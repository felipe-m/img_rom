------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : fondo_space_inv_512_384.ppm 
--- Filas    : 384 
--- Columnas : 512 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_fondo_space_inv_512_384 is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(18-1 downto 0);
    dout : out std_logic_vector(9-1 downto 0) 
  );
end ROM_RGB_9b_fondo_space_inv_512_384;


architecture BEHAVIORAL of ROM_RGB_9b_fondo_space_inv_512_384 is
  signal addr_int  : natural range 0 to 2**18-1;
  type memostruct is array (natural range<>) of std_logic_vector(9-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBBB"
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "011010100",
       "010011100",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010100100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110101",
       "001100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "001101101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001110110",
       "010100100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000110110",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "001101101",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001110110",
       "010100100",
       "011010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "010100100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "001011100",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001110101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "010100101",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010011100",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "001100100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "000110110",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "001100100",
       "001101101",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010100100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "010100101",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "001111110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001101101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110101",
       "010011100",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010100",
       "010011100",
       "001110101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010100100",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001110101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010100100",
       "011010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010011100",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010100100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010100",
       "010100100",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001011100",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "010100100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100100",
       "001110101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010100",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "000101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010100101",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "001011100",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010100101",
       "000111111",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000110101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010100100",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010100100",
       "001100101",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "001110110",
       "000111110",
       "000110110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "001110101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010100100",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110101",
       "001100101",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001110101",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001110101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001110101",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001110101",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010100100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110101",
       "001100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "001110101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111000011",
       "110001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "001011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001110101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010100100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "000110110",
       "000111110",
       "000111111",
       "000111110",
       "000111110",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010010100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "001100100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "110001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010100101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010100",
       "010011100",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "001001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010100100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "100001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "100001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "110001011",
       "111000011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "101001011",
       "101001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "001011100",
       "001011100",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "110001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010100100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001110110",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "101001011",
       "101001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001110101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "011001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100001011",
       "001001011",
       "010001011",
       "001001011",
       "010001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111000011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001110110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110101",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "001100101",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111000011",
       "111000011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "011001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010100101",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010100101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001110101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101000011",
       "010010011",
       "001001011",
       "010001011",
       "001001011",
       "100001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "011001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "101001011",
       "101001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "001110101",
       "001110101",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "101000011",
       "001010011",
       "010001011",
       "010001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111001011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "000110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "110000011",
       "111000011",
       "101000011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "001011100",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010100100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "001010011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001111110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "011010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111001011",
       "111001011",
       "011001011",
       "001001011",
       "100001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111000011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "001100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "010100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "011001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "100001011",
       "001010011",
       "010001011",
       "010001011",
       "001010011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "111001011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100100",
       "001110101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "001010011",
       "100001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "001001011",
       "001001011",
       "001001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "110001011",
       "110001011",
       "110001011",
       "010001011",
       "010001011",
       "011001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010100100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111000011",
       "111000011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "011010100",
       "001100101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "100001011",
       "001010011",
       "010001011",
       "010001011",
       "001010011",
       "011001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "000110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001101101",
       "010010100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "101001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100001011",
       "001001011",
       "010001011",
       "001001011",
       "010001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "001001011",
       "010001011",
       "001001011",
       "011001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100001011",
       "011001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "011010100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "101000011",
       "001010011",
       "101001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "011011100",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010010011",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010010011",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "011001011",
       "001010011",
       "010001011",
       "010001011",
       "011001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "001001011",
       "010001011",
       "001001011",
       "100001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111000011",
       "110001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "001100101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "110001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "110001011",
       "011001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "110001011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000101101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011011100",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111000011",
       "111000011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111110",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110001011",
       "001001011",
       "010001011",
       "010001011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "100001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111000011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "000110110",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "001010011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "101001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "100001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "010010100",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "110000011",
       "110000011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "001110101",
       "000111111",
       "000111110",
       "000111110",
       "001100100",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011011100",
       "001100101",
       "000111111",
       "000111110",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "100001011",
       "001010011",
       "010001011",
       "010001011",
       "001010011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "001010011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100001011",
       "001001011",
       "010001011",
       "001001011",
       "010001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "001001011",
       "010001011",
       "001001011",
       "011001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100001011",
       "011001011",
       "010001011",
       "010001011",
       "001010011",
       "100001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011011100",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "011001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "010010100",
       "010001011",
       "010001011",
       "001010011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "001101101",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "011001011",
       "010001011",
       "010001011",
       "001010011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101001011",
       "001001011",
       "010001011",
       "001001011",
       "010001011",
       "011001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "010010011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "011001011",
       "001010011",
       "011001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100001011",
       "011001011",
       "001001011",
       "010001011",
       "001001011",
       "100001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100001011",
       "010001011",
       "001001011",
       "010001011",
       "001001011",
       "100001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "101000011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "011001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010100100",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111000011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "101000011",
       "001010011",
       "010001011",
       "010001011",
       "011001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110001011",
       "100001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "011001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "101000011",
       "001010011",
       "010001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100001011",
       "001010011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100100",
       "000111111",
       "000111111",
       "000111111",
       "010100101",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "110000011",
       "110000011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "011001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100100",
       "000111110",
       "000111111",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011011100",
       "000110110",
       "000111111",
       "000111110",
       "000111111",
       "010011100",
       "010001011",
       "010001011",
       "001001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "100001011",
       "010001011",
       "010001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010010100",
       "001111110",
       "000111111",
       "000111111",
       "000111110",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "110000011",
       "111000011",
       "101001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "001110101",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011010100",
       "001110110",
       "000111111",
       "000111111",
       "001110110",
       "010010011",
       "010001011",
       "010001011",
       "001001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "011001011",
       "001010011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "001100101",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "001100100",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "101001011",
       "001001011",
       "010001011",
       "001001011",
       "010001011",
       "011001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "100001011",
       "001001011",
       "010001011",
       "001001011",
       "010001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "001100100",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "010001011",
       "001001011",
       "010001011",
       "001010011",
       "100001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "110001011",
       "111000011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100100",
       "011010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "001100100",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "011001011",
       "001010011",
       "010001011",
       "100001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "101000011",
       "001010011",
       "101001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010100100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "001100101",
       "000111111",
       "000111110",
       "000111111",
       "001100100",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "011001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "001100100",
       "010001011",
       "010001011",
       "001001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001100100",
       "000111111",
       "000111110",
       "000111111",
       "001100101",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "001111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010100100",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011010100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "010010011",
       "010001011",
       "010001011",
       "001001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010100100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011011100",
       "000110110",
       "000111111",
       "000111110",
       "000111111",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "001100101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "010100100",
       "010011100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "010100100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "001100100",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010011100",
       "001110101",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "001101101",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010010100",
       "010100100",
       "000111111",
       "000111110",
       "000111111",
       "000110110",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "100001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010010011",
       "001110110",
       "000111111",
       "000111110",
       "000111111",
       "001100101",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010100100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010100100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "011001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "001110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "010100101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "010001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010100101",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "100001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001100100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "110001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "000111110",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001100100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "101001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100100",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "000110110",
       "010100100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011011100",
       "001100100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "100001011",
       "110001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100001011",
       "011001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001011100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011011100",
       "001011100",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "010001011",
       "011001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001101101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "000110110",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001100101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "001110110",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "100010011",
       "101010100",
       "011010011",
       "011010011",
       "010010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "011010100",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010011100",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011010100",
       "010011100",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "001100100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "001100100",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "001101101",
       "001101101",
       "010100100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100100",
       "001101101",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "100010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "011010011",
       "101010100",
       "010010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "010011100",
       "001110101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001110110",
       "001110110",
       "001110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "110001011",
       "110001011",
       "110001011",
       "110001011",
       "101001011",
       "110001011",
       "101010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "010011100",
       "001101101",
       "001110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "001101101",
       "001100100",
       "010011100",
       "011010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "110001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "011010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010011100",
       "010011100",
       "001100101",
       "001101101",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "001101101",
       "001101101",
       "010100100",
       "010011100",
       "010011100",
       "011010011",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010100101",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "101010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "011010011",
       "101010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "001101101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "001101101",
       "001101101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "010100100",
       "010100100",
       "010100100",
       "010100100",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110001011",
       "101010011",
       "110001011",
       "100001011",
       "101001011",
       "101010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "001100101",
       "001101101",
       "001110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001101101",
       "001101101",
       "001100100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "101001011",
       "110001011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "101010100",
       "100010011",
       "010010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010100",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011011",
       "010010011",
       "010010100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "001101101",
       "001110101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "001100100",
       "010011100",
       "011011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "011010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "001110101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "001110110",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "101010011",
       "011001011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "001101101",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001110110",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110001011",
       "100001011",
       "110001011",
       "011010011",
       "011010011",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "101010100",
       "011010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001100101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101110",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "101001011",
       "101001011",
       "100001011",
       "011010011",
       "100010100",
       "100010011",
       "011010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001100100",
       "001110110",
       "000111110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010101101",
       "011100101",
       "010100101",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001100101",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010101101",
       "011100101",
       "010100101",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "011001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "101010011",
       "010010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101110",
       "011100101",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "101001011",
       "101001011",
       "101001011",
       "010010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "011100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110001011",
       "100001011",
       "011010011",
       "100010011",
       "011010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "011010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101110",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "011010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001101101",
       "000111110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010101101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "110001011",
       "100001011",
       "011010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001100101",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "110001011",
       "011001011",
       "100010100",
       "011010011",
       "100010011",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001100101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "110001011",
       "110001011",
       "100010011",
       "011010011",
       "011010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "100010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "110001011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001100101",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "101001011",
       "011001011",
       "010010011",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100001011",
       "101010011",
       "100010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001101101",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110001011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "011001011",
       "100010011",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001100101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100001011",
       "100010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001101101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "110000011",
       "110000011",
       "110000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "110001011",
       "100010100",
       "011010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001101101",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "100001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101010011",
       "100010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010100100",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011011100",
       "010100101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "011010011",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010100101",
       "011100101",
       "001101110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "001110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "001110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "100001011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010100100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "001110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "001110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000111110",
       "010101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "001101110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100100",
       "010100101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "010101101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "011010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001101101",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "001101101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001101101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001110101",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "001101101",
       "001110110",
       "001100100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "001100101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "001110110",
       "000111111",
       "000111110",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "011001011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100101",
       "010100101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101110",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000110110",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010100100",
       "010100101",
       "010100101",
       "011100101",
       "001101101",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001110110",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010101101",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010101101",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010101101",
       "001110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "010100100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "101001011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "001101110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "010010011",
       "100010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "001101101",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "001101101",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "010101101",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "001101101",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "101001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "001101101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "001101101",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "001101101",
       "001110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "001101101",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001101101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "001110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "000110110",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111110",
       "000110110",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "001101101",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010010100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "001101101",
       "000110110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "001101110",
       "010101101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "001101101",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "001100100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "010101101",
       "001101101",
       "000110110",
       "000110101",
       "000110110",
       "000111110",
       "000111110",
       "000110110",
       "000110101",
       "000110110",
       "000110110",
       "001101101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010101101",
       "000110110",
       "000111110",
       "000111110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "001101101",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "001101101",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "001110101",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "011100101",
       "011100101",
       "011100101",
       "011100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "001101101",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000110110",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010100101",
       "001110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111111",
       "000110110",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "001101110",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "001101101",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000110110",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "010101101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111110",
       "010100101",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "011010011",
       "100010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010101101",
       "001101110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "001110110",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101001011",
       "011010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010101101",
       "001110110",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000110110",
       "001100101",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110001011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010010011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "010100101",
       "010101101",
       "000110110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111111",
       "000111111",
       "000111111",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000110110",
       "001101101",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010010011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "010100101",
       "011100101",
       "011100101",
       "010101101",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000110110",
       "001101101",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010100101",
       "010100100",
       "010100101",
       "010100101",
       "010100101",
       "001101110",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000110110",
       "000111110",
       "000111110",
       "000110110",
       "000110110",
       "000110110",
       "001101101",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "011010011",
       "011010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011011",
       "001100101",
       "001101101",
       "001101101",
       "000110110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000111110",
       "000110110",
       "001101101",
       "001101101",
       "001101101",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "001100101",
       "001101101",
       "001100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "011011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "110101100",
       "110100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "110101100",
       "110100100",
       "101100100",
       "101011100",
       "100011100",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "101001011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "011010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "011011011",
       "101011100",
       "110100100",
       "110100100",
       "110101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "110101100",
       "110100100",
       "101011100",
       "011011100",
       "011011100",
       "011011100",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "011010011",
       "011011100",
       "100011100",
       "110101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "110100100",
       "100011011",
       "011011100",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "011010011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "100011011",
       "100011100",
       "100100100",
       "110101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "110101100",
       "100011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "011010011",
       "101010100",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "011011100",
       "101011100",
       "110101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "101100100",
       "101011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "101100100",
       "011011100",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "101100100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "101011100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "101100100",
       "011011100",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "101100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "101100100",
       "110011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "101100100",
       "110100100",
       "110100100",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100100100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "100010100",
       "100010011",
       "100010011",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "101100100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100100100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101011100",
       "101011100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "100100100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100011100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "110000011",
       "110000011",
       "110000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100011100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110100100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100011100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "100011100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "100011100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010011100",
       "100100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "100010100",
       "100100100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "110100100",
       "111101100",
       "110101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110100100",
       "010010100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "101100100",
       "110100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "110100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101001011",
       "100010011",
       "100010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "110101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011010100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "011011011",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111001011",
       "110001011",
       "111001011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "011001011",
       "101001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "011001011",
       "011001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "011001011",
       "100000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "110000011",
       "110000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "110100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "011001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010001011",
       "110000011",
       "110000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "011001011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "100001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "100011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "011001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "110000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001001011",
       "100001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "100001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "100001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "100001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "110101100",
       "111101100",
       "111101100",
       "110101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "110101100",
       "110101100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "110101100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "110011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "110000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "100001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "100001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "100001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "101000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "011001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "100011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "110001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "011001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "100001011",
       "001001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "110101100",
       "110100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111001011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "101000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "101000011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "110001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "101000011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "110000011",
       "101001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "010001011",
       "011001011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "100001011",
       "011001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "001010011",
       "011001011",
       "111000011",
       "110000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "110000011",
       "111000011",
       "011001011",
       "001010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "011011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "101001011",
       "110000011",
       "101000011",
       "101000011",
       "101000011",
       "101000011",
       "101000011",
       "110000011",
       "110001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100011",
       "010010100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010010100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "110101100",
       "110101100",
       "110100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "110100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "100100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110100100",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110101100",
       "011011011",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "011011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "101011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110100100",
       "010010011",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110100100",
       "010010011",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "110100100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111101100",
       "011011100",
       "010010100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "110101100",
       "011011100",
       "010010100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "100011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111101100",
       "101011100",
       "010010100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "110101100",
       "100011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "101100100",
       "010010100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "101100100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111110100",
       "111110100",
       "111110100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110100100",
       "101011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110100100",
       "011011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "101100100",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110100100",
       "011011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "100011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "101100100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "101100100",
       "011011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "110100100",
       "101011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "101100100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110101100",
       "110100100",
       "100011011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101011100",
       "101100100",
       "110100100",
       "110100100",
       "110100100",
       "110100100",
       "101100100",
       "101100100",
       "110100100",
       "110100100",
       "110100100",
       "110100100",
       "110100100",
       "110100100",
       "101100100",
       "110100100",
       "101100100",
       "100100100",
       "101100100",
       "100011100",
       "010011100",
       "010011100",
       "101100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110100100",
       "101011100",
       "101011100",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101011100",
       "101011100",
       "101011100",
       "101010100",
       "101011100",
       "101011100",
       "100011100",
       "100011100",
       "100011100",
       "100011100",
       "100011100",
       "101100100",
       "100011100",
       "100011100",
       "100011100",
       "100011100",
       "100011100",
       "100011100",
       "100011100",
       "100100100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "110100100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "110100100",
       "101011100",
       "101010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "110101100",
       "111101100",
       "111101100",
       "110100100",
       "101011100",
       "101011100",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011011100",
       "101011100",
       "101011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "011010100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010100",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100010100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010100",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "100010011",
       "100010011",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "011010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "111001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "110000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "101010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "101010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111000011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111001011",
       "111000011",
       "110001011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "100010011",
       "011010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010011100",
       "010011100",
       "010011100",
       "010010011",
       "010001011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010010011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011",
       "010001011"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

