---   Background Pattern table COLOR PLANE 1
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: nova_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_NOVA_BG_PLN1 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_NOVA_BG_PLN1;

architecture BEHAVIORAL of ROM_PTABLE_NOVA_BG_PLN1 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table COLOR PLANE 1
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Background 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000011", --    2 -  0x2  :    3 - 0x3
    "00000001", --    3 -  0x3  :    1 - 0x1
    "00000001", --    4 -  0x4  :    1 - 0x1
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000011", --    6 -  0x6  :    3 - 0x3
    "00000001", --    7 -  0x7  :    1 - 0x1
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Background 0x1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00111000", --   10 -  0xa  :   56 - 0x38
    "10110100", --   11 -  0xb  :  180 - 0xb4
    "10101000", --   12 -  0xc  :  168 - 0xa8
    "11010100", --   13 -  0xd  :  212 - 0xd4
    "01110100", --   14 -  0xe  :  116 - 0x74
    "01111110", --   15 -  0xf  :  126 - 0x7e
    "00111000", --   16 - 0x10  :   56 - 0x38 -- Background 0x2
    "01111000", --   17 - 0x11  :  120 - 0x78
    "01111100", --   18 - 0x12  :  124 - 0x7c
    "01111110", --   19 - 0x13  :  126 - 0x7e
    "01111110", --   20 - 0x14  :  126 - 0x7e
    "01111110", --   21 - 0x15  :  126 - 0x7e
    "00111110", --   22 - 0x16  :   62 - 0x3e
    "00011110", --   23 - 0x17  :   30 - 0x1e
    "11110110", --   24 - 0x18  :  246 - 0xf6 -- Background 0x3
    "11110000", --   25 - 0x19  :  240 - 0xf0
    "00111000", --   26 - 0x1a  :   56 - 0x38
    "11010000", --   27 - 0x1b  :  208 - 0xd0
    "11100000", --   28 - 0x1c  :  224 - 0xe0
    "01110000", --   29 - 0x1d  :  112 - 0x70
    "10111000", --   30 - 0x1e  :  184 - 0xb8
    "01000000", --   31 - 0x1f  :   64 - 0x40
    "00011100", --   32 - 0x20  :   28 - 0x1c -- Background 0x4
    "00011100", --   33 - 0x21  :   28 - 0x1c
    "00011110", --   34 - 0x22  :   30 - 0x1e
    "00011111", --   35 - 0x23  :   31 - 0x1f
    "00001100", --   36 - 0x24  :   12 - 0xc
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "10101000", --   40 - 0x28  :  168 - 0xa8 -- Background 0x5
    "01010000", --   41 - 0x29  :   80 - 0x50
    "10101000", --   42 - 0x2a  :  168 - 0xa8
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "01100000", --   44 - 0x2c  :   96 - 0x60
    "01100000", --   45 - 0x2d  :   96 - 0x60
    "01110000", --   46 - 0x2e  :  112 - 0x70
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00011100", --   48 - 0x30  :   28 - 0x1c -- Background 0x6
    "00011100", --   49 - 0x31  :   28 - 0x1c
    "00011110", --   50 - 0x32  :   30 - 0x1e
    "00011111", --   51 - 0x33  :   31 - 0x1f
    "00001100", --   52 - 0x34  :   12 - 0xc
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000001", --   54 - 0x36  :    1 - 0x1
    "00000000", --   55 - 0x37  :    0 - 0x0
    "10101000", --   56 - 0x38  :  168 - 0xa8 -- Background 0x7
    "01010000", --   57 - 0x39  :   80 - 0x50
    "10101000", --   58 - 0x3a  :  168 - 0xa8
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "01011000", --   60 - 0x3c  :   88 - 0x58
    "11011000", --   61 - 0x3d  :  216 - 0xd8
    "10001100", --   62 - 0x3e  :  140 - 0x8c
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00011100", --   64 - 0x40  :   28 - 0x1c -- Background 0x8
    "00011100", --   65 - 0x41  :   28 - 0x1c
    "00011110", --   66 - 0x42  :   30 - 0x1e
    "00011111", --   67 - 0x43  :   31 - 0x1f
    "00001100", --   68 - 0x44  :   12 - 0xc
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "10101000", --   72 - 0x48  :  168 - 0xa8 -- Background 0x9
    "01010100", --   73 - 0x49  :   84 - 0x54
    "10101000", --   74 - 0x4a  :  168 - 0xa8
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "01101110", --   76 - 0x4c  :  110 - 0x6e
    "11000000", --   77 - 0x4d  :  192 - 0xc0
    "10000000", --   78 - 0x4e  :  128 - 0x80
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00011100", --   80 - 0x50  :   28 - 0x1c -- Background 0xa
    "00011100", --   81 - 0x51  :   28 - 0x1c
    "00011110", --   82 - 0x52  :   30 - 0x1e
    "00011111", --   83 - 0x53  :   31 - 0x1f
    "00001100", --   84 - 0x54  :   12 - 0xc
    "00000001", --   85 - 0x55  :    1 - 0x1
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "10101000", --   88 - 0x58  :  168 - 0xa8 -- Background 0xb
    "01010100", --   89 - 0x59  :   84 - 0x54
    "10101000", --   90 - 0x5a  :  168 - 0xa8
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "11011000", --   92 - 0x5c  :  216 - 0xd8
    "11011100", --   93 - 0x5d  :  220 - 0xdc
    "00001100", --   94 - 0x5e  :   12 - 0xc
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "11110110", --   96 - 0x60  :  246 - 0xf6 -- Background 0xc
    "11110000", --   97 - 0x61  :  240 - 0xf0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "11111100", --   99 - 0x63  :  252 - 0xfc
    "11111000", --  100 - 0x64  :  248 - 0xf8
    "00000000", --  101 - 0x65  :    0 - 0x0
    "10101000", --  102 - 0x66  :  168 - 0xa8
    "01010100", --  103 - 0x67  :   84 - 0x54
    "00111000", --  104 - 0x68  :   56 - 0x38 -- Background 0xd
    "01111000", --  105 - 0x69  :  120 - 0x78
    "01111100", --  106 - 0x6a  :  124 - 0x7c
    "01111101", --  107 - 0x6b  :  125 - 0x7d
    "01111101", --  108 - 0x6c  :  125 - 0x7d
    "01111011", --  109 - 0x6d  :  123 - 0x7b
    "00111011", --  110 - 0x6e  :   59 - 0x3b
    "00011011", --  111 - 0x6f  :   27 - 0x1b
    "11110110", --  112 - 0x70  :  246 - 0xf6 -- Background 0xe
    "11110000", --  113 - 0x71  :  240 - 0xf0
    "01111000", --  114 - 0x72  :  120 - 0x78
    "01110000", --  115 - 0x73  :  112 - 0x70
    "10100000", --  116 - 0x74  :  160 - 0xa0
    "10010000", --  117 - 0x75  :  144 - 0x90
    "00101000", --  118 - 0x76  :   40 - 0x28
    "01010100", --  119 - 0x77  :   84 - 0x54
    "00000000", --  120 - 0x78  :    0 - 0x0 -- Background 0xf
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000011", --  122 - 0x7a  :    3 - 0x3
    "00000001", --  123 - 0x7b  :    1 - 0x1
    "00000001", --  124 - 0x7c  :    1 - 0x1
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000011", --  126 - 0x7e  :    3 - 0x3
    "00000001", --  127 - 0x7f  :    1 - 0x1
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Background 0x10
    "00000011", --  129 - 0x81  :    3 - 0x3
    "00001111", --  130 - 0x82  :   15 - 0xf
    "00001111", --  131 - 0x83  :   15 - 0xf
    "00001111", --  132 - 0x84  :   15 - 0xf
    "00011111", --  133 - 0x85  :   31 - 0x1f
    "00011111", --  134 - 0x86  :   31 - 0x1f
    "00011110", --  135 - 0x87  :   30 - 0x1e
    "00110110", --  136 - 0x88  :   54 - 0x36 -- Background 0x11
    "10110000", --  137 - 0x89  :  176 - 0xb0
    "10111000", --  138 - 0x8a  :  184 - 0xb8
    "10010000", --  139 - 0x8b  :  144 - 0x90
    "10100000", --  140 - 0x8c  :  160 - 0xa0
    "01110000", --  141 - 0x8d  :  112 - 0x70
    "00111000", --  142 - 0x8e  :   56 - 0x38
    "01000000", --  143 - 0x8f  :   64 - 0x40
    "00011100", --  144 - 0x90  :   28 - 0x1c -- Background 0x12
    "00011100", --  145 - 0x91  :   28 - 0x1c
    "00011110", --  146 - 0x92  :   30 - 0x1e
    "00011111", --  147 - 0x93  :   31 - 0x1f
    "00001100", --  148 - 0x94  :   12 - 0xc
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- Background 0x13
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000011", --  155 - 0x9b  :    3 - 0x3
    "00000111", --  156 - 0x9c  :    7 - 0x7
    "00001111", --  157 - 0x9d  :   15 - 0xf
    "00001111", --  158 - 0x9e  :   15 - 0xf
    "00011111", --  159 - 0x9f  :   31 - 0x1f
    "11110110", --  160 - 0xa0  :  246 - 0xf6 -- Background 0x14
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "11111000", --  162 - 0xa2  :  248 - 0xf8
    "11111110", --  163 - 0xa3  :  254 - 0xfe
    "11111110", --  164 - 0xa4  :  254 - 0xfe
    "11111110", --  165 - 0xa5  :  254 - 0xfe
    "11111000", --  166 - 0xa6  :  248 - 0xf8
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000011", --  168 - 0xa8  :    3 - 0x3 -- Background 0x15
    "00000011", --  169 - 0xa9  :    3 - 0x3
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000011", --  171 - 0xab  :    3 - 0x3
    "00000011", --  172 - 0xac  :    3 - 0x3
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00001111", --  174 - 0xae  :   15 - 0xf
    "00111111", --  175 - 0xaf  :   63 - 0x3f
    "11011000", --  176 - 0xb0  :  216 - 0xd8 -- Background 0x16
    "11000000", --  177 - 0xb1  :  192 - 0xc0
    "11100000", --  178 - 0xb2  :  224 - 0xe0
    "01000000", --  179 - 0xb3  :   64 - 0x40
    "10000000", --  180 - 0xb4  :  128 - 0x80
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "11100000", --  182 - 0xb6  :  224 - 0xe0
    "11111100", --  183 - 0xb7  :  252 - 0xfc
    "01111111", --  184 - 0xb8  :  127 - 0x7f -- Background 0x17
    "01111111", --  185 - 0xb9  :  127 - 0x7f
    "01111111", --  186 - 0xba  :  127 - 0x7f
    "01111100", --  187 - 0xbb  :  124 - 0x7c
    "00110000", --  188 - 0xbc  :   48 - 0x30
    "00000001", --  189 - 0xbd  :    1 - 0x1
    "00000001", --  190 - 0xbe  :    1 - 0x1
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "11111100", --  192 - 0xc0  :  252 - 0xfc -- Background 0x18
    "11111110", --  193 - 0xc1  :  254 - 0xfe
    "11111100", --  194 - 0xc2  :  252 - 0xfc
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00000000", --  196 - 0xc4  :    0 - 0x0
    "10000000", --  197 - 0xc5  :  128 - 0x80
    "11000000", --  198 - 0xc6  :  192 - 0xc0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000111", --  200 - 0xc8  :    7 - 0x7 -- Background 0x19
    "00000111", --  201 - 0xc9  :    7 - 0x7
    "00000001", --  202 - 0xca  :    1 - 0x1
    "00000110", --  203 - 0xcb  :    6 - 0x6
    "00000111", --  204 - 0xcc  :    7 - 0x7
    "00000110", --  205 - 0xcd  :    6 - 0x6
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00001111", --  207 - 0xcf  :   15 - 0xf
    "10110000", --  208 - 0xd0  :  176 - 0xb0 -- Background 0x1a
    "10000000", --  209 - 0xd1  :  128 - 0x80
    "11000000", --  210 - 0xd2  :  192 - 0xc0
    "10000000", --  211 - 0xd3  :  128 - 0x80
    "00000000", --  212 - 0xd4  :    0 - 0x0
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "11100000", --  215 - 0xd7  :  224 - 0xe0
    "00111111", --  216 - 0xd8  :   63 - 0x3f -- Background 0x1b
    "00111111", --  217 - 0xd9  :   63 - 0x3f
    "01111111", --  218 - 0xda  :  127 - 0x7f
    "01111111", --  219 - 0xdb  :  127 - 0x7f
    "00111111", --  220 - 0xdc  :   63 - 0x3f
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000011", --  222 - 0xde  :    3 - 0x3
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "11111111", --  224 - 0xe0  :  255 - 0xff -- Background 0x1c
    "11111111", --  225 - 0xe1  :  255 - 0xff
    "11111111", --  226 - 0xe2  :  255 - 0xff
    "11111111", --  227 - 0xe3  :  255 - 0xff
    "11111111", --  228 - 0xe4  :  255 - 0xff
    "00000000", --  229 - 0xe5  :    0 - 0x0
    "10000000", --  230 - 0xe6  :  128 - 0x80
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- Background 0x1d
    "11000000", --  233 - 0xe9  :  192 - 0xc0
    "11000000", --  234 - 0xea  :  192 - 0xc0
    "11000000", --  235 - 0xeb  :  192 - 0xc0
    "10000000", --  236 - 0xec  :  128 - 0x80
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "11100000", --  240 - 0xf0  :  224 - 0xe0 -- Background 0x1e
    "10011100", --  241 - 0xf1  :  156 - 0x9c
    "00111000", --  242 - 0xf2  :   56 - 0x38
    "11100000", --  243 - 0xf3  :  224 - 0xe0
    "11001000", --  244 - 0xf4  :  200 - 0xc8
    "00010100", --  245 - 0xf5  :   20 - 0x14
    "10101000", --  246 - 0xf6  :  168 - 0xa8
    "01010100", --  247 - 0xf7  :   84 - 0x54
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- Background 0x1f
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00111000", --  250 - 0xfa  :   56 - 0x38
    "10110100", --  251 - 0xfb  :  180 - 0xb4
    "10101000", --  252 - 0xfc  :  168 - 0xa8
    "11010100", --  253 - 0xfd  :  212 - 0xd4
    "01110100", --  254 - 0xfe  :  116 - 0x74
    "00011110", --  255 - 0xff  :   30 - 0x1e
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Background 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00001100", --  258 - 0x102  :   12 - 0xc
    "00000111", --  259 - 0x103  :    7 - 0x7
    "00001111", --  260 - 0x104  :   15 - 0xf
    "00000111", --  261 - 0x105  :    7 - 0x7
    "00001111", --  262 - 0x106  :   15 - 0xf
    "00001111", --  263 - 0x107  :   15 - 0xf
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Background 0x21
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00110000", --  266 - 0x10a  :   48 - 0x30
    "11100000", --  267 - 0x10b  :  224 - 0xe0
    "11110000", --  268 - 0x10c  :  240 - 0xf0
    "11100000", --  269 - 0x10d  :  224 - 0xe0
    "11110000", --  270 - 0x10e  :  240 - 0xf0
    "11110000", --  271 - 0x10f  :  240 - 0xf0
    "00000111", --  272 - 0x110  :    7 - 0x7 -- Background 0x22
    "00000011", --  273 - 0x111  :    3 - 0x3
    "00011000", --  274 - 0x112  :   24 - 0x18
    "00010101", --  275 - 0x113  :   21 - 0x15
    "00000010", --  276 - 0x114  :    2 - 0x2
    "00000101", --  277 - 0x115  :    5 - 0x5
    "00000010", --  278 - 0x116  :    2 - 0x2
    "00000100", --  279 - 0x117  :    4 - 0x4
    "11100000", --  280 - 0x118  :  224 - 0xe0 -- Background 0x23
    "11000000", --  281 - 0x119  :  192 - 0xc0
    "00111100", --  282 - 0x11a  :   60 - 0x3c
    "01111100", --  283 - 0x11b  :  124 - 0x7c
    "01111100", --  284 - 0x11c  :  124 - 0x7c
    "01111100", --  285 - 0x11d  :  124 - 0x7c
    "11101100", --  286 - 0x11e  :  236 - 0xec
    "11100000", --  287 - 0x11f  :  224 - 0xe0
    "00000010", --  288 - 0x120  :    2 - 0x2 -- Background 0x24
    "00000101", --  289 - 0x121  :    5 - 0x5
    "00001011", --  290 - 0x122  :   11 - 0xb
    "00001011", --  291 - 0x123  :   11 - 0xb
    "00001101", --  292 - 0x124  :   13 - 0xd
    "00011000", --  293 - 0x125  :   24 - 0x18
    "00111000", --  294 - 0x126  :   56 - 0x38
    "00000000", --  295 - 0x127  :    0 - 0x0
    "11100000", --  296 - 0x128  :  224 - 0xe0 -- Background 0x25
    "11100000", --  297 - 0x129  :  224 - 0xe0
    "11100000", --  298 - 0x12a  :  224 - 0xe0
    "11010000", --  299 - 0x12b  :  208 - 0xd0
    "10111000", --  300 - 0x12c  :  184 - 0xb8
    "00111000", --  301 - 0x12d  :   56 - 0x38
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Background 0x26
    "00000000", --  305 - 0x131  :    0 - 0x0
    "00000000", --  306 - 0x132  :    0 - 0x0
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "00000000", --  309 - 0x135  :    0 - 0x0
    "00000000", --  310 - 0x136  :    0 - 0x0
    "00000000", --  311 - 0x137  :    0 - 0x0
    "00000000", --  312 - 0x138  :    0 - 0x0 -- Background 0x27
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Background 0x28
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "00000000", --  324 - 0x144  :    0 - 0x0
    "00000000", --  325 - 0x145  :    0 - 0x0
    "00000000", --  326 - 0x146  :    0 - 0x0
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00011111", --  328 - 0x148  :   31 - 0x1f -- Background 0x29
    "00011111", --  329 - 0x149  :   31 - 0x1f
    "00011111", --  330 - 0x14a  :   31 - 0x1f
    "00011111", --  331 - 0x14b  :   31 - 0x1f
    "00001100", --  332 - 0x14c  :   12 - 0xc
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000001", --  334 - 0x14e  :    1 - 0x1
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00011111", --  336 - 0x150  :   31 - 0x1f -- Background 0x2a
    "00011111", --  337 - 0x151  :   31 - 0x1f
    "00011111", --  338 - 0x152  :   31 - 0x1f
    "00011111", --  339 - 0x153  :   31 - 0x1f
    "00001100", --  340 - 0x154  :   12 - 0xc
    "00000000", --  341 - 0x155  :    0 - 0x0
    "00000000", --  342 - 0x156  :    0 - 0x0
    "00000000", --  343 - 0x157  :    0 - 0x0
    "00000000", --  344 - 0x158  :    0 - 0x0 -- Background 0x2b
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Background 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0 -- Background 0x2d
    "01111110", --  361 - 0x169  :  126 - 0x7e
    "01000010", --  362 - 0x16a  :   66 - 0x42
    "01000010", --  363 - 0x16b  :   66 - 0x42
    "01000010", --  364 - 0x16c  :   66 - 0x42
    "01000010", --  365 - 0x16d  :   66 - 0x42
    "01111110", --  366 - 0x16e  :  126 - 0x7e
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Background 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "01100110", --  376 - 0x178  :  102 - 0x66 -- Background 0x2f
    "01100000", --  377 - 0x179  :   96 - 0x60
    "01101000", --  378 - 0x17a  :  104 - 0x68
    "11100000", --  379 - 0x17b  :  224 - 0xe0
    "11000000", --  380 - 0x17c  :  192 - 0xc0
    "00010000", --  381 - 0x17d  :   16 - 0x10
    "00101000", --  382 - 0x17e  :   40 - 0x28
    "01010000", --  383 - 0x17f  :   80 - 0x50
    "11110110", --  384 - 0x180  :  246 - 0xf6 -- Background 0x30
    "11110000", --  385 - 0x181  :  240 - 0xf0
    "00111000", --  386 - 0x182  :   56 - 0x38
    "11010000", --  387 - 0x183  :  208 - 0xd0
    "11000000", --  388 - 0x184  :  192 - 0xc0
    "11111000", --  389 - 0x185  :  248 - 0xf8
    "01111000", --  390 - 0x186  :  120 - 0x78
    "00000000", --  391 - 0x187  :    0 - 0x0
    "11110110", --  392 - 0x188  :  246 - 0xf6 -- Background 0x31
    "11110000", --  393 - 0x189  :  240 - 0xf0
    "00111000", --  394 - 0x18a  :   56 - 0x38
    "11010000", --  395 - 0x18b  :  208 - 0xd0
    "11000000", --  396 - 0x18c  :  192 - 0xc0
    "11100000", --  397 - 0x18d  :  224 - 0xe0
    "01111000", --  398 - 0x18e  :  120 - 0x78
    "00111000", --  399 - 0x18f  :   56 - 0x38
    "11110110", --  400 - 0x190  :  246 - 0xf6 -- Background 0x32
    "11110000", --  401 - 0x191  :  240 - 0xf0
    "00111000", --  402 - 0x192  :   56 - 0x38
    "11000000", --  403 - 0x193  :  192 - 0xc0
    "11011000", --  404 - 0x194  :  216 - 0xd8
    "11111000", --  405 - 0x195  :  248 - 0xf8
    "01100000", --  406 - 0x196  :   96 - 0x60
    "00010000", --  407 - 0x197  :   16 - 0x10
    "00011100", --  408 - 0x198  :   28 - 0x1c -- Background 0x33
    "00011100", --  409 - 0x199  :   28 - 0x1c
    "00011110", --  410 - 0x19a  :   30 - 0x1e
    "00011111", --  411 - 0x19b  :   31 - 0x1f
    "00001100", --  412 - 0x19c  :   12 - 0xc
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "10000000", --  416 - 0x1a0  :  128 - 0x80 -- Background 0x34
    "01010000", --  417 - 0x1a1  :   80 - 0x50
    "10101000", --  418 - 0x1a2  :  168 - 0xa8
    "00000000", --  419 - 0x1a3  :    0 - 0x0
    "01011000", --  420 - 0x1a4  :   88 - 0x58
    "11011000", --  421 - 0x1a5  :  216 - 0xd8
    "11101100", --  422 - 0x1a6  :  236 - 0xec
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "00011100", --  424 - 0x1a8  :   28 - 0x1c -- Background 0x35
    "00011100", --  425 - 0x1a9  :   28 - 0x1c
    "00011110", --  426 - 0x1aa  :   30 - 0x1e
    "00011111", --  427 - 0x1ab  :   31 - 0x1f
    "00001100", --  428 - 0x1ac  :   12 - 0xc
    "00000001", --  429 - 0x1ad  :    1 - 0x1
    "00000001", --  430 - 0x1ae  :    1 - 0x1
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "10101000", --  432 - 0x1b0  :  168 - 0xa8 -- Background 0x36
    "01010000", --  433 - 0x1b1  :   80 - 0x50
    "10101000", --  434 - 0x1b2  :  168 - 0xa8
    "00000000", --  435 - 0x1b3  :    0 - 0x0
    "01011000", --  436 - 0x1b4  :   88 - 0x58
    "11001110", --  437 - 0x1b5  :  206 - 0xce
    "10000110", --  438 - 0x1b6  :  134 - 0x86
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "10101000", --  440 - 0x1b8  :  168 - 0xa8 -- Background 0x37
    "01010000", --  441 - 0x1b9  :   80 - 0x50
    "10101000", --  442 - 0x1ba  :  168 - 0xa8
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "01011000", --  444 - 0x1bc  :   88 - 0x58
    "11011000", --  445 - 0x1bd  :  216 - 0xd8
    "11101100", --  446 - 0x1be  :  236 - 0xec
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Background 0x38
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "00000000", --  453 - 0x1c5  :    0 - 0x0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- Background 0x39
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Background 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "00000000", --  467 - 0x1d3  :    0 - 0x0
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "00000000", --  469 - 0x1d5  :    0 - 0x0
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Background 0x3b
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Background 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "00000000", --  485 - 0x1e5  :    0 - 0x0
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Background 0x3d
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Background 0x3e
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00000000", --  500 - 0x1f4  :    0 - 0x0
    "00000000", --  501 - 0x1f5  :    0 - 0x0
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- Background 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00111100", --  512 - 0x200  :   60 - 0x3c -- Background 0x40
    "01111100", --  513 - 0x201  :  124 - 0x7c
    "11100110", --  514 - 0x202  :  230 - 0xe6
    "11101110", --  515 - 0x203  :  238 - 0xee
    "11110110", --  516 - 0x204  :  246 - 0xf6
    "11100110", --  517 - 0x205  :  230 - 0xe6
    "00111100", --  518 - 0x206  :   60 - 0x3c
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00111000", --  520 - 0x208  :   56 - 0x38 -- Background 0x41
    "01111000", --  521 - 0x209  :  120 - 0x78
    "00111000", --  522 - 0x20a  :   56 - 0x38
    "00111000", --  523 - 0x20b  :   56 - 0x38
    "00111000", --  524 - 0x20c  :   56 - 0x38
    "00111000", --  525 - 0x20d  :   56 - 0x38
    "00111000", --  526 - 0x20e  :   56 - 0x38
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "01111100", --  528 - 0x210  :  124 - 0x7c -- Background 0x42
    "11111110", --  529 - 0x211  :  254 - 0xfe
    "11100110", --  530 - 0x212  :  230 - 0xe6
    "00011110", --  531 - 0x213  :   30 - 0x1e
    "01111100", --  532 - 0x214  :  124 - 0x7c
    "11100000", --  533 - 0x215  :  224 - 0xe0
    "11111110", --  534 - 0x216  :  254 - 0xfe
    "00000000", --  535 - 0x217  :    0 - 0x0
    "01111100", --  536 - 0x218  :  124 - 0x7c -- Background 0x43
    "11111100", --  537 - 0x219  :  252 - 0xfc
    "11100110", --  538 - 0x21a  :  230 - 0xe6
    "00011100", --  539 - 0x21b  :   28 - 0x1c
    "01100110", --  540 - 0x21c  :  102 - 0x66
    "11101110", --  541 - 0x21d  :  238 - 0xee
    "11111100", --  542 - 0x21e  :  252 - 0xfc
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00001100", --  544 - 0x220  :   12 - 0xc -- Background 0x44
    "00011100", --  545 - 0x221  :   28 - 0x1c
    "00111100", --  546 - 0x222  :   60 - 0x3c
    "01111100", --  547 - 0x223  :  124 - 0x7c
    "11101100", --  548 - 0x224  :  236 - 0xec
    "11111110", --  549 - 0x225  :  254 - 0xfe
    "00001100", --  550 - 0x226  :   12 - 0xc
    "00000000", --  551 - 0x227  :    0 - 0x0
    "11111110", --  552 - 0x228  :  254 - 0xfe -- Background 0x45
    "11111110", --  553 - 0x229  :  254 - 0xfe
    "11100000", --  554 - 0x22a  :  224 - 0xe0
    "11111110", --  555 - 0x22b  :  254 - 0xfe
    "00000110", --  556 - 0x22c  :    6 - 0x6
    "11101110", --  557 - 0x22d  :  238 - 0xee
    "11111100", --  558 - 0x22e  :  252 - 0xfc
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00111100", --  560 - 0x230  :   60 - 0x3c -- Background 0x46
    "01111100", --  561 - 0x231  :  124 - 0x7c
    "11100000", --  562 - 0x232  :  224 - 0xe0
    "11111110", --  563 - 0x233  :  254 - 0xfe
    "11100110", --  564 - 0x234  :  230 - 0xe6
    "11101110", --  565 - 0x235  :  238 - 0xee
    "00111100", --  566 - 0x236  :   60 - 0x3c
    "00000000", --  567 - 0x237  :    0 - 0x0
    "11111110", --  568 - 0x238  :  254 - 0xfe -- Background 0x47
    "11111100", --  569 - 0x239  :  252 - 0xfc
    "00001100", --  570 - 0x23a  :   12 - 0xc
    "00111000", --  571 - 0x23b  :   56 - 0x38
    "00111000", --  572 - 0x23c  :   56 - 0x38
    "01110000", --  573 - 0x23d  :  112 - 0x70
    "01110000", --  574 - 0x23e  :  112 - 0x70
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00111110", --  576 - 0x240  :   62 - 0x3e -- Background 0x48
    "01111100", --  577 - 0x241  :  124 - 0x7c
    "11100110", --  578 - 0x242  :  230 - 0xe6
    "10111100", --  579 - 0x243  :  188 - 0xbc
    "11100110", --  580 - 0x244  :  230 - 0xe6
    "11101110", --  581 - 0x245  :  238 - 0xee
    "00111100", --  582 - 0x246  :   60 - 0x3c
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00111100", --  584 - 0x248  :   60 - 0x3c -- Background 0x49
    "01111100", --  585 - 0x249  :  124 - 0x7c
    "11100110", --  586 - 0x24a  :  230 - 0xe6
    "11101110", --  587 - 0x24b  :  238 - 0xee
    "11111110", --  588 - 0x24c  :  254 - 0xfe
    "10000110", --  589 - 0x24d  :  134 - 0x86
    "01111100", --  590 - 0x24e  :  124 - 0x7c
    "01000000", --  591 - 0x24f  :   64 - 0x40
    "11101110", --  592 - 0x250  :  238 - 0xee -- Background 0x4a
    "11101110", --  593 - 0x251  :  238 - 0xee
    "11101110", --  594 - 0x252  :  238 - 0xee
    "11101110", --  595 - 0x253  :  238 - 0xee
    "11101110", --  596 - 0x254  :  238 - 0xee
    "11101110", --  597 - 0x255  :  238 - 0xee
    "11101110", --  598 - 0x256  :  238 - 0xee
    "10001000", --  599 - 0x257  :  136 - 0x88
    "11100000", --  600 - 0x258  :  224 - 0xe0 -- Background 0x4b
    "11100000", --  601 - 0x259  :  224 - 0xe0
    "11100000", --  602 - 0x25a  :  224 - 0xe0
    "11100000", --  603 - 0x25b  :  224 - 0xe0
    "11100000", --  604 - 0x25c  :  224 - 0xe0
    "11100000", --  605 - 0x25d  :  224 - 0xe0
    "11100000", --  606 - 0x25e  :  224 - 0xe0
    "10000000", --  607 - 0x25f  :  128 - 0x80
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Background 0x4c
    "01111111", --  609 - 0x261  :  127 - 0x7f
    "01111111", --  610 - 0x262  :  127 - 0x7f
    "01111111", --  611 - 0x263  :  127 - 0x7f
    "01111111", --  612 - 0x264  :  127 - 0x7f
    "01111111", --  613 - 0x265  :  127 - 0x7f
    "01111111", --  614 - 0x266  :  127 - 0x7f
    "01111111", --  615 - 0x267  :  127 - 0x7f
    "01111111", --  616 - 0x268  :  127 - 0x7f -- Background 0x4d
    "01111111", --  617 - 0x269  :  127 - 0x7f
    "01111111", --  618 - 0x26a  :  127 - 0x7f
    "01111111", --  619 - 0x26b  :  127 - 0x7f
    "01111111", --  620 - 0x26c  :  127 - 0x7f
    "01111111", --  621 - 0x26d  :  127 - 0x7f
    "01111111", --  622 - 0x26e  :  127 - 0x7f
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Background 0x4e
    "11111110", --  625 - 0x271  :  254 - 0xfe
    "11111110", --  626 - 0x272  :  254 - 0xfe
    "11111110", --  627 - 0x273  :  254 - 0xfe
    "11111110", --  628 - 0x274  :  254 - 0xfe
    "11111110", --  629 - 0x275  :  254 - 0xfe
    "11111110", --  630 - 0x276  :  254 - 0xfe
    "11111110", --  631 - 0x277  :  254 - 0xfe
    "11111110", --  632 - 0x278  :  254 - 0xfe -- Background 0x4f
    "11111110", --  633 - 0x279  :  254 - 0xfe
    "11111110", --  634 - 0x27a  :  254 - 0xfe
    "11111110", --  635 - 0x27b  :  254 - 0xfe
    "11111110", --  636 - 0x27c  :  254 - 0xfe
    "11111110", --  637 - 0x27d  :  254 - 0xfe
    "11111110", --  638 - 0x27e  :  254 - 0xfe
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Background 0x50
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Background 0x51
    "00010000", --  649 - 0x289  :   16 - 0x10
    "00010000", --  650 - 0x28a  :   16 - 0x10
    "01111100", --  651 - 0x28b  :  124 - 0x7c
    "00111000", --  652 - 0x28c  :   56 - 0x38
    "00111000", --  653 - 0x28d  :   56 - 0x38
    "01101100", --  654 - 0x28e  :  108 - 0x6c
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Background 0x52
    "00010000", --  657 - 0x291  :   16 - 0x10
    "00010000", --  658 - 0x292  :   16 - 0x10
    "01111100", --  659 - 0x293  :  124 - 0x7c
    "00111000", --  660 - 0x294  :   56 - 0x38
    "00111000", --  661 - 0x295  :   56 - 0x38
    "01101100", --  662 - 0x296  :  108 - 0x6c
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Background 0x53
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "11111111", --  672 - 0x2a0  :  255 - 0xff -- Background 0x54
    "11111111", --  673 - 0x2a1  :  255 - 0xff
    "11111111", --  674 - 0x2a2  :  255 - 0xff
    "11111111", --  675 - 0x2a3  :  255 - 0xff
    "11111111", --  676 - 0x2a4  :  255 - 0xff
    "11111111", --  677 - 0x2a5  :  255 - 0xff
    "11111111", --  678 - 0x2a6  :  255 - 0xff
    "11111111", --  679 - 0x2a7  :  255 - 0xff
    "11111111", --  680 - 0x2a8  :  255 - 0xff -- Background 0x55
    "11111111", --  681 - 0x2a9  :  255 - 0xff
    "11111111", --  682 - 0x2aa  :  255 - 0xff
    "11111111", --  683 - 0x2ab  :  255 - 0xff
    "11111111", --  684 - 0x2ac  :  255 - 0xff
    "11111111", --  685 - 0x2ad  :  255 - 0xff
    "11111111", --  686 - 0x2ae  :  255 - 0xff
    "11111111", --  687 - 0x2af  :  255 - 0xff
    "00000010", --  688 - 0x2b0  :    2 - 0x2 -- Background 0x56
    "00000101", --  689 - 0x2b1  :    5 - 0x5
    "10101010", --  690 - 0x2b2  :  170 - 0xaa
    "01010001", --  691 - 0x2b3  :   81 - 0x51
    "10101010", --  692 - 0x2b4  :  170 - 0xaa
    "01010001", --  693 - 0x2b5  :   81 - 0x51
    "10100010", --  694 - 0x2b6  :  162 - 0xa2
    "00000100", --  695 - 0x2b7  :    4 - 0x4
    "00001000", --  696 - 0x2b8  :    8 - 0x8 -- Background 0x57
    "01010101", --  697 - 0x2b9  :   85 - 0x55
    "00101010", --  698 - 0x2ba  :   42 - 0x2a
    "01010101", --  699 - 0x2bb  :   85 - 0x55
    "00101010", --  700 - 0x2bc  :   42 - 0x2a
    "01000101", --  701 - 0x2bd  :   69 - 0x45
    "00001010", --  702 - 0x2be  :   10 - 0xa
    "00010000", --  703 - 0x2bf  :   16 - 0x10
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Background 0x58
    "00111111", --  705 - 0x2c1  :   63 - 0x3f
    "01011111", --  706 - 0x2c2  :   95 - 0x5f
    "01101111", --  707 - 0x2c3  :  111 - 0x6f
    "01110000", --  708 - 0x2c4  :  112 - 0x70
    "01110111", --  709 - 0x2c5  :  119 - 0x77
    "01110111", --  710 - 0x2c6  :  119 - 0x77
    "01110111", --  711 - 0x2c7  :  119 - 0x77
    "01110111", --  712 - 0x2c8  :  119 - 0x77 -- Background 0x59
    "01110111", --  713 - 0x2c9  :  119 - 0x77
    "01110111", --  714 - 0x2ca  :  119 - 0x77
    "01110000", --  715 - 0x2cb  :  112 - 0x70
    "01101111", --  716 - 0x2cc  :  111 - 0x6f
    "01011111", --  717 - 0x2cd  :   95 - 0x5f
    "00010101", --  718 - 0x2ce  :   21 - 0x15
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Background 0x5a
    "11111100", --  721 - 0x2d1  :  252 - 0xfc
    "11111000", --  722 - 0x2d2  :  248 - 0xf8
    "11110110", --  723 - 0x2d3  :  246 - 0xf6
    "00001100", --  724 - 0x2d4  :   12 - 0xc
    "11101110", --  725 - 0x2d5  :  238 - 0xee
    "11101100", --  726 - 0x2d6  :  236 - 0xec
    "11101110", --  727 - 0x2d7  :  238 - 0xee
    "11101100", --  728 - 0x2d8  :  236 - 0xec -- Background 0x5b
    "11101110", --  729 - 0x2d9  :  238 - 0xee
    "11101100", --  730 - 0x2da  :  236 - 0xec
    "00001110", --  731 - 0x2db  :   14 - 0xe
    "11110100", --  732 - 0x2dc  :  244 - 0xf4
    "11111010", --  733 - 0x2dd  :  250 - 0xfa
    "01010100", --  734 - 0x2de  :   84 - 0x54
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Background 0x5c
    "00011100", --  737 - 0x2e1  :   28 - 0x1c
    "00111110", --  738 - 0x2e2  :   62 - 0x3e
    "00111110", --  739 - 0x2e3  :   62 - 0x3e
    "00111110", --  740 - 0x2e4  :   62 - 0x3e
    "00011100", --  741 - 0x2e5  :   28 - 0x1c
    "00011100", --  742 - 0x2e6  :   28 - 0x1c
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- Background 0x5d
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Background 0x5e
    "00010100", --  753 - 0x2f1  :   20 - 0x14
    "00110110", --  754 - 0x2f2  :   54 - 0x36
    "00111110", --  755 - 0x2f3  :   62 - 0x3e
    "00111110", --  756 - 0x2f4  :   62 - 0x3e
    "00011100", --  757 - 0x2f5  :   28 - 0x1c
    "00001000", --  758 - 0x2f6  :    8 - 0x8
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- Background 0x5f
    "00010100", --  761 - 0x2f9  :   20 - 0x14
    "00011100", --  762 - 0x2fa  :   28 - 0x1c
    "00011100", --  763 - 0x2fb  :   28 - 0x1c
    "00011100", --  764 - 0x2fc  :   28 - 0x1c
    "00011100", --  765 - 0x2fd  :   28 - 0x1c
    "00011100", --  766 - 0x2fe  :   28 - 0x1c
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Background 0x60
    "01111111", --  769 - 0x301  :  127 - 0x7f
    "01111111", --  770 - 0x302  :  127 - 0x7f
    "01111111", --  771 - 0x303  :  127 - 0x7f
    "01111111", --  772 - 0x304  :  127 - 0x7f
    "01111111", --  773 - 0x305  :  127 - 0x7f
    "00101010", --  774 - 0x306  :   42 - 0x2a
    "00000000", --  775 - 0x307  :    0 - 0x0
    "00000000", --  776 - 0x308  :    0 - 0x0 -- Background 0x61
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11111111", --  778 - 0x30a  :  255 - 0xff
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "11111111", --  780 - 0x30c  :  255 - 0xff
    "11111111", --  781 - 0x30d  :  255 - 0xff
    "10101010", --  782 - 0x30e  :  170 - 0xaa
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Background 0x62
    "11111110", --  785 - 0x311  :  254 - 0xfe
    "11111110", --  786 - 0x312  :  254 - 0xfe
    "11111110", --  787 - 0x313  :  254 - 0xfe
    "11111110", --  788 - 0x314  :  254 - 0xfe
    "11111110", --  789 - 0x315  :  254 - 0xfe
    "10101010", --  790 - 0x316  :  170 - 0xaa
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0 -- Background 0x63
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Background 0x64
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000001", --  802 - 0x322  :    1 - 0x1
    "00000001", --  803 - 0x323  :    1 - 0x1
    "00000011", --  804 - 0x324  :    3 - 0x3
    "00000011", --  805 - 0x325  :    3 - 0x3
    "00000111", --  806 - 0x326  :    7 - 0x7
    "00000111", --  807 - 0x327  :    7 - 0x7
    "00001111", --  808 - 0x328  :   15 - 0xf -- Background 0x65
    "00001111", --  809 - 0x329  :   15 - 0xf
    "00011111", --  810 - 0x32a  :   31 - 0x1f
    "00011111", --  811 - 0x32b  :   31 - 0x1f
    "00111111", --  812 - 0x32c  :   63 - 0x3f
    "00111111", --  813 - 0x32d  :   63 - 0x3f
    "01010101", --  814 - 0x32e  :   85 - 0x55
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Background 0x66
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000000", --  818 - 0x332  :    0 - 0x0
    "10000000", --  819 - 0x333  :  128 - 0x80
    "01000000", --  820 - 0x334  :   64 - 0x40
    "10000000", --  821 - 0x335  :  128 - 0x80
    "11000000", --  822 - 0x336  :  192 - 0xc0
    "11100000", --  823 - 0x337  :  224 - 0xe0
    "11010000", --  824 - 0x338  :  208 - 0xd0 -- Background 0x67
    "11100000", --  825 - 0x339  :  224 - 0xe0
    "11110000", --  826 - 0x33a  :  240 - 0xf0
    "11101000", --  827 - 0x33b  :  232 - 0xe8
    "11110100", --  828 - 0x33c  :  244 - 0xf4
    "11111000", --  829 - 0x33d  :  248 - 0xf8
    "01010100", --  830 - 0x33e  :   84 - 0x54
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Background 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Background 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Background 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0 -- Background 0x6b
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Background 0x6c
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "00000000", --  868 - 0x364  :    0 - 0x0
    "00000000", --  869 - 0x365  :    0 - 0x0
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Background 0x6d
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Background 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00000000", --  888 - 0x378  :    0 - 0x0 -- Background 0x6f
    "00000000", --  889 - 0x379  :    0 - 0x0
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Background 0x70
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0 -- Background 0x71
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Background 0x72
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0 -- Background 0x73
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Background 0x74
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- Background 0x75
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Background 0x76
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- Background 0x77
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Background 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Background 0x79
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Background 0x7a
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Background 0x7b
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Background 0x7c
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Background 0x7d
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- Background 0x7f
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Background 0x80
    "00000011", -- 1025 - 0x401  :    3 - 0x3
    "00001111", -- 1026 - 0x402  :   15 - 0xf
    "00011111", -- 1027 - 0x403  :   31 - 0x1f
    "00011111", -- 1028 - 0x404  :   31 - 0x1f
    "00111111", -- 1029 - 0x405  :   63 - 0x3f
    "00111111", -- 1030 - 0x406  :   63 - 0x3f
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00000000", -- 1032 - 0x408  :    0 - 0x0 -- Background 0x81
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Background 0x82
    "11000000", -- 1041 - 0x411  :  192 - 0xc0
    "11110000", -- 1042 - 0x412  :  240 - 0xf0
    "11110000", -- 1043 - 0x413  :  240 - 0xf0
    "11101100", -- 1044 - 0x414  :  236 - 0xec
    "11100000", -- 1045 - 0x415  :  224 - 0xe0
    "11111100", -- 1046 - 0x416  :  252 - 0xfc
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- Background 0x83
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "11100000", -- 1054 - 0x41e  :  224 - 0xe0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- Background 0x84
    "00000011", -- 1057 - 0x421  :    3 - 0x3
    "00001111", -- 1058 - 0x422  :   15 - 0xf
    "00011111", -- 1059 - 0x423  :   31 - 0x1f
    "00011111", -- 1060 - 0x424  :   31 - 0x1f
    "00111111", -- 1061 - 0x425  :   63 - 0x3f
    "00111111", -- 1062 - 0x426  :   63 - 0x3f
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0 -- Background 0x85
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00001000", -- 1069 - 0x42d  :    8 - 0x8
    "00001110", -- 1070 - 0x42e  :   14 - 0xe
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Background 0x86
    "11000000", -- 1073 - 0x431  :  192 - 0xc0
    "11110000", -- 1074 - 0x432  :  240 - 0xf0
    "11110000", -- 1075 - 0x433  :  240 - 0xf0
    "11101100", -- 1076 - 0x434  :  236 - 0xec
    "11100000", -- 1077 - 0x435  :  224 - 0xe0
    "11111100", -- 1078 - 0x436  :  252 - 0xfc
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- Background 0x87
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000110", -- 1085 - 0x43d  :    6 - 0x6
    "00001100", -- 1086 - 0x43e  :   12 - 0xc
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Background 0x88
    "00000011", -- 1089 - 0x441  :    3 - 0x3
    "00000011", -- 1090 - 0x442  :    3 - 0x3
    "00000100", -- 1091 - 0x443  :    4 - 0x4
    "00001111", -- 1092 - 0x444  :   15 - 0xf
    "00011111", -- 1093 - 0x445  :   31 - 0x1f
    "01101111", -- 1094 - 0x446  :  111 - 0x6f
    "01101111", -- 1095 - 0x447  :  111 - 0x6f
    "01101111", -- 1096 - 0x448  :  111 - 0x6f -- Background 0x89
    "01101111", -- 1097 - 0x449  :  111 - 0x6f
    "00011111", -- 1098 - 0x44a  :   31 - 0x1f
    "00001111", -- 1099 - 0x44b  :   15 - 0xf
    "00000100", -- 1100 - 0x44c  :    4 - 0x4
    "00000011", -- 1101 - 0x44d  :    3 - 0x3
    "00000011", -- 1102 - 0x44e  :    3 - 0x3
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Background 0x8a
    "00000000", -- 1105 - 0x451  :    0 - 0x0
    "00011000", -- 1106 - 0x452  :   24 - 0x18
    "00110111", -- 1107 - 0x453  :   55 - 0x37
    "00101111", -- 1108 - 0x454  :   47 - 0x2f
    "00011111", -- 1109 - 0x455  :   31 - 0x1f
    "00011111", -- 1110 - 0x456  :   31 - 0x1f
    "00011111", -- 1111 - 0x457  :   31 - 0x1f
    "00011111", -- 1112 - 0x458  :   31 - 0x1f -- Background 0x8b
    "00011111", -- 1113 - 0x459  :   31 - 0x1f
    "00011111", -- 1114 - 0x45a  :   31 - 0x1f
    "00101111", -- 1115 - 0x45b  :   47 - 0x2f
    "00110111", -- 1116 - 0x45c  :   55 - 0x37
    "00011000", -- 1117 - 0x45d  :   24 - 0x18
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Background 0x8c
    "00000011", -- 1121 - 0x461  :    3 - 0x3
    "00000001", -- 1122 - 0x462  :    1 - 0x1
    "00011001", -- 1123 - 0x463  :   25 - 0x19
    "00111001", -- 1124 - 0x464  :   57 - 0x39
    "00011011", -- 1125 - 0x465  :   27 - 0x1b
    "00001111", -- 1126 - 0x466  :   15 - 0xf
    "00001111", -- 1127 - 0x467  :   15 - 0xf
    "01111111", -- 1128 - 0x468  :  127 - 0x7f -- Background 0x8d
    "01111111", -- 1129 - 0x469  :  127 - 0x7f
    "00111111", -- 1130 - 0x46a  :   63 - 0x3f
    "00010111", -- 1131 - 0x46b  :   23 - 0x17
    "00000110", -- 1132 - 0x46c  :    6 - 0x6
    "00000100", -- 1133 - 0x46d  :    4 - 0x4
    "00000111", -- 1134 - 0x46e  :    7 - 0x7
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0 -- Background 0x8e
    "11000000", -- 1137 - 0x471  :  192 - 0xc0
    "11110000", -- 1138 - 0x472  :  240 - 0xf0
    "10111000", -- 1139 - 0x473  :  184 - 0xb8
    "10011100", -- 1140 - 0x474  :  156 - 0x9c
    "11111100", -- 1141 - 0x475  :  252 - 0xfc
    "11111110", -- 1142 - 0x476  :  254 - 0xfe
    "11000000", -- 1143 - 0x477  :  192 - 0xc0
    "11111110", -- 1144 - 0x478  :  254 - 0xfe -- Background 0x8f
    "11111110", -- 1145 - 0x479  :  254 - 0xfe
    "11111000", -- 1146 - 0x47a  :  248 - 0xf8
    "11110000", -- 1147 - 0x47b  :  240 - 0xf0
    "11000000", -- 1148 - 0x47c  :  192 - 0xc0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "10000000", -- 1151 - 0x47f  :  128 - 0x80
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Background 0x90
    "00000001", -- 1153 - 0x481  :    1 - 0x1
    "00001001", -- 1154 - 0x482  :    9 - 0x9
    "00011001", -- 1155 - 0x483  :   25 - 0x19
    "00011100", -- 1156 - 0x484  :   28 - 0x1c
    "00001101", -- 1157 - 0x485  :   13 - 0xd
    "00001111", -- 1158 - 0x486  :   15 - 0xf
    "00101111", -- 1159 - 0x487  :   47 - 0x2f
    "01111111", -- 1160 - 0x488  :  127 - 0x7f -- Background 0x91
    "01111111", -- 1161 - 0x489  :  127 - 0x7f
    "00111111", -- 1162 - 0x48a  :   63 - 0x3f
    "00011011", -- 1163 - 0x48b  :   27 - 0x1b
    "00000011", -- 1164 - 0x48c  :    3 - 0x3
    "00000011", -- 1165 - 0x48d  :    3 - 0x3
    "00000001", -- 1166 - 0x48e  :    1 - 0x1
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0 -- Background 0x92
    "11000000", -- 1169 - 0x491  :  192 - 0xc0
    "11110000", -- 1170 - 0x492  :  240 - 0xf0
    "11011000", -- 1171 - 0x493  :  216 - 0xd8
    "11001100", -- 1172 - 0x494  :  204 - 0xcc
    "11111100", -- 1173 - 0x495  :  252 - 0xfc
    "11111110", -- 1174 - 0x496  :  254 - 0xfe
    "11100000", -- 1175 - 0x497  :  224 - 0xe0
    "11111110", -- 1176 - 0x498  :  254 - 0xfe -- Background 0x93
    "11111110", -- 1177 - 0x499  :  254 - 0xfe
    "11111000", -- 1178 - 0x49a  :  248 - 0xf8
    "01110000", -- 1179 - 0x49b  :  112 - 0x70
    "01000000", -- 1180 - 0x49c  :   64 - 0x40
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "11000000", -- 1182 - 0x49e  :  192 - 0xc0
    "00100000", -- 1183 - 0x49f  :   32 - 0x20
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- Background 0x94
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00001100", -- 1186 - 0x4a2  :   12 - 0xc
    "00001110", -- 1187 - 0x4a3  :   14 - 0xe
    "00000110", -- 1188 - 0x4a4  :    6 - 0x6
    "00100110", -- 1189 - 0x4a5  :   38 - 0x26
    "00110111", -- 1190 - 0x4a6  :   55 - 0x37
    "00110011", -- 1191 - 0x4a7  :   51 - 0x33
    "01111111", -- 1192 - 0x4a8  :  127 - 0x7f -- Background 0x95
    "01111111", -- 1193 - 0x4a9  :  127 - 0x7f
    "00111111", -- 1194 - 0x4aa  :   63 - 0x3f
    "00011111", -- 1195 - 0x4ab  :   31 - 0x1f
    "00001110", -- 1196 - 0x4ac  :   14 - 0xe
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0 -- Background 0x96
    "11000000", -- 1201 - 0x4b1  :  192 - 0xc0
    "11110000", -- 1202 - 0x4b2  :  240 - 0xf0
    "01101000", -- 1203 - 0x4b3  :  104 - 0x68
    "01100100", -- 1204 - 0x4b4  :  100 - 0x64
    "11111100", -- 1205 - 0x4b5  :  252 - 0xfc
    "11111110", -- 1206 - 0x4b6  :  254 - 0xfe
    "11110000", -- 1207 - 0x4b7  :  240 - 0xf0
    "11111111", -- 1208 - 0x4b8  :  255 - 0xff -- Background 0x97
    "11111110", -- 1209 - 0x4b9  :  254 - 0xfe
    "11111100", -- 1210 - 0x4ba  :  252 - 0xfc
    "10110000", -- 1211 - 0x4bb  :  176 - 0xb0
    "11000000", -- 1212 - 0x4bc  :  192 - 0xc0
    "11000000", -- 1213 - 0x4bd  :  192 - 0xc0
    "01110000", -- 1214 - 0x4be  :  112 - 0x70
    "00001000", -- 1215 - 0x4bf  :    8 - 0x8
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- Background 0x98
    "00000001", -- 1217 - 0x4c1  :    1 - 0x1
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000000", -- 1219 - 0x4c3  :    0 - 0x0
    "00000000", -- 1220 - 0x4c4  :    0 - 0x0
    "00000000", -- 1221 - 0x4c5  :    0 - 0x0
    "00000001", -- 1222 - 0x4c6  :    1 - 0x1
    "00000011", -- 1223 - 0x4c7  :    3 - 0x3
    "00000111", -- 1224 - 0x4c8  :    7 - 0x7 -- Background 0x99
    "00010111", -- 1225 - 0x4c9  :   23 - 0x17
    "00101111", -- 1226 - 0x4ca  :   47 - 0x2f
    "00011110", -- 1227 - 0x4cb  :   30 - 0x1e
    "00010001", -- 1228 - 0x4cc  :   17 - 0x11
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000001", -- 1230 - 0x4ce  :    1 - 0x1
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Background 0x9a
    "00010000", -- 1233 - 0x4d1  :   16 - 0x10
    "01111000", -- 1234 - 0x4d2  :  120 - 0x78
    "01110100", -- 1235 - 0x4d3  :  116 - 0x74
    "11111110", -- 1236 - 0x4d4  :  254 - 0xfe
    "11111000", -- 1237 - 0x4d5  :  248 - 0xf8
    "11111100", -- 1238 - 0x4d6  :  252 - 0xfc
    "11111000", -- 1239 - 0x4d7  :  248 - 0xf8
    "11111000", -- 1240 - 0x4d8  :  248 - 0xf8 -- Background 0x9b
    "11010000", -- 1241 - 0x4d9  :  208 - 0xd0
    "00110000", -- 1242 - 0x4da  :   48 - 0x30
    "01100000", -- 1243 - 0x4db  :   96 - 0x60
    "10000000", -- 1244 - 0x4dc  :  128 - 0x80
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0 -- Background 0x9c
    "00000001", -- 1249 - 0x4e1  :    1 - 0x1
    "00000000", -- 1250 - 0x4e2  :    0 - 0x0
    "00000000", -- 1251 - 0x4e3  :    0 - 0x0
    "00000000", -- 1252 - 0x4e4  :    0 - 0x0
    "00000000", -- 1253 - 0x4e5  :    0 - 0x0
    "00000001", -- 1254 - 0x4e6  :    1 - 0x1
    "00000011", -- 1255 - 0x4e7  :    3 - 0x3
    "00000111", -- 1256 - 0x4e8  :    7 - 0x7 -- Background 0x9d
    "00010111", -- 1257 - 0x4e9  :   23 - 0x17
    "00101111", -- 1258 - 0x4ea  :   47 - 0x2f
    "00011110", -- 1259 - 0x4eb  :   30 - 0x1e
    "00010000", -- 1260 - 0x4ec  :   16 - 0x10
    "00000100", -- 1261 - 0x4ed  :    4 - 0x4
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0 -- Background 0x9e
    "00010000", -- 1265 - 0x4f1  :   16 - 0x10
    "01111000", -- 1266 - 0x4f2  :  120 - 0x78
    "01110100", -- 1267 - 0x4f3  :  116 - 0x74
    "11111110", -- 1268 - 0x4f4  :  254 - 0xfe
    "11111000", -- 1269 - 0x4f5  :  248 - 0xf8
    "11111100", -- 1270 - 0x4f6  :  252 - 0xfc
    "11111000", -- 1271 - 0x4f7  :  248 - 0xf8
    "11111000", -- 1272 - 0x4f8  :  248 - 0xf8 -- Background 0x9f
    "11010000", -- 1273 - 0x4f9  :  208 - 0xd0
    "00110000", -- 1274 - 0x4fa  :   48 - 0x30
    "11000000", -- 1275 - 0x4fb  :  192 - 0xc0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- Background 0xa0
    "00000011", -- 1281 - 0x501  :    3 - 0x3
    "00001111", -- 1282 - 0x502  :   15 - 0xf
    "00011111", -- 1283 - 0x503  :   31 - 0x1f
    "00111111", -- 1284 - 0x504  :   63 - 0x3f
    "00111111", -- 1285 - 0x505  :   63 - 0x3f
    "01111111", -- 1286 - 0x506  :  127 - 0x7f
    "01111111", -- 1287 - 0x507  :  127 - 0x7f
    "01111111", -- 1288 - 0x508  :  127 - 0x7f -- Background 0xa1
    "01111111", -- 1289 - 0x509  :  127 - 0x7f
    "00111111", -- 1290 - 0x50a  :   63 - 0x3f
    "00111111", -- 1291 - 0x50b  :   63 - 0x3f
    "00011111", -- 1292 - 0x50c  :   31 - 0x1f
    "00000101", -- 1293 - 0x50d  :    5 - 0x5
    "00000010", -- 1294 - 0x50e  :    2 - 0x2
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00000000", -- 1296 - 0x510  :    0 - 0x0 -- Background 0xa2
    "11000000", -- 1297 - 0x511  :  192 - 0xc0
    "11110000", -- 1298 - 0x512  :  240 - 0xf0
    "11111000", -- 1299 - 0x513  :  248 - 0xf8
    "11111000", -- 1300 - 0x514  :  248 - 0xf8
    "11111100", -- 1301 - 0x515  :  252 - 0xfc
    "11111010", -- 1302 - 0x516  :  250 - 0xfa
    "11111100", -- 1303 - 0x517  :  252 - 0xfc
    "11111010", -- 1304 - 0x518  :  250 - 0xfa -- Background 0xa3
    "11110100", -- 1305 - 0x519  :  244 - 0xf4
    "11101000", -- 1306 - 0x51a  :  232 - 0xe8
    "11010100", -- 1307 - 0x51b  :  212 - 0xd4
    "10101000", -- 1308 - 0x51c  :  168 - 0xa8
    "01010000", -- 1309 - 0x51d  :   80 - 0x50
    "10000000", -- 1310 - 0x51e  :  128 - 0x80
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Background 0xa4
    "00000000", -- 1313 - 0x521  :    0 - 0x0
    "00000000", -- 1314 - 0x522  :    0 - 0x0
    "00001110", -- 1315 - 0x523  :   14 - 0xe
    "00000000", -- 1316 - 0x524  :    0 - 0x0
    "00001010", -- 1317 - 0x525  :   10 - 0xa
    "01001010", -- 1318 - 0x526  :   74 - 0x4a
    "01100000", -- 1319 - 0x527  :   96 - 0x60
    "01111111", -- 1320 - 0x528  :  127 - 0x7f -- Background 0xa5
    "01111000", -- 1321 - 0x529  :  120 - 0x78
    "00110111", -- 1322 - 0x52a  :   55 - 0x37
    "00111011", -- 1323 - 0x52b  :   59 - 0x3b
    "00111100", -- 1324 - 0x52c  :   60 - 0x3c
    "00011111", -- 1325 - 0x52d  :   31 - 0x1f
    "00000111", -- 1326 - 0x52e  :    7 - 0x7
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Background 0xa6
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "01110000", -- 1331 - 0x533  :  112 - 0x70
    "00000000", -- 1332 - 0x534  :    0 - 0x0
    "01010000", -- 1333 - 0x535  :   80 - 0x50
    "01010010", -- 1334 - 0x536  :   82 - 0x52
    "00000110", -- 1335 - 0x537  :    6 - 0x6
    "11111100", -- 1336 - 0x538  :  252 - 0xfc -- Background 0xa7
    "00011010", -- 1337 - 0x539  :   26 - 0x1a
    "11101100", -- 1338 - 0x53a  :  236 - 0xec
    "11011000", -- 1339 - 0x53b  :  216 - 0xd8
    "00110100", -- 1340 - 0x53c  :   52 - 0x34
    "11101000", -- 1341 - 0x53d  :  232 - 0xe8
    "11000000", -- 1342 - 0x53e  :  192 - 0xc0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Background 0xa8
    "00000000", -- 1345 - 0x541  :    0 - 0x0
    "00000000", -- 1346 - 0x542  :    0 - 0x0
    "00001110", -- 1347 - 0x543  :   14 - 0xe
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00001110", -- 1349 - 0x545  :   14 - 0xe
    "01001010", -- 1350 - 0x546  :   74 - 0x4a
    "01100000", -- 1351 - 0x547  :   96 - 0x60
    "01111111", -- 1352 - 0x548  :  127 - 0x7f -- Background 0xa9
    "01111100", -- 1353 - 0x549  :  124 - 0x7c
    "01111011", -- 1354 - 0x54a  :  123 - 0x7b
    "01110111", -- 1355 - 0x54b  :  119 - 0x77
    "01111000", -- 1356 - 0x54c  :  120 - 0x78
    "01111111", -- 1357 - 0x54d  :  127 - 0x7f
    "01111111", -- 1358 - 0x54e  :  127 - 0x7f
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Background 0xaa
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "01110000", -- 1363 - 0x553  :  112 - 0x70
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "01110000", -- 1365 - 0x555  :  112 - 0x70
    "01010010", -- 1366 - 0x556  :   82 - 0x52
    "00000110", -- 1367 - 0x557  :    6 - 0x6
    "11111100", -- 1368 - 0x558  :  252 - 0xfc -- Background 0xab
    "00111010", -- 1369 - 0x559  :   58 - 0x3a
    "11011100", -- 1370 - 0x55a  :  220 - 0xdc
    "11101010", -- 1371 - 0x55b  :  234 - 0xea
    "00011100", -- 1372 - 0x55c  :   28 - 0x1c
    "11111010", -- 1373 - 0x55d  :  250 - 0xfa
    "11110100", -- 1374 - 0x55e  :  244 - 0xf4
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Background 0xac
    "00000011", -- 1377 - 0x561  :    3 - 0x3
    "00001111", -- 1378 - 0x562  :   15 - 0xf
    "00001111", -- 1379 - 0x563  :   15 - 0xf
    "00011111", -- 1380 - 0x564  :   31 - 0x1f
    "01011111", -- 1381 - 0x565  :   95 - 0x5f
    "01010000", -- 1382 - 0x566  :   80 - 0x50
    "00010000", -- 1383 - 0x567  :   16 - 0x10
    "00000000", -- 1384 - 0x568  :    0 - 0x0 -- Background 0xad
    "11111010", -- 1385 - 0x569  :  250 - 0xfa
    "11111010", -- 1386 - 0x56a  :  250 - 0xfa
    "11111010", -- 1387 - 0x56b  :  250 - 0xfa
    "10111010", -- 1388 - 0x56c  :  186 - 0xba
    "10011010", -- 1389 - 0x56d  :  154 - 0x9a
    "00001010", -- 1390 - 0x56e  :   10 - 0xa
    "00000010", -- 1391 - 0x56f  :    2 - 0x2
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Background 0xae
    "00000011", -- 1393 - 0x571  :    3 - 0x3
    "00001111", -- 1394 - 0x572  :   15 - 0xf
    "00001111", -- 1395 - 0x573  :   15 - 0xf
    "00011111", -- 1396 - 0x574  :   31 - 0x1f
    "01011111", -- 1397 - 0x575  :   95 - 0x5f
    "01010000", -- 1398 - 0x576  :   80 - 0x50
    "00010111", -- 1399 - 0x577  :   23 - 0x17
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Background 0xaf
    "11111010", -- 1401 - 0x579  :  250 - 0xfa
    "11111010", -- 1402 - 0x57a  :  250 - 0xfa
    "11111010", -- 1403 - 0x57b  :  250 - 0xfa
    "00111010", -- 1404 - 0x57c  :   58 - 0x3a
    "01011010", -- 1405 - 0x57d  :   90 - 0x5a
    "01101010", -- 1406 - 0x57e  :  106 - 0x6a
    "11110010", -- 1407 - 0x57f  :  242 - 0xf2
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Background 0xb0
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "00000011", -- 1410 - 0x582  :    3 - 0x3
    "00001111", -- 1411 - 0x583  :   15 - 0xf
    "00111011", -- 1412 - 0x584  :   59 - 0x3b
    "00111111", -- 1413 - 0x585  :   63 - 0x3f
    "01101111", -- 1414 - 0x586  :  111 - 0x6f
    "01111101", -- 1415 - 0x587  :  125 - 0x7d
    "00001111", -- 1416 - 0x588  :   15 - 0xf -- Background 0xb1
    "01110000", -- 1417 - 0x589  :  112 - 0x70
    "01111111", -- 1418 - 0x58a  :  127 - 0x7f
    "00001111", -- 1419 - 0x58b  :   15 - 0xf
    "01110000", -- 1420 - 0x58c  :  112 - 0x70
    "01111111", -- 1421 - 0x58d  :  127 - 0x7f
    "00001111", -- 1422 - 0x58e  :   15 - 0xf
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "00000000", -- 1424 - 0x590  :    0 - 0x0 -- Background 0xb2
    "00000000", -- 1425 - 0x591  :    0 - 0x0
    "11000000", -- 1426 - 0x592  :  192 - 0xc0
    "11110000", -- 1427 - 0x593  :  240 - 0xf0
    "10111100", -- 1428 - 0x594  :  188 - 0xbc
    "11110100", -- 1429 - 0x595  :  244 - 0xf4
    "11111110", -- 1430 - 0x596  :  254 - 0xfe
    "11011110", -- 1431 - 0x597  :  222 - 0xde
    "11110000", -- 1432 - 0x598  :  240 - 0xf0 -- Background 0xb3
    "00001110", -- 1433 - 0x599  :   14 - 0xe
    "11111110", -- 1434 - 0x59a  :  254 - 0xfe
    "11110000", -- 1435 - 0x59b  :  240 - 0xf0
    "00001110", -- 1436 - 0x59c  :   14 - 0xe
    "11111110", -- 1437 - 0x59d  :  254 - 0xfe
    "11110000", -- 1438 - 0x59e  :  240 - 0xf0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0 -- Background 0xb4
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "00000011", -- 1442 - 0x5a2  :    3 - 0x3
    "00001111", -- 1443 - 0x5a3  :   15 - 0xf
    "00111011", -- 1444 - 0x5a4  :   59 - 0x3b
    "00111111", -- 1445 - 0x5a5  :   63 - 0x3f
    "01101111", -- 1446 - 0x5a6  :  111 - 0x6f
    "01111101", -- 1447 - 0x5a7  :  125 - 0x7d
    "00001111", -- 1448 - 0x5a8  :   15 - 0xf -- Background 0xb5
    "01110000", -- 1449 - 0x5a9  :  112 - 0x70
    "01111111", -- 1450 - 0x5aa  :  127 - 0x7f
    "00001111", -- 1451 - 0x5ab  :   15 - 0xf
    "01110000", -- 1452 - 0x5ac  :  112 - 0x70
    "01111111", -- 1453 - 0x5ad  :  127 - 0x7f
    "00001111", -- 1454 - 0x5ae  :   15 - 0xf
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Background 0xb6
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "11000000", -- 1458 - 0x5b2  :  192 - 0xc0
    "11110000", -- 1459 - 0x5b3  :  240 - 0xf0
    "10111100", -- 1460 - 0x5b4  :  188 - 0xbc
    "11110100", -- 1461 - 0x5b5  :  244 - 0xf4
    "11111110", -- 1462 - 0x5b6  :  254 - 0xfe
    "11011110", -- 1463 - 0x5b7  :  222 - 0xde
    "11110000", -- 1464 - 0x5b8  :  240 - 0xf0 -- Background 0xb7
    "00001110", -- 1465 - 0x5b9  :   14 - 0xe
    "11111110", -- 1466 - 0x5ba  :  254 - 0xfe
    "11110000", -- 1467 - 0x5bb  :  240 - 0xf0
    "00001110", -- 1468 - 0x5bc  :   14 - 0xe
    "11111110", -- 1469 - 0x5bd  :  254 - 0xfe
    "11110000", -- 1470 - 0x5be  :  240 - 0xf0
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Background 0xb8
    "00000000", -- 1473 - 0x5c1  :    0 - 0x0
    "00000011", -- 1474 - 0x5c2  :    3 - 0x3
    "00001111", -- 1475 - 0x5c3  :   15 - 0xf
    "00111011", -- 1476 - 0x5c4  :   59 - 0x3b
    "00111111", -- 1477 - 0x5c5  :   63 - 0x3f
    "01101111", -- 1478 - 0x5c6  :  111 - 0x6f
    "01111101", -- 1479 - 0x5c7  :  125 - 0x7d
    "00001111", -- 1480 - 0x5c8  :   15 - 0xf -- Background 0xb9
    "00100000", -- 1481 - 0x5c9  :   32 - 0x20
    "01010101", -- 1482 - 0x5ca  :   85 - 0x55
    "00001010", -- 1483 - 0x5cb  :   10 - 0xa
    "01110000", -- 1484 - 0x5cc  :  112 - 0x70
    "01111111", -- 1485 - 0x5cd  :  127 - 0x7f
    "00001111", -- 1486 - 0x5ce  :   15 - 0xf
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Background 0xba
    "00000000", -- 1489 - 0x5d1  :    0 - 0x0
    "11000000", -- 1490 - 0x5d2  :  192 - 0xc0
    "11110000", -- 1491 - 0x5d3  :  240 - 0xf0
    "10111100", -- 1492 - 0x5d4  :  188 - 0xbc
    "11110100", -- 1493 - 0x5d5  :  244 - 0xf4
    "11111110", -- 1494 - 0x5d6  :  254 - 0xfe
    "11011110", -- 1495 - 0x5d7  :  222 - 0xde
    "11110000", -- 1496 - 0x5d8  :  240 - 0xf0 -- Background 0xbb
    "00001010", -- 1497 - 0x5d9  :   10 - 0xa
    "01010100", -- 1498 - 0x5da  :   84 - 0x54
    "10100000", -- 1499 - 0x5db  :  160 - 0xa0
    "00001110", -- 1500 - 0x5dc  :   14 - 0xe
    "11111110", -- 1501 - 0x5dd  :  254 - 0xfe
    "11110000", -- 1502 - 0x5de  :  240 - 0xf0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Background 0xbc
    "01110011", -- 1505 - 0x5e1  :  115 - 0x73
    "01111011", -- 1506 - 0x5e2  :  123 - 0x7b
    "01111111", -- 1507 - 0x5e3  :  127 - 0x7f
    "00111111", -- 1508 - 0x5e4  :   63 - 0x3f
    "00011100", -- 1509 - 0x5e5  :   28 - 0x1c
    "01111011", -- 1510 - 0x5e6  :  123 - 0x7b
    "01111011", -- 1511 - 0x5e7  :  123 - 0x7b
    "01111011", -- 1512 - 0x5e8  :  123 - 0x7b -- Background 0xbd
    "01111011", -- 1513 - 0x5e9  :  123 - 0x7b
    "00011100", -- 1514 - 0x5ea  :   28 - 0x1c
    "00111111", -- 1515 - 0x5eb  :   63 - 0x3f
    "01111111", -- 1516 - 0x5ec  :  127 - 0x7f
    "01111011", -- 1517 - 0x5ed  :  123 - 0x7b
    "01110011", -- 1518 - 0x5ee  :  115 - 0x73
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Background 0xbe
    "11001110", -- 1521 - 0x5f1  :  206 - 0xce
    "11011110", -- 1522 - 0x5f2  :  222 - 0xde
    "11111110", -- 1523 - 0x5f3  :  254 - 0xfe
    "11111100", -- 1524 - 0x5f4  :  252 - 0xfc
    "00111000", -- 1525 - 0x5f5  :   56 - 0x38
    "11011110", -- 1526 - 0x5f6  :  222 - 0xde
    "11011110", -- 1527 - 0x5f7  :  222 - 0xde
    "11011110", -- 1528 - 0x5f8  :  222 - 0xde -- Background 0xbf
    "11011110", -- 1529 - 0x5f9  :  222 - 0xde
    "00111000", -- 1530 - 0x5fa  :   56 - 0x38
    "11111100", -- 1531 - 0x5fb  :  252 - 0xfc
    "11111110", -- 1532 - 0x5fc  :  254 - 0xfe
    "11011110", -- 1533 - 0x5fd  :  222 - 0xde
    "11001110", -- 1534 - 0x5fe  :  206 - 0xce
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "01000000", -- 1538 - 0x602  :   64 - 0x40
    "01100000", -- 1539 - 0x603  :   96 - 0x60
    "01100001", -- 1540 - 0x604  :   97 - 0x61
    "00000010", -- 1541 - 0x605  :    2 - 0x2
    "00000010", -- 1542 - 0x606  :    2 - 0x2
    "00000111", -- 1543 - 0x607  :    7 - 0x7
    "00000111", -- 1544 - 0x608  :    7 - 0x7 -- Background 0xc1
    "00000100", -- 1545 - 0x609  :    4 - 0x4
    "00000111", -- 1546 - 0x60a  :    7 - 0x7
    "00000001", -- 1547 - 0x60b  :    1 - 0x1
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00010000", -- 1549 - 0x60d  :   16 - 0x10
    "00101000", -- 1550 - 0x60e  :   40 - 0x28
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000010", -- 1554 - 0x612  :    2 - 0x2
    "00000110", -- 1555 - 0x613  :    6 - 0x6
    "11100110", -- 1556 - 0x614  :  230 - 0xe6
    "10100000", -- 1557 - 0x615  :  160 - 0xa0
    "10100000", -- 1558 - 0x616  :  160 - 0xa0
    "11110000", -- 1559 - 0x617  :  240 - 0xf0
    "11110000", -- 1560 - 0x618  :  240 - 0xf0 -- Background 0xc3
    "00110000", -- 1561 - 0x619  :   48 - 0x30
    "11000000", -- 1562 - 0x61a  :  192 - 0xc0
    "10000000", -- 1563 - 0x61b  :  128 - 0x80
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00001000", -- 1565 - 0x61d  :    8 - 0x8
    "00010100", -- 1566 - 0x61e  :   20 - 0x14
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Background 0xc4
    "00000101", -- 1569 - 0x621  :    5 - 0x5
    "00000111", -- 1570 - 0x622  :    7 - 0x7
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000001", -- 1575 - 0x627  :    1 - 0x1
    "00000010", -- 1576 - 0x628  :    2 - 0x2 -- Background 0xc5
    "00000111", -- 1577 - 0x629  :    7 - 0x7
    "00100111", -- 1578 - 0x62a  :   39 - 0x27
    "01010011", -- 1579 - 0x62b  :   83 - 0x53
    "00000000", -- 1580 - 0x62c  :    0 - 0x0
    "00000010", -- 1581 - 0x62d  :    2 - 0x2
    "00000101", -- 1582 - 0x62e  :    5 - 0x5
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "00000000", -- 1584 - 0x630  :    0 - 0x0 -- Background 0xc6
    "00000000", -- 1585 - 0x631  :    0 - 0x0
    "00000000", -- 1586 - 0x632  :    0 - 0x0
    "00000000", -- 1587 - 0x633  :    0 - 0x0
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "01100000", -- 1589 - 0x635  :   96 - 0x60
    "11011000", -- 1590 - 0x636  :  216 - 0xd8
    "10110000", -- 1591 - 0x637  :  176 - 0xb0
    "11101000", -- 1592 - 0x638  :  232 - 0xe8 -- Background 0xc7
    "01111000", -- 1593 - 0x639  :  120 - 0x78
    "10110110", -- 1594 - 0x63a  :  182 - 0xb6
    "11100100", -- 1595 - 0x63b  :  228 - 0xe4
    "00000110", -- 1596 - 0x63c  :    6 - 0x6
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Background 0xc8
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "01000000", -- 1602 - 0x642  :   64 - 0x40
    "00100000", -- 1603 - 0x643  :   32 - 0x20
    "01000000", -- 1604 - 0x644  :   64 - 0x40
    "00000111", -- 1605 - 0x645  :    7 - 0x7
    "00000101", -- 1606 - 0x646  :    5 - 0x5
    "00001101", -- 1607 - 0x647  :   13 - 0xd
    "00001101", -- 1608 - 0x648  :   13 - 0xd -- Background 0xc9
    "00000101", -- 1609 - 0x649  :    5 - 0x5
    "00000011", -- 1610 - 0x64a  :    3 - 0x3
    "01000011", -- 1611 - 0x64b  :   67 - 0x43
    "00100000", -- 1612 - 0x64c  :   32 - 0x20
    "01000000", -- 1613 - 0x64d  :   64 - 0x40
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Background 0xca
    "00011100", -- 1617 - 0x651  :   28 - 0x1c
    "00011000", -- 1618 - 0x652  :   24 - 0x18
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "10000000", -- 1621 - 0x655  :  128 - 0x80
    "11100000", -- 1622 - 0x656  :  224 - 0xe0
    "10010000", -- 1623 - 0x657  :  144 - 0x90
    "11110000", -- 1624 - 0x658  :  240 - 0xf0 -- Background 0xcb
    "10010000", -- 1625 - 0x659  :  144 - 0x90
    "11110000", -- 1626 - 0x65a  :  240 - 0xf0
    "10000000", -- 1627 - 0x65b  :  128 - 0x80
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00011000", -- 1629 - 0x65d  :   24 - 0x18
    "00011100", -- 1630 - 0x65e  :   28 - 0x1c
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Background 0xcc
    "00001000", -- 1633 - 0x661  :    8 - 0x8
    "00000100", -- 1634 - 0x662  :    4 - 0x4
    "00001000", -- 1635 - 0x663  :    8 - 0x8
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "01000110", -- 1637 - 0x665  :   70 - 0x46
    "00101111", -- 1638 - 0x666  :   47 - 0x2f
    "01001110", -- 1639 - 0x667  :   78 - 0x4e
    "00001101", -- 1640 - 0x668  :   13 - 0xd -- Background 0xcd
    "00001011", -- 1641 - 0x669  :   11 - 0xb
    "00001111", -- 1642 - 0x66a  :   15 - 0xf
    "00000110", -- 1643 - 0x66b  :    6 - 0x6
    "00000011", -- 1644 - 0x66c  :    3 - 0x3
    "00011100", -- 1645 - 0x66d  :   28 - 0x1c
    "00010100", -- 1646 - 0x66e  :   20 - 0x14
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Background 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000110", -- 1653 - 0x675  :    6 - 0x6
    "00000100", -- 1654 - 0x676  :    4 - 0x4
    "10000110", -- 1655 - 0x677  :  134 - 0x86
    "11000000", -- 1656 - 0x678  :  192 - 0xc0 -- Background 0xcf
    "01100000", -- 1657 - 0x679  :   96 - 0x60
    "10100000", -- 1658 - 0x67a  :  160 - 0xa0
    "11000000", -- 1659 - 0x67b  :  192 - 0xc0
    "01000000", -- 1660 - 0x67c  :   64 - 0x40
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Background 0xd0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000100", -- 1668 - 0x684  :    4 - 0x4
    "00001110", -- 1669 - 0x685  :   14 - 0xe
    "00111111", -- 1670 - 0x686  :   63 - 0x3f
    "00111001", -- 1671 - 0x687  :   57 - 0x39
    "01110000", -- 1672 - 0x688  :  112 - 0x70 -- Background 0xd1
    "01111000", -- 1673 - 0x689  :  120 - 0x78
    "00111111", -- 1674 - 0x68a  :   63 - 0x3f
    "00111111", -- 1675 - 0x68b  :   63 - 0x3f
    "00000011", -- 1676 - 0x68c  :    3 - 0x3
    "00001100", -- 1677 - 0x68d  :   12 - 0xc
    "00001110", -- 1678 - 0x68e  :   14 - 0xe
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00000000", -- 1680 - 0x690  :    0 - 0x0 -- Background 0xd2
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00001000", -- 1683 - 0x693  :    8 - 0x8
    "11011000", -- 1684 - 0x694  :  216 - 0xd8
    "11111100", -- 1685 - 0x695  :  252 - 0xfc
    "11111100", -- 1686 - 0x696  :  252 - 0xfc
    "10011100", -- 1687 - 0x697  :  156 - 0x9c
    "00001100", -- 1688 - 0x698  :   12 - 0xc -- Background 0xd3
    "10011100", -- 1689 - 0x699  :  156 - 0x9c
    "11111000", -- 1690 - 0x69a  :  248 - 0xf8
    "01111000", -- 1691 - 0x69b  :  120 - 0x78
    "10001000", -- 1692 - 0x69c  :  136 - 0x88
    "00110000", -- 1693 - 0x69d  :   48 - 0x30
    "00111000", -- 1694 - 0x69e  :   56 - 0x38
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000001", -- 1700 - 0x6a4  :    1 - 0x1
    "00001011", -- 1701 - 0x6a5  :   11 - 0xb
    "00011111", -- 1702 - 0x6a6  :   31 - 0x1f
    "00111001", -- 1703 - 0x6a7  :   57 - 0x39
    "01110000", -- 1704 - 0x6a8  :  112 - 0x70 -- Background 0xd5
    "01111000", -- 1705 - 0x6a9  :  120 - 0x78
    "00111111", -- 1706 - 0x6aa  :   63 - 0x3f
    "00111111", -- 1707 - 0x6ab  :   63 - 0x3f
    "00000011", -- 1708 - 0x6ac  :    3 - 0x3
    "00111000", -- 1709 - 0x6ad  :   56 - 0x38
    "00011100", -- 1710 - 0x6ae  :   28 - 0x1c
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "11000000", -- 1715 - 0x6b3  :  192 - 0xc0
    "11001000", -- 1716 - 0x6b4  :  200 - 0xc8
    "11111000", -- 1717 - 0x6b5  :  248 - 0xf8
    "11111100", -- 1718 - 0x6b6  :  252 - 0xfc
    "10011100", -- 1719 - 0x6b7  :  156 - 0x9c
    "00001100", -- 1720 - 0x6b8  :   12 - 0xc -- Background 0xd7
    "10011100", -- 1721 - 0x6b9  :  156 - 0x9c
    "11111000", -- 1722 - 0x6ba  :  248 - 0xf8
    "01111000", -- 1723 - 0x6bb  :  120 - 0x78
    "11100010", -- 1724 - 0x6bc  :  226 - 0xe2
    "00011110", -- 1725 - 0x6bd  :   30 - 0x1e
    "00001100", -- 1726 - 0x6be  :   12 - 0xc
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Background 0xd8
    "00110000", -- 1729 - 0x6c1  :   48 - 0x30
    "00111100", -- 1730 - 0x6c2  :   60 - 0x3c
    "01111100", -- 1731 - 0x6c3  :  124 - 0x7c
    "01111100", -- 1732 - 0x6c4  :  124 - 0x7c
    "00111110", -- 1733 - 0x6c5  :   62 - 0x3e
    "00011100", -- 1734 - 0x6c6  :   28 - 0x1c
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0 -- Background 0xd9
    "00001110", -- 1737 - 0x6c9  :   14 - 0xe
    "00111110", -- 1738 - 0x6ca  :   62 - 0x3e
    "01111110", -- 1739 - 0x6cb  :  126 - 0x7e
    "01111110", -- 1740 - 0x6cc  :  126 - 0x7e
    "00111100", -- 1741 - 0x6cd  :   60 - 0x3c
    "00001100", -- 1742 - 0x6ce  :   12 - 0xc
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Background 0xda
    "00100000", -- 1745 - 0x6d1  :   32 - 0x20
    "01111110", -- 1746 - 0x6d2  :  126 - 0x7e
    "01111110", -- 1747 - 0x6d3  :  126 - 0x7e
    "01111110", -- 1748 - 0x6d4  :  126 - 0x7e
    "00111100", -- 1749 - 0x6d5  :   60 - 0x3c
    "00111000", -- 1750 - 0x6d6  :   56 - 0x38
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0 -- Background 0xdb
    "00011100", -- 1753 - 0x6d9  :   28 - 0x1c
    "00111110", -- 1754 - 0x6da  :   62 - 0x3e
    "01111110", -- 1755 - 0x6db  :  126 - 0x7e
    "01111110", -- 1756 - 0x6dc  :  126 - 0x7e
    "00111100", -- 1757 - 0x6dd  :   60 - 0x3c
    "00010000", -- 1758 - 0x6de  :   16 - 0x10
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000001", -- 1763 - 0x6e3  :    1 - 0x1
    "00000011", -- 1764 - 0x6e4  :    3 - 0x3
    "00000001", -- 1765 - 0x6e5  :    1 - 0x1
    "00000001", -- 1766 - 0x6e6  :    1 - 0x1
    "00001111", -- 1767 - 0x6e7  :   15 - 0xf
    "00000111", -- 1768 - 0x6e8  :    7 - 0x7 -- Background 0xdd
    "00000111", -- 1769 - 0x6e9  :    7 - 0x7
    "00000111", -- 1770 - 0x6ea  :    7 - 0x7
    "00011111", -- 1771 - 0x6eb  :   31 - 0x1f
    "00001111", -- 1772 - 0x6ec  :   15 - 0xf
    "00000111", -- 1773 - 0x6ed  :    7 - 0x7
    "00000011", -- 1774 - 0x6ee  :    3 - 0x3
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0 -- Background 0xde
    "00000000", -- 1777 - 0x6f1  :    0 - 0x0
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00000000", -- 1779 - 0x6f3  :    0 - 0x0
    "10000000", -- 1780 - 0x6f4  :  128 - 0x80
    "10000000", -- 1781 - 0x6f5  :  128 - 0x80
    "10010000", -- 1782 - 0x6f6  :  144 - 0x90
    "11110000", -- 1783 - 0x6f7  :  240 - 0xf0
    "11100000", -- 1784 - 0x6f8  :  224 - 0xe0 -- Background 0xdf
    "11100000", -- 1785 - 0x6f9  :  224 - 0xe0
    "11110000", -- 1786 - 0x6fa  :  240 - 0xf0
    "11110000", -- 1787 - 0x6fb  :  240 - 0xf0
    "11100000", -- 1788 - 0x6fc  :  224 - 0xe0
    "11000000", -- 1789 - 0x6fd  :  192 - 0xc0
    "11000000", -- 1790 - 0x6fe  :  192 - 0xc0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00001111", -- 1792 - 0x700  :   15 - 0xf -- Background 0xe0
    "00011111", -- 1793 - 0x701  :   31 - 0x1f
    "00011111", -- 1794 - 0x702  :   31 - 0x1f
    "00111111", -- 1795 - 0x703  :   63 - 0x3f
    "01111111", -- 1796 - 0x704  :  127 - 0x7f
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "11111111", -- 1798 - 0x706  :  255 - 0xff
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "11111111", -- 1800 - 0x708  :  255 - 0xff -- Background 0xe1
    "11111111", -- 1801 - 0x709  :  255 - 0xff
    "01111111", -- 1802 - 0x70a  :  127 - 0x7f
    "00111111", -- 1803 - 0x70b  :   63 - 0x3f
    "00111111", -- 1804 - 0x70c  :   63 - 0x3f
    "00011111", -- 1805 - 0x70d  :   31 - 0x1f
    "00001111", -- 1806 - 0x70e  :   15 - 0xf
    "00000111", -- 1807 - 0x70f  :    7 - 0x7
    "11111110", -- 1808 - 0x710  :  254 - 0xfe -- Background 0xe2
    "11111111", -- 1809 - 0x711  :  255 - 0xff
    "11111111", -- 1810 - 0x712  :  255 - 0xff
    "00001111", -- 1811 - 0x713  :   15 - 0xf
    "10111111", -- 1812 - 0x714  :  191 - 0xbf
    "10100011", -- 1813 - 0x715  :  163 - 0xa3
    "11110111", -- 1814 - 0x716  :  247 - 0xf7
    "11110111", -- 1815 - 0x717  :  247 - 0xf7
    "11111111", -- 1816 - 0x718  :  255 - 0xff -- Background 0xe3
    "11111111", -- 1817 - 0x719  :  255 - 0xff
    "00111111", -- 1818 - 0x71a  :   63 - 0x3f
    "00011111", -- 1819 - 0x71b  :   31 - 0x1f
    "11111110", -- 1820 - 0x71c  :  254 - 0xfe
    "11111100", -- 1821 - 0x71d  :  252 - 0xfc
    "11111000", -- 1822 - 0x71e  :  248 - 0xf8
    "11110000", -- 1823 - 0x71f  :  240 - 0xf0
    "00001111", -- 1824 - 0x720  :   15 - 0xf -- Background 0xe4
    "00011111", -- 1825 - 0x721  :   31 - 0x1f
    "00011111", -- 1826 - 0x722  :   31 - 0x1f
    "00111111", -- 1827 - 0x723  :   63 - 0x3f
    "01111111", -- 1828 - 0x724  :  127 - 0x7f
    "11111111", -- 1829 - 0x725  :  255 - 0xff
    "11111111", -- 1830 - 0x726  :  255 - 0xff
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "11111111", -- 1832 - 0x728  :  255 - 0xff -- Background 0xe5
    "11111111", -- 1833 - 0x729  :  255 - 0xff
    "01111110", -- 1834 - 0x72a  :  126 - 0x7e
    "00111111", -- 1835 - 0x72b  :   63 - 0x3f
    "00111111", -- 1836 - 0x72c  :   63 - 0x3f
    "00011111", -- 1837 - 0x72d  :   31 - 0x1f
    "00001111", -- 1838 - 0x72e  :   15 - 0xf
    "00000111", -- 1839 - 0x72f  :    7 - 0x7
    "11111110", -- 1840 - 0x730  :  254 - 0xfe -- Background 0xe6
    "11111111", -- 1841 - 0x731  :  255 - 0xff
    "11111111", -- 1842 - 0x732  :  255 - 0xff
    "11100011", -- 1843 - 0x733  :  227 - 0xe3
    "00010111", -- 1844 - 0x734  :   23 - 0x17
    "10110111", -- 1845 - 0x735  :  183 - 0xb7
    "10111111", -- 1846 - 0x736  :  191 - 0xbf
    "11111111", -- 1847 - 0x737  :  255 - 0xff
    "11111111", -- 1848 - 0x738  :  255 - 0xff -- Background 0xe7
    "11111111", -- 1849 - 0x739  :  255 - 0xff
    "00111111", -- 1850 - 0x73a  :   63 - 0x3f
    "00001111", -- 1851 - 0x73b  :   15 - 0xf
    "00001110", -- 1852 - 0x73c  :   14 - 0xe
    "11111100", -- 1853 - 0x73d  :  252 - 0xfc
    "11111000", -- 1854 - 0x73e  :  248 - 0xf8
    "11110000", -- 1855 - 0x73f  :  240 - 0xf0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Background 0xe8
    "00000101", -- 1857 - 0x741  :    5 - 0x5
    "00000111", -- 1858 - 0x742  :    7 - 0x7
    "00000011", -- 1859 - 0x743  :    3 - 0x3
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0 -- Background 0xe9
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000011", -- 1872 - 0x750  :    3 - 0x3 -- Background 0xea
    "10011110", -- 1873 - 0x751  :  158 - 0x9e
    "00001110", -- 1874 - 0x752  :   14 - 0xe
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- Background 0xeb
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Background 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000100", -- 1892 - 0x764  :    4 - 0x4
    "00001110", -- 1893 - 0x765  :   14 - 0xe
    "00001111", -- 1894 - 0x766  :   15 - 0xf
    "00001011", -- 1895 - 0x767  :   11 - 0xb
    "00001111", -- 1896 - 0x768  :   15 - 0xf -- Background 0xed
    "00001100", -- 1897 - 0x769  :   12 - 0xc
    "00001111", -- 1898 - 0x76a  :   15 - 0xf
    "00001111", -- 1899 - 0x76b  :   15 - 0xf
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "01111111", -- 1901 - 0x76d  :  127 - 0x7f
    "11010101", -- 1902 - 0x76e  :  213 - 0xd5
    "01111111", -- 1903 - 0x76f  :  127 - 0x7f
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Background 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00100000", -- 1908 - 0x774  :   32 - 0x20
    "01110000", -- 1909 - 0x775  :  112 - 0x70
    "11110000", -- 1910 - 0x776  :  240 - 0xf0
    "11100000", -- 1911 - 0x777  :  224 - 0xe0
    "11110000", -- 1912 - 0x778  :  240 - 0xf0 -- Background 0xef
    "00110000", -- 1913 - 0x779  :   48 - 0x30
    "11110000", -- 1914 - 0x77a  :  240 - 0xf0
    "11110000", -- 1915 - 0x77b  :  240 - 0xf0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "11111110", -- 1917 - 0x77d  :  254 - 0xfe
    "01010101", -- 1918 - 0x77e  :   85 - 0x55
    "11111110", -- 1919 - 0x77f  :  254 - 0xfe
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000100", -- 1924 - 0x784  :    4 - 0x4
    "00001110", -- 1925 - 0x785  :   14 - 0xe
    "00001111", -- 1926 - 0x786  :   15 - 0xf
    "00001011", -- 1927 - 0x787  :   11 - 0xb
    "00001111", -- 1928 - 0x788  :   15 - 0xf -- Background 0xf1
    "00001100", -- 1929 - 0x789  :   12 - 0xc
    "00001111", -- 1930 - 0x78a  :   15 - 0xf
    "00001111", -- 1931 - 0x78b  :   15 - 0xf
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "01111111", -- 1933 - 0x78d  :  127 - 0x7f
    "10101010", -- 1934 - 0x78e  :  170 - 0xaa
    "01111111", -- 1935 - 0x78f  :  127 - 0x7f
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Background 0xf2
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00100000", -- 1940 - 0x794  :   32 - 0x20
    "01110000", -- 1941 - 0x795  :  112 - 0x70
    "11110000", -- 1942 - 0x796  :  240 - 0xf0
    "11100000", -- 1943 - 0x797  :  224 - 0xe0
    "11110000", -- 1944 - 0x798  :  240 - 0xf0 -- Background 0xf3
    "00110000", -- 1945 - 0x799  :   48 - 0x30
    "11110000", -- 1946 - 0x79a  :  240 - 0xf0
    "11110000", -- 1947 - 0x79b  :  240 - 0xf0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "11111110", -- 1949 - 0x79d  :  254 - 0xfe
    "10101011", -- 1950 - 0x79e  :  171 - 0xab
    "11111110", -- 1951 - 0x79f  :  254 - 0xfe
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Background 0xf4
    "00010101", -- 1953 - 0x7a1  :   21 - 0x15
    "00001010", -- 1954 - 0x7a2  :   10 - 0xa
    "00000101", -- 1955 - 0x7a3  :    5 - 0x5
    "00000010", -- 1956 - 0x7a4  :    2 - 0x2
    "00000101", -- 1957 - 0x7a5  :    5 - 0x5
    "00000111", -- 1958 - 0x7a6  :    7 - 0x7
    "00000111", -- 1959 - 0x7a7  :    7 - 0x7
    "00111100", -- 1960 - 0x7a8  :   60 - 0x3c -- Background 0xf5
    "01111011", -- 1961 - 0x7a9  :  123 - 0x7b
    "01111011", -- 1962 - 0x7aa  :  123 - 0x7b
    "01111111", -- 1963 - 0x7ab  :  127 - 0x7f
    "01111110", -- 1964 - 0x7ac  :  126 - 0x7e
    "01111111", -- 1965 - 0x7ad  :  127 - 0x7f
    "00111110", -- 1966 - 0x7ae  :   62 - 0x3e
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Background 0xf6
    "01010000", -- 1969 - 0x7b1  :   80 - 0x50
    "10100000", -- 1970 - 0x7b2  :  160 - 0xa0
    "01000000", -- 1971 - 0x7b3  :   64 - 0x40
    "10100000", -- 1972 - 0x7b4  :  160 - 0xa0
    "01000000", -- 1973 - 0x7b5  :   64 - 0x40
    "11100000", -- 1974 - 0x7b6  :  224 - 0xe0
    "11100000", -- 1975 - 0x7b7  :  224 - 0xe0
    "01111000", -- 1976 - 0x7b8  :  120 - 0x78 -- Background 0xf7
    "10111100", -- 1977 - 0x7b9  :  188 - 0xbc
    "10111000", -- 1978 - 0x7ba  :  184 - 0xb8
    "10111110", -- 1979 - 0x7bb  :  190 - 0xbe
    "01111100", -- 1980 - 0x7bc  :  124 - 0x7c
    "11111110", -- 1981 - 0x7bd  :  254 - 0xfe
    "01111000", -- 1982 - 0x7be  :  120 - 0x78
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000011", -- 1984 - 0x7c0  :    3 - 0x3 -- Background 0xf8
    "00000011", -- 1985 - 0x7c1  :    3 - 0x3
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000011", -- 1987 - 0x7c3  :    3 - 0x3
    "00000111", -- 1988 - 0x7c4  :    7 - 0x7
    "00000110", -- 1989 - 0x7c5  :    6 - 0x6
    "00000111", -- 1990 - 0x7c6  :    7 - 0x7
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- Background 0xf9
    "00011111", -- 1993 - 0x7c9  :   31 - 0x1f
    "00011111", -- 1994 - 0x7ca  :   31 - 0x1f
    "00001111", -- 1995 - 0x7cb  :   15 - 0xf
    "00000011", -- 1996 - 0x7cc  :    3 - 0x3
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "11100000", -- 2000 - 0x7d0  :  224 - 0xe0 -- Background 0xfa
    "11100000", -- 2001 - 0x7d1  :  224 - 0xe0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00110000", -- 2003 - 0x7d3  :   48 - 0x30
    "01110000", -- 2004 - 0x7d4  :  112 - 0x70
    "01100000", -- 2005 - 0x7d5  :   96 - 0x60
    "01110000", -- 2006 - 0x7d6  :  112 - 0x70
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- Background 0xfb
    "11111000", -- 2009 - 0x7d9  :  248 - 0xf8
    "11111000", -- 2010 - 0x7da  :  248 - 0xf8
    "11110000", -- 2011 - 0x7db  :  240 - 0xf0
    "11000000", -- 2012 - 0x7dc  :  192 - 0xc0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00111000", -- 2016 - 0x7e0  :   56 - 0x38 -- Background 0xfc
    "00111000", -- 2017 - 0x7e1  :   56 - 0x38
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "01111100", -- 2019 - 0x7e3  :  124 - 0x7c
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00111000", -- 2021 - 0x7e5  :   56 - 0x38
    "00111000", -- 2022 - 0x7e6  :   56 - 0x38
    "01111100", -- 2023 - 0x7e7  :  124 - 0x7c
    "01111100", -- 2024 - 0x7e8  :  124 - 0x7c -- Background 0xfd
    "01111100", -- 2025 - 0x7e9  :  124 - 0x7c
    "01111100", -- 2026 - 0x7ea  :  124 - 0x7c
    "00111000", -- 2027 - 0x7eb  :   56 - 0x38
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "01111100", -- 2029 - 0x7ed  :  124 - 0x7c
    "01111100", -- 2030 - 0x7ee  :  124 - 0x7c
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Background 0xfe
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00010001", -- 2034 - 0x7f2  :   17 - 0x11
    "11010111", -- 2035 - 0x7f3  :  215 - 0xd7
    "11010111", -- 2036 - 0x7f4  :  215 - 0xd7
    "11010111", -- 2037 - 0x7f5  :  215 - 0xd7
    "00010001", -- 2038 - 0x7f6  :   17 - 0x11
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Background 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "11100110", -- 2042 - 0x7fa  :  230 - 0xe6
    "11110110", -- 2043 - 0x7fb  :  246 - 0xf6
    "11110110", -- 2044 - 0x7fc  :  246 - 0xf6
    "11110110", -- 2045 - 0x7fd  :  246 - 0xf6
    "11100110", -- 2046 - 0x7fe  :  230 - 0xe6
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
