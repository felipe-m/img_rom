--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables

---  Original memory dump file name: smario_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_SMARIO is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(13-1 downto 0);  --8192 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_SMARIO;

architecture BEHAVIORAL of ROM_PTABLE_SMARIO is
  signal addr_int  : natural range 0 to 2**13-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant nametable_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
    "00000011", --    0 -  0x0  :    3 - 0x3
    "00001111", --    1 -  0x1  :   15 - 0xf
    "00011111", --    2 -  0x2  :   31 - 0x1f
    "00011111", --    3 -  0x3  :   31 - 0x1f
    "00011100", --    4 -  0x4  :   28 - 0x1c
    "00100100", --    5 -  0x5  :   36 - 0x24
    "00100110", --    6 -  0x6  :   38 - 0x26
    "01100110", --    7 -  0x7  :  102 - 0x66
    "00000000", --    8 -  0x8  :    0 - 0x0
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00011111", --   12 -  0xc  :   31 - 0x1f
    "00111111", --   13 -  0xd  :   63 - 0x3f
    "00111111", --   14 -  0xe  :   63 - 0x3f
    "01111111", --   15 -  0xf  :  127 - 0x7f
    "11100000", --   16 - 0x10  :  224 - 0xe0
    "11000000", --   17 - 0x11  :  192 - 0xc0
    "10000000", --   18 - 0x12  :  128 - 0x80
    "11111100", --   19 - 0x13  :  252 - 0xfc
    "10000000", --   20 - 0x14  :  128 - 0x80
    "11000000", --   21 - 0x15  :  192 - 0xc0
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00100000", --   23 - 0x17  :   32 - 0x20
    "00000000", --   24 - 0x18  :    0 - 0x0
    "00100000", --   25 - 0x19  :   32 - 0x20
    "01100000", --   26 - 0x1a  :   96 - 0x60
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "11110000", --   28 - 0x1c  :  240 - 0xf0
    "11111100", --   29 - 0x1d  :  252 - 0xfc
    "11111110", --   30 - 0x1e  :  254 - 0xfe
    "11111110", --   31 - 0x1f  :  254 - 0xfe
    "01100000", --   32 - 0x20  :   96 - 0x60
    "01110000", --   33 - 0x21  :  112 - 0x70
    "00011000", --   34 - 0x22  :   24 - 0x18
    "00000111", --   35 - 0x23  :    7 - 0x7
    "00001111", --   36 - 0x24  :   15 - 0xf
    "00011111", --   37 - 0x25  :   31 - 0x1f
    "00111111", --   38 - 0x26  :   63 - 0x3f
    "01111111", --   39 - 0x27  :  127 - 0x7f
    "01111111", --   40 - 0x28  :  127 - 0x7f
    "01111111", --   41 - 0x29  :  127 - 0x7f
    "00011111", --   42 - 0x2a  :   31 - 0x1f
    "00000111", --   43 - 0x2b  :    7 - 0x7
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00011110", --   45 - 0x2d  :   30 - 0x1e
    "00111111", --   46 - 0x2e  :   63 - 0x3f
    "01111111", --   47 - 0x2f  :  127 - 0x7f
    "11111100", --   48 - 0x30  :  252 - 0xfc
    "01111100", --   49 - 0x31  :  124 - 0x7c
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00000000", --   51 - 0x33  :    0 - 0x0
    "11100000", --   52 - 0x34  :  224 - 0xe0
    "11110000", --   53 - 0x35  :  240 - 0xf0
    "11111000", --   54 - 0x36  :  248 - 0xf8
    "11111000", --   55 - 0x37  :  248 - 0xf8
    "11111100", --   56 - 0x38  :  252 - 0xfc
    "11111100", --   57 - 0x39  :  252 - 0xfc
    "11111000", --   58 - 0x3a  :  248 - 0xf8
    "11000000", --   59 - 0x3b  :  192 - 0xc0
    "11000010", --   60 - 0x3c  :  194 - 0xc2
    "01100111", --   61 - 0x3d  :  103 - 0x67
    "00101111", --   62 - 0x3e  :   47 - 0x2f
    "00110111", --   63 - 0x3f  :   55 - 0x37
    "01111111", --   64 - 0x40  :  127 - 0x7f
    "01111111", --   65 - 0x41  :  127 - 0x7f
    "11111111", --   66 - 0x42  :  255 - 0xff
    "11111111", --   67 - 0x43  :  255 - 0xff
    "00000111", --   68 - 0x44  :    7 - 0x7
    "00000111", --   69 - 0x45  :    7 - 0x7
    "00001111", --   70 - 0x46  :   15 - 0xf
    "00001111", --   71 - 0x47  :   15 - 0xf
    "01111111", --   72 - 0x48  :  127 - 0x7f
    "01111110", --   73 - 0x49  :  126 - 0x7e
    "11111100", --   74 - 0x4a  :  252 - 0xfc
    "11110000", --   75 - 0x4b  :  240 - 0xf0
    "11111000", --   76 - 0x4c  :  248 - 0xf8
    "11111000", --   77 - 0x4d  :  248 - 0xf8
    "11110000", --   78 - 0x4e  :  240 - 0xf0
    "01110000", --   79 - 0x4f  :  112 - 0x70
    "11111101", --   80 - 0x50  :  253 - 0xfd
    "11111110", --   81 - 0x51  :  254 - 0xfe
    "10110100", --   82 - 0x52  :  180 - 0xb4
    "11111000", --   83 - 0x53  :  248 - 0xf8
    "11111000", --   84 - 0x54  :  248 - 0xf8
    "11111001", --   85 - 0x55  :  249 - 0xf9
    "11111011", --   86 - 0x56  :  251 - 0xfb
    "11111111", --   87 - 0x57  :  255 - 0xff
    "00110111", --   88 - 0x58  :   55 - 0x37
    "00110110", --   89 - 0x59  :   54 - 0x36
    "01011100", --   90 - 0x5a  :   92 - 0x5c
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000001", --   93 - 0x5d  :    1 - 0x1
    "00000011", --   94 - 0x5e  :    3 - 0x3
    "00011111", --   95 - 0x5f  :   31 - 0x1f
    "00011111", --   96 - 0x60  :   31 - 0x1f
    "00111111", --   97 - 0x61  :   63 - 0x3f
    "11111111", --   98 - 0x62  :  255 - 0xff
    "11111111", --   99 - 0x63  :  255 - 0xff
    "11111100", --  100 - 0x64  :  252 - 0xfc
    "01110000", --  101 - 0x65  :  112 - 0x70
    "01110000", --  102 - 0x66  :  112 - 0x70
    "00111000", --  103 - 0x67  :   56 - 0x38
    "00001000", --  104 - 0x68  :    8 - 0x8
    "00100100", --  105 - 0x69  :   36 - 0x24
    "11100011", --  106 - 0x6a  :  227 - 0xe3
    "11110000", --  107 - 0x6b  :  240 - 0xf0
    "11111000", --  108 - 0x6c  :  248 - 0xf8
    "01110000", --  109 - 0x6d  :  112 - 0x70
    "01110000", --  110 - 0x6e  :  112 - 0x70
    "00111000", --  111 - 0x6f  :   56 - 0x38
    "11111111", --  112 - 0x70  :  255 - 0xff
    "11111111", --  113 - 0x71  :  255 - 0xff
    "11111111", --  114 - 0x72  :  255 - 0xff
    "00011111", --  115 - 0x73  :   31 - 0x1f
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00011111", --  120 - 0x78  :   31 - 0x1f
    "00011111", --  121 - 0x79  :   31 - 0x1f
    "00011111", --  122 - 0x7a  :   31 - 0x1f
    "00011111", --  123 - 0x7b  :   31 - 0x1f
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000001", --  130 - 0x82  :    1 - 0x1
    "00000111", --  131 - 0x83  :    7 - 0x7
    "00001111", --  132 - 0x84  :   15 - 0xf
    "00001111", --  133 - 0x85  :   15 - 0xf
    "00001110", --  134 - 0x86  :   14 - 0xe
    "00010010", --  135 - 0x87  :   18 - 0x12
    "00000000", --  136 - 0x88  :    0 - 0x0
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00001111", --  142 - 0x8e  :   15 - 0xf
    "00011111", --  143 - 0x8f  :   31 - 0x1f
    "00000000", --  144 - 0x90  :    0 - 0x0
    "00000000", --  145 - 0x91  :    0 - 0x0
    "11110000", --  146 - 0x92  :  240 - 0xf0
    "11100000", --  147 - 0x93  :  224 - 0xe0
    "11000000", --  148 - 0x94  :  192 - 0xc0
    "11111110", --  149 - 0x95  :  254 - 0xfe
    "01000000", --  150 - 0x96  :   64 - 0x40
    "01100000", --  151 - 0x97  :   96 - 0x60
    "00000000", --  152 - 0x98  :    0 - 0x0
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00010000", --  155 - 0x9b  :   16 - 0x10
    "00110000", --  156 - 0x9c  :   48 - 0x30
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "11111000", --  158 - 0x9e  :  248 - 0xf8
    "11111110", --  159 - 0x9f  :  254 - 0xfe
    "00010011", --  160 - 0xa0  :   19 - 0x13
    "00110011", --  161 - 0xa1  :   51 - 0x33
    "00110000", --  162 - 0xa2  :   48 - 0x30
    "00011000", --  163 - 0xa3  :   24 - 0x18
    "00000100", --  164 - 0xa4  :    4 - 0x4
    "00001111", --  165 - 0xa5  :   15 - 0xf
    "00011111", --  166 - 0xa6  :   31 - 0x1f
    "00011111", --  167 - 0xa7  :   31 - 0x1f
    "00011111", --  168 - 0xa8  :   31 - 0x1f
    "00111111", --  169 - 0xa9  :   63 - 0x3f
    "00111111", --  170 - 0xaa  :   63 - 0x3f
    "00011111", --  171 - 0xab  :   31 - 0x1f
    "00000111", --  172 - 0xac  :    7 - 0x7
    "00001000", --  173 - 0xad  :    8 - 0x8
    "00010111", --  174 - 0xae  :   23 - 0x17
    "00010111", --  175 - 0xaf  :   23 - 0x17
    "00000000", --  176 - 0xb0  :    0 - 0x0
    "00010000", --  177 - 0xb1  :   16 - 0x10
    "01111110", --  178 - 0xb2  :  126 - 0x7e
    "00111110", --  179 - 0xb3  :   62 - 0x3e
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "11000000", --  182 - 0xb6  :  192 - 0xc0
    "11100000", --  183 - 0xb7  :  224 - 0xe0
    "11111111", --  184 - 0xb8  :  255 - 0xff
    "11111111", --  185 - 0xb9  :  255 - 0xff
    "11111110", --  186 - 0xba  :  254 - 0xfe
    "11111110", --  187 - 0xbb  :  254 - 0xfe
    "11111100", --  188 - 0xbc  :  252 - 0xfc
    "11100000", --  189 - 0xbd  :  224 - 0xe0
    "01000000", --  190 - 0xbe  :   64 - 0x40
    "10100000", --  191 - 0xbf  :  160 - 0xa0
    "00111111", --  192 - 0xc0  :   63 - 0x3f
    "00111111", --  193 - 0xc1  :   63 - 0x3f
    "00111111", --  194 - 0xc2  :   63 - 0x3f
    "00011111", --  195 - 0xc3  :   31 - 0x1f
    "00011111", --  196 - 0xc4  :   31 - 0x1f
    "00011111", --  197 - 0xc5  :   31 - 0x1f
    "00011111", --  198 - 0xc6  :   31 - 0x1f
    "00011111", --  199 - 0xc7  :   31 - 0x1f
    "00110111", --  200 - 0xc8  :   55 - 0x37
    "00100111", --  201 - 0xc9  :   39 - 0x27
    "00100011", --  202 - 0xca  :   35 - 0x23
    "00000011", --  203 - 0xcb  :    3 - 0x3
    "00000001", --  204 - 0xcc  :    1 - 0x1
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "11110000", --  208 - 0xd0  :  240 - 0xf0
    "11110000", --  209 - 0xd1  :  240 - 0xf0
    "11110000", --  210 - 0xd2  :  240 - 0xf0
    "11111000", --  211 - 0xd3  :  248 - 0xf8
    "11111000", --  212 - 0xd4  :  248 - 0xf8
    "11111000", --  213 - 0xd5  :  248 - 0xf8
    "11111000", --  214 - 0xd6  :  248 - 0xf8
    "11111000", --  215 - 0xd7  :  248 - 0xf8
    "11001100", --  216 - 0xd8  :  204 - 0xcc
    "11111111", --  217 - 0xd9  :  255 - 0xff
    "11111111", --  218 - 0xda  :  255 - 0xff
    "11111111", --  219 - 0xdb  :  255 - 0xff
    "11111111", --  220 - 0xdc  :  255 - 0xff
    "01110000", --  221 - 0xdd  :  112 - 0x70
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00001000", --  223 - 0xdf  :    8 - 0x8
    "11111111", --  224 - 0xe0  :  255 - 0xff
    "11111111", --  225 - 0xe1  :  255 - 0xff
    "11111111", --  226 - 0xe2  :  255 - 0xff
    "11111110", --  227 - 0xe3  :  254 - 0xfe
    "11110000", --  228 - 0xe4  :  240 - 0xf0
    "11000000", --  229 - 0xe5  :  192 - 0xc0
    "10000000", --  230 - 0xe6  :  128 - 0x80
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "11110000", --  232 - 0xe8  :  240 - 0xf0
    "11110000", --  233 - 0xe9  :  240 - 0xf0
    "11110000", --  234 - 0xea  :  240 - 0xf0
    "11110000", --  235 - 0xeb  :  240 - 0xf0
    "11110000", --  236 - 0xec  :  240 - 0xf0
    "11000000", --  237 - 0xed  :  192 - 0xc0
    "10000000", --  238 - 0xee  :  128 - 0x80
    "00000000", --  239 - 0xef  :    0 - 0x0
    "11111100", --  240 - 0xf0  :  252 - 0xfc
    "11111100", --  241 - 0xf1  :  252 - 0xfc
    "11111000", --  242 - 0xf2  :  248 - 0xf8
    "01111000", --  243 - 0xf3  :  120 - 0x78
    "01111000", --  244 - 0xf4  :  120 - 0x78
    "01111000", --  245 - 0xf5  :  120 - 0x78
    "01111110", --  246 - 0xf6  :  126 - 0x7e
    "01111110", --  247 - 0xf7  :  126 - 0x7e
    "00010000", --  248 - 0xf8  :   16 - 0x10
    "01100000", --  249 - 0xf9  :   96 - 0x60
    "10000000", --  250 - 0xfa  :  128 - 0x80
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "01111000", --  252 - 0xfc  :  120 - 0x78
    "01111000", --  253 - 0xfd  :  120 - 0x78
    "01111110", --  254 - 0xfe  :  126 - 0x7e
    "01111110", --  255 - 0xff  :  126 - 0x7e
    "00000000", --  256 - 0x100  :    0 - 0x0
    "00000011", --  257 - 0x101  :    3 - 0x3
    "00001111", --  258 - 0x102  :   15 - 0xf
    "00011111", --  259 - 0x103  :   31 - 0x1f
    "00011111", --  260 - 0x104  :   31 - 0x1f
    "00011100", --  261 - 0x105  :   28 - 0x1c
    "00100100", --  262 - 0x106  :   36 - 0x24
    "00100110", --  263 - 0x107  :   38 - 0x26
    "00000000", --  264 - 0x108  :    0 - 0x0
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00011111", --  269 - 0x10d  :   31 - 0x1f
    "00111111", --  270 - 0x10e  :   63 - 0x3f
    "00111111", --  271 - 0x10f  :   63 - 0x3f
    "00000000", --  272 - 0x110  :    0 - 0x0
    "11100000", --  273 - 0x111  :  224 - 0xe0
    "11000000", --  274 - 0x112  :  192 - 0xc0
    "10000000", --  275 - 0x113  :  128 - 0x80
    "11111100", --  276 - 0x114  :  252 - 0xfc
    "10000000", --  277 - 0x115  :  128 - 0x80
    "11000000", --  278 - 0x116  :  192 - 0xc0
    "00000000", --  279 - 0x117  :    0 - 0x0
    "00000000", --  280 - 0x118  :    0 - 0x0
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00100000", --  282 - 0x11a  :   32 - 0x20
    "01100000", --  283 - 0x11b  :   96 - 0x60
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "11110000", --  285 - 0x11d  :  240 - 0xf0
    "11111100", --  286 - 0x11e  :  252 - 0xfc
    "11111110", --  287 - 0x11f  :  254 - 0xfe
    "01100110", --  288 - 0x120  :  102 - 0x66
    "01100000", --  289 - 0x121  :   96 - 0x60
    "00110000", --  290 - 0x122  :   48 - 0x30
    "00011000", --  291 - 0x123  :   24 - 0x18
    "00001111", --  292 - 0x124  :   15 - 0xf
    "00011111", --  293 - 0x125  :   31 - 0x1f
    "00111111", --  294 - 0x126  :   63 - 0x3f
    "00111111", --  295 - 0x127  :   63 - 0x3f
    "01111111", --  296 - 0x128  :  127 - 0x7f
    "01111111", --  297 - 0x129  :  127 - 0x7f
    "00111111", --  298 - 0x12a  :   63 - 0x3f
    "00011111", --  299 - 0x12b  :   31 - 0x1f
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00010110", --  301 - 0x12d  :   22 - 0x16
    "00101111", --  302 - 0x12e  :   47 - 0x2f
    "00101111", --  303 - 0x12f  :   47 - 0x2f
    "00100000", --  304 - 0x130  :   32 - 0x20
    "11111100", --  305 - 0x131  :  252 - 0xfc
    "01111100", --  306 - 0x132  :  124 - 0x7c
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "11100000", --  309 - 0x135  :  224 - 0xe0
    "11100000", --  310 - 0x136  :  224 - 0xe0
    "11110000", --  311 - 0x137  :  240 - 0xf0
    "11111110", --  312 - 0x138  :  254 - 0xfe
    "11111100", --  313 - 0x139  :  252 - 0xfc
    "11111100", --  314 - 0x13a  :  252 - 0xfc
    "11111000", --  315 - 0x13b  :  248 - 0xf8
    "11000000", --  316 - 0x13c  :  192 - 0xc0
    "01100000", --  317 - 0x13d  :   96 - 0x60
    "00100000", --  318 - 0x13e  :   32 - 0x20
    "00110000", --  319 - 0x13f  :   48 - 0x30
    "00111111", --  320 - 0x140  :   63 - 0x3f
    "00111111", --  321 - 0x141  :   63 - 0x3f
    "00111111", --  322 - 0x142  :   63 - 0x3f
    "00111111", --  323 - 0x143  :   63 - 0x3f
    "00111111", --  324 - 0x144  :   63 - 0x3f
    "00111111", --  325 - 0x145  :   63 - 0x3f
    "00111111", --  326 - 0x146  :   63 - 0x3f
    "00011111", --  327 - 0x147  :   31 - 0x1f
    "00101111", --  328 - 0x148  :   47 - 0x2f
    "00101111", --  329 - 0x149  :   47 - 0x2f
    "00101111", --  330 - 0x14a  :   47 - 0x2f
    "00001111", --  331 - 0x14b  :   15 - 0xf
    "00000111", --  332 - 0x14c  :    7 - 0x7
    "00000011", --  333 - 0x14d  :    3 - 0x3
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "11110000", --  336 - 0x150  :  240 - 0xf0
    "10010000", --  337 - 0x151  :  144 - 0x90
    "00000000", --  338 - 0x152  :    0 - 0x0
    "00001000", --  339 - 0x153  :    8 - 0x8
    "00001100", --  340 - 0x154  :   12 - 0xc
    "00011100", --  341 - 0x155  :   28 - 0x1c
    "11111100", --  342 - 0x156  :  252 - 0xfc
    "11111000", --  343 - 0x157  :  248 - 0xf8
    "00010000", --  344 - 0x158  :   16 - 0x10
    "11110000", --  345 - 0x159  :  240 - 0xf0
    "11110000", --  346 - 0x15a  :  240 - 0xf0
    "11110000", --  347 - 0x15b  :  240 - 0xf0
    "11110000", --  348 - 0x15c  :  240 - 0xf0
    "11100000", --  349 - 0x15d  :  224 - 0xe0
    "11000000", --  350 - 0x15e  :  192 - 0xc0
    "11100000", --  351 - 0x15f  :  224 - 0xe0
    "00001111", --  352 - 0x160  :   15 - 0xf
    "00001111", --  353 - 0x161  :   15 - 0xf
    "00000111", --  354 - 0x162  :    7 - 0x7
    "00000111", --  355 - 0x163  :    7 - 0x7
    "00000111", --  356 - 0x164  :    7 - 0x7
    "00001111", --  357 - 0x165  :   15 - 0xf
    "00001111", --  358 - 0x166  :   15 - 0xf
    "00000011", --  359 - 0x167  :    3 - 0x3
    "00000001", --  360 - 0x168  :    1 - 0x1
    "00000011", --  361 - 0x169  :    3 - 0x3
    "00000001", --  362 - 0x16a  :    1 - 0x1
    "00000100", --  363 - 0x16b  :    4 - 0x4
    "00000111", --  364 - 0x16c  :    7 - 0x7
    "00001111", --  365 - 0x16d  :   15 - 0xf
    "00001111", --  366 - 0x16e  :   15 - 0xf
    "00000011", --  367 - 0x16f  :    3 - 0x3
    "11111000", --  368 - 0x170  :  248 - 0xf8
    "11110000", --  369 - 0x171  :  240 - 0xf0
    "11100000", --  370 - 0x172  :  224 - 0xe0
    "11110000", --  371 - 0x173  :  240 - 0xf0
    "10110000", --  372 - 0x174  :  176 - 0xb0
    "10000000", --  373 - 0x175  :  128 - 0x80
    "11100000", --  374 - 0x176  :  224 - 0xe0
    "11100000", --  375 - 0x177  :  224 - 0xe0
    "11111000", --  376 - 0x178  :  248 - 0xf8
    "11110000", --  377 - 0x179  :  240 - 0xf0
    "11100000", --  378 - 0x17a  :  224 - 0xe0
    "01110000", --  379 - 0x17b  :  112 - 0x70
    "10110000", --  380 - 0x17c  :  176 - 0xb0
    "10000000", --  381 - 0x17d  :  128 - 0x80
    "11100000", --  382 - 0x17e  :  224 - 0xe0
    "11100000", --  383 - 0x17f  :  224 - 0xe0
    "00000011", --  384 - 0x180  :    3 - 0x3
    "00111111", --  385 - 0x181  :   63 - 0x3f
    "01111111", --  386 - 0x182  :  127 - 0x7f
    "00011001", --  387 - 0x183  :   25 - 0x19
    "00001001", --  388 - 0x184  :    9 - 0x9
    "00001001", --  389 - 0x185  :    9 - 0x9
    "00101000", --  390 - 0x186  :   40 - 0x28
    "01011100", --  391 - 0x187  :   92 - 0x5c
    "00000000", --  392 - 0x188  :    0 - 0x0
    "00110000", --  393 - 0x189  :   48 - 0x30
    "01110000", --  394 - 0x18a  :  112 - 0x70
    "01111111", --  395 - 0x18b  :  127 - 0x7f
    "11111111", --  396 - 0x18c  :  255 - 0xff
    "11111111", --  397 - 0x18d  :  255 - 0xff
    "11110111", --  398 - 0x18e  :  247 - 0xf7
    "11110011", --  399 - 0x18f  :  243 - 0xf3
    "11111000", --  400 - 0x190  :  248 - 0xf8
    "11100000", --  401 - 0x191  :  224 - 0xe0
    "11100000", --  402 - 0x192  :  224 - 0xe0
    "11111100", --  403 - 0x193  :  252 - 0xfc
    "00100110", --  404 - 0x194  :   38 - 0x26
    "00110000", --  405 - 0x195  :   48 - 0x30
    "10000000", --  406 - 0x196  :  128 - 0x80
    "00010000", --  407 - 0x197  :   16 - 0x10
    "00000000", --  408 - 0x198  :    0 - 0x0
    "00011000", --  409 - 0x199  :   24 - 0x18
    "00010000", --  410 - 0x19a  :   16 - 0x10
    "00000000", --  411 - 0x19b  :    0 - 0x0
    "11111000", --  412 - 0x19c  :  248 - 0xf8
    "11111000", --  413 - 0x19d  :  248 - 0xf8
    "11111110", --  414 - 0x19e  :  254 - 0xfe
    "11111111", --  415 - 0x19f  :  255 - 0xff
    "00111110", --  416 - 0x1a0  :   62 - 0x3e
    "00011110", --  417 - 0x1a1  :   30 - 0x1e
    "00111111", --  418 - 0x1a2  :   63 - 0x3f
    "00111000", --  419 - 0x1a3  :   56 - 0x38
    "00110000", --  420 - 0x1a4  :   48 - 0x30
    "00110000", --  421 - 0x1a5  :   48 - 0x30
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "00111010", --  423 - 0x1a7  :   58 - 0x3a
    "11100111", --  424 - 0x1a8  :  231 - 0xe7
    "00001111", --  425 - 0x1a9  :   15 - 0xf
    "00001111", --  426 - 0x1aa  :   15 - 0xf
    "00011111", --  427 - 0x1ab  :   31 - 0x1f
    "00011111", --  428 - 0x1ac  :   31 - 0x1f
    "00011111", --  429 - 0x1ad  :   31 - 0x1f
    "00001111", --  430 - 0x1ae  :   15 - 0xf
    "00000111", --  431 - 0x1af  :    7 - 0x7
    "01111000", --  432 - 0x1b0  :  120 - 0x78
    "00011110", --  433 - 0x1b1  :   30 - 0x1e
    "10000000", --  434 - 0x1b2  :  128 - 0x80
    "11111110", --  435 - 0x1b3  :  254 - 0xfe
    "01111110", --  436 - 0x1b4  :  126 - 0x7e
    "01111110", --  437 - 0x1b5  :  126 - 0x7e
    "01111111", --  438 - 0x1b6  :  127 - 0x7f
    "01111111", --  439 - 0x1b7  :  127 - 0x7f
    "11111111", --  440 - 0x1b8  :  255 - 0xff
    "11111110", --  441 - 0x1b9  :  254 - 0xfe
    "11111100", --  442 - 0x1ba  :  252 - 0xfc
    "11000110", --  443 - 0x1bb  :  198 - 0xc6
    "10001110", --  444 - 0x1bc  :  142 - 0x8e
    "11101110", --  445 - 0x1bd  :  238 - 0xee
    "11111111", --  446 - 0x1be  :  255 - 0xff
    "11111111", --  447 - 0x1bf  :  255 - 0xff
    "00111100", --  448 - 0x1c0  :   60 - 0x3c
    "00111111", --  449 - 0x1c1  :   63 - 0x3f
    "00011111", --  450 - 0x1c2  :   31 - 0x1f
    "00001111", --  451 - 0x1c3  :   15 - 0xf
    "00000111", --  452 - 0x1c4  :    7 - 0x7
    "00111111", --  453 - 0x1c5  :   63 - 0x3f
    "00100001", --  454 - 0x1c6  :   33 - 0x21
    "00100000", --  455 - 0x1c7  :   32 - 0x20
    "00000011", --  456 - 0x1c8  :    3 - 0x3
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00001110", --  459 - 0x1cb  :   14 - 0xe
    "00000111", --  460 - 0x1cc  :    7 - 0x7
    "00111111", --  461 - 0x1cd  :   63 - 0x3f
    "00111111", --  462 - 0x1ce  :   63 - 0x3f
    "00111111", --  463 - 0x1cf  :   63 - 0x3f
    "11111111", --  464 - 0x1d0  :  255 - 0xff
    "11111111", --  465 - 0x1d1  :  255 - 0xff
    "11111111", --  466 - 0x1d2  :  255 - 0xff
    "11111110", --  467 - 0x1d3  :  254 - 0xfe
    "11111110", --  468 - 0x1d4  :  254 - 0xfe
    "11111110", --  469 - 0x1d5  :  254 - 0xfe
    "11111100", --  470 - 0x1d6  :  252 - 0xfc
    "01110000", --  471 - 0x1d7  :  112 - 0x70
    "11111111", --  472 - 0x1d8  :  255 - 0xff
    "01111111", --  473 - 0x1d9  :  127 - 0x7f
    "00111111", --  474 - 0x1da  :   63 - 0x3f
    "00001110", --  475 - 0x1db  :   14 - 0xe
    "11000000", --  476 - 0x1dc  :  192 - 0xc0
    "11000000", --  477 - 0x1dd  :  192 - 0xc0
    "11100000", --  478 - 0x1de  :  224 - 0xe0
    "11100000", --  479 - 0x1df  :  224 - 0xe0
    "00001111", --  480 - 0x1e0  :   15 - 0xf
    "10011111", --  481 - 0x1e1  :  159 - 0x9f
    "11001111", --  482 - 0x1e2  :  207 - 0xcf
    "11111111", --  483 - 0x1e3  :  255 - 0xff
    "01111111", --  484 - 0x1e4  :  127 - 0x7f
    "00111111", --  485 - 0x1e5  :   63 - 0x3f
    "00011110", --  486 - 0x1e6  :   30 - 0x1e
    "00001110", --  487 - 0x1e7  :   14 - 0xe
    "00000000", --  488 - 0x1e8  :    0 - 0x0
    "10000000", --  489 - 0x1e9  :  128 - 0x80
    "11001000", --  490 - 0x1ea  :  200 - 0xc8
    "11111110", --  491 - 0x1eb  :  254 - 0xfe
    "01111111", --  492 - 0x1ec  :  127 - 0x7f
    "00111111", --  493 - 0x1ed  :   63 - 0x3f
    "00011110", --  494 - 0x1ee  :   30 - 0x1e
    "00001110", --  495 - 0x1ef  :   14 - 0xe
    "00100000", --  496 - 0x1f0  :   32 - 0x20
    "11000000", --  497 - 0x1f1  :  192 - 0xc0
    "10000000", --  498 - 0x1f2  :  128 - 0x80
    "10000000", --  499 - 0x1f3  :  128 - 0x80
    "00000000", --  500 - 0x1f4  :    0 - 0x0
    "00000000", --  501 - 0x1f5  :    0 - 0x0
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "11100000", --  504 - 0x1f8  :  224 - 0xe0
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000011", --  514 - 0x202  :    3 - 0x3
    "00001111", --  515 - 0x203  :   15 - 0xf
    "00011111", --  516 - 0x204  :   31 - 0x1f
    "00011111", --  517 - 0x205  :   31 - 0x1f
    "00011100", --  518 - 0x206  :   28 - 0x1c
    "00100100", --  519 - 0x207  :   36 - 0x24
    "00000000", --  520 - 0x208  :    0 - 0x0
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00011111", --  526 - 0x20e  :   31 - 0x1f
    "00111111", --  527 - 0x20f  :   63 - 0x3f
    "00000000", --  528 - 0x210  :    0 - 0x0
    "00000100", --  529 - 0x211  :    4 - 0x4
    "11100110", --  530 - 0x212  :  230 - 0xe6
    "11100000", --  531 - 0x213  :  224 - 0xe0
    "11111111", --  532 - 0x214  :  255 - 0xff
    "11111111", --  533 - 0x215  :  255 - 0xff
    "10001111", --  534 - 0x216  :  143 - 0x8f
    "10000011", --  535 - 0x217  :  131 - 0x83
    "00001110", --  536 - 0x218  :   14 - 0xe
    "00011111", --  537 - 0x219  :   31 - 0x1f
    "00011111", --  538 - 0x21a  :   31 - 0x1f
    "00011111", --  539 - 0x21b  :   31 - 0x1f
    "00011111", --  540 - 0x21c  :   31 - 0x1f
    "00000011", --  541 - 0x21d  :    3 - 0x3
    "11111111", --  542 - 0x21e  :  255 - 0xff
    "11111111", --  543 - 0x21f  :  255 - 0xff
    "00100110", --  544 - 0x220  :   38 - 0x26
    "00100110", --  545 - 0x221  :   38 - 0x26
    "01100000", --  546 - 0x222  :   96 - 0x60
    "01111000", --  547 - 0x223  :  120 - 0x78
    "00011000", --  548 - 0x224  :   24 - 0x18
    "00001111", --  549 - 0x225  :   15 - 0xf
    "01111111", --  550 - 0x226  :  127 - 0x7f
    "11111111", --  551 - 0x227  :  255 - 0xff
    "00111111", --  552 - 0x228  :   63 - 0x3f
    "00111111", --  553 - 0x229  :   63 - 0x3f
    "01111111", --  554 - 0x22a  :  127 - 0x7f
    "01111111", --  555 - 0x22b  :  127 - 0x7f
    "00011111", --  556 - 0x22c  :   31 - 0x1f
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "01111110", --  558 - 0x22e  :  126 - 0x7e
    "11111111", --  559 - 0x22f  :  255 - 0xff
    "00000001", --  560 - 0x230  :    1 - 0x1
    "00100001", --  561 - 0x231  :   33 - 0x21
    "11111110", --  562 - 0x232  :  254 - 0xfe
    "01111010", --  563 - 0x233  :  122 - 0x7a
    "00000110", --  564 - 0x234  :    6 - 0x6
    "11111110", --  565 - 0x235  :  254 - 0xfe
    "11111100", --  566 - 0x236  :  252 - 0xfc
    "11111100", --  567 - 0x237  :  252 - 0xfc
    "11111111", --  568 - 0x238  :  255 - 0xff
    "11111111", --  569 - 0x239  :  255 - 0xff
    "11111110", --  570 - 0x23a  :  254 - 0xfe
    "11111110", --  571 - 0x23b  :  254 - 0xfe
    "11111110", --  572 - 0x23c  :  254 - 0xfe
    "11011110", --  573 - 0x23d  :  222 - 0xde
    "01011100", --  574 - 0x23e  :   92 - 0x5c
    "01101100", --  575 - 0x23f  :  108 - 0x6c
    "11111111", --  576 - 0x240  :  255 - 0xff
    "11001111", --  577 - 0x241  :  207 - 0xcf
    "10000111", --  578 - 0x242  :  135 - 0x87
    "00000111", --  579 - 0x243  :    7 - 0x7
    "00000111", --  580 - 0x244  :    7 - 0x7
    "00001111", --  581 - 0x245  :   15 - 0xf
    "00011111", --  582 - 0x246  :   31 - 0x1f
    "00011111", --  583 - 0x247  :   31 - 0x1f
    "11111111", --  584 - 0x248  :  255 - 0xff
    "11111111", --  585 - 0x249  :  255 - 0xff
    "11111110", --  586 - 0x24a  :  254 - 0xfe
    "11111100", --  587 - 0x24b  :  252 - 0xfc
    "11111000", --  588 - 0x24c  :  248 - 0xf8
    "10110000", --  589 - 0x24d  :  176 - 0xb0
    "01100000", --  590 - 0x24e  :   96 - 0x60
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "11111000", --  592 - 0x250  :  248 - 0xf8
    "11111000", --  593 - 0x251  :  248 - 0xf8
    "11110000", --  594 - 0x252  :  240 - 0xf0
    "10111000", --  595 - 0x253  :  184 - 0xb8
    "11111000", --  596 - 0x254  :  248 - 0xf8
    "11111001", --  597 - 0x255  :  249 - 0xf9
    "11111011", --  598 - 0x256  :  251 - 0xfb
    "11111111", --  599 - 0x257  :  255 - 0xff
    "00101000", --  600 - 0x258  :   40 - 0x28
    "00110000", --  601 - 0x259  :   48 - 0x30
    "00011000", --  602 - 0x25a  :   24 - 0x18
    "01000000", --  603 - 0x25b  :   64 - 0x40
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000001", --  605 - 0x25d  :    1 - 0x1
    "00000011", --  606 - 0x25e  :    3 - 0x3
    "00001111", --  607 - 0x25f  :   15 - 0xf
    "00011111", --  608 - 0x260  :   31 - 0x1f
    "11111111", --  609 - 0x261  :  255 - 0xff
    "11111111", --  610 - 0x262  :  255 - 0xff
    "11111111", --  611 - 0x263  :  255 - 0xff
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111110", --  613 - 0x265  :  254 - 0xfe
    "11000000", --  614 - 0x266  :  192 - 0xc0
    "10000000", --  615 - 0x267  :  128 - 0x80
    "00010000", --  616 - 0x268  :   16 - 0x10
    "11101100", --  617 - 0x269  :  236 - 0xec
    "11100011", --  618 - 0x26a  :  227 - 0xe3
    "11100000", --  619 - 0x26b  :  224 - 0xe0
    "11100000", --  620 - 0x26c  :  224 - 0xe0
    "11100000", --  621 - 0x26d  :  224 - 0xe0
    "11000000", --  622 - 0x26e  :  192 - 0xc0
    "10000000", --  623 - 0x26f  :  128 - 0x80
    "11111111", --  624 - 0x270  :  255 - 0xff
    "11111111", --  625 - 0x271  :  255 - 0xff
    "11111111", --  626 - 0x272  :  255 - 0xff
    "00111111", --  627 - 0x273  :   63 - 0x3f
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000000", --  629 - 0x275  :    0 - 0x0
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00001111", --  632 - 0x278  :   15 - 0xf
    "00001111", --  633 - 0x279  :   15 - 0xf
    "00001111", --  634 - 0x27a  :   15 - 0xf
    "00001111", --  635 - 0x27b  :   15 - 0xf
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00010011", --  640 - 0x280  :   19 - 0x13
    "00110011", --  641 - 0x281  :   51 - 0x33
    "00110000", --  642 - 0x282  :   48 - 0x30
    "00011000", --  643 - 0x283  :   24 - 0x18
    "00000100", --  644 - 0x284  :    4 - 0x4
    "00001111", --  645 - 0x285  :   15 - 0xf
    "00011111", --  646 - 0x286  :   31 - 0x1f
    "00011111", --  647 - 0x287  :   31 - 0x1f
    "00011111", --  648 - 0x288  :   31 - 0x1f
    "00111111", --  649 - 0x289  :   63 - 0x3f
    "00111111", --  650 - 0x28a  :   63 - 0x3f
    "00011111", --  651 - 0x28b  :   31 - 0x1f
    "00000111", --  652 - 0x28c  :    7 - 0x7
    "00001001", --  653 - 0x28d  :    9 - 0x9
    "00010011", --  654 - 0x28e  :   19 - 0x13
    "00010111", --  655 - 0x28f  :   23 - 0x17
    "00000000", --  656 - 0x290  :    0 - 0x0
    "00010000", --  657 - 0x291  :   16 - 0x10
    "01111110", --  658 - 0x292  :  126 - 0x7e
    "00110000", --  659 - 0x293  :   48 - 0x30
    "11100000", --  660 - 0x294  :  224 - 0xe0
    "11110000", --  661 - 0x295  :  240 - 0xf0
    "11110000", --  662 - 0x296  :  240 - 0xf0
    "11100000", --  663 - 0x297  :  224 - 0xe0
    "11111111", --  664 - 0x298  :  255 - 0xff
    "11111111", --  665 - 0x299  :  255 - 0xff
    "11111110", --  666 - 0x29a  :  254 - 0xfe
    "11111111", --  667 - 0x29b  :  255 - 0xff
    "11111110", --  668 - 0x29c  :  254 - 0xfe
    "11111100", --  669 - 0x29d  :  252 - 0xfc
    "11111000", --  670 - 0x29e  :  248 - 0xf8
    "11100000", --  671 - 0x29f  :  224 - 0xe0
    "00011111", --  672 - 0x2a0  :   31 - 0x1f
    "00011111", --  673 - 0x2a1  :   31 - 0x1f
    "00001111", --  674 - 0x2a2  :   15 - 0xf
    "00001111", --  675 - 0x2a3  :   15 - 0xf
    "00001111", --  676 - 0x2a4  :   15 - 0xf
    "00011111", --  677 - 0x2a5  :   31 - 0x1f
    "00011111", --  678 - 0x2a6  :   31 - 0x1f
    "00011111", --  679 - 0x2a7  :   31 - 0x1f
    "00010111", --  680 - 0x2a8  :   23 - 0x17
    "00010111", --  681 - 0x2a9  :   23 - 0x17
    "00000011", --  682 - 0x2aa  :    3 - 0x3
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "00000000", --  686 - 0x2ae  :    0 - 0x0
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "11110000", --  688 - 0x2b0  :  240 - 0xf0
    "11110000", --  689 - 0x2b1  :  240 - 0xf0
    "11111000", --  690 - 0x2b2  :  248 - 0xf8
    "11111000", --  691 - 0x2b3  :  248 - 0xf8
    "10111000", --  692 - 0x2b4  :  184 - 0xb8
    "11111000", --  693 - 0x2b5  :  248 - 0xf8
    "11111000", --  694 - 0x2b6  :  248 - 0xf8
    "11111000", --  695 - 0x2b7  :  248 - 0xf8
    "11010000", --  696 - 0x2b8  :  208 - 0xd0
    "10010000", --  697 - 0x2b9  :  144 - 0x90
    "00011000", --  698 - 0x2ba  :   24 - 0x18
    "00001000", --  699 - 0x2bb  :    8 - 0x8
    "01000000", --  700 - 0x2bc  :   64 - 0x40
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00111111", --  704 - 0x2c0  :   63 - 0x3f
    "11111111", --  705 - 0x2c1  :  255 - 0xff
    "11111111", --  706 - 0x2c2  :  255 - 0xff
    "11111111", --  707 - 0x2c3  :  255 - 0xff
    "11110110", --  708 - 0x2c4  :  246 - 0xf6
    "11000110", --  709 - 0x2c5  :  198 - 0xc6
    "10000100", --  710 - 0x2c6  :  132 - 0x84
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00110000", --  712 - 0x2c8  :   48 - 0x30
    "11110000", --  713 - 0x2c9  :  240 - 0xf0
    "11110000", --  714 - 0x2ca  :  240 - 0xf0
    "11110001", --  715 - 0x2cb  :  241 - 0xf1
    "11110110", --  716 - 0x2cc  :  246 - 0xf6
    "11000110", --  717 - 0x2cd  :  198 - 0xc6
    "10000100", --  718 - 0x2ce  :  132 - 0x84
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "11110000", --  720 - 0x2d0  :  240 - 0xf0
    "11100000", --  721 - 0x2d1  :  224 - 0xe0
    "10000000", --  722 - 0x2d2  :  128 - 0x80
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00011111", --  736 - 0x2e0  :   31 - 0x1f
    "00011111", --  737 - 0x2e1  :   31 - 0x1f
    "00111111", --  738 - 0x2e2  :   63 - 0x3f
    "00111111", --  739 - 0x2e3  :   63 - 0x3f
    "00011111", --  740 - 0x2e4  :   31 - 0x1f
    "00001111", --  741 - 0x2e5  :   15 - 0xf
    "00001111", --  742 - 0x2e6  :   15 - 0xf
    "00011111", --  743 - 0x2e7  :   31 - 0x1f
    "00011111", --  744 - 0x2e8  :   31 - 0x1f
    "00011111", --  745 - 0x2e9  :   31 - 0x1f
    "00111111", --  746 - 0x2ea  :   63 - 0x3f
    "00111110", --  747 - 0x2eb  :   62 - 0x3e
    "01111100", --  748 - 0x2ec  :  124 - 0x7c
    "01111000", --  749 - 0x2ed  :  120 - 0x78
    "11110000", --  750 - 0x2ee  :  240 - 0xf0
    "11100000", --  751 - 0x2ef  :  224 - 0xe0
    "11110000", --  752 - 0x2f0  :  240 - 0xf0
    "11110000", --  753 - 0x2f1  :  240 - 0xf0
    "11111000", --  754 - 0x2f2  :  248 - 0xf8
    "11111000", --  755 - 0x2f3  :  248 - 0xf8
    "10111000", --  756 - 0x2f4  :  184 - 0xb8
    "11111000", --  757 - 0x2f5  :  248 - 0xf8
    "11111000", --  758 - 0x2f6  :  248 - 0xf8
    "11110000", --  759 - 0x2f7  :  240 - 0xf0
    "10110000", --  760 - 0x2f8  :  176 - 0xb0
    "10010000", --  761 - 0x2f9  :  144 - 0x90
    "00011000", --  762 - 0x2fa  :   24 - 0x18
    "00001000", --  763 - 0x2fb  :    8 - 0x8
    "01000000", --  764 - 0x2fc  :   64 - 0x40
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "11100000", --  768 - 0x300  :  224 - 0xe0
    "11110000", --  769 - 0x301  :  240 - 0xf0
    "11110000", --  770 - 0x302  :  240 - 0xf0
    "11110000", --  771 - 0x303  :  240 - 0xf0
    "11110000", --  772 - 0x304  :  240 - 0xf0
    "11110000", --  773 - 0x305  :  240 - 0xf0
    "11111000", --  774 - 0x306  :  248 - 0xf8
    "11110000", --  775 - 0x307  :  240 - 0xf0
    "11000000", --  776 - 0x308  :  192 - 0xc0
    "11100000", --  777 - 0x309  :  224 - 0xe0
    "11111100", --  778 - 0x30a  :  252 - 0xfc
    "11111110", --  779 - 0x30b  :  254 - 0xfe
    "11111111", --  780 - 0x30c  :  255 - 0xff
    "01111111", --  781 - 0x30d  :  127 - 0x7f
    "00000011", --  782 - 0x30e  :    3 - 0x3
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00011111", --  784 - 0x310  :   31 - 0x1f
    "00011111", --  785 - 0x311  :   31 - 0x1f
    "00011111", --  786 - 0x312  :   31 - 0x1f
    "00111111", --  787 - 0x313  :   63 - 0x3f
    "00111110", --  788 - 0x314  :   62 - 0x3e
    "00111100", --  789 - 0x315  :   60 - 0x3c
    "00111000", --  790 - 0x316  :   56 - 0x38
    "00011000", --  791 - 0x317  :   24 - 0x18
    "00000000", --  792 - 0x318  :    0 - 0x0
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00010000", --  794 - 0x31a  :   16 - 0x10
    "00111000", --  795 - 0x31b  :   56 - 0x38
    "00111110", --  796 - 0x31c  :   62 - 0x3e
    "00111100", --  797 - 0x31d  :   60 - 0x3c
    "00111000", --  798 - 0x31e  :   56 - 0x38
    "00011000", --  799 - 0x31f  :   24 - 0x18
    "00000000", --  800 - 0x320  :    0 - 0x0
    "00000011", --  801 - 0x321  :    3 - 0x3
    "00000111", --  802 - 0x322  :    7 - 0x7
    "00000111", --  803 - 0x323  :    7 - 0x7
    "00001010", --  804 - 0x324  :   10 - 0xa
    "00001011", --  805 - 0x325  :   11 - 0xb
    "00001100", --  806 - 0x326  :   12 - 0xc
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000111", --  811 - 0x32b  :    7 - 0x7
    "00001111", --  812 - 0x32c  :   15 - 0xf
    "00001111", --  813 - 0x32d  :   15 - 0xf
    "00001111", --  814 - 0x32e  :   15 - 0xf
    "00000011", --  815 - 0x32f  :    3 - 0x3
    "00000000", --  816 - 0x330  :    0 - 0x0
    "11100000", --  817 - 0x331  :  224 - 0xe0
    "11111100", --  818 - 0x332  :  252 - 0xfc
    "00100000", --  819 - 0x333  :   32 - 0x20
    "00100000", --  820 - 0x334  :   32 - 0x20
    "00010000", --  821 - 0x335  :   16 - 0x10
    "00111100", --  822 - 0x336  :   60 - 0x3c
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000000", --  824 - 0x338  :    0 - 0x0
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "11110000", --  827 - 0x33b  :  240 - 0xf0
    "11111100", --  828 - 0x33c  :  252 - 0xfc
    "11111110", --  829 - 0x33d  :  254 - 0xfe
    "11111100", --  830 - 0x33e  :  252 - 0xfc
    "11111000", --  831 - 0x33f  :  248 - 0xf8
    "00000111", --  832 - 0x340  :    7 - 0x7
    "00000111", --  833 - 0x341  :    7 - 0x7
    "00000111", --  834 - 0x342  :    7 - 0x7
    "00011111", --  835 - 0x343  :   31 - 0x1f
    "00011111", --  836 - 0x344  :   31 - 0x1f
    "00111110", --  837 - 0x345  :   62 - 0x3e
    "00100001", --  838 - 0x346  :   33 - 0x21
    "00000001", --  839 - 0x347  :    1 - 0x1
    "00000111", --  840 - 0x348  :    7 - 0x7
    "00001111", --  841 - 0x349  :   15 - 0xf
    "00011011", --  842 - 0x34a  :   27 - 0x1b
    "00011000", --  843 - 0x34b  :   24 - 0x18
    "00010000", --  844 - 0x34c  :   16 - 0x10
    "00110000", --  845 - 0x34d  :   48 - 0x30
    "00100001", --  846 - 0x34e  :   33 - 0x21
    "00000001", --  847 - 0x34f  :    1 - 0x1
    "11100000", --  848 - 0x350  :  224 - 0xe0
    "11100000", --  849 - 0x351  :  224 - 0xe0
    "11100000", --  850 - 0x352  :  224 - 0xe0
    "11110000", --  851 - 0x353  :  240 - 0xf0
    "11110000", --  852 - 0x354  :  240 - 0xf0
    "11100000", --  853 - 0x355  :  224 - 0xe0
    "11000000", --  854 - 0x356  :  192 - 0xc0
    "11100000", --  855 - 0x357  :  224 - 0xe0
    "10101000", --  856 - 0x358  :  168 - 0xa8
    "11111100", --  857 - 0x359  :  252 - 0xfc
    "11111000", --  858 - 0x35a  :  248 - 0xf8
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "11000000", --  862 - 0x35e  :  192 - 0xc0
    "11100000", --  863 - 0x35f  :  224 - 0xe0
    "00000111", --  864 - 0x360  :    7 - 0x7
    "00001111", --  865 - 0x361  :   15 - 0xf
    "00001110", --  866 - 0x362  :   14 - 0xe
    "00010100", --  867 - 0x363  :   20 - 0x14
    "00010110", --  868 - 0x364  :   22 - 0x16
    "00011000", --  869 - 0x365  :   24 - 0x18
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00111111", --  871 - 0x367  :   63 - 0x3f
    "00000000", --  872 - 0x368  :    0 - 0x0
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00001111", --  874 - 0x36a  :   15 - 0xf
    "00011111", --  875 - 0x36b  :   31 - 0x1f
    "00011111", --  876 - 0x36c  :   31 - 0x1f
    "00011111", --  877 - 0x36d  :   31 - 0x1f
    "00000111", --  878 - 0x36e  :    7 - 0x7
    "00111100", --  879 - 0x36f  :   60 - 0x3c
    "11000000", --  880 - 0x370  :  192 - 0xc0
    "11111000", --  881 - 0x371  :  248 - 0xf8
    "01000000", --  882 - 0x372  :   64 - 0x40
    "01000000", --  883 - 0x373  :   64 - 0x40
    "00100000", --  884 - 0x374  :   32 - 0x20
    "01111000", --  885 - 0x375  :  120 - 0x78
    "00000000", --  886 - 0x376  :    0 - 0x0
    "11000000", --  887 - 0x377  :  192 - 0xc0
    "00000000", --  888 - 0x378  :    0 - 0x0
    "00000000", --  889 - 0x379  :    0 - 0x0
    "11100000", --  890 - 0x37a  :  224 - 0xe0
    "11111000", --  891 - 0x37b  :  248 - 0xf8
    "11111100", --  892 - 0x37c  :  252 - 0xfc
    "11111000", --  893 - 0x37d  :  248 - 0xf8
    "11110000", --  894 - 0x37e  :  240 - 0xf0
    "11000000", --  895 - 0x37f  :  192 - 0xc0
    "00111111", --  896 - 0x380  :   63 - 0x3f
    "00001110", --  897 - 0x381  :   14 - 0xe
    "00001111", --  898 - 0x382  :   15 - 0xf
    "00011111", --  899 - 0x383  :   31 - 0x1f
    "00111111", --  900 - 0x384  :   63 - 0x3f
    "01111100", --  901 - 0x385  :  124 - 0x7c
    "01110000", --  902 - 0x386  :  112 - 0x70
    "00111000", --  903 - 0x387  :   56 - 0x38
    "11111100", --  904 - 0x388  :  252 - 0xfc
    "11101101", --  905 - 0x389  :  237 - 0xed
    "11000000", --  906 - 0x38a  :  192 - 0xc0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "01100000", --  909 - 0x38d  :   96 - 0x60
    "01110000", --  910 - 0x38e  :  112 - 0x70
    "00111000", --  911 - 0x38f  :   56 - 0x38
    "11110000", --  912 - 0x390  :  240 - 0xf0
    "11111000", --  913 - 0x391  :  248 - 0xf8
    "11100100", --  914 - 0x392  :  228 - 0xe4
    "11111100", --  915 - 0x393  :  252 - 0xfc
    "11111100", --  916 - 0x394  :  252 - 0xfc
    "01111100", --  917 - 0x395  :  124 - 0x7c
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "01111110", --  920 - 0x398  :  126 - 0x7e
    "00011110", --  921 - 0x399  :   30 - 0x1e
    "00000100", --  922 - 0x39a  :    4 - 0x4
    "00001100", --  923 - 0x39b  :   12 - 0xc
    "00001100", --  924 - 0x39c  :   12 - 0xc
    "00001100", --  925 - 0x39d  :   12 - 0xc
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000111", --  928 - 0x3a0  :    7 - 0x7
    "00001111", --  929 - 0x3a1  :   15 - 0xf
    "00001110", --  930 - 0x3a2  :   14 - 0xe
    "00010100", --  931 - 0x3a3  :   20 - 0x14
    "00010110", --  932 - 0x3a4  :   22 - 0x16
    "00011000", --  933 - 0x3a5  :   24 - 0x18
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00001111", --  935 - 0x3a7  :   15 - 0xf
    "00000000", --  936 - 0x3a8  :    0 - 0x0
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00001111", --  938 - 0x3aa  :   15 - 0xf
    "00011111", --  939 - 0x3ab  :   31 - 0x1f
    "00011111", --  940 - 0x3ac  :   31 - 0x1f
    "00011111", --  941 - 0x3ad  :   31 - 0x1f
    "00000111", --  942 - 0x3ae  :    7 - 0x7
    "00001101", --  943 - 0x3af  :   13 - 0xd
    "00011111", --  944 - 0x3b0  :   31 - 0x1f
    "00011111", --  945 - 0x3b1  :   31 - 0x1f
    "00011111", --  946 - 0x3b2  :   31 - 0x1f
    "00011100", --  947 - 0x3b3  :   28 - 0x1c
    "00001100", --  948 - 0x3b4  :   12 - 0xc
    "00000111", --  949 - 0x3b5  :    7 - 0x7
    "00000111", --  950 - 0x3b6  :    7 - 0x7
    "00000111", --  951 - 0x3b7  :    7 - 0x7
    "00011110", --  952 - 0x3b8  :   30 - 0x1e
    "00011100", --  953 - 0x3b9  :   28 - 0x1c
    "00011110", --  954 - 0x3ba  :   30 - 0x1e
    "00001111", --  955 - 0x3bb  :   15 - 0xf
    "00000111", --  956 - 0x3bc  :    7 - 0x7
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000111", --  958 - 0x3be  :    7 - 0x7
    "00000111", --  959 - 0x3bf  :    7 - 0x7
    "11100000", --  960 - 0x3c0  :  224 - 0xe0
    "01100000", --  961 - 0x3c1  :   96 - 0x60
    "11110000", --  962 - 0x3c2  :  240 - 0xf0
    "01110000", --  963 - 0x3c3  :  112 - 0x70
    "11100000", --  964 - 0x3c4  :  224 - 0xe0
    "11100000", --  965 - 0x3c5  :  224 - 0xe0
    "11110000", --  966 - 0x3c6  :  240 - 0xf0
    "10000000", --  967 - 0x3c7  :  128 - 0x80
    "01100000", --  968 - 0x3c8  :   96 - 0x60
    "10010000", --  969 - 0x3c9  :  144 - 0x90
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "10000000", --  971 - 0x3cb  :  128 - 0x80
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "11100000", --  973 - 0x3cd  :  224 - 0xe0
    "11110000", --  974 - 0x3ce  :  240 - 0xf0
    "10000000", --  975 - 0x3cf  :  128 - 0x80
    "00000111", --  976 - 0x3d0  :    7 - 0x7
    "00011111", --  977 - 0x3d1  :   31 - 0x1f
    "00111111", --  978 - 0x3d2  :   63 - 0x3f
    "00010010", --  979 - 0x3d3  :   18 - 0x12
    "00010011", --  980 - 0x3d4  :   19 - 0x13
    "00001000", --  981 - 0x3d5  :    8 - 0x8
    "00011111", --  982 - 0x3d6  :   31 - 0x1f
    "00110001", --  983 - 0x3d7  :   49 - 0x31
    "00000000", --  984 - 0x3d8  :    0 - 0x0
    "00010000", --  985 - 0x3d9  :   16 - 0x10
    "00111111", --  986 - 0x3da  :   63 - 0x3f
    "01111111", --  987 - 0x3db  :  127 - 0x7f
    "01111111", --  988 - 0x3dc  :  127 - 0x7f
    "00111111", --  989 - 0x3dd  :   63 - 0x3f
    "00000011", --  990 - 0x3de  :    3 - 0x3
    "00001111", --  991 - 0x3df  :   15 - 0xf
    "11000000", --  992 - 0x3e0  :  192 - 0xc0
    "11110000", --  993 - 0x3e1  :  240 - 0xf0
    "01000000", --  994 - 0x3e2  :   64 - 0x40
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00110000", --  996 - 0x3e4  :   48 - 0x30
    "00011000", --  997 - 0x3e5  :   24 - 0x18
    "11000000", --  998 - 0x3e6  :  192 - 0xc0
    "11111000", --  999 - 0x3e7  :  248 - 0xf8
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "11100000", -- 1002 - 0x3ea  :  224 - 0xe0
    "11111000", -- 1003 - 0x3eb  :  248 - 0xf8
    "11111100", -- 1004 - 0x3ec  :  252 - 0xfc
    "11111000", -- 1005 - 0x3ed  :  248 - 0xf8
    "10110000", -- 1006 - 0x3ee  :  176 - 0xb0
    "00111000", -- 1007 - 0x3ef  :   56 - 0x38
    "00110001", -- 1008 - 0x3f0  :   49 - 0x31
    "00111001", -- 1009 - 0x3f1  :   57 - 0x39
    "00011111", -- 1010 - 0x3f2  :   31 - 0x1f
    "00011111", -- 1011 - 0x3f3  :   31 - 0x1f
    "00001111", -- 1012 - 0x3f4  :   15 - 0xf
    "01011111", -- 1013 - 0x3f5  :   95 - 0x5f
    "01111110", -- 1014 - 0x3f6  :  126 - 0x7e
    "00111100", -- 1015 - 0x3f7  :   60 - 0x3c
    "00011111", -- 1016 - 0x3f8  :   31 - 0x1f
    "00000111", -- 1017 - 0x3f9  :    7 - 0x7
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00001110", -- 1019 - 0x3fb  :   14 - 0xe
    "00001111", -- 1020 - 0x3fc  :   15 - 0xf
    "01010011", -- 1021 - 0x3fd  :   83 - 0x53
    "01111100", -- 1022 - 0x3fe  :  124 - 0x7c
    "00111100", -- 1023 - 0x3ff  :   60 - 0x3c
    "11111000", -- 1024 - 0x400  :  248 - 0xf8
    "11111000", -- 1025 - 0x401  :  248 - 0xf8
    "11110000", -- 1026 - 0x402  :  240 - 0xf0
    "11100000", -- 1027 - 0x403  :  224 - 0xe0
    "11100000", -- 1028 - 0x404  :  224 - 0xe0
    "11000000", -- 1029 - 0x405  :  192 - 0xc0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "11111000", -- 1032 - 0x408  :  248 - 0xf8
    "11111000", -- 1033 - 0x409  :  248 - 0xf8
    "11110000", -- 1034 - 0x40a  :  240 - 0xf0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "10000000", -- 1037 - 0x40d  :  128 - 0x80
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0
    "11100000", -- 1041 - 0x411  :  224 - 0xe0
    "11111100", -- 1042 - 0x412  :  252 - 0xfc
    "00100111", -- 1043 - 0x413  :   39 - 0x27
    "00100111", -- 1044 - 0x414  :   39 - 0x27
    "00010001", -- 1045 - 0x415  :   17 - 0x11
    "00111110", -- 1046 - 0x416  :   62 - 0x3e
    "00000100", -- 1047 - 0x417  :    4 - 0x4
    "00000111", -- 1048 - 0x418  :    7 - 0x7
    "00000111", -- 1049 - 0x419  :    7 - 0x7
    "00000011", -- 1050 - 0x41a  :    3 - 0x3
    "11110111", -- 1051 - 0x41b  :  247 - 0xf7
    "11111111", -- 1052 - 0x41c  :  255 - 0xff
    "11111111", -- 1053 - 0x41d  :  255 - 0xff
    "11111110", -- 1054 - 0x41e  :  254 - 0xfe
    "11111100", -- 1055 - 0x41f  :  252 - 0xfc
    "00111111", -- 1056 - 0x420  :   63 - 0x3f
    "01111111", -- 1057 - 0x421  :  127 - 0x7f
    "00111111", -- 1058 - 0x422  :   63 - 0x3f
    "00001111", -- 1059 - 0x423  :   15 - 0xf
    "00011111", -- 1060 - 0x424  :   31 - 0x1f
    "00111111", -- 1061 - 0x425  :   63 - 0x3f
    "01111111", -- 1062 - 0x426  :  127 - 0x7f
    "01001111", -- 1063 - 0x427  :   79 - 0x4f
    "00111110", -- 1064 - 0x428  :   62 - 0x3e
    "01111111", -- 1065 - 0x429  :  127 - 0x7f
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "11100010", -- 1067 - 0x42b  :  226 - 0xe2
    "01010000", -- 1068 - 0x42c  :   80 - 0x50
    "00111000", -- 1069 - 0x42d  :   56 - 0x38
    "01110000", -- 1070 - 0x42e  :  112 - 0x70
    "01000000", -- 1071 - 0x42f  :   64 - 0x40
    "11111000", -- 1072 - 0x430  :  248 - 0xf8
    "11111001", -- 1073 - 0x431  :  249 - 0xf9
    "11111001", -- 1074 - 0x432  :  249 - 0xf9
    "10110111", -- 1075 - 0x433  :  183 - 0xb7
    "11111111", -- 1076 - 0x434  :  255 - 0xff
    "11111111", -- 1077 - 0x435  :  255 - 0xff
    "11100000", -- 1078 - 0x436  :  224 - 0xe0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "11101000", -- 1080 - 0x438  :  232 - 0xe8
    "01110001", -- 1081 - 0x439  :  113 - 0x71
    "00000001", -- 1082 - 0x43a  :    1 - 0x1
    "01001011", -- 1083 - 0x43b  :   75 - 0x4b
    "00000011", -- 1084 - 0x43c  :    3 - 0x3
    "00000011", -- 1085 - 0x43d  :    3 - 0x3
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000111", -- 1088 - 0x440  :    7 - 0x7
    "00000111", -- 1089 - 0x441  :    7 - 0x7
    "00001111", -- 1090 - 0x442  :   15 - 0xf
    "00111111", -- 1091 - 0x443  :   63 - 0x3f
    "00111111", -- 1092 - 0x444  :   63 - 0x3f
    "00111111", -- 1093 - 0x445  :   63 - 0x3f
    "00100110", -- 1094 - 0x446  :   38 - 0x26
    "00000100", -- 1095 - 0x447  :    4 - 0x4
    "00000101", -- 1096 - 0x448  :    5 - 0x5
    "00000011", -- 1097 - 0x449  :    3 - 0x3
    "00000001", -- 1098 - 0x44a  :    1 - 0x1
    "00110000", -- 1099 - 0x44b  :   48 - 0x30
    "00110000", -- 1100 - 0x44c  :   48 - 0x30
    "00110000", -- 1101 - 0x44d  :   48 - 0x30
    "00100110", -- 1102 - 0x44e  :   38 - 0x26
    "00000100", -- 1103 - 0x44f  :    4 - 0x4
    "11110000", -- 1104 - 0x450  :  240 - 0xf0
    "11110000", -- 1105 - 0x451  :  240 - 0xf0
    "11110000", -- 1106 - 0x452  :  240 - 0xf0
    "11100000", -- 1107 - 0x453  :  224 - 0xe0
    "11000000", -- 1108 - 0x454  :  192 - 0xc0
    "00000000", -- 1109 - 0x455  :    0 - 0x0
    "00000000", -- 1110 - 0x456  :    0 - 0x0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "11111110", -- 1112 - 0x458  :  254 - 0xfe
    "11111100", -- 1113 - 0x459  :  252 - 0xfc
    "11100000", -- 1114 - 0x45a  :  224 - 0xe0
    "00000000", -- 1115 - 0x45b  :    0 - 0x0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00000000", -- 1117 - 0x45d  :    0 - 0x0
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000111", -- 1120 - 0x460  :    7 - 0x7
    "00000111", -- 1121 - 0x461  :    7 - 0x7
    "00001111", -- 1122 - 0x462  :   15 - 0xf
    "00011111", -- 1123 - 0x463  :   31 - 0x1f
    "00111111", -- 1124 - 0x464  :   63 - 0x3f
    "00001111", -- 1125 - 0x465  :   15 - 0xf
    "00011100", -- 1126 - 0x466  :   28 - 0x1c
    "00011000", -- 1127 - 0x467  :   24 - 0x18
    "00000101", -- 1128 - 0x468  :    5 - 0x5
    "00000011", -- 1129 - 0x469  :    3 - 0x3
    "00000001", -- 1130 - 0x46a  :    1 - 0x1
    "00010000", -- 1131 - 0x46b  :   16 - 0x10
    "00110000", -- 1132 - 0x46c  :   48 - 0x30
    "00001100", -- 1133 - 0x46d  :   12 - 0xc
    "00011100", -- 1134 - 0x46e  :   28 - 0x1c
    "00011000", -- 1135 - 0x46f  :   24 - 0x18
    "11100000", -- 1136 - 0x470  :  224 - 0xe0
    "11100000", -- 1137 - 0x471  :  224 - 0xe0
    "11100000", -- 1138 - 0x472  :  224 - 0xe0
    "11100000", -- 1139 - 0x473  :  224 - 0xe0
    "11000000", -- 1140 - 0x474  :  192 - 0xc0
    "10000000", -- 1141 - 0x475  :  128 - 0x80
    "00000000", -- 1142 - 0x476  :    0 - 0x0
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "11000000", -- 1144 - 0x478  :  192 - 0xc0
    "11100000", -- 1145 - 0x479  :  224 - 0xe0
    "11110000", -- 1146 - 0x47a  :  240 - 0xf0
    "01111000", -- 1147 - 0x47b  :  120 - 0x78
    "00011000", -- 1148 - 0x47c  :   24 - 0x18
    "00001000", -- 1149 - 0x47d  :    8 - 0x8
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000111", -- 1152 - 0x480  :    7 - 0x7
    "00001111", -- 1153 - 0x481  :   15 - 0xf
    "00011111", -- 1154 - 0x482  :   31 - 0x1f
    "00001111", -- 1155 - 0x483  :   15 - 0xf
    "00111111", -- 1156 - 0x484  :   63 - 0x3f
    "00001111", -- 1157 - 0x485  :   15 - 0xf
    "00011100", -- 1158 - 0x486  :   28 - 0x1c
    "00011000", -- 1159 - 0x487  :   24 - 0x18
    "00000111", -- 1160 - 0x488  :    7 - 0x7
    "00001111", -- 1161 - 0x489  :   15 - 0xf
    "00111110", -- 1162 - 0x48a  :   62 - 0x3e
    "01111100", -- 1163 - 0x48b  :  124 - 0x7c
    "00110000", -- 1164 - 0x48c  :   48 - 0x30
    "00001100", -- 1165 - 0x48d  :   12 - 0xc
    "00011100", -- 1166 - 0x48e  :   28 - 0x1c
    "00011000", -- 1167 - 0x48f  :   24 - 0x18
    "11100000", -- 1168 - 0x490  :  224 - 0xe0
    "11100000", -- 1169 - 0x491  :  224 - 0xe0
    "11100000", -- 1170 - 0x492  :  224 - 0xe0
    "01000000", -- 1171 - 0x493  :   64 - 0x40
    "11000000", -- 1172 - 0x494  :  192 - 0xc0
    "10000000", -- 1173 - 0x495  :  128 - 0x80
    "00000000", -- 1174 - 0x496  :    0 - 0x0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "01100000", -- 1176 - 0x498  :   96 - 0x60
    "01100000", -- 1177 - 0x499  :   96 - 0x60
    "01100000", -- 1178 - 0x49a  :   96 - 0x60
    "10000000", -- 1179 - 0x49b  :  128 - 0x80
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "01111111", -- 1184 - 0x4a0  :  127 - 0x7f
    "11111111", -- 1185 - 0x4a1  :  255 - 0xff
    "11111111", -- 1186 - 0x4a2  :  255 - 0xff
    "11111011", -- 1187 - 0x4a3  :  251 - 0xfb
    "00001111", -- 1188 - 0x4a4  :   15 - 0xf
    "00001111", -- 1189 - 0x4a5  :   15 - 0xf
    "00001111", -- 1190 - 0x4a6  :   15 - 0xf
    "00011111", -- 1191 - 0x4a7  :   31 - 0x1f
    "01110011", -- 1192 - 0x4a8  :  115 - 0x73
    "11110011", -- 1193 - 0x4a9  :  243 - 0xf3
    "11110000", -- 1194 - 0x4aa  :  240 - 0xf0
    "11110100", -- 1195 - 0x4ab  :  244 - 0xf4
    "11110000", -- 1196 - 0x4ac  :  240 - 0xf0
    "11110000", -- 1197 - 0x4ad  :  240 - 0xf0
    "01110000", -- 1198 - 0x4ae  :  112 - 0x70
    "01100000", -- 1199 - 0x4af  :   96 - 0x60
    "00111111", -- 1200 - 0x4b0  :   63 - 0x3f
    "01111110", -- 1201 - 0x4b1  :  126 - 0x7e
    "01111100", -- 1202 - 0x4b2  :  124 - 0x7c
    "01111100", -- 1203 - 0x4b3  :  124 - 0x7c
    "00111100", -- 1204 - 0x4b4  :   60 - 0x3c
    "00111100", -- 1205 - 0x4b5  :   60 - 0x3c
    "11111100", -- 1206 - 0x4b6  :  252 - 0xfc
    "11111100", -- 1207 - 0x4b7  :  252 - 0xfc
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "00111100", -- 1212 - 0x4bc  :   60 - 0x3c
    "00111100", -- 1213 - 0x4bd  :   60 - 0x3c
    "11111100", -- 1214 - 0x4be  :  252 - 0xfc
    "11111100", -- 1215 - 0x4bf  :  252 - 0xfc
    "01100000", -- 1216 - 0x4c0  :   96 - 0x60
    "01110000", -- 1217 - 0x4c1  :  112 - 0x70
    "00011000", -- 1218 - 0x4c2  :   24 - 0x18
    "00001000", -- 1219 - 0x4c3  :    8 - 0x8
    "00001111", -- 1220 - 0x4c4  :   15 - 0xf
    "00011111", -- 1221 - 0x4c5  :   31 - 0x1f
    "00111111", -- 1222 - 0x4c6  :   63 - 0x3f
    "01111111", -- 1223 - 0x4c7  :  127 - 0x7f
    "01111111", -- 1224 - 0x4c8  :  127 - 0x7f
    "01111111", -- 1225 - 0x4c9  :  127 - 0x7f
    "00011111", -- 1226 - 0x4ca  :   31 - 0x1f
    "00000111", -- 1227 - 0x4cb  :    7 - 0x7
    "00001011", -- 1228 - 0x4cc  :   11 - 0xb
    "00011011", -- 1229 - 0x4cd  :   27 - 0x1b
    "00111011", -- 1230 - 0x4ce  :   59 - 0x3b
    "01111011", -- 1231 - 0x4cf  :  123 - 0x7b
    "11111100", -- 1232 - 0x4d0  :  252 - 0xfc
    "01111100", -- 1233 - 0x4d1  :  124 - 0x7c
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00100000", -- 1235 - 0x4d3  :   32 - 0x20
    "11110000", -- 1236 - 0x4d4  :  240 - 0xf0
    "11111000", -- 1237 - 0x4d5  :  248 - 0xf8
    "11111100", -- 1238 - 0x4d6  :  252 - 0xfc
    "11111110", -- 1239 - 0x4d7  :  254 - 0xfe
    "11111100", -- 1240 - 0x4d8  :  252 - 0xfc
    "11111100", -- 1241 - 0x4d9  :  252 - 0xfc
    "11111000", -- 1242 - 0x4da  :  248 - 0xf8
    "11100000", -- 1243 - 0x4db  :  224 - 0xe0
    "11010000", -- 1244 - 0x4dc  :  208 - 0xd0
    "11011000", -- 1245 - 0x4dd  :  216 - 0xd8
    "11011100", -- 1246 - 0x4de  :  220 - 0xdc
    "11011110", -- 1247 - 0x4df  :  222 - 0xde
    "00001011", -- 1248 - 0x4e0  :   11 - 0xb
    "00001111", -- 1249 - 0x4e1  :   15 - 0xf
    "00011111", -- 1250 - 0x4e2  :   31 - 0x1f
    "00011110", -- 1251 - 0x4e3  :   30 - 0x1e
    "00111100", -- 1252 - 0x4e4  :   60 - 0x3c
    "00111100", -- 1253 - 0x4e5  :   60 - 0x3c
    "00111100", -- 1254 - 0x4e6  :   60 - 0x3c
    "01111100", -- 1255 - 0x4e7  :  124 - 0x7c
    "11000100", -- 1256 - 0x4e8  :  196 - 0xc4
    "11100000", -- 1257 - 0x4e9  :  224 - 0xe0
    "11100000", -- 1258 - 0x4ea  :  224 - 0xe0
    "01000000", -- 1259 - 0x4eb  :   64 - 0x40
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00111100", -- 1261 - 0x4ed  :   60 - 0x3c
    "00111100", -- 1262 - 0x4ee  :   60 - 0x3c
    "01111100", -- 1263 - 0x4ef  :  124 - 0x7c
    "00011111", -- 1264 - 0x4f0  :   31 - 0x1f
    "00111111", -- 1265 - 0x4f1  :   63 - 0x3f
    "00001101", -- 1266 - 0x4f2  :   13 - 0xd
    "00000111", -- 1267 - 0x4f3  :    7 - 0x7
    "00001111", -- 1268 - 0x4f4  :   15 - 0xf
    "00001110", -- 1269 - 0x4f5  :   14 - 0xe
    "00011100", -- 1270 - 0x4f6  :   28 - 0x1c
    "00111100", -- 1271 - 0x4f7  :   60 - 0x3c
    "00011101", -- 1272 - 0x4f8  :   29 - 0x1d
    "00111100", -- 1273 - 0x4f9  :   60 - 0x3c
    "00111010", -- 1274 - 0x4fa  :   58 - 0x3a
    "00111000", -- 1275 - 0x4fb  :   56 - 0x38
    "00110000", -- 1276 - 0x4fc  :   48 - 0x30
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00011100", -- 1278 - 0x4fe  :   28 - 0x1c
    "00111100", -- 1279 - 0x4ff  :   60 - 0x3c
    "00000000", -- 1280 - 0x500  :    0 - 0x0
    "00000000", -- 1281 - 0x501  :    0 - 0x0
    "00000000", -- 1282 - 0x502  :    0 - 0x0
    "00000000", -- 1283 - 0x503  :    0 - 0x0
    "00000000", -- 1284 - 0x504  :    0 - 0x0
    "00000000", -- 1285 - 0x505  :    0 - 0x0
    "00000000", -- 1286 - 0x506  :    0 - 0x0
    "00000000", -- 1287 - 0x507  :    0 - 0x0
    "00100010", -- 1288 - 0x508  :   34 - 0x22
    "01010101", -- 1289 - 0x509  :   85 - 0x55
    "01010101", -- 1290 - 0x50a  :   85 - 0x55
    "01010101", -- 1291 - 0x50b  :   85 - 0x55
    "01010101", -- 1292 - 0x50c  :   85 - 0x55
    "01010101", -- 1293 - 0x50d  :   85 - 0x55
    "01110111", -- 1294 - 0x50e  :  119 - 0x77
    "00100010", -- 1295 - 0x50f  :   34 - 0x22
    "00000000", -- 1296 - 0x510  :    0 - 0x0
    "00000111", -- 1297 - 0x511  :    7 - 0x7
    "00011111", -- 1298 - 0x512  :   31 - 0x1f
    "11111111", -- 1299 - 0x513  :  255 - 0xff
    "00000111", -- 1300 - 0x514  :    7 - 0x7
    "00011111", -- 1301 - 0x515  :   31 - 0x1f
    "00001111", -- 1302 - 0x516  :   15 - 0xf
    "00000110", -- 1303 - 0x517  :    6 - 0x6
    "00000000", -- 1304 - 0x518  :    0 - 0x0
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "00000000", -- 1306 - 0x51a  :    0 - 0x0
    "00000000", -- 1307 - 0x51b  :    0 - 0x0
    "00000000", -- 1308 - 0x51c  :    0 - 0x0
    "00000000", -- 1309 - 0x51d  :    0 - 0x0
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00111111", -- 1312 - 0x520  :   63 - 0x3f
    "11111111", -- 1313 - 0x521  :  255 - 0xff
    "11111111", -- 1314 - 0x522  :  255 - 0xff
    "11111111", -- 1315 - 0x523  :  255 - 0xff
    "11111111", -- 1316 - 0x524  :  255 - 0xff
    "11111111", -- 1317 - 0x525  :  255 - 0xff
    "11111011", -- 1318 - 0x526  :  251 - 0xfb
    "01110110", -- 1319 - 0x527  :  118 - 0x76
    "00000000", -- 1320 - 0x528  :    0 - 0x0
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "11001111", -- 1322 - 0x52a  :  207 - 0xcf
    "00000111", -- 1323 - 0x52b  :    7 - 0x7
    "01111111", -- 1324 - 0x52c  :  127 - 0x7f
    "00000000", -- 1325 - 0x52d  :    0 - 0x0
    "00000000", -- 1326 - 0x52e  :    0 - 0x0
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00100000", -- 1328 - 0x530  :   32 - 0x20
    "11111000", -- 1329 - 0x531  :  248 - 0xf8
    "11111111", -- 1330 - 0x532  :  255 - 0xff
    "11000011", -- 1331 - 0x533  :  195 - 0xc3
    "11111101", -- 1332 - 0x534  :  253 - 0xfd
    "11111110", -- 1333 - 0x535  :  254 - 0xfe
    "11110000", -- 1334 - 0x536  :  240 - 0xf0
    "01000000", -- 1335 - 0x537  :   64 - 0x40
    "00000000", -- 1336 - 0x538  :    0 - 0x0
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "00111100", -- 1338 - 0x53a  :   60 - 0x3c
    "11111100", -- 1339 - 0x53b  :  252 - 0xfc
    "11111110", -- 1340 - 0x53c  :  254 - 0xfe
    "11100000", -- 1341 - 0x53d  :  224 - 0xe0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "01000000", -- 1344 - 0x540  :   64 - 0x40
    "11100000", -- 1345 - 0x541  :  224 - 0xe0
    "01000000", -- 1346 - 0x542  :   64 - 0x40
    "01000000", -- 1347 - 0x543  :   64 - 0x40
    "01000001", -- 1348 - 0x544  :   65 - 0x41
    "01000001", -- 1349 - 0x545  :   65 - 0x41
    "01001111", -- 1350 - 0x546  :   79 - 0x4f
    "01000111", -- 1351 - 0x547  :   71 - 0x47
    "01000000", -- 1352 - 0x548  :   64 - 0x40
    "11100000", -- 1353 - 0x549  :  224 - 0xe0
    "01000000", -- 1354 - 0x54a  :   64 - 0x40
    "00111111", -- 1355 - 0x54b  :   63 - 0x3f
    "00111110", -- 1356 - 0x54c  :   62 - 0x3e
    "00111110", -- 1357 - 0x54d  :   62 - 0x3e
    "00110000", -- 1358 - 0x54e  :   48 - 0x30
    "00111000", -- 1359 - 0x54f  :   56 - 0x38
    "00000000", -- 1360 - 0x550  :    0 - 0x0
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "11100000", -- 1366 - 0x556  :  224 - 0xe0
    "11000000", -- 1367 - 0x557  :  192 - 0xc0
    "00000000", -- 1368 - 0x558  :    0 - 0x0
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "11111000", -- 1371 - 0x55b  :  248 - 0xf8
    "11111000", -- 1372 - 0x55c  :  248 - 0xf8
    "11111000", -- 1373 - 0x55d  :  248 - 0xf8
    "00011000", -- 1374 - 0x55e  :   24 - 0x18
    "00111000", -- 1375 - 0x55f  :   56 - 0x38
    "01000011", -- 1376 - 0x560  :   67 - 0x43
    "01000110", -- 1377 - 0x561  :   70 - 0x46
    "01000100", -- 1378 - 0x562  :   68 - 0x44
    "01000000", -- 1379 - 0x563  :   64 - 0x40
    "01000000", -- 1380 - 0x564  :   64 - 0x40
    "01000000", -- 1381 - 0x565  :   64 - 0x40
    "01000000", -- 1382 - 0x566  :   64 - 0x40
    "01000000", -- 1383 - 0x567  :   64 - 0x40
    "00111100", -- 1384 - 0x568  :   60 - 0x3c
    "00111001", -- 1385 - 0x569  :   57 - 0x39
    "00111011", -- 1386 - 0x56a  :   59 - 0x3b
    "00111111", -- 1387 - 0x56b  :   63 - 0x3f
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "10000000", -- 1392 - 0x570  :  128 - 0x80
    "11000000", -- 1393 - 0x571  :  192 - 0xc0
    "01000000", -- 1394 - 0x572  :   64 - 0x40
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000000", -- 1396 - 0x574  :    0 - 0x0
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "01111000", -- 1400 - 0x578  :  120 - 0x78
    "00111000", -- 1401 - 0x579  :   56 - 0x38
    "10111000", -- 1402 - 0x57a  :  184 - 0xb8
    "11111000", -- 1403 - 0x57b  :  248 - 0xf8
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "00110001", -- 1408 - 0x580  :   49 - 0x31
    "00110000", -- 1409 - 0x581  :   48 - 0x30
    "00111000", -- 1410 - 0x582  :   56 - 0x38
    "01111100", -- 1411 - 0x583  :  124 - 0x7c
    "01111111", -- 1412 - 0x584  :  127 - 0x7f
    "11111111", -- 1413 - 0x585  :  255 - 0xff
    "11111111", -- 1414 - 0x586  :  255 - 0xff
    "11111011", -- 1415 - 0x587  :  251 - 0xfb
    "00111111", -- 1416 - 0x588  :   63 - 0x3f
    "00111111", -- 1417 - 0x589  :   63 - 0x3f
    "00001111", -- 1418 - 0x58a  :   15 - 0xf
    "01110111", -- 1419 - 0x58b  :  119 - 0x77
    "01110111", -- 1420 - 0x58c  :  119 - 0x77
    "11110111", -- 1421 - 0x58d  :  247 - 0xf7
    "11110111", -- 1422 - 0x58e  :  247 - 0xf7
    "11110111", -- 1423 - 0x58f  :  247 - 0xf7
    "00010000", -- 1424 - 0x590  :   16 - 0x10
    "01111110", -- 1425 - 0x591  :  126 - 0x7e
    "00111110", -- 1426 - 0x592  :   62 - 0x3e
    "00000000", -- 1427 - 0x593  :    0 - 0x0
    "00011110", -- 1428 - 0x594  :   30 - 0x1e
    "11111110", -- 1429 - 0x595  :  254 - 0xfe
    "11111111", -- 1430 - 0x596  :  255 - 0xff
    "11111111", -- 1431 - 0x597  :  255 - 0xff
    "11111111", -- 1432 - 0x598  :  255 - 0xff
    "11111110", -- 1433 - 0x599  :  254 - 0xfe
    "11111110", -- 1434 - 0x59a  :  254 - 0xfe
    "11111110", -- 1435 - 0x59b  :  254 - 0xfe
    "11111010", -- 1436 - 0x59c  :  250 - 0xfa
    "11111010", -- 1437 - 0x59d  :  250 - 0xfa
    "11110011", -- 1438 - 0x59e  :  243 - 0xf3
    "11100111", -- 1439 - 0x59f  :  231 - 0xe7
    "11111111", -- 1440 - 0x5a0  :  255 - 0xff
    "11111111", -- 1441 - 0x5a1  :  255 - 0xff
    "11100011", -- 1442 - 0x5a2  :  227 - 0xe3
    "11000011", -- 1443 - 0x5a3  :  195 - 0xc3
    "10000111", -- 1444 - 0x5a4  :  135 - 0x87
    "01001000", -- 1445 - 0x5a5  :   72 - 0x48
    "00111100", -- 1446 - 0x5a6  :   60 - 0x3c
    "11111100", -- 1447 - 0x5a7  :  252 - 0xfc
    "11110000", -- 1448 - 0x5a8  :  240 - 0xf0
    "11111000", -- 1449 - 0x5a9  :  248 - 0xf8
    "11111100", -- 1450 - 0x5aa  :  252 - 0xfc
    "01111100", -- 1451 - 0x5ab  :  124 - 0x7c
    "01111000", -- 1452 - 0x5ac  :  120 - 0x78
    "00111000", -- 1453 - 0x5ad  :   56 - 0x38
    "00111100", -- 1454 - 0x5ae  :   60 - 0x3c
    "11111100", -- 1455 - 0x5af  :  252 - 0xfc
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0
    "11111111", -- 1457 - 0x5b1  :  255 - 0xff
    "11000011", -- 1458 - 0x5b2  :  195 - 0xc3
    "10000011", -- 1459 - 0x5b3  :  131 - 0x83
    "10000011", -- 1460 - 0x5b4  :  131 - 0x83
    "11111111", -- 1461 - 0x5b5  :  255 - 0xff
    "11111111", -- 1462 - 0x5b6  :  255 - 0xff
    "11111111", -- 1463 - 0x5b7  :  255 - 0xff
    "11111111", -- 1464 - 0x5b8  :  255 - 0xff
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "11000011", -- 1466 - 0x5ba  :  195 - 0xc3
    "10000001", -- 1467 - 0x5bb  :  129 - 0x81
    "10000001", -- 1468 - 0x5bc  :  129 - 0x81
    "11000011", -- 1469 - 0x5bd  :  195 - 0xc3
    "11111111", -- 1470 - 0x5be  :  255 - 0xff
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00011111", -- 1472 - 0x5c0  :   31 - 0x1f
    "00011111", -- 1473 - 0x5c1  :   31 - 0x1f
    "00001111", -- 1474 - 0x5c2  :   15 - 0xf
    "00000111", -- 1475 - 0x5c3  :    7 - 0x7
    "00000001", -- 1476 - 0x5c4  :    1 - 0x1
    "00000000", -- 1477 - 0x5c5  :    0 - 0x0
    "00000000", -- 1478 - 0x5c6  :    0 - 0x0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "00000000", -- 1482 - 0x5ca  :    0 - 0x0
    "00000000", -- 1483 - 0x5cb  :    0 - 0x0
    "00000000", -- 1484 - 0x5cc  :    0 - 0x0
    "00000000", -- 1485 - 0x5cd  :    0 - 0x0
    "00000000", -- 1486 - 0x5ce  :    0 - 0x0
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "11110000", -- 1488 - 0x5d0  :  240 - 0xf0
    "11111011", -- 1489 - 0x5d1  :  251 - 0xfb
    "11111111", -- 1490 - 0x5d2  :  255 - 0xff
    "11111111", -- 1491 - 0x5d3  :  255 - 0xff
    "11111110", -- 1492 - 0x5d4  :  254 - 0xfe
    "00111110", -- 1493 - 0x5d5  :   62 - 0x3e
    "00001100", -- 1494 - 0x5d6  :   12 - 0xc
    "00000100", -- 1495 - 0x5d7  :    4 - 0x4
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0
    "00001011", -- 1497 - 0x5d9  :   11 - 0xb
    "00011111", -- 1498 - 0x5da  :   31 - 0x1f
    "00011111", -- 1499 - 0x5db  :   31 - 0x1f
    "00011110", -- 1500 - 0x5dc  :   30 - 0x1e
    "00111110", -- 1501 - 0x5dd  :   62 - 0x3e
    "00001100", -- 1502 - 0x5de  :   12 - 0xc
    "00000100", -- 1503 - 0x5df  :    4 - 0x4
    "00011111", -- 1504 - 0x5e0  :   31 - 0x1f
    "00011111", -- 1505 - 0x5e1  :   31 - 0x1f
    "00001111", -- 1506 - 0x5e2  :   15 - 0xf
    "00001111", -- 1507 - 0x5e3  :   15 - 0xf
    "00000111", -- 1508 - 0x5e4  :    7 - 0x7
    "00000000", -- 1509 - 0x5e5  :    0 - 0x0
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00000000", -- 1514 - 0x5ea  :    0 - 0x0
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "00000000", -- 1516 - 0x5ec  :    0 - 0x0
    "00000000", -- 1517 - 0x5ed  :    0 - 0x0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "11111011", -- 1520 - 0x5f0  :  251 - 0xfb
    "11111111", -- 1521 - 0x5f1  :  255 - 0xff
    "11111111", -- 1522 - 0x5f2  :  255 - 0xff
    "11111111", -- 1523 - 0x5f3  :  255 - 0xff
    "11111111", -- 1524 - 0x5f4  :  255 - 0xff
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000011", -- 1528 - 0x5f8  :    3 - 0x3
    "00001111", -- 1529 - 0x5f9  :   15 - 0xf
    "00001111", -- 1530 - 0x5fa  :   15 - 0xf
    "00001111", -- 1531 - 0x5fb  :   15 - 0xf
    "00001111", -- 1532 - 0x5fc  :   15 - 0xf
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0
    "00011000", -- 1537 - 0x601  :   24 - 0x18
    "00111100", -- 1538 - 0x602  :   60 - 0x3c
    "01111110", -- 1539 - 0x603  :  126 - 0x7e
    "01101110", -- 1540 - 0x604  :  110 - 0x6e
    "11011111", -- 1541 - 0x605  :  223 - 0xdf
    "11011111", -- 1542 - 0x606  :  223 - 0xdf
    "11011111", -- 1543 - 0x607  :  223 - 0xdf
    "00000000", -- 1544 - 0x608  :    0 - 0x0
    "00011000", -- 1545 - 0x609  :   24 - 0x18
    "00111100", -- 1546 - 0x60a  :   60 - 0x3c
    "01111110", -- 1547 - 0x60b  :  126 - 0x7e
    "01110110", -- 1548 - 0x60c  :  118 - 0x76
    "11111011", -- 1549 - 0x60d  :  251 - 0xfb
    "11111011", -- 1550 - 0x60e  :  251 - 0xfb
    "11111011", -- 1551 - 0x60f  :  251 - 0xfb
    "00000000", -- 1552 - 0x610  :    0 - 0x0
    "00011000", -- 1553 - 0x611  :   24 - 0x18
    "00011000", -- 1554 - 0x612  :   24 - 0x18
    "00111100", -- 1555 - 0x613  :   60 - 0x3c
    "00111100", -- 1556 - 0x614  :   60 - 0x3c
    "00111100", -- 1557 - 0x615  :   60 - 0x3c
    "00111100", -- 1558 - 0x616  :   60 - 0x3c
    "00011100", -- 1559 - 0x617  :   28 - 0x1c
    "00000000", -- 1560 - 0x618  :    0 - 0x0
    "00010000", -- 1561 - 0x619  :   16 - 0x10
    "00010000", -- 1562 - 0x61a  :   16 - 0x10
    "00100000", -- 1563 - 0x61b  :   32 - 0x20
    "00100000", -- 1564 - 0x61c  :   32 - 0x20
    "00100000", -- 1565 - 0x61d  :   32 - 0x20
    "00100000", -- 1566 - 0x61e  :   32 - 0x20
    "00100000", -- 1567 - 0x61f  :   32 - 0x20
    "00000000", -- 1568 - 0x620  :    0 - 0x0
    "00001000", -- 1569 - 0x621  :    8 - 0x8
    "00001000", -- 1570 - 0x622  :    8 - 0x8
    "00001000", -- 1571 - 0x623  :    8 - 0x8
    "00001000", -- 1572 - 0x624  :    8 - 0x8
    "00001000", -- 1573 - 0x625  :    8 - 0x8
    "00001000", -- 1574 - 0x626  :    8 - 0x8
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0
    "00001000", -- 1577 - 0x629  :    8 - 0x8
    "00001000", -- 1578 - 0x62a  :    8 - 0x8
    "00001000", -- 1579 - 0x62b  :    8 - 0x8
    "00001000", -- 1580 - 0x62c  :    8 - 0x8
    "00001000", -- 1581 - 0x62d  :    8 - 0x8
    "00001000", -- 1582 - 0x62e  :    8 - 0x8
    "00001000", -- 1583 - 0x62f  :    8 - 0x8
    "00000000", -- 1584 - 0x630  :    0 - 0x0
    "00001000", -- 1585 - 0x631  :    8 - 0x8
    "00001000", -- 1586 - 0x632  :    8 - 0x8
    "00000100", -- 1587 - 0x633  :    4 - 0x4
    "00000100", -- 1588 - 0x634  :    4 - 0x4
    "00000100", -- 1589 - 0x635  :    4 - 0x4
    "00000100", -- 1590 - 0x636  :    4 - 0x4
    "00000100", -- 1591 - 0x637  :    4 - 0x4
    "00000000", -- 1592 - 0x638  :    0 - 0x0
    "00010000", -- 1593 - 0x639  :   16 - 0x10
    "00010000", -- 1594 - 0x63a  :   16 - 0x10
    "00111000", -- 1595 - 0x63b  :   56 - 0x38
    "00111000", -- 1596 - 0x63c  :   56 - 0x38
    "00111000", -- 1597 - 0x63d  :   56 - 0x38
    "00111000", -- 1598 - 0x63e  :   56 - 0x38
    "00111000", -- 1599 - 0x63f  :   56 - 0x38
    "00111100", -- 1600 - 0x640  :   60 - 0x3c
    "01111110", -- 1601 - 0x641  :  126 - 0x7e
    "01110111", -- 1602 - 0x642  :  119 - 0x77
    "11111011", -- 1603 - 0x643  :  251 - 0xfb
    "10011111", -- 1604 - 0x644  :  159 - 0x9f
    "01011111", -- 1605 - 0x645  :   95 - 0x5f
    "10001110", -- 1606 - 0x646  :  142 - 0x8e
    "00100000", -- 1607 - 0x647  :   32 - 0x20
    "00000000", -- 1608 - 0x648  :    0 - 0x0
    "00011000", -- 1609 - 0x649  :   24 - 0x18
    "00111100", -- 1610 - 0x64a  :   60 - 0x3c
    "00001110", -- 1611 - 0x64b  :   14 - 0xe
    "00001110", -- 1612 - 0x64c  :   14 - 0xe
    "00000100", -- 1613 - 0x64d  :    4 - 0x4
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "01011100", -- 1616 - 0x650  :   92 - 0x5c
    "00101110", -- 1617 - 0x651  :   46 - 0x2e
    "10001111", -- 1618 - 0x652  :  143 - 0x8f
    "00111111", -- 1619 - 0x653  :   63 - 0x3f
    "01111011", -- 1620 - 0x654  :  123 - 0x7b
    "01110111", -- 1621 - 0x655  :  119 - 0x77
    "01111110", -- 1622 - 0x656  :  126 - 0x7e
    "00111100", -- 1623 - 0x657  :   60 - 0x3c
    "00000000", -- 1624 - 0x658  :    0 - 0x0
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000100", -- 1626 - 0x65a  :    4 - 0x4
    "00000110", -- 1627 - 0x65b  :    6 - 0x6
    "00011110", -- 1628 - 0x65c  :   30 - 0x1e
    "00111100", -- 1629 - 0x65d  :   60 - 0x3c
    "00011000", -- 1630 - 0x65e  :   24 - 0x18
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00010011", -- 1632 - 0x660  :   19 - 0x13
    "01001111", -- 1633 - 0x661  :   79 - 0x4f
    "00111111", -- 1634 - 0x662  :   63 - 0x3f
    "10111111", -- 1635 - 0x663  :  191 - 0xbf
    "00111111", -- 1636 - 0x664  :   63 - 0x3f
    "01111010", -- 1637 - 0x665  :  122 - 0x7a
    "11111000", -- 1638 - 0x666  :  248 - 0xf8
    "11111000", -- 1639 - 0x667  :  248 - 0xf8
    "00000000", -- 1640 - 0x668  :    0 - 0x0
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000001", -- 1642 - 0x66a  :    1 - 0x1
    "00001010", -- 1643 - 0x66b  :   10 - 0xa
    "00010111", -- 1644 - 0x66c  :   23 - 0x17
    "00001111", -- 1645 - 0x66d  :   15 - 0xf
    "00101111", -- 1646 - 0x66e  :   47 - 0x2f
    "00011111", -- 1647 - 0x66f  :   31 - 0x1f
    "00000000", -- 1648 - 0x670  :    0 - 0x0
    "00001000", -- 1649 - 0x671  :    8 - 0x8
    "00000101", -- 1650 - 0x672  :    5 - 0x5
    "00001111", -- 1651 - 0x673  :   15 - 0xf
    "00101111", -- 1652 - 0x674  :   47 - 0x2f
    "00011101", -- 1653 - 0x675  :   29 - 0x1d
    "00011100", -- 1654 - 0x676  :   28 - 0x1c
    "00111100", -- 1655 - 0x677  :   60 - 0x3c
    "00000000", -- 1656 - 0x678  :    0 - 0x0
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000101", -- 1660 - 0x67c  :    5 - 0x5
    "00000111", -- 1661 - 0x67d  :    7 - 0x7
    "00001111", -- 1662 - 0x67e  :   15 - 0xf
    "00000111", -- 1663 - 0x67f  :    7 - 0x7
    "00000000", -- 1664 - 0x680  :    0 - 0x0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000010", -- 1668 - 0x684  :    2 - 0x2
    "00001011", -- 1669 - 0x685  :   11 - 0xb
    "00000111", -- 1670 - 0x686  :    7 - 0x7
    "00001111", -- 1671 - 0x687  :   15 - 0xf
    "00000000", -- 1672 - 0x688  :    0 - 0x0
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000001", -- 1678 - 0x68e  :    1 - 0x1
    "00000011", -- 1679 - 0x68f  :    3 - 0x3
    "00000000", -- 1680 - 0x690  :    0 - 0x0
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00001000", -- 1685 - 0x695  :    8 - 0x8
    "00000100", -- 1686 - 0x696  :    4 - 0x4
    "00000100", -- 1687 - 0x697  :    4 - 0x4
    "00000000", -- 1688 - 0x698  :    0 - 0x0
    "01100000", -- 1689 - 0x699  :   96 - 0x60
    "11110000", -- 1690 - 0x69a  :  240 - 0xf0
    "11111000", -- 1691 - 0x69b  :  248 - 0xf8
    "01111100", -- 1692 - 0x69c  :  124 - 0x7c
    "00111110", -- 1693 - 0x69d  :   62 - 0x3e
    "01111110", -- 1694 - 0x69e  :  126 - 0x7e
    "01111111", -- 1695 - 0x69f  :  127 - 0x7f
    "00000010", -- 1696 - 0x6a0  :    2 - 0x2
    "00000010", -- 1697 - 0x6a1  :    2 - 0x2
    "00000010", -- 1698 - 0x6a2  :    2 - 0x2
    "00000101", -- 1699 - 0x6a3  :    5 - 0x5
    "01110001", -- 1700 - 0x6a4  :  113 - 0x71
    "01111111", -- 1701 - 0x6a5  :  127 - 0x7f
    "01111111", -- 1702 - 0x6a6  :  127 - 0x7f
    "01111111", -- 1703 - 0x6a7  :  127 - 0x7f
    "00111111", -- 1704 - 0x6a8  :   63 - 0x3f
    "01011111", -- 1705 - 0x6a9  :   95 - 0x5f
    "01111111", -- 1706 - 0x6aa  :  127 - 0x7f
    "00111110", -- 1707 - 0x6ab  :   62 - 0x3e
    "00001110", -- 1708 - 0x6ac  :   14 - 0xe
    "00001010", -- 1709 - 0x6ad  :   10 - 0xa
    "01010001", -- 1710 - 0x6ae  :   81 - 0x51
    "00100000", -- 1711 - 0x6af  :   32 - 0x20
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "00000000", -- 1715 - 0x6b3  :    0 - 0x0
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000100", -- 1719 - 0x6b7  :    4 - 0x4
    "00000000", -- 1720 - 0x6b8  :    0 - 0x0
    "00000000", -- 1721 - 0x6b9  :    0 - 0x0
    "00000000", -- 1722 - 0x6ba  :    0 - 0x0
    "00000000", -- 1723 - 0x6bb  :    0 - 0x0
    "00000000", -- 1724 - 0x6bc  :    0 - 0x0
    "00000000", -- 1725 - 0x6bd  :    0 - 0x0
    "00001110", -- 1726 - 0x6be  :   14 - 0xe
    "00011111", -- 1727 - 0x6bf  :   31 - 0x1f
    "00000010", -- 1728 - 0x6c0  :    2 - 0x2
    "00000010", -- 1729 - 0x6c1  :    2 - 0x2
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000001", -- 1731 - 0x6c3  :    1 - 0x1
    "00010011", -- 1732 - 0x6c4  :   19 - 0x13
    "00111111", -- 1733 - 0x6c5  :   63 - 0x3f
    "01111111", -- 1734 - 0x6c6  :  127 - 0x7f
    "01111111", -- 1735 - 0x6c7  :  127 - 0x7f
    "00111111", -- 1736 - 0x6c8  :   63 - 0x3f
    "01111111", -- 1737 - 0x6c9  :  127 - 0x7f
    "01111111", -- 1738 - 0x6ca  :  127 - 0x7f
    "11111110", -- 1739 - 0x6cb  :  254 - 0xfe
    "11101100", -- 1740 - 0x6cc  :  236 - 0xec
    "11001010", -- 1741 - 0x6cd  :  202 - 0xca
    "01010001", -- 1742 - 0x6ce  :   81 - 0x51
    "00100000", -- 1743 - 0x6cf  :   32 - 0x20
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0
    "01000000", -- 1745 - 0x6d1  :   64 - 0x40
    "01100000", -- 1746 - 0x6d2  :   96 - 0x60
    "01110000", -- 1747 - 0x6d3  :  112 - 0x70
    "01110011", -- 1748 - 0x6d4  :  115 - 0x73
    "00100111", -- 1749 - 0x6d5  :   39 - 0x27
    "00001111", -- 1750 - 0x6d6  :   15 - 0xf
    "00011111", -- 1751 - 0x6d7  :   31 - 0x1f
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0
    "01000000", -- 1753 - 0x6d9  :   64 - 0x40
    "01100011", -- 1754 - 0x6da  :   99 - 0x63
    "01110111", -- 1755 - 0x6db  :  119 - 0x77
    "01111100", -- 1756 - 0x6dc  :  124 - 0x7c
    "00111000", -- 1757 - 0x6dd  :   56 - 0x38
    "11111000", -- 1758 - 0x6de  :  248 - 0xf8
    "11100100", -- 1759 - 0x6df  :  228 - 0xe4
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000011", -- 1764 - 0x6e4  :    3 - 0x3
    "00000111", -- 1765 - 0x6e5  :    7 - 0x7
    "00001111", -- 1766 - 0x6e6  :   15 - 0xf
    "00011111", -- 1767 - 0x6e7  :   31 - 0x1f
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000011", -- 1770 - 0x6ea  :    3 - 0x3
    "00000111", -- 1771 - 0x6eb  :    7 - 0x7
    "00001100", -- 1772 - 0x6ec  :   12 - 0xc
    "00011000", -- 1773 - 0x6ed  :   24 - 0x18
    "11111000", -- 1774 - 0x6ee  :  248 - 0xf8
    "11100100", -- 1775 - 0x6ef  :  228 - 0xe4
    "01111111", -- 1776 - 0x6f0  :  127 - 0x7f
    "01111111", -- 1777 - 0x6f1  :  127 - 0x7f
    "00111111", -- 1778 - 0x6f2  :   63 - 0x3f
    "00111111", -- 1779 - 0x6f3  :   63 - 0x3f
    "00011111", -- 1780 - 0x6f4  :   31 - 0x1f
    "00011111", -- 1781 - 0x6f5  :   31 - 0x1f
    "00001111", -- 1782 - 0x6f6  :   15 - 0xf
    "00000111", -- 1783 - 0x6f7  :    7 - 0x7
    "00000011", -- 1784 - 0x6f8  :    3 - 0x3
    "01000100", -- 1785 - 0x6f9  :   68 - 0x44
    "00101000", -- 1786 - 0x6fa  :   40 - 0x28
    "00010000", -- 1787 - 0x6fb  :   16 - 0x10
    "00001000", -- 1788 - 0x6fc  :    8 - 0x8
    "00000100", -- 1789 - 0x6fd  :    4 - 0x4
    "00000011", -- 1790 - 0x6fe  :    3 - 0x3
    "00000100", -- 1791 - 0x6ff  :    4 - 0x4
    "00000011", -- 1792 - 0x700  :    3 - 0x3
    "00000111", -- 1793 - 0x701  :    7 - 0x7
    "00001111", -- 1794 - 0x702  :   15 - 0xf
    "00011111", -- 1795 - 0x703  :   31 - 0x1f
    "00111111", -- 1796 - 0x704  :   63 - 0x3f
    "01110111", -- 1797 - 0x705  :  119 - 0x77
    "01110111", -- 1798 - 0x706  :  119 - 0x77
    "11110101", -- 1799 - 0x707  :  245 - 0xf5
    "00000011", -- 1800 - 0x708  :    3 - 0x3
    "00000111", -- 1801 - 0x709  :    7 - 0x7
    "00001111", -- 1802 - 0x70a  :   15 - 0xf
    "00011111", -- 1803 - 0x70b  :   31 - 0x1f
    "00100111", -- 1804 - 0x70c  :   39 - 0x27
    "01111011", -- 1805 - 0x70d  :  123 - 0x7b
    "01111000", -- 1806 - 0x70e  :  120 - 0x78
    "11111011", -- 1807 - 0x70f  :  251 - 0xfb
    "11000000", -- 1808 - 0x710  :  192 - 0xc0
    "11100000", -- 1809 - 0x711  :  224 - 0xe0
    "11110000", -- 1810 - 0x712  :  240 - 0xf0
    "11111000", -- 1811 - 0x713  :  248 - 0xf8
    "11111100", -- 1812 - 0x714  :  252 - 0xfc
    "11101110", -- 1813 - 0x715  :  238 - 0xee
    "11101110", -- 1814 - 0x716  :  238 - 0xee
    "10101111", -- 1815 - 0x717  :  175 - 0xaf
    "11000000", -- 1816 - 0x718  :  192 - 0xc0
    "11100000", -- 1817 - 0x719  :  224 - 0xe0
    "11110000", -- 1818 - 0x71a  :  240 - 0xf0
    "11111000", -- 1819 - 0x71b  :  248 - 0xf8
    "11100100", -- 1820 - 0x71c  :  228 - 0xe4
    "11011110", -- 1821 - 0x71d  :  222 - 0xde
    "00011110", -- 1822 - 0x71e  :   30 - 0x1e
    "11011111", -- 1823 - 0x71f  :  223 - 0xdf
    "11110001", -- 1824 - 0x720  :  241 - 0xf1
    "11111111", -- 1825 - 0x721  :  255 - 0xff
    "01111000", -- 1826 - 0x722  :  120 - 0x78
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000000", -- 1828 - 0x724  :    0 - 0x0
    "00011000", -- 1829 - 0x725  :   24 - 0x18
    "00011100", -- 1830 - 0x726  :   28 - 0x1c
    "00001110", -- 1831 - 0x727  :   14 - 0xe
    "11111111", -- 1832 - 0x728  :  255 - 0xff
    "11111111", -- 1833 - 0x729  :  255 - 0xff
    "01111111", -- 1834 - 0x72a  :  127 - 0x7f
    "00001111", -- 1835 - 0x72b  :   15 - 0xf
    "00001111", -- 1836 - 0x72c  :   15 - 0xf
    "00000111", -- 1837 - 0x72d  :    7 - 0x7
    "00000011", -- 1838 - 0x72e  :    3 - 0x3
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "10001111", -- 1840 - 0x730  :  143 - 0x8f
    "11111111", -- 1841 - 0x731  :  255 - 0xff
    "00011110", -- 1842 - 0x732  :   30 - 0x1e
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00001100", -- 1844 - 0x734  :   12 - 0xc
    "00111110", -- 1845 - 0x735  :   62 - 0x3e
    "01111110", -- 1846 - 0x736  :  126 - 0x7e
    "01111100", -- 1847 - 0x737  :  124 - 0x7c
    "11111111", -- 1848 - 0x738  :  255 - 0xff
    "11111111", -- 1849 - 0x739  :  255 - 0xff
    "11111110", -- 1850 - 0x73a  :  254 - 0xfe
    "11110000", -- 1851 - 0x73b  :  240 - 0xf0
    "11110000", -- 1852 - 0x73c  :  240 - 0xf0
    "11000000", -- 1853 - 0x73d  :  192 - 0xc0
    "10000000", -- 1854 - 0x73e  :  128 - 0x80
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00011000", -- 1866 - 0x74a  :   24 - 0x18
    "00100100", -- 1867 - 0x74b  :   36 - 0x24
    "00100100", -- 1868 - 0x74c  :   36 - 0x24
    "00011000", -- 1869 - 0x74d  :   24 - 0x18
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0
    "00000010", -- 1873 - 0x751  :    2 - 0x2
    "01000001", -- 1874 - 0x752  :   65 - 0x41
    "01000001", -- 1875 - 0x753  :   65 - 0x41
    "01100001", -- 1876 - 0x754  :   97 - 0x61
    "00110011", -- 1877 - 0x755  :   51 - 0x33
    "00000110", -- 1878 - 0x756  :    6 - 0x6
    "00111100", -- 1879 - 0x757  :   60 - 0x3c
    "00111100", -- 1880 - 0x758  :   60 - 0x3c
    "01111110", -- 1881 - 0x759  :  126 - 0x7e
    "11111111", -- 1882 - 0x75a  :  255 - 0xff
    "11111111", -- 1883 - 0x75b  :  255 - 0xff
    "11111111", -- 1884 - 0x75c  :  255 - 0xff
    "11111111", -- 1885 - 0x75d  :  255 - 0xff
    "01111110", -- 1886 - 0x75e  :  126 - 0x7e
    "00111100", -- 1887 - 0x75f  :   60 - 0x3c
    "00000011", -- 1888 - 0x760  :    3 - 0x3
    "00000111", -- 1889 - 0x761  :    7 - 0x7
    "00001111", -- 1890 - 0x762  :   15 - 0xf
    "00011111", -- 1891 - 0x763  :   31 - 0x1f
    "00111111", -- 1892 - 0x764  :   63 - 0x3f
    "01111111", -- 1893 - 0x765  :  127 - 0x7f
    "01111111", -- 1894 - 0x766  :  127 - 0x7f
    "11111111", -- 1895 - 0x767  :  255 - 0xff
    "00000011", -- 1896 - 0x768  :    3 - 0x3
    "00000111", -- 1897 - 0x769  :    7 - 0x7
    "00001111", -- 1898 - 0x76a  :   15 - 0xf
    "00011111", -- 1899 - 0x76b  :   31 - 0x1f
    "00111111", -- 1900 - 0x76c  :   63 - 0x3f
    "01100011", -- 1901 - 0x76d  :   99 - 0x63
    "01000001", -- 1902 - 0x76e  :   65 - 0x41
    "11000001", -- 1903 - 0x76f  :  193 - 0xc1
    "11000000", -- 1904 - 0x770  :  192 - 0xc0
    "11100000", -- 1905 - 0x771  :  224 - 0xe0
    "11110000", -- 1906 - 0x772  :  240 - 0xf0
    "11111000", -- 1907 - 0x773  :  248 - 0xf8
    "11111100", -- 1908 - 0x774  :  252 - 0xfc
    "11111110", -- 1909 - 0x775  :  254 - 0xfe
    "11111110", -- 1910 - 0x776  :  254 - 0xfe
    "11111111", -- 1911 - 0x777  :  255 - 0xff
    "11000000", -- 1912 - 0x778  :  192 - 0xc0
    "10000000", -- 1913 - 0x779  :  128 - 0x80
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "10001100", -- 1916 - 0x77c  :  140 - 0x8c
    "11111110", -- 1917 - 0x77d  :  254 - 0xfe
    "11111110", -- 1918 - 0x77e  :  254 - 0xfe
    "11110011", -- 1919 - 0x77f  :  243 - 0xf3
    "11111111", -- 1920 - 0x780  :  255 - 0xff
    "11111111", -- 1921 - 0x781  :  255 - 0xff
    "11111111", -- 1922 - 0x782  :  255 - 0xff
    "01111000", -- 1923 - 0x783  :  120 - 0x78
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "11000001", -- 1928 - 0x788  :  193 - 0xc1
    "11100011", -- 1929 - 0x789  :  227 - 0xe3
    "11111111", -- 1930 - 0x78a  :  255 - 0xff
    "01000111", -- 1931 - 0x78b  :   71 - 0x47
    "00001111", -- 1932 - 0x78c  :   15 - 0xf
    "00001111", -- 1933 - 0x78d  :   15 - 0xf
    "00001111", -- 1934 - 0x78e  :   15 - 0xf
    "00000111", -- 1935 - 0x78f  :    7 - 0x7
    "11111111", -- 1936 - 0x790  :  255 - 0xff
    "11111111", -- 1937 - 0x791  :  255 - 0xff
    "11111111", -- 1938 - 0x792  :  255 - 0xff
    "00011110", -- 1939 - 0x793  :   30 - 0x1e
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00100000", -- 1941 - 0x795  :   32 - 0x20
    "00100000", -- 1942 - 0x796  :   32 - 0x20
    "01000000", -- 1943 - 0x797  :   64 - 0x40
    "11110001", -- 1944 - 0x798  :  241 - 0xf1
    "11111001", -- 1945 - 0x799  :  249 - 0xf9
    "11111111", -- 1946 - 0x79a  :  255 - 0xff
    "11100010", -- 1947 - 0x79b  :  226 - 0xe2
    "11110000", -- 1948 - 0x79c  :  240 - 0xf0
    "11110000", -- 1949 - 0x79d  :  240 - 0xf0
    "11110000", -- 1950 - 0x79e  :  240 - 0xf0
    "11100000", -- 1951 - 0x79f  :  224 - 0xe0
    "00010110", -- 1952 - 0x7a0  :   22 - 0x16
    "00011111", -- 1953 - 0x7a1  :   31 - 0x1f
    "00111111", -- 1954 - 0x7a2  :   63 - 0x3f
    "01111111", -- 1955 - 0x7a3  :  127 - 0x7f
    "00111101", -- 1956 - 0x7a4  :   61 - 0x3d
    "00011101", -- 1957 - 0x7a5  :   29 - 0x1d
    "00111111", -- 1958 - 0x7a6  :   63 - 0x3f
    "00011111", -- 1959 - 0x7a7  :   31 - 0x1f
    "00010110", -- 1960 - 0x7a8  :   22 - 0x16
    "00011111", -- 1961 - 0x7a9  :   31 - 0x1f
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000101", -- 1964 - 0x7ac  :    5 - 0x5
    "00001101", -- 1965 - 0x7ad  :   13 - 0xd
    "00111111", -- 1966 - 0x7ae  :   63 - 0x3f
    "00011111", -- 1967 - 0x7af  :   31 - 0x1f
    "10000000", -- 1968 - 0x7b0  :  128 - 0x80
    "10000000", -- 1969 - 0x7b1  :  128 - 0x80
    "11000000", -- 1970 - 0x7b2  :  192 - 0xc0
    "11100000", -- 1971 - 0x7b3  :  224 - 0xe0
    "11110000", -- 1972 - 0x7b4  :  240 - 0xf0
    "11110000", -- 1973 - 0x7b5  :  240 - 0xf0
    "11110000", -- 1974 - 0x7b6  :  240 - 0xf0
    "11111000", -- 1975 - 0x7b7  :  248 - 0xf8
    "10000000", -- 1976 - 0x7b8  :  128 - 0x80
    "10000000", -- 1977 - 0x7b9  :  128 - 0x80
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "10100000", -- 1981 - 0x7bd  :  160 - 0xa0
    "10100000", -- 1982 - 0x7be  :  160 - 0xa0
    "11100000", -- 1983 - 0x7bf  :  224 - 0xe0
    "00111100", -- 1984 - 0x7c0  :   60 - 0x3c
    "11111010", -- 1985 - 0x7c1  :  250 - 0xfa
    "10110001", -- 1986 - 0x7c2  :  177 - 0xb1
    "01110010", -- 1987 - 0x7c3  :  114 - 0x72
    "11110010", -- 1988 - 0x7c4  :  242 - 0xf2
    "11011011", -- 1989 - 0x7c5  :  219 - 0xdb
    "11011111", -- 1990 - 0x7c6  :  223 - 0xdf
    "01011111", -- 1991 - 0x7c7  :   95 - 0x5f
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0
    "00000100", -- 1993 - 0x7c9  :    4 - 0x4
    "01001110", -- 1994 - 0x7ca  :   78 - 0x4e
    "10001100", -- 1995 - 0x7cb  :  140 - 0x8c
    "00001100", -- 1996 - 0x7cc  :   12 - 0xc
    "01111111", -- 1997 - 0x7cd  :  127 - 0x7f
    "11111111", -- 1998 - 0x7ce  :  255 - 0xff
    "11111111", -- 1999 - 0x7cf  :  255 - 0xff
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000001", -- 2003 - 0x7d3  :    1 - 0x1
    "00000001", -- 2004 - 0x7d4  :    1 - 0x1
    "00000001", -- 2005 - 0x7d5  :    1 - 0x1
    "00000110", -- 2006 - 0x7d6  :    6 - 0x6
    "00011110", -- 2007 - 0x7d7  :   30 - 0x1e
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000001", -- 2014 - 0x7de  :    1 - 0x1
    "00000001", -- 2015 - 0x7df  :    1 - 0x1
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "11111111", -- 2024 - 0x7e8  :  255 - 0xff
    "01111111", -- 2025 - 0x7e9  :  127 - 0x7f
    "00111111", -- 2026 - 0x7ea  :   63 - 0x3f
    "00011111", -- 2027 - 0x7eb  :   31 - 0x1f
    "00001111", -- 2028 - 0x7ec  :   15 - 0xf
    "00000111", -- 2029 - 0x7ed  :    7 - 0x7
    "00000011", -- 2030 - 0x7ee  :    3 - 0x3
    "00000001", -- 2031 - 0x7ef  :    1 - 0x1
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0
    "01111100", -- 2033 - 0x7f1  :  124 - 0x7c
    "11010110", -- 2034 - 0x7f2  :  214 - 0xd6
    "10010010", -- 2035 - 0x7f3  :  146 - 0x92
    "10111010", -- 2036 - 0x7f4  :  186 - 0xba
    "11101110", -- 2037 - 0x7f5  :  238 - 0xee
    "11111110", -- 2038 - 0x7f6  :  254 - 0xfe
    "00111000", -- 2039 - 0x7f7  :   56 - 0x38
    "11111111", -- 2040 - 0x7f8  :  255 - 0xff
    "10000011", -- 2041 - 0x7f9  :  131 - 0x83
    "00101001", -- 2042 - 0x7fa  :   41 - 0x29
    "01101101", -- 2043 - 0x7fb  :  109 - 0x6d
    "01000101", -- 2044 - 0x7fc  :   69 - 0x45
    "00010001", -- 2045 - 0x7fd  :   17 - 0x11
    "00000001", -- 2046 - 0x7fe  :    1 - 0x1
    "11000111", -- 2047 - 0x7ff  :  199 - 0xc7
    "00000000", -- 2048 - 0x800  :    0 - 0x0
    "00010101", -- 2049 - 0x801  :   21 - 0x15
    "00111111", -- 2050 - 0x802  :   63 - 0x3f
    "01100010", -- 2051 - 0x803  :   98 - 0x62
    "01011111", -- 2052 - 0x804  :   95 - 0x5f
    "11111111", -- 2053 - 0x805  :  255 - 0xff
    "10011111", -- 2054 - 0x806  :  159 - 0x9f
    "01111101", -- 2055 - 0x807  :  125 - 0x7d
    "00001000", -- 2056 - 0x808  :    8 - 0x8
    "00001000", -- 2057 - 0x809  :    8 - 0x8
    "00000010", -- 2058 - 0x80a  :    2 - 0x2
    "00011111", -- 2059 - 0x80b  :   31 - 0x1f
    "00100010", -- 2060 - 0x80c  :   34 - 0x22
    "00000010", -- 2061 - 0x80d  :    2 - 0x2
    "00000010", -- 2062 - 0x80e  :    2 - 0x2
    "00000000", -- 2063 - 0x80f  :    0 - 0x0
    "00000000", -- 2064 - 0x810  :    0 - 0x0
    "00000000", -- 2065 - 0x811  :    0 - 0x0
    "00000000", -- 2066 - 0x812  :    0 - 0x0
    "00000000", -- 2067 - 0x813  :    0 - 0x0
    "00000000", -- 2068 - 0x814  :    0 - 0x0
    "00000000", -- 2069 - 0x815  :    0 - 0x0
    "00000000", -- 2070 - 0x816  :    0 - 0x0
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "00001000", -- 2072 - 0x818  :    8 - 0x8
    "00001000", -- 2073 - 0x819  :    8 - 0x8
    "00001000", -- 2074 - 0x81a  :    8 - 0x8
    "00001000", -- 2075 - 0x81b  :    8 - 0x8
    "00001000", -- 2076 - 0x81c  :    8 - 0x8
    "00001000", -- 2077 - 0x81d  :    8 - 0x8
    "00001000", -- 2078 - 0x81e  :    8 - 0x8
    "00001000", -- 2079 - 0x81f  :    8 - 0x8
    "00101111", -- 2080 - 0x820  :   47 - 0x2f
    "00011110", -- 2081 - 0x821  :   30 - 0x1e
    "00101111", -- 2082 - 0x822  :   47 - 0x2f
    "00101111", -- 2083 - 0x823  :   47 - 0x2f
    "00101111", -- 2084 - 0x824  :   47 - 0x2f
    "00010101", -- 2085 - 0x825  :   21 - 0x15
    "00001101", -- 2086 - 0x826  :   13 - 0xd
    "00001110", -- 2087 - 0x827  :   14 - 0xe
    "00010000", -- 2088 - 0x828  :   16 - 0x10
    "00011110", -- 2089 - 0x829  :   30 - 0x1e
    "00010000", -- 2090 - 0x82a  :   16 - 0x10
    "01010000", -- 2091 - 0x82b  :   80 - 0x50
    "00010000", -- 2092 - 0x82c  :   16 - 0x10
    "00001000", -- 2093 - 0x82d  :    8 - 0x8
    "00000000", -- 2094 - 0x82e  :    0 - 0x0
    "00000000", -- 2095 - 0x82f  :    0 - 0x0
    "00000000", -- 2096 - 0x830  :    0 - 0x0
    "00000000", -- 2097 - 0x831  :    0 - 0x0
    "00000000", -- 2098 - 0x832  :    0 - 0x0
    "00000000", -- 2099 - 0x833  :    0 - 0x0
    "00000000", -- 2100 - 0x834  :    0 - 0x0
    "00000000", -- 2101 - 0x835  :    0 - 0x0
    "00000000", -- 2102 - 0x836  :    0 - 0x0
    "00000000", -- 2103 - 0x837  :    0 - 0x0
    "00000000", -- 2104 - 0x838  :    0 - 0x0
    "00000000", -- 2105 - 0x839  :    0 - 0x0
    "00000000", -- 2106 - 0x83a  :    0 - 0x0
    "11111110", -- 2107 - 0x83b  :  254 - 0xfe
    "00000000", -- 2108 - 0x83c  :    0 - 0x0
    "00000000", -- 2109 - 0x83d  :    0 - 0x0
    "00000000", -- 2110 - 0x83e  :    0 - 0x0
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "00011100", -- 2112 - 0x840  :   28 - 0x1c
    "00111110", -- 2113 - 0x841  :   62 - 0x3e
    "01111111", -- 2114 - 0x842  :  127 - 0x7f
    "11111111", -- 2115 - 0x843  :  255 - 0xff
    "11111111", -- 2116 - 0x844  :  255 - 0xff
    "11111110", -- 2117 - 0x845  :  254 - 0xfe
    "01111100", -- 2118 - 0x846  :  124 - 0x7c
    "00111000", -- 2119 - 0x847  :   56 - 0x38
    "00011100", -- 2120 - 0x848  :   28 - 0x1c
    "00101010", -- 2121 - 0x849  :   42 - 0x2a
    "01110111", -- 2122 - 0x84a  :  119 - 0x77
    "11101110", -- 2123 - 0x84b  :  238 - 0xee
    "11011101", -- 2124 - 0x84c  :  221 - 0xdd
    "10101010", -- 2125 - 0x84d  :  170 - 0xaa
    "01110100", -- 2126 - 0x84e  :  116 - 0x74
    "00101000", -- 2127 - 0x84f  :   40 - 0x28
    "00000000", -- 2128 - 0x850  :    0 - 0x0
    "11111111", -- 2129 - 0x851  :  255 - 0xff
    "11111111", -- 2130 - 0x852  :  255 - 0xff
    "11111111", -- 2131 - 0x853  :  255 - 0xff
    "11111111", -- 2132 - 0x854  :  255 - 0xff
    "11111111", -- 2133 - 0x855  :  255 - 0xff
    "11111111", -- 2134 - 0x856  :  255 - 0xff
    "11111111", -- 2135 - 0x857  :  255 - 0xff
    "11111111", -- 2136 - 0x858  :  255 - 0xff
    "11111110", -- 2137 - 0x859  :  254 - 0xfe
    "11111110", -- 2138 - 0x85a  :  254 - 0xfe
    "00000000", -- 2139 - 0x85b  :    0 - 0x0
    "11101111", -- 2140 - 0x85c  :  239 - 0xef
    "11101111", -- 2141 - 0x85d  :  239 - 0xef
    "11101111", -- 2142 - 0x85e  :  239 - 0xef
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "11111111", -- 2144 - 0x860  :  255 - 0xff
    "11111111", -- 2145 - 0x861  :  255 - 0xff
    "11111111", -- 2146 - 0x862  :  255 - 0xff
    "11111111", -- 2147 - 0x863  :  255 - 0xff
    "11111111", -- 2148 - 0x864  :  255 - 0xff
    "11111111", -- 2149 - 0x865  :  255 - 0xff
    "11111111", -- 2150 - 0x866  :  255 - 0xff
    "11111111", -- 2151 - 0x867  :  255 - 0xff
    "11111110", -- 2152 - 0x868  :  254 - 0xfe
    "11111110", -- 2153 - 0x869  :  254 - 0xfe
    "11111110", -- 2154 - 0x86a  :  254 - 0xfe
    "00000000", -- 2155 - 0x86b  :    0 - 0x0
    "11101111", -- 2156 - 0x86c  :  239 - 0xef
    "11101111", -- 2157 - 0x86d  :  239 - 0xef
    "11101111", -- 2158 - 0x86e  :  239 - 0xef
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "01111111", -- 2160 - 0x870  :  127 - 0x7f
    "11111111", -- 2161 - 0x871  :  255 - 0xff
    "11111111", -- 2162 - 0x872  :  255 - 0xff
    "11111111", -- 2163 - 0x873  :  255 - 0xff
    "11111111", -- 2164 - 0x874  :  255 - 0xff
    "11111111", -- 2165 - 0x875  :  255 - 0xff
    "11111111", -- 2166 - 0x876  :  255 - 0xff
    "11111111", -- 2167 - 0x877  :  255 - 0xff
    "00000000", -- 2168 - 0x878  :    0 - 0x0
    "01111111", -- 2169 - 0x879  :  127 - 0x7f
    "01011111", -- 2170 - 0x87a  :   95 - 0x5f
    "01111111", -- 2171 - 0x87b  :  127 - 0x7f
    "01111111", -- 2172 - 0x87c  :  127 - 0x7f
    "01111111", -- 2173 - 0x87d  :  127 - 0x7f
    "01111111", -- 2174 - 0x87e  :  127 - 0x7f
    "01111111", -- 2175 - 0x87f  :  127 - 0x7f
    "01101000", -- 2176 - 0x880  :  104 - 0x68
    "01001110", -- 2177 - 0x881  :   78 - 0x4e
    "11100000", -- 2178 - 0x882  :  224 - 0xe0
    "11100000", -- 2179 - 0x883  :  224 - 0xe0
    "11100000", -- 2180 - 0x884  :  224 - 0xe0
    "11110000", -- 2181 - 0x885  :  240 - 0xf0
    "11111000", -- 2182 - 0x886  :  248 - 0xf8
    "11111100", -- 2183 - 0x887  :  252 - 0xfc
    "10111000", -- 2184 - 0x888  :  184 - 0xb8
    "10011110", -- 2185 - 0x889  :  158 - 0x9e
    "10000000", -- 2186 - 0x88a  :  128 - 0x80
    "11000000", -- 2187 - 0x88b  :  192 - 0xc0
    "11100000", -- 2188 - 0x88c  :  224 - 0xe0
    "11110000", -- 2189 - 0x88d  :  240 - 0xf0
    "11111000", -- 2190 - 0x88e  :  248 - 0xf8
    "01111100", -- 2191 - 0x88f  :  124 - 0x7c
    "00111111", -- 2192 - 0x890  :   63 - 0x3f
    "01011100", -- 2193 - 0x891  :   92 - 0x5c
    "00111001", -- 2194 - 0x892  :   57 - 0x39
    "00111011", -- 2195 - 0x893  :   59 - 0x3b
    "10111011", -- 2196 - 0x894  :  187 - 0xbb
    "11111001", -- 2197 - 0x895  :  249 - 0xf9
    "11111100", -- 2198 - 0x896  :  252 - 0xfc
    "11111110", -- 2199 - 0x897  :  254 - 0xfe
    "00000000", -- 2200 - 0x898  :    0 - 0x0
    "00100011", -- 2201 - 0x899  :   35 - 0x23
    "01010111", -- 2202 - 0x89a  :   87 - 0x57
    "01001111", -- 2203 - 0x89b  :   79 - 0x4f
    "01010111", -- 2204 - 0x89c  :   87 - 0x57
    "00100111", -- 2205 - 0x89d  :   39 - 0x27
    "11000011", -- 2206 - 0x89e  :  195 - 0xc3
    "00100001", -- 2207 - 0x89f  :   33 - 0x21
    "11000000", -- 2208 - 0x8a0  :  192 - 0xc0
    "11110000", -- 2209 - 0x8a1  :  240 - 0xf0
    "11110000", -- 2210 - 0x8a2  :  240 - 0xf0
    "11110000", -- 2211 - 0x8a3  :  240 - 0xf0
    "11110000", -- 2212 - 0x8a4  :  240 - 0xf0
    "11100000", -- 2213 - 0x8a5  :  224 - 0xe0
    "11000000", -- 2214 - 0x8a6  :  192 - 0xc0
    "00000000", -- 2215 - 0x8a7  :    0 - 0x0
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0
    "00110000", -- 2217 - 0x8a9  :   48 - 0x30
    "01110000", -- 2218 - 0x8aa  :  112 - 0x70
    "01110000", -- 2219 - 0x8ab  :  112 - 0x70
    "11110000", -- 2220 - 0x8ac  :  240 - 0xf0
    "11100000", -- 2221 - 0x8ad  :  224 - 0xe0
    "11000000", -- 2222 - 0x8ae  :  192 - 0xc0
    "00000000", -- 2223 - 0x8af  :    0 - 0x0
    "11111110", -- 2224 - 0x8b0  :  254 - 0xfe
    "11111100", -- 2225 - 0x8b1  :  252 - 0xfc
    "01100001", -- 2226 - 0x8b2  :   97 - 0x61
    "00001111", -- 2227 - 0x8b3  :   15 - 0xf
    "11111111", -- 2228 - 0x8b4  :  255 - 0xff
    "11111110", -- 2229 - 0x8b5  :  254 - 0xfe
    "11110000", -- 2230 - 0x8b6  :  240 - 0xf0
    "11100000", -- 2231 - 0x8b7  :  224 - 0xe0
    "00010011", -- 2232 - 0x8b8  :   19 - 0x13
    "00001111", -- 2233 - 0x8b9  :   15 - 0xf
    "00011110", -- 2234 - 0x8ba  :   30 - 0x1e
    "11110000", -- 2235 - 0x8bb  :  240 - 0xf0
    "11111100", -- 2236 - 0x8bc  :  252 - 0xfc
    "11111000", -- 2237 - 0x8bd  :  248 - 0xf8
    "11110000", -- 2238 - 0x8be  :  240 - 0xf0
    "11100000", -- 2239 - 0x8bf  :  224 - 0xe0
    "01101110", -- 2240 - 0x8c0  :  110 - 0x6e
    "01000000", -- 2241 - 0x8c1  :   64 - 0x40
    "11100000", -- 2242 - 0x8c2  :  224 - 0xe0
    "11100000", -- 2243 - 0x8c3  :  224 - 0xe0
    "11100000", -- 2244 - 0x8c4  :  224 - 0xe0
    "11100000", -- 2245 - 0x8c5  :  224 - 0xe0
    "11100000", -- 2246 - 0x8c6  :  224 - 0xe0
    "11000000", -- 2247 - 0x8c7  :  192 - 0xc0
    "10111110", -- 2248 - 0x8c8  :  190 - 0xbe
    "10010000", -- 2249 - 0x8c9  :  144 - 0x90
    "10000000", -- 2250 - 0x8ca  :  128 - 0x80
    "11000000", -- 2251 - 0x8cb  :  192 - 0xc0
    "11000000", -- 2252 - 0x8cc  :  192 - 0xc0
    "10000000", -- 2253 - 0x8cd  :  128 - 0x80
    "00000000", -- 2254 - 0x8ce  :    0 - 0x0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "00000001", -- 2256 - 0x8d0  :    1 - 0x1
    "00000001", -- 2257 - 0x8d1  :    1 - 0x1
    "00000011", -- 2258 - 0x8d2  :    3 - 0x3
    "00000011", -- 2259 - 0x8d3  :    3 - 0x3
    "00000111", -- 2260 - 0x8d4  :    7 - 0x7
    "01111111", -- 2261 - 0x8d5  :  127 - 0x7f
    "01111111", -- 2262 - 0x8d6  :  127 - 0x7f
    "00111111", -- 2263 - 0x8d7  :   63 - 0x3f
    "00000001", -- 2264 - 0x8d8  :    1 - 0x1
    "00000001", -- 2265 - 0x8d9  :    1 - 0x1
    "00000011", -- 2266 - 0x8da  :    3 - 0x3
    "00000011", -- 2267 - 0x8db  :    3 - 0x3
    "00000111", -- 2268 - 0x8dc  :    7 - 0x7
    "01111111", -- 2269 - 0x8dd  :  127 - 0x7f
    "01111101", -- 2270 - 0x8de  :  125 - 0x7d
    "00111101", -- 2271 - 0x8df  :   61 - 0x3d
    "00000110", -- 2272 - 0x8e0  :    6 - 0x6
    "00000111", -- 2273 - 0x8e1  :    7 - 0x7
    "00111111", -- 2274 - 0x8e2  :   63 - 0x3f
    "00111100", -- 2275 - 0x8e3  :   60 - 0x3c
    "00011001", -- 2276 - 0x8e4  :   25 - 0x19
    "01111011", -- 2277 - 0x8e5  :  123 - 0x7b
    "01111111", -- 2278 - 0x8e6  :  127 - 0x7f
    "00111111", -- 2279 - 0x8e7  :   63 - 0x3f
    "00000110", -- 2280 - 0x8e8  :    6 - 0x6
    "00000100", -- 2281 - 0x8e9  :    4 - 0x4
    "00110000", -- 2282 - 0x8ea  :   48 - 0x30
    "00100011", -- 2283 - 0x8eb  :   35 - 0x23
    "00000110", -- 2284 - 0x8ec  :    6 - 0x6
    "01100100", -- 2285 - 0x8ed  :  100 - 0x64
    "01100000", -- 2286 - 0x8ee  :   96 - 0x60
    "00000000", -- 2287 - 0x8ef  :    0 - 0x0
    "00111111", -- 2288 - 0x8f0  :   63 - 0x3f
    "01111111", -- 2289 - 0x8f1  :  127 - 0x7f
    "01111111", -- 2290 - 0x8f2  :  127 - 0x7f
    "00011111", -- 2291 - 0x8f3  :   31 - 0x1f
    "00111111", -- 2292 - 0x8f4  :   63 - 0x3f
    "00111111", -- 2293 - 0x8f5  :   63 - 0x3f
    "00000111", -- 2294 - 0x8f6  :    7 - 0x7
    "00000110", -- 2295 - 0x8f7  :    6 - 0x6
    "00000000", -- 2296 - 0x8f8  :    0 - 0x0
    "01100000", -- 2297 - 0x8f9  :   96 - 0x60
    "01100000", -- 2298 - 0x8fa  :   96 - 0x60
    "00000000", -- 2299 - 0x8fb  :    0 - 0x0
    "00100000", -- 2300 - 0x8fc  :   32 - 0x20
    "00110000", -- 2301 - 0x8fd  :   48 - 0x30
    "00000100", -- 2302 - 0x8fe  :    4 - 0x4
    "00000110", -- 2303 - 0x8ff  :    6 - 0x6
    "00000011", -- 2304 - 0x900  :    3 - 0x3
    "00000111", -- 2305 - 0x901  :    7 - 0x7
    "00001111", -- 2306 - 0x902  :   15 - 0xf
    "00001111", -- 2307 - 0x903  :   15 - 0xf
    "00001111", -- 2308 - 0x904  :   15 - 0xf
    "00001111", -- 2309 - 0x905  :   15 - 0xf
    "00000111", -- 2310 - 0x906  :    7 - 0x7
    "00000011", -- 2311 - 0x907  :    3 - 0x3
    "00000000", -- 2312 - 0x908  :    0 - 0x0
    "00000001", -- 2313 - 0x909  :    1 - 0x1
    "00000001", -- 2314 - 0x90a  :    1 - 0x1
    "00000000", -- 2315 - 0x90b  :    0 - 0x0
    "00000000", -- 2316 - 0x90c  :    0 - 0x0
    "00000000", -- 2317 - 0x90d  :    0 - 0x0
    "00000000", -- 2318 - 0x90e  :    0 - 0x0
    "00000000", -- 2319 - 0x90f  :    0 - 0x0
    "11111000", -- 2320 - 0x910  :  248 - 0xf8
    "11111000", -- 2321 - 0x911  :  248 - 0xf8
    "11111000", -- 2322 - 0x912  :  248 - 0xf8
    "10100000", -- 2323 - 0x913  :  160 - 0xa0
    "11100001", -- 2324 - 0x914  :  225 - 0xe1
    "11111111", -- 2325 - 0x915  :  255 - 0xff
    "11111111", -- 2326 - 0x916  :  255 - 0xff
    "11111111", -- 2327 - 0x917  :  255 - 0xff
    "11111110", -- 2328 - 0x918  :  254 - 0xfe
    "11111111", -- 2329 - 0x919  :  255 - 0xff
    "11111111", -- 2330 - 0x91a  :  255 - 0xff
    "01000000", -- 2331 - 0x91b  :   64 - 0x40
    "00000001", -- 2332 - 0x91c  :    1 - 0x1
    "00000011", -- 2333 - 0x91d  :    3 - 0x3
    "00000011", -- 2334 - 0x91e  :    3 - 0x3
    "00000011", -- 2335 - 0x91f  :    3 - 0x3
    "00001111", -- 2336 - 0x920  :   15 - 0xf
    "00001111", -- 2337 - 0x921  :   15 - 0xf
    "00001111", -- 2338 - 0x922  :   15 - 0xf
    "00011111", -- 2339 - 0x923  :   31 - 0x1f
    "00011111", -- 2340 - 0x924  :   31 - 0x1f
    "00011111", -- 2341 - 0x925  :   31 - 0x1f
    "00001111", -- 2342 - 0x926  :   15 - 0xf
    "00000111", -- 2343 - 0x927  :    7 - 0x7
    "00000001", -- 2344 - 0x928  :    1 - 0x1
    "00000001", -- 2345 - 0x929  :    1 - 0x1
    "00000000", -- 2346 - 0x92a  :    0 - 0x0
    "00000000", -- 2347 - 0x92b  :    0 - 0x0
    "00000000", -- 2348 - 0x92c  :    0 - 0x0
    "00000000", -- 2349 - 0x92d  :    0 - 0x0
    "00000000", -- 2350 - 0x92e  :    0 - 0x0
    "00000000", -- 2351 - 0x92f  :    0 - 0x0
    "11100000", -- 2352 - 0x930  :  224 - 0xe0
    "11111000", -- 2353 - 0x931  :  248 - 0xf8
    "11111000", -- 2354 - 0x932  :  248 - 0xf8
    "11111000", -- 2355 - 0x933  :  248 - 0xf8
    "11111111", -- 2356 - 0x934  :  255 - 0xff
    "11111110", -- 2357 - 0x935  :  254 - 0xfe
    "11110000", -- 2358 - 0x936  :  240 - 0xf0
    "11000000", -- 2359 - 0x937  :  192 - 0xc0
    "11100000", -- 2360 - 0x938  :  224 - 0xe0
    "11111110", -- 2361 - 0x939  :  254 - 0xfe
    "11111111", -- 2362 - 0x93a  :  255 - 0xff
    "01111111", -- 2363 - 0x93b  :  127 - 0x7f
    "00000011", -- 2364 - 0x93c  :    3 - 0x3
    "00000010", -- 2365 - 0x93d  :    2 - 0x2
    "00000000", -- 2366 - 0x93e  :    0 - 0x0
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000001", -- 2368 - 0x940  :    1 - 0x1
    "00001111", -- 2369 - 0x941  :   15 - 0xf
    "00001111", -- 2370 - 0x942  :   15 - 0xf
    "00011111", -- 2371 - 0x943  :   31 - 0x1f
    "00111001", -- 2372 - 0x944  :   57 - 0x39
    "00110011", -- 2373 - 0x945  :   51 - 0x33
    "00110111", -- 2374 - 0x946  :   55 - 0x37
    "01111111", -- 2375 - 0x947  :  127 - 0x7f
    "00000001", -- 2376 - 0x948  :    1 - 0x1
    "00001101", -- 2377 - 0x949  :   13 - 0xd
    "00001000", -- 2378 - 0x94a  :    8 - 0x8
    "00000000", -- 2379 - 0x94b  :    0 - 0x0
    "00110110", -- 2380 - 0x94c  :   54 - 0x36
    "00101100", -- 2381 - 0x94d  :   44 - 0x2c
    "00001000", -- 2382 - 0x94e  :    8 - 0x8
    "01100000", -- 2383 - 0x94f  :   96 - 0x60
    "01111111", -- 2384 - 0x950  :  127 - 0x7f
    "00111111", -- 2385 - 0x951  :   63 - 0x3f
    "00111111", -- 2386 - 0x952  :   63 - 0x3f
    "00111111", -- 2387 - 0x953  :   63 - 0x3f
    "00011111", -- 2388 - 0x954  :   31 - 0x1f
    "00001111", -- 2389 - 0x955  :   15 - 0xf
    "00001111", -- 2390 - 0x956  :   15 - 0xf
    "00000001", -- 2391 - 0x957  :    1 - 0x1
    "01100000", -- 2392 - 0x958  :   96 - 0x60
    "00000000", -- 2393 - 0x959  :    0 - 0x0
    "00100000", -- 2394 - 0x95a  :   32 - 0x20
    "00110000", -- 2395 - 0x95b  :   48 - 0x30
    "00000000", -- 2396 - 0x95c  :    0 - 0x0
    "00001000", -- 2397 - 0x95d  :    8 - 0x8
    "00001101", -- 2398 - 0x95e  :   13 - 0xd
    "00000001", -- 2399 - 0x95f  :    1 - 0x1
    "00000000", -- 2400 - 0x960  :    0 - 0x0
    "00000000", -- 2401 - 0x961  :    0 - 0x0
    "00000011", -- 2402 - 0x962  :    3 - 0x3
    "00000011", -- 2403 - 0x963  :    3 - 0x3
    "01000111", -- 2404 - 0x964  :   71 - 0x47
    "01100111", -- 2405 - 0x965  :  103 - 0x67
    "01110111", -- 2406 - 0x966  :  119 - 0x77
    "01110111", -- 2407 - 0x967  :  119 - 0x77
    "00000001", -- 2408 - 0x968  :    1 - 0x1
    "00000001", -- 2409 - 0x969  :    1 - 0x1
    "00000011", -- 2410 - 0x96a  :    3 - 0x3
    "01000011", -- 2411 - 0x96b  :   67 - 0x43
    "01100111", -- 2412 - 0x96c  :  103 - 0x67
    "01110111", -- 2413 - 0x96d  :  119 - 0x77
    "01111011", -- 2414 - 0x96e  :  123 - 0x7b
    "01111000", -- 2415 - 0x96f  :  120 - 0x78
    "00000000", -- 2416 - 0x970  :    0 - 0x0
    "00000000", -- 2417 - 0x971  :    0 - 0x0
    "00000000", -- 2418 - 0x972  :    0 - 0x0
    "00000000", -- 2419 - 0x973  :    0 - 0x0
    "10001000", -- 2420 - 0x974  :  136 - 0x88
    "10011000", -- 2421 - 0x975  :  152 - 0x98
    "11111000", -- 2422 - 0x976  :  248 - 0xf8
    "11110000", -- 2423 - 0x977  :  240 - 0xf0
    "00000000", -- 2424 - 0x978  :    0 - 0x0
    "00000000", -- 2425 - 0x979  :    0 - 0x0
    "10000000", -- 2426 - 0x97a  :  128 - 0x80
    "10000100", -- 2427 - 0x97b  :  132 - 0x84
    "11001100", -- 2428 - 0x97c  :  204 - 0xcc
    "11011100", -- 2429 - 0x97d  :  220 - 0xdc
    "10111100", -- 2430 - 0x97e  :  188 - 0xbc
    "00111100", -- 2431 - 0x97f  :   60 - 0x3c
    "01111110", -- 2432 - 0x980  :  126 - 0x7e
    "01111111", -- 2433 - 0x981  :  127 - 0x7f
    "11111111", -- 2434 - 0x982  :  255 - 0xff
    "00011111", -- 2435 - 0x983  :   31 - 0x1f
    "00000111", -- 2436 - 0x984  :    7 - 0x7
    "00110000", -- 2437 - 0x985  :   48 - 0x30
    "00011100", -- 2438 - 0x986  :   28 - 0x1c
    "00001100", -- 2439 - 0x987  :   12 - 0xc
    "00110011", -- 2440 - 0x988  :   51 - 0x33
    "00000111", -- 2441 - 0x989  :    7 - 0x7
    "00000111", -- 2442 - 0x98a  :    7 - 0x7
    "11100011", -- 2443 - 0x98b  :  227 - 0xe3
    "00111000", -- 2444 - 0x98c  :   56 - 0x38
    "00111111", -- 2445 - 0x98d  :   63 - 0x3f
    "00011100", -- 2446 - 0x98e  :   28 - 0x1c
    "00001100", -- 2447 - 0x98f  :   12 - 0xc
    "01111110", -- 2448 - 0x990  :  126 - 0x7e
    "00111000", -- 2449 - 0x991  :   56 - 0x38
    "11110110", -- 2450 - 0x992  :  246 - 0xf6
    "11101101", -- 2451 - 0x993  :  237 - 0xed
    "11011111", -- 2452 - 0x994  :  223 - 0xdf
    "00111000", -- 2453 - 0x995  :   56 - 0x38
    "01110000", -- 2454 - 0x996  :  112 - 0x70
    "01100000", -- 2455 - 0x997  :   96 - 0x60
    "10011000", -- 2456 - 0x998  :  152 - 0x98
    "11000111", -- 2457 - 0x999  :  199 - 0xc7
    "11001000", -- 2458 - 0x99a  :  200 - 0xc8
    "10010010", -- 2459 - 0x99b  :  146 - 0x92
    "00110000", -- 2460 - 0x99c  :   48 - 0x30
    "11111000", -- 2461 - 0x99d  :  248 - 0xf8
    "01110000", -- 2462 - 0x99e  :  112 - 0x70
    "01100000", -- 2463 - 0x99f  :   96 - 0x60
    "00000000", -- 2464 - 0x9a0  :    0 - 0x0
    "00000000", -- 2465 - 0x9a1  :    0 - 0x0
    "00000000", -- 2466 - 0x9a2  :    0 - 0x0
    "00000011", -- 2467 - 0x9a3  :    3 - 0x3
    "00000011", -- 2468 - 0x9a4  :    3 - 0x3
    "01000111", -- 2469 - 0x9a5  :   71 - 0x47
    "01100111", -- 2470 - 0x9a6  :  103 - 0x67
    "01110111", -- 2471 - 0x9a7  :  119 - 0x77
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0
    "00000001", -- 2473 - 0x9a9  :    1 - 0x1
    "00000001", -- 2474 - 0x9aa  :    1 - 0x1
    "00000011", -- 2475 - 0x9ab  :    3 - 0x3
    "01000011", -- 2476 - 0x9ac  :   67 - 0x43
    "01100111", -- 2477 - 0x9ad  :  103 - 0x67
    "01110111", -- 2478 - 0x9ae  :  119 - 0x77
    "01111011", -- 2479 - 0x9af  :  123 - 0x7b
    "00000000", -- 2480 - 0x9b0  :    0 - 0x0
    "00000000", -- 2481 - 0x9b1  :    0 - 0x0
    "00000000", -- 2482 - 0x9b2  :    0 - 0x0
    "00000000", -- 2483 - 0x9b3  :    0 - 0x0
    "00000000", -- 2484 - 0x9b4  :    0 - 0x0
    "10001000", -- 2485 - 0x9b5  :  136 - 0x88
    "10011000", -- 2486 - 0x9b6  :  152 - 0x98
    "11111000", -- 2487 - 0x9b7  :  248 - 0xf8
    "00000000", -- 2488 - 0x9b8  :    0 - 0x0
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "00000000", -- 2490 - 0x9ba  :    0 - 0x0
    "10000000", -- 2491 - 0x9bb  :  128 - 0x80
    "10000100", -- 2492 - 0x9bc  :  132 - 0x84
    "11001100", -- 2493 - 0x9bd  :  204 - 0xcc
    "11011100", -- 2494 - 0x9be  :  220 - 0xdc
    "10111100", -- 2495 - 0x9bf  :  188 - 0xbc
    "01110111", -- 2496 - 0x9c0  :  119 - 0x77
    "01111110", -- 2497 - 0x9c1  :  126 - 0x7e
    "01111111", -- 2498 - 0x9c2  :  127 - 0x7f
    "11111111", -- 2499 - 0x9c3  :  255 - 0xff
    "00011111", -- 2500 - 0x9c4  :   31 - 0x1f
    "00000111", -- 2501 - 0x9c5  :    7 - 0x7
    "01110000", -- 2502 - 0x9c6  :  112 - 0x70
    "11110000", -- 2503 - 0x9c7  :  240 - 0xf0
    "01111000", -- 2504 - 0x9c8  :  120 - 0x78
    "00110011", -- 2505 - 0x9c9  :   51 - 0x33
    "00000111", -- 2506 - 0x9ca  :    7 - 0x7
    "00000111", -- 2507 - 0x9cb  :    7 - 0x7
    "11100011", -- 2508 - 0x9cc  :  227 - 0xe3
    "00111000", -- 2509 - 0x9cd  :   56 - 0x38
    "01111111", -- 2510 - 0x9ce  :  127 - 0x7f
    "11110000", -- 2511 - 0x9cf  :  240 - 0xf0
    "11110000", -- 2512 - 0x9d0  :  240 - 0xf0
    "01111110", -- 2513 - 0x9d1  :  126 - 0x7e
    "00111000", -- 2514 - 0x9d2  :   56 - 0x38
    "11110110", -- 2515 - 0x9d3  :  246 - 0xf6
    "11101101", -- 2516 - 0x9d4  :  237 - 0xed
    "11011111", -- 2517 - 0x9d5  :  223 - 0xdf
    "00111000", -- 2518 - 0x9d6  :   56 - 0x38
    "00111100", -- 2519 - 0x9d7  :   60 - 0x3c
    "00111100", -- 2520 - 0x9d8  :   60 - 0x3c
    "10011000", -- 2521 - 0x9d9  :  152 - 0x98
    "11000111", -- 2522 - 0x9da  :  199 - 0xc7
    "11001000", -- 2523 - 0x9db  :  200 - 0xc8
    "10010010", -- 2524 - 0x9dc  :  146 - 0x92
    "00110000", -- 2525 - 0x9dd  :   48 - 0x30
    "11111000", -- 2526 - 0x9de  :  248 - 0xf8
    "00111100", -- 2527 - 0x9df  :   60 - 0x3c
    "00000011", -- 2528 - 0x9e0  :    3 - 0x3
    "00000111", -- 2529 - 0x9e1  :    7 - 0x7
    "00001010", -- 2530 - 0x9e2  :   10 - 0xa
    "00011010", -- 2531 - 0x9e3  :   26 - 0x1a
    "00011100", -- 2532 - 0x9e4  :   28 - 0x1c
    "00011110", -- 2533 - 0x9e5  :   30 - 0x1e
    "00001011", -- 2534 - 0x9e6  :   11 - 0xb
    "00001000", -- 2535 - 0x9e7  :    8 - 0x8
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0
    "00010000", -- 2537 - 0x9e9  :   16 - 0x10
    "01111111", -- 2538 - 0x9ea  :  127 - 0x7f
    "01111111", -- 2539 - 0x9eb  :  127 - 0x7f
    "01111111", -- 2540 - 0x9ec  :  127 - 0x7f
    "00011111", -- 2541 - 0x9ed  :   31 - 0x1f
    "00001111", -- 2542 - 0x9ee  :   15 - 0xf
    "00001111", -- 2543 - 0x9ef  :   15 - 0xf
    "00011100", -- 2544 - 0x9f0  :   28 - 0x1c
    "00111111", -- 2545 - 0x9f1  :   63 - 0x3f
    "00111111", -- 2546 - 0x9f2  :   63 - 0x3f
    "00111101", -- 2547 - 0x9f3  :   61 - 0x3d
    "00111111", -- 2548 - 0x9f4  :   63 - 0x3f
    "00011111", -- 2549 - 0x9f5  :   31 - 0x1f
    "00000000", -- 2550 - 0x9f6  :    0 - 0x0
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "00000011", -- 2552 - 0x9f8  :    3 - 0x3
    "00110011", -- 2553 - 0x9f9  :   51 - 0x33
    "00111001", -- 2554 - 0x9fa  :   57 - 0x39
    "00111010", -- 2555 - 0x9fb  :   58 - 0x3a
    "00111000", -- 2556 - 0x9fc  :   56 - 0x38
    "00011000", -- 2557 - 0x9fd  :   24 - 0x18
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00000000", -- 2560 - 0xa00  :    0 - 0x0
    "00000000", -- 2561 - 0xa01  :    0 - 0x0
    "00000100", -- 2562 - 0xa02  :    4 - 0x4
    "01001100", -- 2563 - 0xa03  :   76 - 0x4c
    "01001110", -- 2564 - 0xa04  :   78 - 0x4e
    "01001110", -- 2565 - 0xa05  :   78 - 0x4e
    "01000110", -- 2566 - 0xa06  :   70 - 0x46
    "01101111", -- 2567 - 0xa07  :  111 - 0x6f
    "00010000", -- 2568 - 0xa08  :   16 - 0x10
    "00111000", -- 2569 - 0xa09  :   56 - 0x38
    "00111100", -- 2570 - 0xa0a  :   60 - 0x3c
    "01110100", -- 2571 - 0xa0b  :  116 - 0x74
    "01110110", -- 2572 - 0xa0c  :  118 - 0x76
    "01110110", -- 2573 - 0xa0d  :  118 - 0x76
    "01111110", -- 2574 - 0xa0e  :  126 - 0x7e
    "01111101", -- 2575 - 0xa0f  :  125 - 0x7d
    "00000000", -- 2576 - 0xa10  :    0 - 0x0
    "00011111", -- 2577 - 0xa11  :   31 - 0x1f
    "00111111", -- 2578 - 0xa12  :   63 - 0x3f
    "00111111", -- 2579 - 0xa13  :   63 - 0x3f
    "01001111", -- 2580 - 0xa14  :   79 - 0x4f
    "01011111", -- 2581 - 0xa15  :   95 - 0x5f
    "01111111", -- 2582 - 0xa16  :  127 - 0x7f
    "01111111", -- 2583 - 0xa17  :  127 - 0x7f
    "00000000", -- 2584 - 0xa18  :    0 - 0x0
    "00000000", -- 2585 - 0xa19  :    0 - 0x0
    "00010001", -- 2586 - 0xa1a  :   17 - 0x11
    "00001010", -- 2587 - 0xa1b  :   10 - 0xa
    "00110100", -- 2588 - 0xa1c  :   52 - 0x34
    "00101010", -- 2589 - 0xa1d  :   42 - 0x2a
    "01010001", -- 2590 - 0xa1e  :   81 - 0x51
    "00100000", -- 2591 - 0xa1f  :   32 - 0x20
    "01111111", -- 2592 - 0xa20  :  127 - 0x7f
    "01100111", -- 2593 - 0xa21  :  103 - 0x67
    "10100011", -- 2594 - 0xa22  :  163 - 0xa3
    "10110000", -- 2595 - 0xa23  :  176 - 0xb0
    "11011000", -- 2596 - 0xa24  :  216 - 0xd8
    "11011110", -- 2597 - 0xa25  :  222 - 0xde
    "11011100", -- 2598 - 0xa26  :  220 - 0xdc
    "11001000", -- 2599 - 0xa27  :  200 - 0xc8
    "01111111", -- 2600 - 0xa28  :  127 - 0x7f
    "01100111", -- 2601 - 0xa29  :  103 - 0x67
    "01100011", -- 2602 - 0xa2a  :   99 - 0x63
    "01110000", -- 2603 - 0xa2b  :  112 - 0x70
    "00111000", -- 2604 - 0xa2c  :   56 - 0x38
    "00111110", -- 2605 - 0xa2d  :   62 - 0x3e
    "01111100", -- 2606 - 0xa2e  :  124 - 0x7c
    "10111000", -- 2607 - 0xa2f  :  184 - 0xb8
    "01111111", -- 2608 - 0xa30  :  127 - 0x7f
    "01111111", -- 2609 - 0xa31  :  127 - 0x7f
    "01111111", -- 2610 - 0xa32  :  127 - 0x7f
    "00011111", -- 2611 - 0xa33  :   31 - 0x1f
    "01000111", -- 2612 - 0xa34  :   71 - 0x47
    "01110000", -- 2613 - 0xa35  :  112 - 0x70
    "01110000", -- 2614 - 0xa36  :  112 - 0x70
    "00111001", -- 2615 - 0xa37  :   57 - 0x39
    "01010001", -- 2616 - 0xa38  :   81 - 0x51
    "00001010", -- 2617 - 0xa39  :   10 - 0xa
    "00000100", -- 2618 - 0xa3a  :    4 - 0x4
    "11101010", -- 2619 - 0xa3b  :  234 - 0xea
    "01111001", -- 2620 - 0xa3c  :  121 - 0x79
    "01111111", -- 2621 - 0xa3d  :  127 - 0x7f
    "01110000", -- 2622 - 0xa3e  :  112 - 0x70
    "00111001", -- 2623 - 0xa3f  :   57 - 0x39
    "11101000", -- 2624 - 0xa40  :  232 - 0xe8
    "11101000", -- 2625 - 0xa41  :  232 - 0xe8
    "11100000", -- 2626 - 0xa42  :  224 - 0xe0
    "11000000", -- 2627 - 0xa43  :  192 - 0xc0
    "00010000", -- 2628 - 0xa44  :   16 - 0x10
    "01110000", -- 2629 - 0xa45  :  112 - 0x70
    "11100000", -- 2630 - 0xa46  :  224 - 0xe0
    "11000000", -- 2631 - 0xa47  :  192 - 0xc0
    "01011000", -- 2632 - 0xa48  :   88 - 0x58
    "00111000", -- 2633 - 0xa49  :   56 - 0x38
    "00010000", -- 2634 - 0xa4a  :   16 - 0x10
    "00110000", -- 2635 - 0xa4b  :   48 - 0x30
    "11110000", -- 2636 - 0xa4c  :  240 - 0xf0
    "11110000", -- 2637 - 0xa4d  :  240 - 0xf0
    "11100000", -- 2638 - 0xa4e  :  224 - 0xe0
    "11000000", -- 2639 - 0xa4f  :  192 - 0xc0
    "00000000", -- 2640 - 0xa50  :    0 - 0x0
    "00000000", -- 2641 - 0xa51  :    0 - 0x0
    "00000000", -- 2642 - 0xa52  :    0 - 0x0
    "00100000", -- 2643 - 0xa53  :   32 - 0x20
    "01100110", -- 2644 - 0xa54  :  102 - 0x66
    "01100110", -- 2645 - 0xa55  :  102 - 0x66
    "01100110", -- 2646 - 0xa56  :  102 - 0x66
    "01100010", -- 2647 - 0xa57  :   98 - 0x62
    "00000000", -- 2648 - 0xa58  :    0 - 0x0
    "00001000", -- 2649 - 0xa59  :    8 - 0x8
    "00011100", -- 2650 - 0xa5a  :   28 - 0x1c
    "00111100", -- 2651 - 0xa5b  :   60 - 0x3c
    "01111010", -- 2652 - 0xa5c  :  122 - 0x7a
    "01111010", -- 2653 - 0xa5d  :  122 - 0x7a
    "01111010", -- 2654 - 0xa5e  :  122 - 0x7a
    "01111110", -- 2655 - 0xa5f  :  126 - 0x7e
    "00000000", -- 2656 - 0xa60  :    0 - 0x0
    "00000000", -- 2657 - 0xa61  :    0 - 0x0
    "00011111", -- 2658 - 0xa62  :   31 - 0x1f
    "00111111", -- 2659 - 0xa63  :   63 - 0x3f
    "01111111", -- 2660 - 0xa64  :  127 - 0x7f
    "01001111", -- 2661 - 0xa65  :   79 - 0x4f
    "01011111", -- 2662 - 0xa66  :   95 - 0x5f
    "01111111", -- 2663 - 0xa67  :  127 - 0x7f
    "00000000", -- 2664 - 0xa68  :    0 - 0x0
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "00000000", -- 2666 - 0xa6a  :    0 - 0x0
    "00010001", -- 2667 - 0xa6b  :   17 - 0x11
    "00001010", -- 2668 - 0xa6c  :   10 - 0xa
    "00110100", -- 2669 - 0xa6d  :   52 - 0x34
    "00101010", -- 2670 - 0xa6e  :   42 - 0x2a
    "01010001", -- 2671 - 0xa6f  :   81 - 0x51
    "01110111", -- 2672 - 0xa70  :  119 - 0x77
    "01111111", -- 2673 - 0xa71  :  127 - 0x7f
    "00111111", -- 2674 - 0xa72  :   63 - 0x3f
    "10110111", -- 2675 - 0xa73  :  183 - 0xb7
    "10110011", -- 2676 - 0xa74  :  179 - 0xb3
    "11011011", -- 2677 - 0xa75  :  219 - 0xdb
    "11011010", -- 2678 - 0xa76  :  218 - 0xda
    "11011000", -- 2679 - 0xa77  :  216 - 0xd8
    "01111111", -- 2680 - 0xa78  :  127 - 0x7f
    "01111101", -- 2681 - 0xa79  :  125 - 0x7d
    "00111111", -- 2682 - 0xa7a  :   63 - 0x3f
    "00110111", -- 2683 - 0xa7b  :   55 - 0x37
    "00110011", -- 2684 - 0xa7c  :   51 - 0x33
    "00111011", -- 2685 - 0xa7d  :   59 - 0x3b
    "00111010", -- 2686 - 0xa7e  :   58 - 0x3a
    "01111000", -- 2687 - 0xa7f  :  120 - 0x78
    "01111111", -- 2688 - 0xa80  :  127 - 0x7f
    "01111111", -- 2689 - 0xa81  :  127 - 0x7f
    "01111111", -- 2690 - 0xa82  :  127 - 0x7f
    "01111111", -- 2691 - 0xa83  :  127 - 0x7f
    "00011111", -- 2692 - 0xa84  :   31 - 0x1f
    "00000111", -- 2693 - 0xa85  :    7 - 0x7
    "01110000", -- 2694 - 0xa86  :  112 - 0x70
    "11110000", -- 2695 - 0xa87  :  240 - 0xf0
    "00100000", -- 2696 - 0xa88  :   32 - 0x20
    "01010001", -- 2697 - 0xa89  :   81 - 0x51
    "00001010", -- 2698 - 0xa8a  :   10 - 0xa
    "00000100", -- 2699 - 0xa8b  :    4 - 0x4
    "11101010", -- 2700 - 0xa8c  :  234 - 0xea
    "00111001", -- 2701 - 0xa8d  :   57 - 0x39
    "01111111", -- 2702 - 0xa8e  :  127 - 0x7f
    "11110000", -- 2703 - 0xa8f  :  240 - 0xf0
    "11001100", -- 2704 - 0xa90  :  204 - 0xcc
    "11101000", -- 2705 - 0xa91  :  232 - 0xe8
    "11101000", -- 2706 - 0xa92  :  232 - 0xe8
    "11100000", -- 2707 - 0xa93  :  224 - 0xe0
    "11000000", -- 2708 - 0xa94  :  192 - 0xc0
    "00011000", -- 2709 - 0xa95  :   24 - 0x18
    "01111100", -- 2710 - 0xa96  :  124 - 0x7c
    "00111110", -- 2711 - 0xa97  :   62 - 0x3e
    "10111100", -- 2712 - 0xa98  :  188 - 0xbc
    "01011000", -- 2713 - 0xa99  :   88 - 0x58
    "00111000", -- 2714 - 0xa9a  :   56 - 0x38
    "00010000", -- 2715 - 0xa9b  :   16 - 0x10
    "00110000", -- 2716 - 0xa9c  :   48 - 0x30
    "11111000", -- 2717 - 0xa9d  :  248 - 0xf8
    "11111100", -- 2718 - 0xa9e  :  252 - 0xfc
    "00111110", -- 2719 - 0xa9f  :   62 - 0x3e
    "00000011", -- 2720 - 0xaa0  :    3 - 0x3
    "00001111", -- 2721 - 0xaa1  :   15 - 0xf
    "00011111", -- 2722 - 0xaa2  :   31 - 0x1f
    "00111111", -- 2723 - 0xaa3  :   63 - 0x3f
    "00111011", -- 2724 - 0xaa4  :   59 - 0x3b
    "00111111", -- 2725 - 0xaa5  :   63 - 0x3f
    "01111111", -- 2726 - 0xaa6  :  127 - 0x7f
    "01111111", -- 2727 - 0xaa7  :  127 - 0x7f
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "00000000", -- 2730 - 0xaaa  :    0 - 0x0
    "00000110", -- 2731 - 0xaab  :    6 - 0x6
    "00001110", -- 2732 - 0xaac  :   14 - 0xe
    "00001100", -- 2733 - 0xaad  :   12 - 0xc
    "00000000", -- 2734 - 0xaae  :    0 - 0x0
    "00000000", -- 2735 - 0xaaf  :    0 - 0x0
    "10000000", -- 2736 - 0xab0  :  128 - 0x80
    "11110000", -- 2737 - 0xab1  :  240 - 0xf0
    "11111000", -- 2738 - 0xab2  :  248 - 0xf8
    "11111100", -- 2739 - 0xab3  :  252 - 0xfc
    "11111110", -- 2740 - 0xab4  :  254 - 0xfe
    "11111110", -- 2741 - 0xab5  :  254 - 0xfe
    "11111111", -- 2742 - 0xab6  :  255 - 0xff
    "11111110", -- 2743 - 0xab7  :  254 - 0xfe
    "00000000", -- 2744 - 0xab8  :    0 - 0x0
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "00000000", -- 2747 - 0xabb  :    0 - 0x0
    "00000000", -- 2748 - 0xabc  :    0 - 0x0
    "00000000", -- 2749 - 0xabd  :    0 - 0x0
    "00001111", -- 2750 - 0xabe  :   15 - 0xf
    "00011000", -- 2751 - 0xabf  :   24 - 0x18
    "01111111", -- 2752 - 0xac0  :  127 - 0x7f
    "01111111", -- 2753 - 0xac1  :  127 - 0x7f
    "01111111", -- 2754 - 0xac2  :  127 - 0x7f
    "01111111", -- 2755 - 0xac3  :  127 - 0x7f
    "11111111", -- 2756 - 0xac4  :  255 - 0xff
    "00001111", -- 2757 - 0xac5  :   15 - 0xf
    "00000011", -- 2758 - 0xac6  :    3 - 0x3
    "00000000", -- 2759 - 0xac7  :    0 - 0x0
    "00000000", -- 2760 - 0xac8  :    0 - 0x0
    "00000000", -- 2761 - 0xac9  :    0 - 0x0
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000000", -- 2763 - 0xacb  :    0 - 0x0
    "11111000", -- 2764 - 0xacc  :  248 - 0xf8
    "00111110", -- 2765 - 0xacd  :   62 - 0x3e
    "00111011", -- 2766 - 0xace  :   59 - 0x3b
    "00011000", -- 2767 - 0xacf  :   24 - 0x18
    "11111110", -- 2768 - 0xad0  :  254 - 0xfe
    "11111011", -- 2769 - 0xad1  :  251 - 0xfb
    "11111111", -- 2770 - 0xad2  :  255 - 0xff
    "11111111", -- 2771 - 0xad3  :  255 - 0xff
    "11110110", -- 2772 - 0xad4  :  246 - 0xf6
    "11100000", -- 2773 - 0xad5  :  224 - 0xe0
    "11000000", -- 2774 - 0xad6  :  192 - 0xc0
    "00000000", -- 2775 - 0xad7  :    0 - 0x0
    "00010000", -- 2776 - 0xad8  :   16 - 0x10
    "00010100", -- 2777 - 0xad9  :   20 - 0x14
    "00010000", -- 2778 - 0xada  :   16 - 0x10
    "00010000", -- 2779 - 0xadb  :   16 - 0x10
    "00111000", -- 2780 - 0xadc  :   56 - 0x38
    "01111000", -- 2781 - 0xadd  :  120 - 0x78
    "11111000", -- 2782 - 0xade  :  248 - 0xf8
    "00110000", -- 2783 - 0xadf  :   48 - 0x30
    "00000000", -- 2784 - 0xae0  :    0 - 0x0
    "00000011", -- 2785 - 0xae1  :    3 - 0x3
    "00001111", -- 2786 - 0xae2  :   15 - 0xf
    "00011111", -- 2787 - 0xae3  :   31 - 0x1f
    "00111111", -- 2788 - 0xae4  :   63 - 0x3f
    "00111011", -- 2789 - 0xae5  :   59 - 0x3b
    "00111111", -- 2790 - 0xae6  :   63 - 0x3f
    "01111111", -- 2791 - 0xae7  :  127 - 0x7f
    "00000000", -- 2792 - 0xae8  :    0 - 0x0
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000000", -- 2794 - 0xaea  :    0 - 0x0
    "00000000", -- 2795 - 0xaeb  :    0 - 0x0
    "00000110", -- 2796 - 0xaec  :    6 - 0x6
    "00001110", -- 2797 - 0xaed  :   14 - 0xe
    "00001100", -- 2798 - 0xaee  :   12 - 0xc
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "00000000", -- 2800 - 0xaf0  :    0 - 0x0
    "11000000", -- 2801 - 0xaf1  :  192 - 0xc0
    "11110000", -- 2802 - 0xaf2  :  240 - 0xf0
    "11111000", -- 2803 - 0xaf3  :  248 - 0xf8
    "11111100", -- 2804 - 0xaf4  :  252 - 0xfc
    "11111110", -- 2805 - 0xaf5  :  254 - 0xfe
    "11111110", -- 2806 - 0xaf6  :  254 - 0xfe
    "11111111", -- 2807 - 0xaf7  :  255 - 0xff
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0
    "00000000", -- 2809 - 0xaf9  :    0 - 0x0
    "00000000", -- 2810 - 0xafa  :    0 - 0x0
    "00000000", -- 2811 - 0xafb  :    0 - 0x0
    "00000000", -- 2812 - 0xafc  :    0 - 0x0
    "00000000", -- 2813 - 0xafd  :    0 - 0x0
    "00000000", -- 2814 - 0xafe  :    0 - 0x0
    "00001111", -- 2815 - 0xaff  :   15 - 0xf
    "01111111", -- 2816 - 0xb00  :  127 - 0x7f
    "01111111", -- 2817 - 0xb01  :  127 - 0x7f
    "01111111", -- 2818 - 0xb02  :  127 - 0x7f
    "01111111", -- 2819 - 0xb03  :  127 - 0x7f
    "01111111", -- 2820 - 0xb04  :  127 - 0x7f
    "11111111", -- 2821 - 0xb05  :  255 - 0xff
    "00001111", -- 2822 - 0xb06  :   15 - 0xf
    "00000011", -- 2823 - 0xb07  :    3 - 0x3
    "00000000", -- 2824 - 0xb08  :    0 - 0x0
    "00000000", -- 2825 - 0xb09  :    0 - 0x0
    "00000000", -- 2826 - 0xb0a  :    0 - 0x0
    "00000000", -- 2827 - 0xb0b  :    0 - 0x0
    "00000000", -- 2828 - 0xb0c  :    0 - 0x0
    "11111000", -- 2829 - 0xb0d  :  248 - 0xf8
    "01111110", -- 2830 - 0xb0e  :  126 - 0x7e
    "11110011", -- 2831 - 0xb0f  :  243 - 0xf3
    "11111110", -- 2832 - 0xb10  :  254 - 0xfe
    "11111110", -- 2833 - 0xb11  :  254 - 0xfe
    "11111011", -- 2834 - 0xb12  :  251 - 0xfb
    "11111111", -- 2835 - 0xb13  :  255 - 0xff
    "11111111", -- 2836 - 0xb14  :  255 - 0xff
    "11110110", -- 2837 - 0xb15  :  246 - 0xf6
    "11100000", -- 2838 - 0xb16  :  224 - 0xe0
    "11000000", -- 2839 - 0xb17  :  192 - 0xc0
    "00011000", -- 2840 - 0xb18  :   24 - 0x18
    "00010000", -- 2841 - 0xb19  :   16 - 0x10
    "00010100", -- 2842 - 0xb1a  :   20 - 0x14
    "00010000", -- 2843 - 0xb1b  :   16 - 0x10
    "00010000", -- 2844 - 0xb1c  :   16 - 0x10
    "00111000", -- 2845 - 0xb1d  :   56 - 0x38
    "01111100", -- 2846 - 0xb1e  :  124 - 0x7c
    "11011110", -- 2847 - 0xb1f  :  222 - 0xde
    "00000000", -- 2848 - 0xb20  :    0 - 0x0
    "00000001", -- 2849 - 0xb21  :    1 - 0x1
    "00000001", -- 2850 - 0xb22  :    1 - 0x1
    "00000001", -- 2851 - 0xb23  :    1 - 0x1
    "00000001", -- 2852 - 0xb24  :    1 - 0x1
    "00000000", -- 2853 - 0xb25  :    0 - 0x0
    "00000000", -- 2854 - 0xb26  :    0 - 0x0
    "00001000", -- 2855 - 0xb27  :    8 - 0x8
    "00000000", -- 2856 - 0xb28  :    0 - 0x0
    "00001101", -- 2857 - 0xb29  :   13 - 0xd
    "00011110", -- 2858 - 0xb2a  :   30 - 0x1e
    "00011110", -- 2859 - 0xb2b  :   30 - 0x1e
    "00011110", -- 2860 - 0xb2c  :   30 - 0x1e
    "00011111", -- 2861 - 0xb2d  :   31 - 0x1f
    "00001111", -- 2862 - 0xb2e  :   15 - 0xf
    "00000111", -- 2863 - 0xb2f  :    7 - 0x7
    "01111000", -- 2864 - 0xb30  :  120 - 0x78
    "11110000", -- 2865 - 0xb31  :  240 - 0xf0
    "11111000", -- 2866 - 0xb32  :  248 - 0xf8
    "11100100", -- 2867 - 0xb33  :  228 - 0xe4
    "11000000", -- 2868 - 0xb34  :  192 - 0xc0
    "11001010", -- 2869 - 0xb35  :  202 - 0xca
    "11001010", -- 2870 - 0xb36  :  202 - 0xca
    "11000000", -- 2871 - 0xb37  :  192 - 0xc0
    "01111000", -- 2872 - 0xb38  :  120 - 0x78
    "11110000", -- 2873 - 0xb39  :  240 - 0xf0
    "00000000", -- 2874 - 0xb3a  :    0 - 0x0
    "00011010", -- 2875 - 0xb3b  :   26 - 0x1a
    "00111111", -- 2876 - 0xb3c  :   63 - 0x3f
    "00110101", -- 2877 - 0xb3d  :   53 - 0x35
    "00110101", -- 2878 - 0xb3e  :   53 - 0x35
    "00111111", -- 2879 - 0xb3f  :   63 - 0x3f
    "00001111", -- 2880 - 0xb40  :   15 - 0xf
    "00011111", -- 2881 - 0xb41  :   31 - 0x1f
    "10011111", -- 2882 - 0xb42  :  159 - 0x9f
    "11111111", -- 2883 - 0xb43  :  255 - 0xff
    "11111111", -- 2884 - 0xb44  :  255 - 0xff
    "01111111", -- 2885 - 0xb45  :  127 - 0x7f
    "01110100", -- 2886 - 0xb46  :  116 - 0x74
    "00100000", -- 2887 - 0xb47  :   32 - 0x20
    "00000000", -- 2888 - 0xb48  :    0 - 0x0
    "00000000", -- 2889 - 0xb49  :    0 - 0x0
    "10000000", -- 2890 - 0xb4a  :  128 - 0x80
    "11100000", -- 2891 - 0xb4b  :  224 - 0xe0
    "11100000", -- 2892 - 0xb4c  :  224 - 0xe0
    "01110000", -- 2893 - 0xb4d  :  112 - 0x70
    "01110011", -- 2894 - 0xb4e  :  115 - 0x73
    "00100001", -- 2895 - 0xb4f  :   33 - 0x21
    "11100100", -- 2896 - 0xb50  :  228 - 0xe4
    "11111111", -- 2897 - 0xb51  :  255 - 0xff
    "11111110", -- 2898 - 0xb52  :  254 - 0xfe
    "11111100", -- 2899 - 0xb53  :  252 - 0xfc
    "10011100", -- 2900 - 0xb54  :  156 - 0x9c
    "00011110", -- 2901 - 0xb55  :   30 - 0x1e
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "00011010", -- 2904 - 0xb58  :   26 - 0x1a
    "00000111", -- 2905 - 0xb59  :    7 - 0x7
    "00001100", -- 2906 - 0xb5a  :   12 - 0xc
    "00011000", -- 2907 - 0xb5b  :   24 - 0x18
    "01111000", -- 2908 - 0xb5c  :  120 - 0x78
    "11111110", -- 2909 - 0xb5d  :  254 - 0xfe
    "11111100", -- 2910 - 0xb5e  :  252 - 0xfc
    "11110000", -- 2911 - 0xb5f  :  240 - 0xf0
    "00000000", -- 2912 - 0xb60  :    0 - 0x0
    "00000001", -- 2913 - 0xb61  :    1 - 0x1
    "00000011", -- 2914 - 0xb62  :    3 - 0x3
    "00000011", -- 2915 - 0xb63  :    3 - 0x3
    "00000111", -- 2916 - 0xb64  :    7 - 0x7
    "00000011", -- 2917 - 0xb65  :    3 - 0x3
    "00000001", -- 2918 - 0xb66  :    1 - 0x1
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "00000000", -- 2920 - 0xb68  :    0 - 0x0
    "00000001", -- 2921 - 0xb69  :    1 - 0x1
    "00000010", -- 2922 - 0xb6a  :    2 - 0x2
    "00000000", -- 2923 - 0xb6b  :    0 - 0x0
    "00111000", -- 2924 - 0xb6c  :   56 - 0x38
    "01111100", -- 2925 - 0xb6d  :  124 - 0x7c
    "01111110", -- 2926 - 0xb6e  :  126 - 0x7e
    "00111111", -- 2927 - 0xb6f  :   63 - 0x3f
    "00000000", -- 2928 - 0xb70  :    0 - 0x0
    "01011111", -- 2929 - 0xb71  :   95 - 0x5f
    "01111111", -- 2930 - 0xb72  :  127 - 0x7f
    "01111111", -- 2931 - 0xb73  :  127 - 0x7f
    "00111111", -- 2932 - 0xb74  :   63 - 0x3f
    "00111111", -- 2933 - 0xb75  :   63 - 0x3f
    "00010100", -- 2934 - 0xb76  :   20 - 0x14
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "00111111", -- 2936 - 0xb78  :   63 - 0x3f
    "01000000", -- 2937 - 0xb79  :   64 - 0x40
    "01100000", -- 2938 - 0xb7a  :   96 - 0x60
    "01100000", -- 2939 - 0xb7b  :   96 - 0x60
    "00100000", -- 2940 - 0xb7c  :   32 - 0x20
    "00110000", -- 2941 - 0xb7d  :   48 - 0x30
    "00010011", -- 2942 - 0xb7e  :   19 - 0x13
    "00000001", -- 2943 - 0xb7f  :    1 - 0x1
    "11000000", -- 2944 - 0xb80  :  192 - 0xc0
    "11100000", -- 2945 - 0xb81  :  224 - 0xe0
    "11110000", -- 2946 - 0xb82  :  240 - 0xf0
    "00110000", -- 2947 - 0xb83  :   48 - 0x30
    "00111000", -- 2948 - 0xb84  :   56 - 0x38
    "00111100", -- 2949 - 0xb85  :   60 - 0x3c
    "00111100", -- 2950 - 0xb86  :   60 - 0x3c
    "11111100", -- 2951 - 0xb87  :  252 - 0xfc
    "11000000", -- 2952 - 0xb88  :  192 - 0xc0
    "11100000", -- 2953 - 0xb89  :  224 - 0xe0
    "00110000", -- 2954 - 0xb8a  :   48 - 0x30
    "11010000", -- 2955 - 0xb8b  :  208 - 0xd0
    "11010000", -- 2956 - 0xb8c  :  208 - 0xd0
    "11010000", -- 2957 - 0xb8d  :  208 - 0xd0
    "11010000", -- 2958 - 0xb8e  :  208 - 0xd0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00000111", -- 2960 - 0xb90  :    7 - 0x7
    "00001111", -- 2961 - 0xb91  :   15 - 0xf
    "00011111", -- 2962 - 0xb92  :   31 - 0x1f
    "00100010", -- 2963 - 0xb93  :   34 - 0x22
    "00100000", -- 2964 - 0xb94  :   32 - 0x20
    "00100101", -- 2965 - 0xb95  :   37 - 0x25
    "00100101", -- 2966 - 0xb96  :   37 - 0x25
    "00011111", -- 2967 - 0xb97  :   31 - 0x1f
    "00000111", -- 2968 - 0xb98  :    7 - 0x7
    "00001111", -- 2969 - 0xb99  :   15 - 0xf
    "00000010", -- 2970 - 0xb9a  :    2 - 0x2
    "00011101", -- 2971 - 0xb9b  :   29 - 0x1d
    "00011111", -- 2972 - 0xb9c  :   31 - 0x1f
    "00011010", -- 2973 - 0xb9d  :   26 - 0x1a
    "00011010", -- 2974 - 0xb9e  :   26 - 0x1a
    "00000010", -- 2975 - 0xb9f  :    2 - 0x2
    "11111110", -- 2976 - 0xba0  :  254 - 0xfe
    "11111110", -- 2977 - 0xba1  :  254 - 0xfe
    "01111110", -- 2978 - 0xba2  :  126 - 0x7e
    "00111010", -- 2979 - 0xba3  :   58 - 0x3a
    "00000010", -- 2980 - 0xba4  :    2 - 0x2
    "00000001", -- 2981 - 0xba5  :    1 - 0x1
    "01000001", -- 2982 - 0xba6  :   65 - 0x41
    "01000001", -- 2983 - 0xba7  :   65 - 0x41
    "00111000", -- 2984 - 0xba8  :   56 - 0x38
    "01111100", -- 2985 - 0xba9  :  124 - 0x7c
    "11111100", -- 2986 - 0xbaa  :  252 - 0xfc
    "11111100", -- 2987 - 0xbab  :  252 - 0xfc
    "11111100", -- 2988 - 0xbac  :  252 - 0xfc
    "11111110", -- 2989 - 0xbad  :  254 - 0xfe
    "10111110", -- 2990 - 0xbae  :  190 - 0xbe
    "10111110", -- 2991 - 0xbaf  :  190 - 0xbe
    "00011111", -- 2992 - 0xbb0  :   31 - 0x1f
    "00111111", -- 2993 - 0xbb1  :   63 - 0x3f
    "01111110", -- 2994 - 0xbb2  :  126 - 0x7e
    "01011100", -- 2995 - 0xbb3  :   92 - 0x5c
    "01000000", -- 2996 - 0xbb4  :   64 - 0x40
    "10000000", -- 2997 - 0xbb5  :  128 - 0x80
    "10000010", -- 2998 - 0xbb6  :  130 - 0x82
    "10000010", -- 2999 - 0xbb7  :  130 - 0x82
    "00011100", -- 3000 - 0xbb8  :   28 - 0x1c
    "00111110", -- 3001 - 0xbb9  :   62 - 0x3e
    "00111111", -- 3002 - 0xbba  :   63 - 0x3f
    "00111111", -- 3003 - 0xbbb  :   63 - 0x3f
    "00111111", -- 3004 - 0xbbc  :   63 - 0x3f
    "01111111", -- 3005 - 0xbbd  :  127 - 0x7f
    "01111101", -- 3006 - 0xbbe  :  125 - 0x7d
    "01111101", -- 3007 - 0xbbf  :  125 - 0x7d
    "10000010", -- 3008 - 0xbc0  :  130 - 0x82
    "10000000", -- 3009 - 0xbc1  :  128 - 0x80
    "10100000", -- 3010 - 0xbc2  :  160 - 0xa0
    "01000100", -- 3011 - 0xbc3  :   68 - 0x44
    "01000011", -- 3012 - 0xbc4  :   67 - 0x43
    "01000000", -- 3013 - 0xbc5  :   64 - 0x40
    "00100001", -- 3014 - 0xbc6  :   33 - 0x21
    "00011110", -- 3015 - 0xbc7  :   30 - 0x1e
    "01111101", -- 3016 - 0xbc8  :  125 - 0x7d
    "01111111", -- 3017 - 0xbc9  :  127 - 0x7f
    "01011111", -- 3018 - 0xbca  :   95 - 0x5f
    "00111011", -- 3019 - 0xbcb  :   59 - 0x3b
    "00111100", -- 3020 - 0xbcc  :   60 - 0x3c
    "00111111", -- 3021 - 0xbcd  :   63 - 0x3f
    "00011110", -- 3022 - 0xbce  :   30 - 0x1e
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00011100", -- 3024 - 0xbd0  :   28 - 0x1c
    "00111111", -- 3025 - 0xbd1  :   63 - 0x3f
    "00111110", -- 3026 - 0xbd2  :   62 - 0x3e
    "00111100", -- 3027 - 0xbd3  :   60 - 0x3c
    "01000000", -- 3028 - 0xbd4  :   64 - 0x40
    "10000000", -- 3029 - 0xbd5  :  128 - 0x80
    "10000010", -- 3030 - 0xbd6  :  130 - 0x82
    "10000010", -- 3031 - 0xbd7  :  130 - 0x82
    "00011100", -- 3032 - 0xbd8  :   28 - 0x1c
    "00111110", -- 3033 - 0xbd9  :   62 - 0x3e
    "00111111", -- 3034 - 0xbda  :   63 - 0x3f
    "00011111", -- 3035 - 0xbdb  :   31 - 0x1f
    "00111111", -- 3036 - 0xbdc  :   63 - 0x3f
    "01111111", -- 3037 - 0xbdd  :  127 - 0x7f
    "01111101", -- 3038 - 0xbde  :  125 - 0x7d
    "01111101", -- 3039 - 0xbdf  :  125 - 0x7d
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0
    "00000000", -- 3041 - 0xbe1  :    0 - 0x0
    "10000000", -- 3042 - 0xbe2  :  128 - 0x80
    "10000000", -- 3043 - 0xbe3  :  128 - 0x80
    "10010010", -- 3044 - 0xbe4  :  146 - 0x92
    "10011101", -- 3045 - 0xbe5  :  157 - 0x9d
    "11000111", -- 3046 - 0xbe6  :  199 - 0xc7
    "11101111", -- 3047 - 0xbe7  :  239 - 0xef
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0
    "00000000", -- 3049 - 0xbe9  :    0 - 0x0
    "00000000", -- 3050 - 0xbea  :    0 - 0x0
    "01100000", -- 3051 - 0xbeb  :   96 - 0x60
    "01100010", -- 3052 - 0xbec  :   98 - 0x62
    "01100101", -- 3053 - 0xbed  :  101 - 0x65
    "00111111", -- 3054 - 0xbee  :   63 - 0x3f
    "00011111", -- 3055 - 0xbef  :   31 - 0x1f
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0
    "00100011", -- 3057 - 0xbf1  :   35 - 0x23
    "00110011", -- 3058 - 0xbf2  :   51 - 0x33
    "00111111", -- 3059 - 0xbf3  :   63 - 0x3f
    "00111111", -- 3060 - 0xbf4  :   63 - 0x3f
    "01111111", -- 3061 - 0xbf5  :  127 - 0x7f
    "01111111", -- 3062 - 0xbf6  :  127 - 0x7f
    "01111111", -- 3063 - 0xbf7  :  127 - 0x7f
    "01110000", -- 3064 - 0xbf8  :  112 - 0x70
    "00111100", -- 3065 - 0xbf9  :   60 - 0x3c
    "00111100", -- 3066 - 0xbfa  :   60 - 0x3c
    "00011000", -- 3067 - 0xbfb  :   24 - 0x18
    "00000000", -- 3068 - 0xbfc  :    0 - 0x0
    "00000000", -- 3069 - 0xbfd  :    0 - 0x0
    "00000010", -- 3070 - 0xbfe  :    2 - 0x2
    "00000111", -- 3071 - 0xbff  :    7 - 0x7
    "11111110", -- 3072 - 0xc00  :  254 - 0xfe
    "11111000", -- 3073 - 0xc01  :  248 - 0xf8
    "10100000", -- 3074 - 0xc02  :  160 - 0xa0
    "00000000", -- 3075 - 0xc03  :    0 - 0x0
    "00000000", -- 3076 - 0xc04  :    0 - 0x0
    "00000000", -- 3077 - 0xc05  :    0 - 0x0
    "10000000", -- 3078 - 0xc06  :  128 - 0x80
    "10000000", -- 3079 - 0xc07  :  128 - 0x80
    "11001111", -- 3080 - 0xc08  :  207 - 0xcf
    "01111010", -- 3081 - 0xc09  :  122 - 0x7a
    "01011010", -- 3082 - 0xc0a  :   90 - 0x5a
    "00010000", -- 3083 - 0xc0b  :   16 - 0x10
    "00000000", -- 3084 - 0xc0c  :    0 - 0x0
    "00000000", -- 3085 - 0xc0d  :    0 - 0x0
    "11000000", -- 3086 - 0xc0e  :  192 - 0xc0
    "10000000", -- 3087 - 0xc0f  :  128 - 0x80
    "01111110", -- 3088 - 0xc10  :  126 - 0x7e
    "01111111", -- 3089 - 0xc11  :  127 - 0x7f
    "01111101", -- 3090 - 0xc12  :  125 - 0x7d
    "00111111", -- 3091 - 0xc13  :   63 - 0x3f
    "00011110", -- 3092 - 0xc14  :   30 - 0x1e
    "10001111", -- 3093 - 0xc15  :  143 - 0x8f
    "10001111", -- 3094 - 0xc16  :  143 - 0x8f
    "00011001", -- 3095 - 0xc17  :   25 - 0x19
    "10000101", -- 3096 - 0xc18  :  133 - 0x85
    "10000100", -- 3097 - 0xc19  :  132 - 0x84
    "10000110", -- 3098 - 0xc1a  :  134 - 0x86
    "11000110", -- 3099 - 0xc1b  :  198 - 0xc6
    "11100111", -- 3100 - 0xc1c  :  231 - 0xe7
    "01110011", -- 3101 - 0xc1d  :  115 - 0x73
    "01110011", -- 3102 - 0xc1e  :  115 - 0x73
    "11100001", -- 3103 - 0xc1f  :  225 - 0xe1
    "11100000", -- 3104 - 0xc20  :  224 - 0xe0
    "00001110", -- 3105 - 0xc21  :   14 - 0xe
    "01110011", -- 3106 - 0xc22  :  115 - 0x73
    "11110011", -- 3107 - 0xc23  :  243 - 0xf3
    "11111001", -- 3108 - 0xc24  :  249 - 0xf9
    "11111001", -- 3109 - 0xc25  :  249 - 0xf9
    "11111000", -- 3110 - 0xc26  :  248 - 0xf8
    "01110000", -- 3111 - 0xc27  :  112 - 0x70
    "10000000", -- 3112 - 0xc28  :  128 - 0x80
    "01001110", -- 3113 - 0xc29  :   78 - 0x4e
    "01110111", -- 3114 - 0xc2a  :  119 - 0x77
    "11110011", -- 3115 - 0xc2b  :  243 - 0xf3
    "11111011", -- 3116 - 0xc2c  :  251 - 0xfb
    "11111001", -- 3117 - 0xc2d  :  249 - 0xf9
    "11111010", -- 3118 - 0xc2e  :  250 - 0xfa
    "01111000", -- 3119 - 0xc2f  :  120 - 0x78
    "00001110", -- 3120 - 0xc30  :   14 - 0xe
    "01100110", -- 3121 - 0xc31  :  102 - 0x66
    "11100010", -- 3122 - 0xc32  :  226 - 0xe2
    "11110110", -- 3123 - 0xc33  :  246 - 0xf6
    "11111111", -- 3124 - 0xc34  :  255 - 0xff
    "11111111", -- 3125 - 0xc35  :  255 - 0xff
    "00011111", -- 3126 - 0xc36  :   31 - 0x1f
    "10011000", -- 3127 - 0xc37  :  152 - 0x98
    "00010001", -- 3128 - 0xc38  :   17 - 0x11
    "00111001", -- 3129 - 0xc39  :   57 - 0x39
    "01111101", -- 3130 - 0xc3a  :  125 - 0x7d
    "00111001", -- 3131 - 0xc3b  :   57 - 0x39
    "00000000", -- 3132 - 0xc3c  :    0 - 0x0
    "00000000", -- 3133 - 0xc3d  :    0 - 0x0
    "11100000", -- 3134 - 0xc3e  :  224 - 0xe0
    "11100111", -- 3135 - 0xc3f  :  231 - 0xe7
    "00000000", -- 3136 - 0xc40  :    0 - 0x0
    "00000000", -- 3137 - 0xc41  :    0 - 0x0
    "00000000", -- 3138 - 0xc42  :    0 - 0x0
    "00000100", -- 3139 - 0xc43  :    4 - 0x4
    "00001111", -- 3140 - 0xc44  :   15 - 0xf
    "00001111", -- 3141 - 0xc45  :   15 - 0xf
    "00011111", -- 3142 - 0xc46  :   31 - 0x1f
    "00000111", -- 3143 - 0xc47  :    7 - 0x7
    "00000000", -- 3144 - 0xc48  :    0 - 0x0
    "00000000", -- 3145 - 0xc49  :    0 - 0x0
    "00000111", -- 3146 - 0xc4a  :    7 - 0x7
    "00000111", -- 3147 - 0xc4b  :    7 - 0x7
    "00010110", -- 3148 - 0xc4c  :   22 - 0x16
    "00010000", -- 3149 - 0xc4d  :   16 - 0x10
    "00000000", -- 3150 - 0xc4e  :    0 - 0x0
    "00111000", -- 3151 - 0xc4f  :   56 - 0x38
    "11110011", -- 3152 - 0xc50  :  243 - 0xf3
    "11100111", -- 3153 - 0xc51  :  231 - 0xe7
    "11101110", -- 3154 - 0xc52  :  238 - 0xee
    "11101100", -- 3155 - 0xc53  :  236 - 0xec
    "11001101", -- 3156 - 0xc54  :  205 - 0xcd
    "11001111", -- 3157 - 0xc55  :  207 - 0xcf
    "11001111", -- 3158 - 0xc56  :  207 - 0xcf
    "11011111", -- 3159 - 0xc57  :  223 - 0xdf
    "11001111", -- 3160 - 0xc58  :  207 - 0xcf
    "00011111", -- 3161 - 0xc59  :   31 - 0x1f
    "00010111", -- 3162 - 0xc5a  :   23 - 0x17
    "00010000", -- 3163 - 0xc5b  :   16 - 0x10
    "00110011", -- 3164 - 0xc5c  :   51 - 0x33
    "00110000", -- 3165 - 0xc5d  :   48 - 0x30
    "00110000", -- 3166 - 0xc5e  :   48 - 0x30
    "00100000", -- 3167 - 0xc5f  :   32 - 0x20
    "00100111", -- 3168 - 0xc60  :   39 - 0x27
    "00111111", -- 3169 - 0xc61  :   63 - 0x3f
    "00111111", -- 3170 - 0xc62  :   63 - 0x3f
    "01111000", -- 3171 - 0xc63  :  120 - 0x78
    "00111100", -- 3172 - 0xc64  :   60 - 0x3c
    "00011111", -- 3173 - 0xc65  :   31 - 0x1f
    "00011111", -- 3174 - 0xc66  :   31 - 0x1f
    "01110011", -- 3175 - 0xc67  :  115 - 0x73
    "00111000", -- 3176 - 0xc68  :   56 - 0x38
    "00110000", -- 3177 - 0xc69  :   48 - 0x30
    "01000000", -- 3178 - 0xc6a  :   64 - 0x40
    "11000111", -- 3179 - 0xc6b  :  199 - 0xc7
    "00000111", -- 3180 - 0xc6c  :    7 - 0x7
    "01100110", -- 3181 - 0xc6d  :  102 - 0x66
    "11100000", -- 3182 - 0xc6e  :  224 - 0xe0
    "01101100", -- 3183 - 0xc6f  :  108 - 0x6c
    "10011111", -- 3184 - 0xc70  :  159 - 0x9f
    "00111110", -- 3185 - 0xc71  :   62 - 0x3e
    "01111100", -- 3186 - 0xc72  :  124 - 0x7c
    "11111100", -- 3187 - 0xc73  :  252 - 0xfc
    "11111000", -- 3188 - 0xc74  :  248 - 0xf8
    "11111000", -- 3189 - 0xc75  :  248 - 0xf8
    "11000000", -- 3190 - 0xc76  :  192 - 0xc0
    "01000000", -- 3191 - 0xc77  :   64 - 0x40
    "01100000", -- 3192 - 0xc78  :   96 - 0x60
    "11000000", -- 3193 - 0xc79  :  192 - 0xc0
    "10000000", -- 3194 - 0xc7a  :  128 - 0x80
    "00000100", -- 3195 - 0xc7b  :    4 - 0x4
    "10011110", -- 3196 - 0xc7c  :  158 - 0x9e
    "11111111", -- 3197 - 0xc7d  :  255 - 0xff
    "11110000", -- 3198 - 0xc7e  :  240 - 0xf0
    "11111000", -- 3199 - 0xc7f  :  248 - 0xf8
    "01111111", -- 3200 - 0xc80  :  127 - 0x7f
    "01111110", -- 3201 - 0xc81  :  126 - 0x7e
    "01111000", -- 3202 - 0xc82  :  120 - 0x78
    "00000001", -- 3203 - 0xc83  :    1 - 0x1
    "00000111", -- 3204 - 0xc84  :    7 - 0x7
    "00011111", -- 3205 - 0xc85  :   31 - 0x1f
    "00111100", -- 3206 - 0xc86  :   60 - 0x3c
    "01111100", -- 3207 - 0xc87  :  124 - 0x7c
    "00100100", -- 3208 - 0xc88  :   36 - 0x24
    "00000001", -- 3209 - 0xc89  :    1 - 0x1
    "00000111", -- 3210 - 0xc8a  :    7 - 0x7
    "11111110", -- 3211 - 0xc8b  :  254 - 0xfe
    "11111111", -- 3212 - 0xc8c  :  255 - 0xff
    "01111111", -- 3213 - 0xc8d  :  127 - 0x7f
    "00111111", -- 3214 - 0xc8e  :   63 - 0x3f
    "01111111", -- 3215 - 0xc8f  :  127 - 0x7f
    "11111100", -- 3216 - 0xc90  :  252 - 0xfc
    "11111000", -- 3217 - 0xc91  :  248 - 0xf8
    "10100000", -- 3218 - 0xc92  :  160 - 0xa0
    "11111110", -- 3219 - 0xc93  :  254 - 0xfe
    "11111100", -- 3220 - 0xc94  :  252 - 0xfc
    "11110000", -- 3221 - 0xc95  :  240 - 0xf0
    "10000000", -- 3222 - 0xc96  :  128 - 0x80
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "11001111", -- 3224 - 0xc98  :  207 - 0xcf
    "01111010", -- 3225 - 0xc99  :  122 - 0x7a
    "00001010", -- 3226 - 0xc9a  :   10 - 0xa
    "11111110", -- 3227 - 0xc9b  :  254 - 0xfe
    "11111100", -- 3228 - 0xc9c  :  252 - 0xfc
    "00000000", -- 3229 - 0xc9d  :    0 - 0x0
    "00000000", -- 3230 - 0xc9e  :    0 - 0x0
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "01111110", -- 3232 - 0xca0  :  126 - 0x7e
    "01111111", -- 3233 - 0xca1  :  127 - 0x7f
    "01111111", -- 3234 - 0xca2  :  127 - 0x7f
    "00111111", -- 3235 - 0xca3  :   63 - 0x3f
    "00011111", -- 3236 - 0xca4  :   31 - 0x1f
    "10001111", -- 3237 - 0xca5  :  143 - 0x8f
    "10001111", -- 3238 - 0xca6  :  143 - 0x8f
    "00011000", -- 3239 - 0xca7  :   24 - 0x18
    "10000101", -- 3240 - 0xca8  :  133 - 0x85
    "10000110", -- 3241 - 0xca9  :  134 - 0x86
    "10000011", -- 3242 - 0xcaa  :  131 - 0x83
    "11000011", -- 3243 - 0xcab  :  195 - 0xc3
    "11100001", -- 3244 - 0xcac  :  225 - 0xe1
    "01110000", -- 3245 - 0xcad  :  112 - 0x70
    "01110000", -- 3246 - 0xcae  :  112 - 0x70
    "11100000", -- 3247 - 0xcaf  :  224 - 0xe0
    "10011111", -- 3248 - 0xcb0  :  159 - 0x9f
    "00111110", -- 3249 - 0xcb1  :   62 - 0x3e
    "01111100", -- 3250 - 0xcb2  :  124 - 0x7c
    "11111000", -- 3251 - 0xcb3  :  248 - 0xf8
    "11111000", -- 3252 - 0xcb4  :  248 - 0xf8
    "00111100", -- 3253 - 0xcb5  :   60 - 0x3c
    "00011000", -- 3254 - 0xcb6  :   24 - 0x18
    "11111000", -- 3255 - 0xcb7  :  248 - 0xf8
    "01100000", -- 3256 - 0xcb8  :   96 - 0x60
    "11000000", -- 3257 - 0xcb9  :  192 - 0xc0
    "10000000", -- 3258 - 0xcba  :  128 - 0x80
    "00000000", -- 3259 - 0xcbb  :    0 - 0x0
    "10011000", -- 3260 - 0xcbc  :  152 - 0x98
    "11111100", -- 3261 - 0xcbd  :  252 - 0xfc
    "11111110", -- 3262 - 0xcbe  :  254 - 0xfe
    "11111111", -- 3263 - 0xcbf  :  255 - 0xff
    "01111111", -- 3264 - 0xcc0  :  127 - 0x7f
    "01111111", -- 3265 - 0xcc1  :  127 - 0x7f
    "01111000", -- 3266 - 0xcc2  :  120 - 0x78
    "00000001", -- 3267 - 0xcc3  :    1 - 0x1
    "00000111", -- 3268 - 0xcc4  :    7 - 0x7
    "00010011", -- 3269 - 0xcc5  :   19 - 0x13
    "11110001", -- 3270 - 0xcc6  :  241 - 0xf1
    "00000011", -- 3271 - 0xcc7  :    3 - 0x3
    "00100100", -- 3272 - 0xcc8  :   36 - 0x24
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000111", -- 3274 - 0xcca  :    7 - 0x7
    "11111110", -- 3275 - 0xccb  :  254 - 0xfe
    "11111111", -- 3276 - 0xccc  :  255 - 0xff
    "01111111", -- 3277 - 0xccd  :  127 - 0x7f
    "11111111", -- 3278 - 0xcce  :  255 - 0xff
    "00000011", -- 3279 - 0xccf  :    3 - 0x3
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00011100", -- 3282 - 0xcd2  :   28 - 0x1c
    "00011101", -- 3283 - 0xcd3  :   29 - 0x1d
    "00011011", -- 3284 - 0xcd4  :   27 - 0x1b
    "11000011", -- 3285 - 0xcd5  :  195 - 0xc3
    "11100011", -- 3286 - 0xcd6  :  227 - 0xe3
    "11100001", -- 3287 - 0xcd7  :  225 - 0xe1
    "00000011", -- 3288 - 0xcd8  :    3 - 0x3
    "00001111", -- 3289 - 0xcd9  :   15 - 0xf
    "00100011", -- 3290 - 0xcda  :   35 - 0x23
    "01100010", -- 3291 - 0xcdb  :   98 - 0x62
    "01100100", -- 3292 - 0xcdc  :  100 - 0x64
    "00111100", -- 3293 - 0xcdd  :   60 - 0x3c
    "00011100", -- 3294 - 0xcde  :   28 - 0x1c
    "00011110", -- 3295 - 0xcdf  :   30 - 0x1e
    "11100000", -- 3296 - 0xce0  :  224 - 0xe0
    "11001101", -- 3297 - 0xce1  :  205 - 0xcd
    "00011101", -- 3298 - 0xce2  :   29 - 0x1d
    "01001111", -- 3299 - 0xce3  :   79 - 0x4f
    "11101110", -- 3300 - 0xce4  :  238 - 0xee
    "11111111", -- 3301 - 0xce5  :  255 - 0xff
    "00111111", -- 3302 - 0xce6  :   63 - 0x3f
    "00111111", -- 3303 - 0xce7  :   63 - 0x3f
    "00011111", -- 3304 - 0xce8  :   31 - 0x1f
    "00111101", -- 3305 - 0xce9  :   61 - 0x3d
    "01101101", -- 3306 - 0xcea  :  109 - 0x6d
    "01001111", -- 3307 - 0xceb  :   79 - 0x4f
    "11101110", -- 3308 - 0xcec  :  238 - 0xee
    "11110011", -- 3309 - 0xced  :  243 - 0xf3
    "00100000", -- 3310 - 0xcee  :   32 - 0x20
    "00000011", -- 3311 - 0xcef  :    3 - 0x3
    "00111111", -- 3312 - 0xcf0  :   63 - 0x3f
    "00111111", -- 3313 - 0xcf1  :   63 - 0x3f
    "00000000", -- 3314 - 0xcf2  :    0 - 0x0
    "00000000", -- 3315 - 0xcf3  :    0 - 0x0
    "01110000", -- 3316 - 0xcf4  :  112 - 0x70
    "10111000", -- 3317 - 0xcf5  :  184 - 0xb8
    "11111100", -- 3318 - 0xcf6  :  252 - 0xfc
    "11111100", -- 3319 - 0xcf7  :  252 - 0xfc
    "00000111", -- 3320 - 0xcf8  :    7 - 0x7
    "00000111", -- 3321 - 0xcf9  :    7 - 0x7
    "00011111", -- 3322 - 0xcfa  :   31 - 0x1f
    "00111111", -- 3323 - 0xcfb  :   63 - 0x3f
    "00001111", -- 3324 - 0xcfc  :   15 - 0xf
    "01000111", -- 3325 - 0xcfd  :   71 - 0x47
    "00000011", -- 3326 - 0xcfe  :    3 - 0x3
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00000111", -- 3328 - 0xd00  :    7 - 0x7
    "00001111", -- 3329 - 0xd01  :   15 - 0xf
    "00011111", -- 3330 - 0xd02  :   31 - 0x1f
    "00111111", -- 3331 - 0xd03  :   63 - 0x3f
    "00111110", -- 3332 - 0xd04  :   62 - 0x3e
    "01111100", -- 3333 - 0xd05  :  124 - 0x7c
    "01111000", -- 3334 - 0xd06  :  120 - 0x78
    "01111000", -- 3335 - 0xd07  :  120 - 0x78
    "00000000", -- 3336 - 0xd08  :    0 - 0x0
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "00000011", -- 3338 - 0xd0a  :    3 - 0x3
    "00000111", -- 3339 - 0xd0b  :    7 - 0x7
    "00001111", -- 3340 - 0xd0c  :   15 - 0xf
    "00001111", -- 3341 - 0xd0d  :   15 - 0xf
    "00011111", -- 3342 - 0xd0e  :   31 - 0x1f
    "00011111", -- 3343 - 0xd0f  :   31 - 0x1f
    "00111111", -- 3344 - 0xd10  :   63 - 0x3f
    "01011100", -- 3345 - 0xd11  :   92 - 0x5c
    "00111001", -- 3346 - 0xd12  :   57 - 0x39
    "00111011", -- 3347 - 0xd13  :   59 - 0x3b
    "10111111", -- 3348 - 0xd14  :  191 - 0xbf
    "11111111", -- 3349 - 0xd15  :  255 - 0xff
    "11111110", -- 3350 - 0xd16  :  254 - 0xfe
    "11111110", -- 3351 - 0xd17  :  254 - 0xfe
    "00000000", -- 3352 - 0xd18  :    0 - 0x0
    "00100011", -- 3353 - 0xd19  :   35 - 0x23
    "01010111", -- 3354 - 0xd1a  :   87 - 0x57
    "01001111", -- 3355 - 0xd1b  :   79 - 0x4f
    "01010111", -- 3356 - 0xd1c  :   87 - 0x57
    "00101111", -- 3357 - 0xd1d  :   47 - 0x2f
    "11011111", -- 3358 - 0xd1e  :  223 - 0xdf
    "00100001", -- 3359 - 0xd1f  :   33 - 0x21
    "11000000", -- 3360 - 0xd20  :  192 - 0xc0
    "11000000", -- 3361 - 0xd21  :  192 - 0xc0
    "10000000", -- 3362 - 0xd22  :  128 - 0x80
    "10000000", -- 3363 - 0xd23  :  128 - 0x80
    "10000000", -- 3364 - 0xd24  :  128 - 0x80
    "10000000", -- 3365 - 0xd25  :  128 - 0x80
    "00000000", -- 3366 - 0xd26  :    0 - 0x0
    "00000000", -- 3367 - 0xd27  :    0 - 0x0
    "00000000", -- 3368 - 0xd28  :    0 - 0x0
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "00000000", -- 3370 - 0xd2a  :    0 - 0x0
    "00000000", -- 3371 - 0xd2b  :    0 - 0x0
    "10000000", -- 3372 - 0xd2c  :  128 - 0x80
    "10000000", -- 3373 - 0xd2d  :  128 - 0x80
    "00000000", -- 3374 - 0xd2e  :    0 - 0x0
    "00000000", -- 3375 - 0xd2f  :    0 - 0x0
    "11111110", -- 3376 - 0xd30  :  254 - 0xfe
    "11111100", -- 3377 - 0xd31  :  252 - 0xfc
    "01100001", -- 3378 - 0xd32  :   97 - 0x61
    "00001111", -- 3379 - 0xd33  :   15 - 0xf
    "01111111", -- 3380 - 0xd34  :  127 - 0x7f
    "00111111", -- 3381 - 0xd35  :   63 - 0x3f
    "00011111", -- 3382 - 0xd36  :   31 - 0x1f
    "00011110", -- 3383 - 0xd37  :   30 - 0x1e
    "00100011", -- 3384 - 0xd38  :   35 - 0x23
    "00001111", -- 3385 - 0xd39  :   15 - 0xf
    "00011110", -- 3386 - 0xd3a  :   30 - 0x1e
    "11110000", -- 3387 - 0xd3b  :  240 - 0xf0
    "00011100", -- 3388 - 0xd3c  :   28 - 0x1c
    "00111111", -- 3389 - 0xd3d  :   63 - 0x3f
    "00011111", -- 3390 - 0xd3e  :   31 - 0x1f
    "00011110", -- 3391 - 0xd3f  :   30 - 0x1e
    "11110000", -- 3392 - 0xd40  :  240 - 0xf0
    "01111000", -- 3393 - 0xd41  :  120 - 0x78
    "11100100", -- 3394 - 0xd42  :  228 - 0xe4
    "11001000", -- 3395 - 0xd43  :  200 - 0xc8
    "11001100", -- 3396 - 0xd44  :  204 - 0xcc
    "10111110", -- 3397 - 0xd45  :  190 - 0xbe
    "10111110", -- 3398 - 0xd46  :  190 - 0xbe
    "00111110", -- 3399 - 0xd47  :   62 - 0x3e
    "00000000", -- 3400 - 0xd48  :    0 - 0x0
    "10000000", -- 3401 - 0xd49  :  128 - 0x80
    "00011000", -- 3402 - 0xd4a  :   24 - 0x18
    "00110000", -- 3403 - 0xd4b  :   48 - 0x30
    "00110100", -- 3404 - 0xd4c  :   52 - 0x34
    "11111110", -- 3405 - 0xd4d  :  254 - 0xfe
    "11111110", -- 3406 - 0xd4e  :  254 - 0xfe
    "11111110", -- 3407 - 0xd4f  :  254 - 0xfe
    "00000000", -- 3408 - 0xd50  :    0 - 0x0
    "00000001", -- 3409 - 0xd51  :    1 - 0x1
    "00000000", -- 3410 - 0xd52  :    0 - 0x0
    "00000111", -- 3411 - 0xd53  :    7 - 0x7
    "00000111", -- 3412 - 0xd54  :    7 - 0x7
    "00000111", -- 3413 - 0xd55  :    7 - 0x7
    "00000111", -- 3414 - 0xd56  :    7 - 0x7
    "00011111", -- 3415 - 0xd57  :   31 - 0x1f
    "00000000", -- 3416 - 0xd58  :    0 - 0x0
    "00000000", -- 3417 - 0xd59  :    0 - 0x0
    "00000001", -- 3418 - 0xd5a  :    1 - 0x1
    "00000100", -- 3419 - 0xd5b  :    4 - 0x4
    "00000110", -- 3420 - 0xd5c  :    6 - 0x6
    "00000110", -- 3421 - 0xd5d  :    6 - 0x6
    "00000111", -- 3422 - 0xd5e  :    7 - 0x7
    "00000111", -- 3423 - 0xd5f  :    7 - 0x7
    "00000000", -- 3424 - 0xd60  :    0 - 0x0
    "00000000", -- 3425 - 0xd61  :    0 - 0x0
    "00001111", -- 3426 - 0xd62  :   15 - 0xf
    "00111111", -- 3427 - 0xd63  :   63 - 0x3f
    "00111111", -- 3428 - 0xd64  :   63 - 0x3f
    "00001111", -- 3429 - 0xd65  :   15 - 0xf
    "00000000", -- 3430 - 0xd66  :    0 - 0x0
    "00000000", -- 3431 - 0xd67  :    0 - 0x0
    "00001111", -- 3432 - 0xd68  :   15 - 0xf
    "00111111", -- 3433 - 0xd69  :   63 - 0x3f
    "01111111", -- 3434 - 0xd6a  :  127 - 0x7f
    "11111000", -- 3435 - 0xd6b  :  248 - 0xf8
    "11111000", -- 3436 - 0xd6c  :  248 - 0xf8
    "01111111", -- 3437 - 0xd6d  :  127 - 0x7f
    "00111111", -- 3438 - 0xd6e  :   63 - 0x3f
    "00001111", -- 3439 - 0xd6f  :   15 - 0xf
    "01111000", -- 3440 - 0xd70  :  120 - 0x78
    "01111100", -- 3441 - 0xd71  :  124 - 0x7c
    "01111110", -- 3442 - 0xd72  :  126 - 0x7e
    "01111111", -- 3443 - 0xd73  :  127 - 0x7f
    "00111111", -- 3444 - 0xd74  :   63 - 0x3f
    "00111111", -- 3445 - 0xd75  :   63 - 0x3f
    "00011011", -- 3446 - 0xd76  :   27 - 0x1b
    "00001001", -- 3447 - 0xd77  :    9 - 0x9
    "00011111", -- 3448 - 0xd78  :   31 - 0x1f
    "00011111", -- 3449 - 0xd79  :   31 - 0x1f
    "00011111", -- 3450 - 0xd7a  :   31 - 0x1f
    "00001011", -- 3451 - 0xd7b  :   11 - 0xb
    "00000001", -- 3452 - 0xd7c  :    1 - 0x1
    "00000001", -- 3453 - 0xd7d  :    1 - 0x1
    "00000000", -- 3454 - 0xd7e  :    0 - 0x0
    "00000000", -- 3455 - 0xd7f  :    0 - 0x0
    "00001100", -- 3456 - 0xd80  :   12 - 0xc
    "00000000", -- 3457 - 0xd81  :    0 - 0x0
    "00000000", -- 3458 - 0xd82  :    0 - 0x0
    "00000000", -- 3459 - 0xd83  :    0 - 0x0
    "00000111", -- 3460 - 0xd84  :    7 - 0x7
    "01111111", -- 3461 - 0xd85  :  127 - 0x7f
    "01111100", -- 3462 - 0xd86  :  124 - 0x7c
    "00000000", -- 3463 - 0xd87  :    0 - 0x0
    "00000011", -- 3464 - 0xd88  :    3 - 0x3
    "00011111", -- 3465 - 0xd89  :   31 - 0x1f
    "00111111", -- 3466 - 0xd8a  :   63 - 0x3f
    "00111111", -- 3467 - 0xd8b  :   63 - 0x3f
    "01111000", -- 3468 - 0xd8c  :  120 - 0x78
    "00000000", -- 3469 - 0xd8d  :    0 - 0x0
    "00000011", -- 3470 - 0xd8e  :    3 - 0x3
    "11111111", -- 3471 - 0xd8f  :  255 - 0xff
    "00000001", -- 3472 - 0xd90  :    1 - 0x1
    "11100001", -- 3473 - 0xd91  :  225 - 0xe1
    "01110001", -- 3474 - 0xd92  :  113 - 0x71
    "01111001", -- 3475 - 0xd93  :  121 - 0x79
    "00111101", -- 3476 - 0xd94  :   61 - 0x3d
    "00111101", -- 3477 - 0xd95  :   61 - 0x3d
    "00011111", -- 3478 - 0xd96  :   31 - 0x1f
    "00000011", -- 3479 - 0xd97  :    3 - 0x3
    "00000000", -- 3480 - 0xd98  :    0 - 0x0
    "00000000", -- 3481 - 0xd99  :    0 - 0x0
    "00000000", -- 3482 - 0xd9a  :    0 - 0x0
    "00000000", -- 3483 - 0xd9b  :    0 - 0x0
    "00000000", -- 3484 - 0xd9c  :    0 - 0x0
    "00000000", -- 3485 - 0xd9d  :    0 - 0x0
    "00000000", -- 3486 - 0xd9e  :    0 - 0x0
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "00111111", -- 3488 - 0xda0  :   63 - 0x3f
    "00111111", -- 3489 - 0xda1  :   63 - 0x3f
    "00011111", -- 3490 - 0xda2  :   31 - 0x1f
    "00011011", -- 3491 - 0xda3  :   27 - 0x1b
    "00110110", -- 3492 - 0xda4  :   54 - 0x36
    "00110000", -- 3493 - 0xda5  :   48 - 0x30
    "01111111", -- 3494 - 0xda6  :  127 - 0x7f
    "00111111", -- 3495 - 0xda7  :   63 - 0x3f
    "00100011", -- 3496 - 0xda8  :   35 - 0x23
    "00100111", -- 3497 - 0xda9  :   39 - 0x27
    "00011111", -- 3498 - 0xdaa  :   31 - 0x1f
    "00000111", -- 3499 - 0xdab  :    7 - 0x7
    "00001111", -- 3500 - 0xdac  :   15 - 0xf
    "00011111", -- 3501 - 0xdad  :   31 - 0x1f
    "01111111", -- 3502 - 0xdae  :  127 - 0x7f
    "00111111", -- 3503 - 0xdaf  :   63 - 0x3f
    "11111000", -- 3504 - 0xdb0  :  248 - 0xf8
    "11111000", -- 3505 - 0xdb1  :  248 - 0xf8
    "11111000", -- 3506 - 0xdb2  :  248 - 0xf8
    "10111000", -- 3507 - 0xdb3  :  184 - 0xb8
    "00011000", -- 3508 - 0xdb4  :   24 - 0x18
    "11011000", -- 3509 - 0xdb5  :  216 - 0xd8
    "11011000", -- 3510 - 0xdb6  :  216 - 0xd8
    "10111000", -- 3511 - 0xdb7  :  184 - 0xb8
    "11100000", -- 3512 - 0xdb8  :  224 - 0xe0
    "10000000", -- 3513 - 0xdb9  :  128 - 0x80
    "10000000", -- 3514 - 0xdba  :  128 - 0x80
    "01000000", -- 3515 - 0xdbb  :   64 - 0x40
    "11100000", -- 3516 - 0xdbc  :  224 - 0xe0
    "11100000", -- 3517 - 0xdbd  :  224 - 0xe0
    "11100000", -- 3518 - 0xdbe  :  224 - 0xe0
    "11000000", -- 3519 - 0xdbf  :  192 - 0xc0
    "00000001", -- 3520 - 0xdc0  :    1 - 0x1
    "00000010", -- 3521 - 0xdc1  :    2 - 0x2
    "00000100", -- 3522 - 0xdc2  :    4 - 0x4
    "00000100", -- 3523 - 0xdc3  :    4 - 0x4
    "00001000", -- 3524 - 0xdc4  :    8 - 0x8
    "00001000", -- 3525 - 0xdc5  :    8 - 0x8
    "00010000", -- 3526 - 0xdc6  :   16 - 0x10
    "00010000", -- 3527 - 0xdc7  :   16 - 0x10
    "00000011", -- 3528 - 0xdc8  :    3 - 0x3
    "00000111", -- 3529 - 0xdc9  :    7 - 0x7
    "00001111", -- 3530 - 0xdca  :   15 - 0xf
    "00011111", -- 3531 - 0xdcb  :   31 - 0x1f
    "00111111", -- 3532 - 0xdcc  :   63 - 0x3f
    "01111111", -- 3533 - 0xdcd  :  127 - 0x7f
    "11111111", -- 3534 - 0xdce  :  255 - 0xff
    "00011111", -- 3535 - 0xdcf  :   31 - 0x1f
    "00000000", -- 3536 - 0xdd0  :    0 - 0x0
    "00001111", -- 3537 - 0xdd1  :   15 - 0xf
    "00010011", -- 3538 - 0xdd2  :   19 - 0x13
    "00001101", -- 3539 - 0xdd3  :   13 - 0xd
    "00001101", -- 3540 - 0xdd4  :   13 - 0xd
    "00010011", -- 3541 - 0xdd5  :   19 - 0x13
    "00001100", -- 3542 - 0xdd6  :   12 - 0xc
    "00100000", -- 3543 - 0xdd7  :   32 - 0x20
    "00011111", -- 3544 - 0xdd8  :   31 - 0x1f
    "00010000", -- 3545 - 0xdd9  :   16 - 0x10
    "00001100", -- 3546 - 0xdda  :   12 - 0xc
    "00010010", -- 3547 - 0xddb  :   18 - 0x12
    "00010010", -- 3548 - 0xddc  :   18 - 0x12
    "00101100", -- 3549 - 0xddd  :   44 - 0x2c
    "00111111", -- 3550 - 0xdde  :   63 - 0x3f
    "00111111", -- 3551 - 0xddf  :   63 - 0x3f
    "00000000", -- 3552 - 0xde0  :    0 - 0x0
    "00100100", -- 3553 - 0xde1  :   36 - 0x24
    "00000000", -- 3554 - 0xde2  :    0 - 0x0
    "00100100", -- 3555 - 0xde3  :   36 - 0x24
    "00000000", -- 3556 - 0xde4  :    0 - 0x0
    "00000100", -- 3557 - 0xde5  :    4 - 0x4
    "00000000", -- 3558 - 0xde6  :    0 - 0x0
    "00000000", -- 3559 - 0xde7  :    0 - 0x0
    "00110111", -- 3560 - 0xde8  :   55 - 0x37
    "00110110", -- 3561 - 0xde9  :   54 - 0x36
    "00110110", -- 3562 - 0xdea  :   54 - 0x36
    "00110110", -- 3563 - 0xdeb  :   54 - 0x36
    "00010110", -- 3564 - 0xdec  :   22 - 0x16
    "00010110", -- 3565 - 0xded  :   22 - 0x16
    "00010010", -- 3566 - 0xdee  :   18 - 0x12
    "00000010", -- 3567 - 0xdef  :    2 - 0x2
    "00001111", -- 3568 - 0xdf0  :   15 - 0xf
    "01000001", -- 3569 - 0xdf1  :   65 - 0x41
    "00000000", -- 3570 - 0xdf2  :    0 - 0x0
    "10001000", -- 3571 - 0xdf3  :  136 - 0x88
    "00000000", -- 3572 - 0xdf4  :    0 - 0x0
    "01000100", -- 3573 - 0xdf5  :   68 - 0x44
    "00000000", -- 3574 - 0xdf6  :    0 - 0x0
    "00000000", -- 3575 - 0xdf7  :    0 - 0x0
    "00010000", -- 3576 - 0xdf8  :   16 - 0x10
    "01111110", -- 3577 - 0xdf9  :  126 - 0x7e
    "11111111", -- 3578 - 0xdfa  :  255 - 0xff
    "11111111", -- 3579 - 0xdfb  :  255 - 0xff
    "11110110", -- 3580 - 0xdfc  :  246 - 0xf6
    "01110110", -- 3581 - 0xdfd  :  118 - 0x76
    "00111010", -- 3582 - 0xdfe  :   58 - 0x3a
    "00011010", -- 3583 - 0xdff  :   26 - 0x1a
    "00111000", -- 3584 - 0xe00  :   56 - 0x38
    "01111100", -- 3585 - 0xe01  :  124 - 0x7c
    "11111110", -- 3586 - 0xe02  :  254 - 0xfe
    "11111110", -- 3587 - 0xe03  :  254 - 0xfe
    "00111011", -- 3588 - 0xe04  :   59 - 0x3b
    "00000011", -- 3589 - 0xe05  :    3 - 0x3
    "00000011", -- 3590 - 0xe06  :    3 - 0x3
    "00000011", -- 3591 - 0xe07  :    3 - 0x3
    "00000000", -- 3592 - 0xe08  :    0 - 0x0
    "00000000", -- 3593 - 0xe09  :    0 - 0x0
    "00111000", -- 3594 - 0xe0a  :   56 - 0x38
    "00000100", -- 3595 - 0xe0b  :    4 - 0x4
    "00000000", -- 3596 - 0xe0c  :    0 - 0x0
    "00000000", -- 3597 - 0xe0d  :    0 - 0x0
    "00000000", -- 3598 - 0xe0e  :    0 - 0x0
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "00000011", -- 3600 - 0xe10  :    3 - 0x3
    "00110011", -- 3601 - 0xe11  :   51 - 0x33
    "01111011", -- 3602 - 0xe12  :  123 - 0x7b
    "01111111", -- 3603 - 0xe13  :  127 - 0x7f
    "11111111", -- 3604 - 0xe14  :  255 - 0xff
    "11111011", -- 3605 - 0xe15  :  251 - 0xfb
    "00000011", -- 3606 - 0xe16  :    3 - 0x3
    "00000011", -- 3607 - 0xe17  :    3 - 0x3
    "00000000", -- 3608 - 0xe18  :    0 - 0x0
    "00000000", -- 3609 - 0xe19  :    0 - 0x0
    "00000000", -- 3610 - 0xe1a  :    0 - 0x0
    "00111000", -- 3611 - 0xe1b  :   56 - 0x38
    "01000000", -- 3612 - 0xe1c  :   64 - 0x40
    "00000000", -- 3613 - 0xe1d  :    0 - 0x0
    "00000000", -- 3614 - 0xe1e  :    0 - 0x0
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "11011100", -- 3616 - 0xe20  :  220 - 0xdc
    "11000000", -- 3617 - 0xe21  :  192 - 0xc0
    "11100000", -- 3618 - 0xe22  :  224 - 0xe0
    "11100000", -- 3619 - 0xe23  :  224 - 0xe0
    "11100000", -- 3620 - 0xe24  :  224 - 0xe0
    "11100000", -- 3621 - 0xe25  :  224 - 0xe0
    "11100000", -- 3622 - 0xe26  :  224 - 0xe0
    "11000000", -- 3623 - 0xe27  :  192 - 0xc0
    "11111100", -- 3624 - 0xe28  :  252 - 0xfc
    "10100000", -- 3625 - 0xe29  :  160 - 0xa0
    "10000000", -- 3626 - 0xe2a  :  128 - 0x80
    "10000000", -- 3627 - 0xe2b  :  128 - 0x80
    "00000000", -- 3628 - 0xe2c  :    0 - 0x0
    "00000000", -- 3629 - 0xe2d  :    0 - 0x0
    "00000000", -- 3630 - 0xe2e  :    0 - 0x0
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "00111111", -- 3632 - 0xe30  :   63 - 0x3f
    "01011111", -- 3633 - 0xe31  :   95 - 0x5f
    "00111111", -- 3634 - 0xe32  :   63 - 0x3f
    "00111111", -- 3635 - 0xe33  :   63 - 0x3f
    "10111011", -- 3636 - 0xe34  :  187 - 0xbb
    "11111000", -- 3637 - 0xe35  :  248 - 0xf8
    "11111110", -- 3638 - 0xe36  :  254 - 0xfe
    "11111110", -- 3639 - 0xe37  :  254 - 0xfe
    "00000111", -- 3640 - 0xe38  :    7 - 0x7
    "00100111", -- 3641 - 0xe39  :   39 - 0x27
    "01010111", -- 3642 - 0xe3a  :   87 - 0x57
    "01001111", -- 3643 - 0xe3b  :   79 - 0x4f
    "01010111", -- 3644 - 0xe3c  :   87 - 0x57
    "00100111", -- 3645 - 0xe3d  :   39 - 0x27
    "11000001", -- 3646 - 0xe3e  :  193 - 0xc1
    "00100001", -- 3647 - 0xe3f  :   33 - 0x21
    "00011111", -- 3648 - 0xe40  :   31 - 0x1f
    "00001111", -- 3649 - 0xe41  :   15 - 0xf
    "00001111", -- 3650 - 0xe42  :   15 - 0xf
    "00011111", -- 3651 - 0xe43  :   31 - 0x1f
    "00011111", -- 3652 - 0xe44  :   31 - 0x1f
    "00011110", -- 3653 - 0xe45  :   30 - 0x1e
    "00111000", -- 3654 - 0xe46  :   56 - 0x38
    "00110000", -- 3655 - 0xe47  :   48 - 0x30
    "00011101", -- 3656 - 0xe48  :   29 - 0x1d
    "00001111", -- 3657 - 0xe49  :   15 - 0xf
    "00001111", -- 3658 - 0xe4a  :   15 - 0xf
    "00011111", -- 3659 - 0xe4b  :   31 - 0x1f
    "00011111", -- 3660 - 0xe4c  :   31 - 0x1f
    "00011110", -- 3661 - 0xe4d  :   30 - 0x1e
    "00111000", -- 3662 - 0xe4e  :   56 - 0x38
    "00110000", -- 3663 - 0xe4f  :   48 - 0x30
    "00000000", -- 3664 - 0xe50  :    0 - 0x0
    "00100000", -- 3665 - 0xe51  :   32 - 0x20
    "01100000", -- 3666 - 0xe52  :   96 - 0x60
    "01100000", -- 3667 - 0xe53  :   96 - 0x60
    "01110000", -- 3668 - 0xe54  :  112 - 0x70
    "11110000", -- 3669 - 0xe55  :  240 - 0xf0
    "11111000", -- 3670 - 0xe56  :  248 - 0xf8
    "11111000", -- 3671 - 0xe57  :  248 - 0xf8
    "00000000", -- 3672 - 0xe58  :    0 - 0x0
    "00000000", -- 3673 - 0xe59  :    0 - 0x0
    "00111000", -- 3674 - 0xe5a  :   56 - 0x38
    "00010000", -- 3675 - 0xe5b  :   16 - 0x10
    "01001100", -- 3676 - 0xe5c  :   76 - 0x4c
    "00011000", -- 3677 - 0xe5d  :   24 - 0x18
    "10000110", -- 3678 - 0xe5e  :  134 - 0x86
    "00100100", -- 3679 - 0xe5f  :   36 - 0x24
    "11111000", -- 3680 - 0xe60  :  248 - 0xf8
    "11111100", -- 3681 - 0xe61  :  252 - 0xfc
    "11111100", -- 3682 - 0xe62  :  252 - 0xfc
    "01111110", -- 3683 - 0xe63  :  126 - 0x7e
    "01111110", -- 3684 - 0xe64  :  126 - 0x7e
    "00111110", -- 3685 - 0xe65  :   62 - 0x3e
    "00011111", -- 3686 - 0xe66  :   31 - 0x1f
    "00000111", -- 3687 - 0xe67  :    7 - 0x7
    "00000000", -- 3688 - 0xe68  :    0 - 0x0
    "01000010", -- 3689 - 0xe69  :   66 - 0x42
    "00001010", -- 3690 - 0xe6a  :   10 - 0xa
    "01000000", -- 3691 - 0xe6b  :   64 - 0x40
    "00010000", -- 3692 - 0xe6c  :   16 - 0x10
    "00000010", -- 3693 - 0xe6d  :    2 - 0x2
    "00001000", -- 3694 - 0xe6e  :    8 - 0x8
    "00000010", -- 3695 - 0xe6f  :    2 - 0x2
    "00000000", -- 3696 - 0xe70  :    0 - 0x0
    "11000000", -- 3697 - 0xe71  :  192 - 0xc0
    "01110000", -- 3698 - 0xe72  :  112 - 0x70
    "10111000", -- 3699 - 0xe73  :  184 - 0xb8
    "11110100", -- 3700 - 0xe74  :  244 - 0xf4
    "11110010", -- 3701 - 0xe75  :  242 - 0xf2
    "11110101", -- 3702 - 0xe76  :  245 - 0xf5
    "01111011", -- 3703 - 0xe77  :  123 - 0x7b
    "00000000", -- 3704 - 0xe78  :    0 - 0x0
    "00000000", -- 3705 - 0xe79  :    0 - 0x0
    "10000000", -- 3706 - 0xe7a  :  128 - 0x80
    "01000000", -- 3707 - 0xe7b  :   64 - 0x40
    "00001000", -- 3708 - 0xe7c  :    8 - 0x8
    "00001100", -- 3709 - 0xe7d  :   12 - 0xc
    "00001010", -- 3710 - 0xe7e  :   10 - 0xa
    "10000100", -- 3711 - 0xe7f  :  132 - 0x84
    "00000000", -- 3712 - 0xe80  :    0 - 0x0
    "11011111", -- 3713 - 0xe81  :  223 - 0xdf
    "00010000", -- 3714 - 0xe82  :   16 - 0x10
    "11111111", -- 3715 - 0xe83  :  255 - 0xff
    "11011111", -- 3716 - 0xe84  :  223 - 0xdf
    "11111111", -- 3717 - 0xe85  :  255 - 0xff
    "11111111", -- 3718 - 0xe86  :  255 - 0xff
    "11111001", -- 3719 - 0xe87  :  249 - 0xf9
    "00000000", -- 3720 - 0xe88  :    0 - 0x0
    "00000000", -- 3721 - 0xe89  :    0 - 0x0
    "11001111", -- 3722 - 0xe8a  :  207 - 0xcf
    "00100000", -- 3723 - 0xe8b  :   32 - 0x20
    "00100000", -- 3724 - 0xe8c  :   32 - 0x20
    "00100000", -- 3725 - 0xe8d  :   32 - 0x20
    "00100110", -- 3726 - 0xe8e  :   38 - 0x26
    "00101110", -- 3727 - 0xe8f  :   46 - 0x2e
    "00011111", -- 3728 - 0xe90  :   31 - 0x1f
    "00011111", -- 3729 - 0xe91  :   31 - 0x1f
    "00111110", -- 3730 - 0xe92  :   62 - 0x3e
    "11111100", -- 3731 - 0xe93  :  252 - 0xfc
    "11111000", -- 3732 - 0xe94  :  248 - 0xf8
    "11110000", -- 3733 - 0xe95  :  240 - 0xf0
    "11000000", -- 3734 - 0xe96  :  192 - 0xc0
    "00000000", -- 3735 - 0xe97  :    0 - 0x0
    "11100000", -- 3736 - 0xe98  :  224 - 0xe0
    "11100000", -- 3737 - 0xe99  :  224 - 0xe0
    "11000000", -- 3738 - 0xe9a  :  192 - 0xc0
    "00000000", -- 3739 - 0xe9b  :    0 - 0x0
    "00000000", -- 3740 - 0xe9c  :    0 - 0x0
    "00000000", -- 3741 - 0xe9d  :    0 - 0x0
    "00000000", -- 3742 - 0xe9e  :    0 - 0x0
    "00000000", -- 3743 - 0xe9f  :    0 - 0x0
    "11111000", -- 3744 - 0xea0  :  248 - 0xf8
    "11111100", -- 3745 - 0xea1  :  252 - 0xfc
    "11111110", -- 3746 - 0xea2  :  254 - 0xfe
    "11111111", -- 3747 - 0xea3  :  255 - 0xff
    "11111111", -- 3748 - 0xea4  :  255 - 0xff
    "11011111", -- 3749 - 0xea5  :  223 - 0xdf
    "11011111", -- 3750 - 0xea6  :  223 - 0xdf
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "00101111", -- 3752 - 0xea8  :   47 - 0x2f
    "00100011", -- 3753 - 0xea9  :   35 - 0x23
    "00100001", -- 3754 - 0xeaa  :   33 - 0x21
    "00100000", -- 3755 - 0xeab  :   32 - 0x20
    "00100000", -- 3756 - 0xeac  :   32 - 0x20
    "00000000", -- 3757 - 0xead  :    0 - 0x0
    "00000000", -- 3758 - 0xeae  :    0 - 0x0
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "11000001", -- 3760 - 0xeb0  :  193 - 0xc1
    "11110001", -- 3761 - 0xeb1  :  241 - 0xf1
    "01111001", -- 3762 - 0xeb2  :  121 - 0x79
    "01111101", -- 3763 - 0xeb3  :  125 - 0x7d
    "00111101", -- 3764 - 0xeb4  :   61 - 0x3d
    "00111111", -- 3765 - 0xeb5  :   63 - 0x3f
    "00011111", -- 3766 - 0xeb6  :   31 - 0x1f
    "00000011", -- 3767 - 0xeb7  :    3 - 0x3
    "11000001", -- 3768 - 0xeb8  :  193 - 0xc1
    "10110001", -- 3769 - 0xeb9  :  177 - 0xb1
    "01011001", -- 3770 - 0xeba  :   89 - 0x59
    "01101101", -- 3771 - 0xebb  :  109 - 0x6d
    "00110101", -- 3772 - 0xebc  :   53 - 0x35
    "00111011", -- 3773 - 0xebd  :   59 - 0x3b
    "00011111", -- 3774 - 0xebe  :   31 - 0x1f
    "00000011", -- 3775 - 0xebf  :    3 - 0x3
    "00000010", -- 3776 - 0xec0  :    2 - 0x2
    "00000110", -- 3777 - 0xec1  :    6 - 0x6
    "00001110", -- 3778 - 0xec2  :   14 - 0xe
    "00001110", -- 3779 - 0xec3  :   14 - 0xe
    "00011110", -- 3780 - 0xec4  :   30 - 0x1e
    "00011110", -- 3781 - 0xec5  :   30 - 0x1e
    "00111110", -- 3782 - 0xec6  :   62 - 0x3e
    "00111110", -- 3783 - 0xec7  :   62 - 0x3e
    "00000000", -- 3784 - 0xec8  :    0 - 0x0
    "00000010", -- 3785 - 0xec9  :    2 - 0x2
    "00000000", -- 3786 - 0xeca  :    0 - 0x0
    "00001000", -- 3787 - 0xecb  :    8 - 0x8
    "00000010", -- 3788 - 0xecc  :    2 - 0x2
    "00000000", -- 3789 - 0xecd  :    0 - 0x0
    "00101000", -- 3790 - 0xece  :   40 - 0x28
    "00000000", -- 3791 - 0xecf  :    0 - 0x0
    "00111110", -- 3792 - 0xed0  :   62 - 0x3e
    "00111110", -- 3793 - 0xed1  :   62 - 0x3e
    "00111110", -- 3794 - 0xed2  :   62 - 0x3e
    "00111110", -- 3795 - 0xed3  :   62 - 0x3e
    "00011110", -- 3796 - 0xed4  :   30 - 0x1e
    "00011110", -- 3797 - 0xed5  :   30 - 0x1e
    "00001110", -- 3798 - 0xed6  :   14 - 0xe
    "00000010", -- 3799 - 0xed7  :    2 - 0x2
    "00000100", -- 3800 - 0xed8  :    4 - 0x4
    "00010000", -- 3801 - 0xed9  :   16 - 0x10
    "00000010", -- 3802 - 0xeda  :    2 - 0x2
    "00010000", -- 3803 - 0xedb  :   16 - 0x10
    "00000100", -- 3804 - 0xedc  :    4 - 0x4
    "00000000", -- 3805 - 0xedd  :    0 - 0x0
    "00001010", -- 3806 - 0xede  :   10 - 0xa
    "00000000", -- 3807 - 0xedf  :    0 - 0x0
    "11000001", -- 3808 - 0xee0  :  193 - 0xc1
    "11110001", -- 3809 - 0xee1  :  241 - 0xf1
    "01111001", -- 3810 - 0xee2  :  121 - 0x79
    "01111101", -- 3811 - 0xee3  :  125 - 0x7d
    "00111101", -- 3812 - 0xee4  :   61 - 0x3d
    "00111111", -- 3813 - 0xee5  :   63 - 0x3f
    "00011111", -- 3814 - 0xee6  :   31 - 0x1f
    "00000011", -- 3815 - 0xee7  :    3 - 0x3
    "11000001", -- 3816 - 0xee8  :  193 - 0xc1
    "10110001", -- 3817 - 0xee9  :  177 - 0xb1
    "01011001", -- 3818 - 0xeea  :   89 - 0x59
    "01101101", -- 3819 - 0xeeb  :  109 - 0x6d
    "00110101", -- 3820 - 0xeec  :   53 - 0x35
    "00111011", -- 3821 - 0xeed  :   59 - 0x3b
    "00011111", -- 3822 - 0xeee  :   31 - 0x1f
    "00000011", -- 3823 - 0xeef  :    3 - 0x3
    "01111100", -- 3824 - 0xef0  :  124 - 0x7c
    "00000000", -- 3825 - 0xef1  :    0 - 0x0
    "00000000", -- 3826 - 0xef2  :    0 - 0x0
    "11111111", -- 3827 - 0xef3  :  255 - 0xff
    "11000011", -- 3828 - 0xef4  :  195 - 0xc3
    "01111111", -- 3829 - 0xef5  :  127 - 0x7f
    "00011111", -- 3830 - 0xef6  :   31 - 0x1f
    "00000011", -- 3831 - 0xef7  :    3 - 0x3
    "00000000", -- 3832 - 0xef8  :    0 - 0x0
    "00001111", -- 3833 - 0xef9  :   15 - 0xf
    "00011111", -- 3834 - 0xefa  :   31 - 0x1f
    "11111111", -- 3835 - 0xefb  :  255 - 0xff
    "11111100", -- 3836 - 0xefc  :  252 - 0xfc
    "01100011", -- 3837 - 0xefd  :   99 - 0x63
    "00011111", -- 3838 - 0xefe  :   31 - 0x1f
    "00000011", -- 3839 - 0xeff  :    3 - 0x3
    "11111111", -- 3840 - 0xf00  :  255 - 0xff
    "11111111", -- 3841 - 0xf01  :  255 - 0xff
    "01111100", -- 3842 - 0xf02  :  124 - 0x7c
    "00000000", -- 3843 - 0xf03  :    0 - 0x0
    "00000000", -- 3844 - 0xf04  :    0 - 0x0
    "01111100", -- 3845 - 0xf05  :  124 - 0x7c
    "11111111", -- 3846 - 0xf06  :  255 - 0xff
    "11111111", -- 3847 - 0xf07  :  255 - 0xff
    "00000000", -- 3848 - 0xf08  :    0 - 0x0
    "00000000", -- 3849 - 0xf09  :    0 - 0x0
    "11111110", -- 3850 - 0xf0a  :  254 - 0xfe
    "11000110", -- 3851 - 0xf0b  :  198 - 0xc6
    "11000110", -- 3852 - 0xf0c  :  198 - 0xc6
    "11111110", -- 3853 - 0xf0d  :  254 - 0xfe
    "00000000", -- 3854 - 0xf0e  :    0 - 0x0
    "00000000", -- 3855 - 0xf0f  :    0 - 0x0
    "11111111", -- 3856 - 0xf10  :  255 - 0xff
    "11111111", -- 3857 - 0xf11  :  255 - 0xff
    "00000000", -- 3858 - 0xf12  :    0 - 0x0
    "00000100", -- 3859 - 0xf13  :    4 - 0x4
    "00001100", -- 3860 - 0xf14  :   12 - 0xc
    "00011000", -- 3861 - 0xf15  :   24 - 0x18
    "00110000", -- 3862 - 0xf16  :   48 - 0x30
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "00000000", -- 3864 - 0xf18  :    0 - 0x0
    "00000000", -- 3865 - 0xf19  :    0 - 0x0
    "00000110", -- 3866 - 0xf1a  :    6 - 0x6
    "00000110", -- 3867 - 0xf1b  :    6 - 0x6
    "00001100", -- 3868 - 0xf1c  :   12 - 0xc
    "00011000", -- 3869 - 0xf1d  :   24 - 0x18
    "01110000", -- 3870 - 0xf1e  :  112 - 0x70
    "01100000", -- 3871 - 0xf1f  :   96 - 0x60
    "11111111", -- 3872 - 0xf20  :  255 - 0xff
    "11111111", -- 3873 - 0xf21  :  255 - 0xff
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000100", -- 3875 - 0xf23  :    4 - 0x4
    "00000100", -- 3876 - 0xf24  :    4 - 0x4
    "00000100", -- 3877 - 0xf25  :    4 - 0x4
    "00001000", -- 3878 - 0xf26  :    8 - 0x8
    "00001000", -- 3879 - 0xf27  :    8 - 0x8
    "00000000", -- 3880 - 0xf28  :    0 - 0x0
    "00000000", -- 3881 - 0xf29  :    0 - 0x0
    "00000110", -- 3882 - 0xf2a  :    6 - 0x6
    "00000110", -- 3883 - 0xf2b  :    6 - 0x6
    "00000100", -- 3884 - 0xf2c  :    4 - 0x4
    "00000100", -- 3885 - 0xf2d  :    4 - 0x4
    "00001000", -- 3886 - 0xf2e  :    8 - 0x8
    "00001000", -- 3887 - 0xf2f  :    8 - 0x8
    "00001000", -- 3888 - 0xf30  :    8 - 0x8
    "00010000", -- 3889 - 0xf31  :   16 - 0x10
    "00010000", -- 3890 - 0xf32  :   16 - 0x10
    "00000000", -- 3891 - 0xf33  :    0 - 0x0
    "00000000", -- 3892 - 0xf34  :    0 - 0x0
    "00010000", -- 3893 - 0xf35  :   16 - 0x10
    "00010000", -- 3894 - 0xf36  :   16 - 0x10
    "00001000", -- 3895 - 0xf37  :    8 - 0x8
    "00001000", -- 3896 - 0xf38  :    8 - 0x8
    "00010000", -- 3897 - 0xf39  :   16 - 0x10
    "00110000", -- 3898 - 0xf3a  :   48 - 0x30
    "00110000", -- 3899 - 0xf3b  :   48 - 0x30
    "00110000", -- 3900 - 0xf3c  :   48 - 0x30
    "00110000", -- 3901 - 0xf3d  :   48 - 0x30
    "00010000", -- 3902 - 0xf3e  :   16 - 0x10
    "00001000", -- 3903 - 0xf3f  :    8 - 0x8
    "01111111", -- 3904 - 0xf40  :  127 - 0x7f
    "00111111", -- 3905 - 0xf41  :   63 - 0x3f
    "00111111", -- 3906 - 0xf42  :   63 - 0x3f
    "00111110", -- 3907 - 0xf43  :   62 - 0x3e
    "00011111", -- 3908 - 0xf44  :   31 - 0x1f
    "00001111", -- 3909 - 0xf45  :   15 - 0xf
    "00000011", -- 3910 - 0xf46  :    3 - 0x3
    "00000000", -- 3911 - 0xf47  :    0 - 0x0
    "00000000", -- 3912 - 0xf48  :    0 - 0x0
    "00000000", -- 3913 - 0xf49  :    0 - 0x0
    "00000001", -- 3914 - 0xf4a  :    1 - 0x1
    "00000011", -- 3915 - 0xf4b  :    3 - 0x3
    "00000001", -- 3916 - 0xf4c  :    1 - 0x1
    "00000000", -- 3917 - 0xf4d  :    0 - 0x0
    "00000000", -- 3918 - 0xf4e  :    0 - 0x0
    "00000000", -- 3919 - 0xf4f  :    0 - 0x0
    "00000011", -- 3920 - 0xf50  :    3 - 0x3
    "00001111", -- 3921 - 0xf51  :   15 - 0xf
    "11111111", -- 3922 - 0xf52  :  255 - 0xff
    "01111111", -- 3923 - 0xf53  :  127 - 0x7f
    "01111111", -- 3924 - 0xf54  :  127 - 0x7f
    "01111111", -- 3925 - 0xf55  :  127 - 0x7f
    "01111111", -- 3926 - 0xf56  :  127 - 0x7f
    "01111111", -- 3927 - 0xf57  :  127 - 0x7f
    "00000011", -- 3928 - 0xf58  :    3 - 0x3
    "00001110", -- 3929 - 0xf59  :   14 - 0xe
    "11111000", -- 3930 - 0xf5a  :  248 - 0xf8
    "00000000", -- 3931 - 0xf5b  :    0 - 0x0
    "00000000", -- 3932 - 0xf5c  :    0 - 0x0
    "00000000", -- 3933 - 0xf5d  :    0 - 0x0
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00000000", -- 3941 - 0xf65  :    0 - 0x0
    "00000000", -- 3942 - 0xf66  :    0 - 0x0
    "00000000", -- 3943 - 0xf67  :    0 - 0x0
    "00100010", -- 3944 - 0xf68  :   34 - 0x22
    "01100101", -- 3945 - 0xf69  :  101 - 0x65
    "00100101", -- 3946 - 0xf6a  :   37 - 0x25
    "00100101", -- 3947 - 0xf6b  :   37 - 0x25
    "00100101", -- 3948 - 0xf6c  :   37 - 0x25
    "00100101", -- 3949 - 0xf6d  :   37 - 0x25
    "01110111", -- 3950 - 0xf6e  :  119 - 0x77
    "01110010", -- 3951 - 0xf6f  :  114 - 0x72
    "00000000", -- 3952 - 0xf70  :    0 - 0x0
    "00000000", -- 3953 - 0xf71  :    0 - 0x0
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00000000", -- 3958 - 0xf76  :    0 - 0x0
    "00000000", -- 3959 - 0xf77  :    0 - 0x0
    "01100010", -- 3960 - 0xf78  :   98 - 0x62
    "10010101", -- 3961 - 0xf79  :  149 - 0x95
    "00010101", -- 3962 - 0xf7a  :   21 - 0x15
    "00100101", -- 3963 - 0xf7b  :   37 - 0x25
    "01000101", -- 3964 - 0xf7c  :   69 - 0x45
    "10000101", -- 3965 - 0xf7d  :  133 - 0x85
    "11110111", -- 3966 - 0xf7e  :  247 - 0xf7
    "11110010", -- 3967 - 0xf7f  :  242 - 0xf2
    "00000000", -- 3968 - 0xf80  :    0 - 0x0
    "00000000", -- 3969 - 0xf81  :    0 - 0x0
    "00000000", -- 3970 - 0xf82  :    0 - 0x0
    "00000000", -- 3971 - 0xf83  :    0 - 0x0
    "00000000", -- 3972 - 0xf84  :    0 - 0x0
    "00000000", -- 3973 - 0xf85  :    0 - 0x0
    "00000000", -- 3974 - 0xf86  :    0 - 0x0
    "00000000", -- 3975 - 0xf87  :    0 - 0x0
    "10100010", -- 3976 - 0xf88  :  162 - 0xa2
    "10100101", -- 3977 - 0xf89  :  165 - 0xa5
    "10100101", -- 3978 - 0xf8a  :  165 - 0xa5
    "10100101", -- 3979 - 0xf8b  :  165 - 0xa5
    "11110101", -- 3980 - 0xf8c  :  245 - 0xf5
    "11110101", -- 3981 - 0xf8d  :  245 - 0xf5
    "00100111", -- 3982 - 0xf8e  :   39 - 0x27
    "00100010", -- 3983 - 0xf8f  :   34 - 0x22
    "00000000", -- 3984 - 0xf90  :    0 - 0x0
    "00000000", -- 3985 - 0xf91  :    0 - 0x0
    "00000000", -- 3986 - 0xf92  :    0 - 0x0
    "00000000", -- 3987 - 0xf93  :    0 - 0x0
    "00000000", -- 3988 - 0xf94  :    0 - 0x0
    "00000000", -- 3989 - 0xf95  :    0 - 0x0
    "00000000", -- 3990 - 0xf96  :    0 - 0x0
    "00000000", -- 3991 - 0xf97  :    0 - 0x0
    "11110010", -- 3992 - 0xf98  :  242 - 0xf2
    "10000101", -- 3993 - 0xf99  :  133 - 0x85
    "10000101", -- 3994 - 0xf9a  :  133 - 0x85
    "11100101", -- 3995 - 0xf9b  :  229 - 0xe5
    "00010101", -- 3996 - 0xf9c  :   21 - 0x15
    "00010101", -- 3997 - 0xf9d  :   21 - 0x15
    "11110111", -- 3998 - 0xf9e  :  247 - 0xf7
    "11100010", -- 3999 - 0xf9f  :  226 - 0xe2
    "00000000", -- 4000 - 0xfa0  :    0 - 0x0
    "00000000", -- 4001 - 0xfa1  :    0 - 0x0
    "00000000", -- 4002 - 0xfa2  :    0 - 0x0
    "00000000", -- 4003 - 0xfa3  :    0 - 0x0
    "00000000", -- 4004 - 0xfa4  :    0 - 0x0
    "00000000", -- 4005 - 0xfa5  :    0 - 0x0
    "00000000", -- 4006 - 0xfa6  :    0 - 0x0
    "00000000", -- 4007 - 0xfa7  :    0 - 0x0
    "01100010", -- 4008 - 0xfa8  :   98 - 0x62
    "10010101", -- 4009 - 0xfa9  :  149 - 0x95
    "01010101", -- 4010 - 0xfaa  :   85 - 0x55
    "01100101", -- 4011 - 0xfab  :  101 - 0x65
    "10110101", -- 4012 - 0xfac  :  181 - 0xb5
    "10010101", -- 4013 - 0xfad  :  149 - 0x95
    "10010111", -- 4014 - 0xfae  :  151 - 0x97
    "01100010", -- 4015 - 0xfaf  :   98 - 0x62
    "00000000", -- 4016 - 0xfb0  :    0 - 0x0
    "00000000", -- 4017 - 0xfb1  :    0 - 0x0
    "00000000", -- 4018 - 0xfb2  :    0 - 0x0
    "00000000", -- 4019 - 0xfb3  :    0 - 0x0
    "00000000", -- 4020 - 0xfb4  :    0 - 0x0
    "00000000", -- 4021 - 0xfb5  :    0 - 0x0
    "00000000", -- 4022 - 0xfb6  :    0 - 0x0
    "00000000", -- 4023 - 0xfb7  :    0 - 0x0
    "00100000", -- 4024 - 0xfb8  :   32 - 0x20
    "01010000", -- 4025 - 0xfb9  :   80 - 0x50
    "01010000", -- 4026 - 0xfba  :   80 - 0x50
    "01010000", -- 4027 - 0xfbb  :   80 - 0x50
    "01010000", -- 4028 - 0xfbc  :   80 - 0x50
    "01010000", -- 4029 - 0xfbd  :   80 - 0x50
    "01110000", -- 4030 - 0xfbe  :  112 - 0x70
    "00100000", -- 4031 - 0xfbf  :   32 - 0x20
    "00000000", -- 4032 - 0xfc0  :    0 - 0x0
    "00000000", -- 4033 - 0xfc1  :    0 - 0x0
    "00000000", -- 4034 - 0xfc2  :    0 - 0x0
    "00000000", -- 4035 - 0xfc3  :    0 - 0x0
    "00000000", -- 4036 - 0xfc4  :    0 - 0x0
    "00000000", -- 4037 - 0xfc5  :    0 - 0x0
    "00000000", -- 4038 - 0xfc6  :    0 - 0x0
    "00000000", -- 4039 - 0xfc7  :    0 - 0x0
    "00000000", -- 4040 - 0xfc8  :    0 - 0x0
    "00000000", -- 4041 - 0xfc9  :    0 - 0x0
    "00000000", -- 4042 - 0xfca  :    0 - 0x0
    "00000000", -- 4043 - 0xfcb  :    0 - 0x0
    "00000000", -- 4044 - 0xfcc  :    0 - 0x0
    "00000000", -- 4045 - 0xfcd  :    0 - 0x0
    "00000000", -- 4046 - 0xfce  :    0 - 0x0
    "00000000", -- 4047 - 0xfcf  :    0 - 0x0
    "00000000", -- 4048 - 0xfd0  :    0 - 0x0
    "00000000", -- 4049 - 0xfd1  :    0 - 0x0
    "00000000", -- 4050 - 0xfd2  :    0 - 0x0
    "00000000", -- 4051 - 0xfd3  :    0 - 0x0
    "00000000", -- 4052 - 0xfd4  :    0 - 0x0
    "00000000", -- 4053 - 0xfd5  :    0 - 0x0
    "00000000", -- 4054 - 0xfd6  :    0 - 0x0
    "00000000", -- 4055 - 0xfd7  :    0 - 0x0
    "01100110", -- 4056 - 0xfd8  :  102 - 0x66
    "11100110", -- 4057 - 0xfd9  :  230 - 0xe6
    "01100110", -- 4058 - 0xfda  :  102 - 0x66
    "01100110", -- 4059 - 0xfdb  :  102 - 0x66
    "01100110", -- 4060 - 0xfdc  :  102 - 0x66
    "01100111", -- 4061 - 0xfdd  :  103 - 0x67
    "11110011", -- 4062 - 0xfde  :  243 - 0xf3
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00000000", -- 4064 - 0xfe0  :    0 - 0x0
    "00000000", -- 4065 - 0xfe1  :    0 - 0x0
    "00000000", -- 4066 - 0xfe2  :    0 - 0x0
    "00000000", -- 4067 - 0xfe3  :    0 - 0x0
    "00000000", -- 4068 - 0xfe4  :    0 - 0x0
    "00000000", -- 4069 - 0xfe5  :    0 - 0x0
    "00000000", -- 4070 - 0xfe6  :    0 - 0x0
    "00000000", -- 4071 - 0xfe7  :    0 - 0x0
    "01011110", -- 4072 - 0xfe8  :   94 - 0x5e
    "01011001", -- 4073 - 0xfe9  :   89 - 0x59
    "01011001", -- 4074 - 0xfea  :   89 - 0x59
    "01011001", -- 4075 - 0xfeb  :   89 - 0x59
    "01011110", -- 4076 - 0xfec  :   94 - 0x5e
    "11011000", -- 4077 - 0xfed  :  216 - 0xd8
    "10011000", -- 4078 - 0xfee  :  152 - 0x98
    "00000000", -- 4079 - 0xfef  :    0 - 0x0
    "00000000", -- 4080 - 0xff0  :    0 - 0x0
    "00000000", -- 4081 - 0xff1  :    0 - 0x0
    "00000000", -- 4082 - 0xff2  :    0 - 0x0
    "00000000", -- 4083 - 0xff3  :    0 - 0x0
    "00000000", -- 4084 - 0xff4  :    0 - 0x0
    "01111100", -- 4085 - 0xff5  :  124 - 0x7c
    "00111000", -- 4086 - 0xff6  :   56 - 0x38
    "00000000", -- 4087 - 0xff7  :    0 - 0x0
    "00000000", -- 4088 - 0xff8  :    0 - 0x0
    "00000000", -- 4089 - 0xff9  :    0 - 0x0
    "00000000", -- 4090 - 0xffa  :    0 - 0x0
    "00000000", -- 4091 - 0xffb  :    0 - 0x0
    "00000000", -- 4092 - 0xffc  :    0 - 0x0
    "00000100", -- 4093 - 0xffd  :    4 - 0x4
    "00001000", -- 4094 - 0xffe  :    8 - 0x8
    "00000000", -- 4095 - 0xfff  :    0 - 0x0
    "00111000", -- 4096 - 0x1000  :   56 - 0x38
    "01001100", -- 4097 - 0x1001  :   76 - 0x4c
    "11000110", -- 4098 - 0x1002  :  198 - 0xc6
    "11000110", -- 4099 - 0x1003  :  198 - 0xc6
    "11000110", -- 4100 - 0x1004  :  198 - 0xc6
    "01100100", -- 4101 - 0x1005  :  100 - 0x64
    "00111000", -- 4102 - 0x1006  :   56 - 0x38
    "00000000", -- 4103 - 0x1007  :    0 - 0x0
    "00000000", -- 4104 - 0x1008  :    0 - 0x0
    "00000000", -- 4105 - 0x1009  :    0 - 0x0
    "00000000", -- 4106 - 0x100a  :    0 - 0x0
    "00000000", -- 4107 - 0x100b  :    0 - 0x0
    "00000000", -- 4108 - 0x100c  :    0 - 0x0
    "00000000", -- 4109 - 0x100d  :    0 - 0x0
    "00000000", -- 4110 - 0x100e  :    0 - 0x0
    "00000000", -- 4111 - 0x100f  :    0 - 0x0
    "00011000", -- 4112 - 0x1010  :   24 - 0x18
    "00111000", -- 4113 - 0x1011  :   56 - 0x38
    "00011000", -- 4114 - 0x1012  :   24 - 0x18
    "00011000", -- 4115 - 0x1013  :   24 - 0x18
    "00011000", -- 4116 - 0x1014  :   24 - 0x18
    "00011000", -- 4117 - 0x1015  :   24 - 0x18
    "01111110", -- 4118 - 0x1016  :  126 - 0x7e
    "00000000", -- 4119 - 0x1017  :    0 - 0x0
    "00000000", -- 4120 - 0x1018  :    0 - 0x0
    "00000000", -- 4121 - 0x1019  :    0 - 0x0
    "00000000", -- 4122 - 0x101a  :    0 - 0x0
    "00000000", -- 4123 - 0x101b  :    0 - 0x0
    "00000000", -- 4124 - 0x101c  :    0 - 0x0
    "00000000", -- 4125 - 0x101d  :    0 - 0x0
    "00000000", -- 4126 - 0x101e  :    0 - 0x0
    "00000000", -- 4127 - 0x101f  :    0 - 0x0
    "01111100", -- 4128 - 0x1020  :  124 - 0x7c
    "11000110", -- 4129 - 0x1021  :  198 - 0xc6
    "00001110", -- 4130 - 0x1022  :   14 - 0xe
    "00111100", -- 4131 - 0x1023  :   60 - 0x3c
    "01111000", -- 4132 - 0x1024  :  120 - 0x78
    "11100000", -- 4133 - 0x1025  :  224 - 0xe0
    "11111110", -- 4134 - 0x1026  :  254 - 0xfe
    "00000000", -- 4135 - 0x1027  :    0 - 0x0
    "00000000", -- 4136 - 0x1028  :    0 - 0x0
    "00000000", -- 4137 - 0x1029  :    0 - 0x0
    "00000000", -- 4138 - 0x102a  :    0 - 0x0
    "00000000", -- 4139 - 0x102b  :    0 - 0x0
    "00000000", -- 4140 - 0x102c  :    0 - 0x0
    "00000000", -- 4141 - 0x102d  :    0 - 0x0
    "00000000", -- 4142 - 0x102e  :    0 - 0x0
    "00000000", -- 4143 - 0x102f  :    0 - 0x0
    "01111110", -- 4144 - 0x1030  :  126 - 0x7e
    "00001100", -- 4145 - 0x1031  :   12 - 0xc
    "00011000", -- 4146 - 0x1032  :   24 - 0x18
    "00111100", -- 4147 - 0x1033  :   60 - 0x3c
    "00000110", -- 4148 - 0x1034  :    6 - 0x6
    "11000110", -- 4149 - 0x1035  :  198 - 0xc6
    "01111100", -- 4150 - 0x1036  :  124 - 0x7c
    "00000000", -- 4151 - 0x1037  :    0 - 0x0
    "00000000", -- 4152 - 0x1038  :    0 - 0x0
    "00000000", -- 4153 - 0x1039  :    0 - 0x0
    "00000000", -- 4154 - 0x103a  :    0 - 0x0
    "00000000", -- 4155 - 0x103b  :    0 - 0x0
    "00000000", -- 4156 - 0x103c  :    0 - 0x0
    "00000000", -- 4157 - 0x103d  :    0 - 0x0
    "00000000", -- 4158 - 0x103e  :    0 - 0x0
    "00000000", -- 4159 - 0x103f  :    0 - 0x0
    "00011100", -- 4160 - 0x1040  :   28 - 0x1c
    "00111100", -- 4161 - 0x1041  :   60 - 0x3c
    "01101100", -- 4162 - 0x1042  :  108 - 0x6c
    "11001100", -- 4163 - 0x1043  :  204 - 0xcc
    "11111110", -- 4164 - 0x1044  :  254 - 0xfe
    "00001100", -- 4165 - 0x1045  :   12 - 0xc
    "00001100", -- 4166 - 0x1046  :   12 - 0xc
    "00000000", -- 4167 - 0x1047  :    0 - 0x0
    "00000000", -- 4168 - 0x1048  :    0 - 0x0
    "00000000", -- 4169 - 0x1049  :    0 - 0x0
    "00000000", -- 4170 - 0x104a  :    0 - 0x0
    "00000000", -- 4171 - 0x104b  :    0 - 0x0
    "00000000", -- 4172 - 0x104c  :    0 - 0x0
    "00000000", -- 4173 - 0x104d  :    0 - 0x0
    "00000000", -- 4174 - 0x104e  :    0 - 0x0
    "00000000", -- 4175 - 0x104f  :    0 - 0x0
    "11111100", -- 4176 - 0x1050  :  252 - 0xfc
    "11000000", -- 4177 - 0x1051  :  192 - 0xc0
    "11111100", -- 4178 - 0x1052  :  252 - 0xfc
    "00000110", -- 4179 - 0x1053  :    6 - 0x6
    "00000110", -- 4180 - 0x1054  :    6 - 0x6
    "11000110", -- 4181 - 0x1055  :  198 - 0xc6
    "01111100", -- 4182 - 0x1056  :  124 - 0x7c
    "00000000", -- 4183 - 0x1057  :    0 - 0x0
    "00000000", -- 4184 - 0x1058  :    0 - 0x0
    "00000000", -- 4185 - 0x1059  :    0 - 0x0
    "00000000", -- 4186 - 0x105a  :    0 - 0x0
    "00000000", -- 4187 - 0x105b  :    0 - 0x0
    "00000000", -- 4188 - 0x105c  :    0 - 0x0
    "00000000", -- 4189 - 0x105d  :    0 - 0x0
    "00000000", -- 4190 - 0x105e  :    0 - 0x0
    "00000000", -- 4191 - 0x105f  :    0 - 0x0
    "00111100", -- 4192 - 0x1060  :   60 - 0x3c
    "01100000", -- 4193 - 0x1061  :   96 - 0x60
    "11000000", -- 4194 - 0x1062  :  192 - 0xc0
    "11111100", -- 4195 - 0x1063  :  252 - 0xfc
    "11000110", -- 4196 - 0x1064  :  198 - 0xc6
    "11000110", -- 4197 - 0x1065  :  198 - 0xc6
    "01111100", -- 4198 - 0x1066  :  124 - 0x7c
    "00000000", -- 4199 - 0x1067  :    0 - 0x0
    "00000000", -- 4200 - 0x1068  :    0 - 0x0
    "00000000", -- 4201 - 0x1069  :    0 - 0x0
    "00000000", -- 4202 - 0x106a  :    0 - 0x0
    "00000000", -- 4203 - 0x106b  :    0 - 0x0
    "00000000", -- 4204 - 0x106c  :    0 - 0x0
    "00000000", -- 4205 - 0x106d  :    0 - 0x0
    "00000000", -- 4206 - 0x106e  :    0 - 0x0
    "00000000", -- 4207 - 0x106f  :    0 - 0x0
    "11111110", -- 4208 - 0x1070  :  254 - 0xfe
    "11000110", -- 4209 - 0x1071  :  198 - 0xc6
    "00001100", -- 4210 - 0x1072  :   12 - 0xc
    "00011000", -- 4211 - 0x1073  :   24 - 0x18
    "00110000", -- 4212 - 0x1074  :   48 - 0x30
    "00110000", -- 4213 - 0x1075  :   48 - 0x30
    "00110000", -- 4214 - 0x1076  :   48 - 0x30
    "00000000", -- 4215 - 0x1077  :    0 - 0x0
    "00000000", -- 4216 - 0x1078  :    0 - 0x0
    "00000000", -- 4217 - 0x1079  :    0 - 0x0
    "00000000", -- 4218 - 0x107a  :    0 - 0x0
    "00000000", -- 4219 - 0x107b  :    0 - 0x0
    "00000000", -- 4220 - 0x107c  :    0 - 0x0
    "00000000", -- 4221 - 0x107d  :    0 - 0x0
    "00000000", -- 4222 - 0x107e  :    0 - 0x0
    "00000000", -- 4223 - 0x107f  :    0 - 0x0
    "01111100", -- 4224 - 0x1080  :  124 - 0x7c
    "11000110", -- 4225 - 0x1081  :  198 - 0xc6
    "11000110", -- 4226 - 0x1082  :  198 - 0xc6
    "01111100", -- 4227 - 0x1083  :  124 - 0x7c
    "11000110", -- 4228 - 0x1084  :  198 - 0xc6
    "11000110", -- 4229 - 0x1085  :  198 - 0xc6
    "01111100", -- 4230 - 0x1086  :  124 - 0x7c
    "00000000", -- 4231 - 0x1087  :    0 - 0x0
    "00000000", -- 4232 - 0x1088  :    0 - 0x0
    "00000000", -- 4233 - 0x1089  :    0 - 0x0
    "00000000", -- 4234 - 0x108a  :    0 - 0x0
    "00000000", -- 4235 - 0x108b  :    0 - 0x0
    "00000000", -- 4236 - 0x108c  :    0 - 0x0
    "00000000", -- 4237 - 0x108d  :    0 - 0x0
    "00000000", -- 4238 - 0x108e  :    0 - 0x0
    "00000000", -- 4239 - 0x108f  :    0 - 0x0
    "01111100", -- 4240 - 0x1090  :  124 - 0x7c
    "11000110", -- 4241 - 0x1091  :  198 - 0xc6
    "11000110", -- 4242 - 0x1092  :  198 - 0xc6
    "01111110", -- 4243 - 0x1093  :  126 - 0x7e
    "00000110", -- 4244 - 0x1094  :    6 - 0x6
    "00001100", -- 4245 - 0x1095  :   12 - 0xc
    "01111000", -- 4246 - 0x1096  :  120 - 0x78
    "00000000", -- 4247 - 0x1097  :    0 - 0x0
    "00000000", -- 4248 - 0x1098  :    0 - 0x0
    "00000000", -- 4249 - 0x1099  :    0 - 0x0
    "00000000", -- 4250 - 0x109a  :    0 - 0x0
    "00000000", -- 4251 - 0x109b  :    0 - 0x0
    "00000000", -- 4252 - 0x109c  :    0 - 0x0
    "00000000", -- 4253 - 0x109d  :    0 - 0x0
    "00000000", -- 4254 - 0x109e  :    0 - 0x0
    "00000000", -- 4255 - 0x109f  :    0 - 0x0
    "00111000", -- 4256 - 0x10a0  :   56 - 0x38
    "01101100", -- 4257 - 0x10a1  :  108 - 0x6c
    "11000110", -- 4258 - 0x10a2  :  198 - 0xc6
    "11000110", -- 4259 - 0x10a3  :  198 - 0xc6
    "11111110", -- 4260 - 0x10a4  :  254 - 0xfe
    "11000110", -- 4261 - 0x10a5  :  198 - 0xc6
    "11000110", -- 4262 - 0x10a6  :  198 - 0xc6
    "00000000", -- 4263 - 0x10a7  :    0 - 0x0
    "00000000", -- 4264 - 0x10a8  :    0 - 0x0
    "00000000", -- 4265 - 0x10a9  :    0 - 0x0
    "00000000", -- 4266 - 0x10aa  :    0 - 0x0
    "00000000", -- 4267 - 0x10ab  :    0 - 0x0
    "00000000", -- 4268 - 0x10ac  :    0 - 0x0
    "00000000", -- 4269 - 0x10ad  :    0 - 0x0
    "00000000", -- 4270 - 0x10ae  :    0 - 0x0
    "00000000", -- 4271 - 0x10af  :    0 - 0x0
    "11111100", -- 4272 - 0x10b0  :  252 - 0xfc
    "11000110", -- 4273 - 0x10b1  :  198 - 0xc6
    "11000110", -- 4274 - 0x10b2  :  198 - 0xc6
    "11111100", -- 4275 - 0x10b3  :  252 - 0xfc
    "11000110", -- 4276 - 0x10b4  :  198 - 0xc6
    "11000110", -- 4277 - 0x10b5  :  198 - 0xc6
    "11111100", -- 4278 - 0x10b6  :  252 - 0xfc
    "00000000", -- 4279 - 0x10b7  :    0 - 0x0
    "00000000", -- 4280 - 0x10b8  :    0 - 0x0
    "00000000", -- 4281 - 0x10b9  :    0 - 0x0
    "00000000", -- 4282 - 0x10ba  :    0 - 0x0
    "00000000", -- 4283 - 0x10bb  :    0 - 0x0
    "00000000", -- 4284 - 0x10bc  :    0 - 0x0
    "00000000", -- 4285 - 0x10bd  :    0 - 0x0
    "00000000", -- 4286 - 0x10be  :    0 - 0x0
    "00000000", -- 4287 - 0x10bf  :    0 - 0x0
    "00111100", -- 4288 - 0x10c0  :   60 - 0x3c
    "01100110", -- 4289 - 0x10c1  :  102 - 0x66
    "11000000", -- 4290 - 0x10c2  :  192 - 0xc0
    "11000000", -- 4291 - 0x10c3  :  192 - 0xc0
    "11000000", -- 4292 - 0x10c4  :  192 - 0xc0
    "01100110", -- 4293 - 0x10c5  :  102 - 0x66
    "00111100", -- 4294 - 0x10c6  :   60 - 0x3c
    "00000000", -- 4295 - 0x10c7  :    0 - 0x0
    "00000000", -- 4296 - 0x10c8  :    0 - 0x0
    "00000000", -- 4297 - 0x10c9  :    0 - 0x0
    "00000000", -- 4298 - 0x10ca  :    0 - 0x0
    "00000000", -- 4299 - 0x10cb  :    0 - 0x0
    "00000000", -- 4300 - 0x10cc  :    0 - 0x0
    "00000000", -- 4301 - 0x10cd  :    0 - 0x0
    "00000000", -- 4302 - 0x10ce  :    0 - 0x0
    "00000000", -- 4303 - 0x10cf  :    0 - 0x0
    "11111000", -- 4304 - 0x10d0  :  248 - 0xf8
    "11001100", -- 4305 - 0x10d1  :  204 - 0xcc
    "11000110", -- 4306 - 0x10d2  :  198 - 0xc6
    "11000110", -- 4307 - 0x10d3  :  198 - 0xc6
    "11000110", -- 4308 - 0x10d4  :  198 - 0xc6
    "11001100", -- 4309 - 0x10d5  :  204 - 0xcc
    "11111000", -- 4310 - 0x10d6  :  248 - 0xf8
    "00000000", -- 4311 - 0x10d7  :    0 - 0x0
    "00000000", -- 4312 - 0x10d8  :    0 - 0x0
    "00000000", -- 4313 - 0x10d9  :    0 - 0x0
    "00000000", -- 4314 - 0x10da  :    0 - 0x0
    "00000000", -- 4315 - 0x10db  :    0 - 0x0
    "00000000", -- 4316 - 0x10dc  :    0 - 0x0
    "00000000", -- 4317 - 0x10dd  :    0 - 0x0
    "00000000", -- 4318 - 0x10de  :    0 - 0x0
    "00000000", -- 4319 - 0x10df  :    0 - 0x0
    "11111110", -- 4320 - 0x10e0  :  254 - 0xfe
    "11000000", -- 4321 - 0x10e1  :  192 - 0xc0
    "11000000", -- 4322 - 0x10e2  :  192 - 0xc0
    "11111100", -- 4323 - 0x10e3  :  252 - 0xfc
    "11000000", -- 4324 - 0x10e4  :  192 - 0xc0
    "11000000", -- 4325 - 0x10e5  :  192 - 0xc0
    "11111110", -- 4326 - 0x10e6  :  254 - 0xfe
    "00000000", -- 4327 - 0x10e7  :    0 - 0x0
    "00000000", -- 4328 - 0x10e8  :    0 - 0x0
    "00000000", -- 4329 - 0x10e9  :    0 - 0x0
    "00000000", -- 4330 - 0x10ea  :    0 - 0x0
    "00000000", -- 4331 - 0x10eb  :    0 - 0x0
    "00000000", -- 4332 - 0x10ec  :    0 - 0x0
    "00000000", -- 4333 - 0x10ed  :    0 - 0x0
    "00000000", -- 4334 - 0x10ee  :    0 - 0x0
    "00000000", -- 4335 - 0x10ef  :    0 - 0x0
    "11111110", -- 4336 - 0x10f0  :  254 - 0xfe
    "11000000", -- 4337 - 0x10f1  :  192 - 0xc0
    "11000000", -- 4338 - 0x10f2  :  192 - 0xc0
    "11111100", -- 4339 - 0x10f3  :  252 - 0xfc
    "11000000", -- 4340 - 0x10f4  :  192 - 0xc0
    "11000000", -- 4341 - 0x10f5  :  192 - 0xc0
    "11000000", -- 4342 - 0x10f6  :  192 - 0xc0
    "00000000", -- 4343 - 0x10f7  :    0 - 0x0
    "00000000", -- 4344 - 0x10f8  :    0 - 0x0
    "00000000", -- 4345 - 0x10f9  :    0 - 0x0
    "00000000", -- 4346 - 0x10fa  :    0 - 0x0
    "00000000", -- 4347 - 0x10fb  :    0 - 0x0
    "00000000", -- 4348 - 0x10fc  :    0 - 0x0
    "00000000", -- 4349 - 0x10fd  :    0 - 0x0
    "00000000", -- 4350 - 0x10fe  :    0 - 0x0
    "00000000", -- 4351 - 0x10ff  :    0 - 0x0
    "00111110", -- 4352 - 0x1100  :   62 - 0x3e
    "01100000", -- 4353 - 0x1101  :   96 - 0x60
    "11000000", -- 4354 - 0x1102  :  192 - 0xc0
    "11001110", -- 4355 - 0x1103  :  206 - 0xce
    "11000110", -- 4356 - 0x1104  :  198 - 0xc6
    "01100110", -- 4357 - 0x1105  :  102 - 0x66
    "00111110", -- 4358 - 0x1106  :   62 - 0x3e
    "00000000", -- 4359 - 0x1107  :    0 - 0x0
    "00000000", -- 4360 - 0x1108  :    0 - 0x0
    "00000000", -- 4361 - 0x1109  :    0 - 0x0
    "00000000", -- 4362 - 0x110a  :    0 - 0x0
    "00000000", -- 4363 - 0x110b  :    0 - 0x0
    "00000000", -- 4364 - 0x110c  :    0 - 0x0
    "00000000", -- 4365 - 0x110d  :    0 - 0x0
    "00000000", -- 4366 - 0x110e  :    0 - 0x0
    "00000000", -- 4367 - 0x110f  :    0 - 0x0
    "11000110", -- 4368 - 0x1110  :  198 - 0xc6
    "11000110", -- 4369 - 0x1111  :  198 - 0xc6
    "11000110", -- 4370 - 0x1112  :  198 - 0xc6
    "11111110", -- 4371 - 0x1113  :  254 - 0xfe
    "11000110", -- 4372 - 0x1114  :  198 - 0xc6
    "11000110", -- 4373 - 0x1115  :  198 - 0xc6
    "11000110", -- 4374 - 0x1116  :  198 - 0xc6
    "00000000", -- 4375 - 0x1117  :    0 - 0x0
    "00000000", -- 4376 - 0x1118  :    0 - 0x0
    "00000000", -- 4377 - 0x1119  :    0 - 0x0
    "00000000", -- 4378 - 0x111a  :    0 - 0x0
    "00000000", -- 4379 - 0x111b  :    0 - 0x0
    "00000000", -- 4380 - 0x111c  :    0 - 0x0
    "00000000", -- 4381 - 0x111d  :    0 - 0x0
    "00000000", -- 4382 - 0x111e  :    0 - 0x0
    "00000000", -- 4383 - 0x111f  :    0 - 0x0
    "01111110", -- 4384 - 0x1120  :  126 - 0x7e
    "00011000", -- 4385 - 0x1121  :   24 - 0x18
    "00011000", -- 4386 - 0x1122  :   24 - 0x18
    "00011000", -- 4387 - 0x1123  :   24 - 0x18
    "00011000", -- 4388 - 0x1124  :   24 - 0x18
    "00011000", -- 4389 - 0x1125  :   24 - 0x18
    "01111110", -- 4390 - 0x1126  :  126 - 0x7e
    "00000000", -- 4391 - 0x1127  :    0 - 0x0
    "00000000", -- 4392 - 0x1128  :    0 - 0x0
    "00000000", -- 4393 - 0x1129  :    0 - 0x0
    "00000000", -- 4394 - 0x112a  :    0 - 0x0
    "00000000", -- 4395 - 0x112b  :    0 - 0x0
    "00000000", -- 4396 - 0x112c  :    0 - 0x0
    "00000000", -- 4397 - 0x112d  :    0 - 0x0
    "00000000", -- 4398 - 0x112e  :    0 - 0x0
    "00000000", -- 4399 - 0x112f  :    0 - 0x0
    "00011110", -- 4400 - 0x1130  :   30 - 0x1e
    "00000110", -- 4401 - 0x1131  :    6 - 0x6
    "00000110", -- 4402 - 0x1132  :    6 - 0x6
    "00000110", -- 4403 - 0x1133  :    6 - 0x6
    "11000110", -- 4404 - 0x1134  :  198 - 0xc6
    "11000110", -- 4405 - 0x1135  :  198 - 0xc6
    "01111100", -- 4406 - 0x1136  :  124 - 0x7c
    "00000000", -- 4407 - 0x1137  :    0 - 0x0
    "00000000", -- 4408 - 0x1138  :    0 - 0x0
    "00000000", -- 4409 - 0x1139  :    0 - 0x0
    "00000000", -- 4410 - 0x113a  :    0 - 0x0
    "00000000", -- 4411 - 0x113b  :    0 - 0x0
    "00000000", -- 4412 - 0x113c  :    0 - 0x0
    "00000000", -- 4413 - 0x113d  :    0 - 0x0
    "00000000", -- 4414 - 0x113e  :    0 - 0x0
    "00000000", -- 4415 - 0x113f  :    0 - 0x0
    "11000110", -- 4416 - 0x1140  :  198 - 0xc6
    "11001100", -- 4417 - 0x1141  :  204 - 0xcc
    "11011000", -- 4418 - 0x1142  :  216 - 0xd8
    "11110000", -- 4419 - 0x1143  :  240 - 0xf0
    "11111000", -- 4420 - 0x1144  :  248 - 0xf8
    "11011100", -- 4421 - 0x1145  :  220 - 0xdc
    "11001110", -- 4422 - 0x1146  :  206 - 0xce
    "00000000", -- 4423 - 0x1147  :    0 - 0x0
    "00000000", -- 4424 - 0x1148  :    0 - 0x0
    "00000000", -- 4425 - 0x1149  :    0 - 0x0
    "00000000", -- 4426 - 0x114a  :    0 - 0x0
    "00000000", -- 4427 - 0x114b  :    0 - 0x0
    "00000000", -- 4428 - 0x114c  :    0 - 0x0
    "00000000", -- 4429 - 0x114d  :    0 - 0x0
    "00000000", -- 4430 - 0x114e  :    0 - 0x0
    "00000000", -- 4431 - 0x114f  :    0 - 0x0
    "01100000", -- 4432 - 0x1150  :   96 - 0x60
    "01100000", -- 4433 - 0x1151  :   96 - 0x60
    "01100000", -- 4434 - 0x1152  :   96 - 0x60
    "01100000", -- 4435 - 0x1153  :   96 - 0x60
    "01100000", -- 4436 - 0x1154  :   96 - 0x60
    "01100000", -- 4437 - 0x1155  :   96 - 0x60
    "01111110", -- 4438 - 0x1156  :  126 - 0x7e
    "00000000", -- 4439 - 0x1157  :    0 - 0x0
    "00000000", -- 4440 - 0x1158  :    0 - 0x0
    "00000000", -- 4441 - 0x1159  :    0 - 0x0
    "00000000", -- 4442 - 0x115a  :    0 - 0x0
    "00000000", -- 4443 - 0x115b  :    0 - 0x0
    "00000000", -- 4444 - 0x115c  :    0 - 0x0
    "00000000", -- 4445 - 0x115d  :    0 - 0x0
    "00000000", -- 4446 - 0x115e  :    0 - 0x0
    "00000000", -- 4447 - 0x115f  :    0 - 0x0
    "11000110", -- 4448 - 0x1160  :  198 - 0xc6
    "11101110", -- 4449 - 0x1161  :  238 - 0xee
    "11111110", -- 4450 - 0x1162  :  254 - 0xfe
    "11111110", -- 4451 - 0x1163  :  254 - 0xfe
    "11010110", -- 4452 - 0x1164  :  214 - 0xd6
    "11000110", -- 4453 - 0x1165  :  198 - 0xc6
    "11000110", -- 4454 - 0x1166  :  198 - 0xc6
    "00000000", -- 4455 - 0x1167  :    0 - 0x0
    "00000000", -- 4456 - 0x1168  :    0 - 0x0
    "00000000", -- 4457 - 0x1169  :    0 - 0x0
    "00000000", -- 4458 - 0x116a  :    0 - 0x0
    "00000000", -- 4459 - 0x116b  :    0 - 0x0
    "00000000", -- 4460 - 0x116c  :    0 - 0x0
    "00000000", -- 4461 - 0x116d  :    0 - 0x0
    "00000000", -- 4462 - 0x116e  :    0 - 0x0
    "00000000", -- 4463 - 0x116f  :    0 - 0x0
    "11000110", -- 4464 - 0x1170  :  198 - 0xc6
    "11100110", -- 4465 - 0x1171  :  230 - 0xe6
    "11110110", -- 4466 - 0x1172  :  246 - 0xf6
    "11111110", -- 4467 - 0x1173  :  254 - 0xfe
    "11011110", -- 4468 - 0x1174  :  222 - 0xde
    "11001110", -- 4469 - 0x1175  :  206 - 0xce
    "11000110", -- 4470 - 0x1176  :  198 - 0xc6
    "00000000", -- 4471 - 0x1177  :    0 - 0x0
    "00000000", -- 4472 - 0x1178  :    0 - 0x0
    "00000000", -- 4473 - 0x1179  :    0 - 0x0
    "00000000", -- 4474 - 0x117a  :    0 - 0x0
    "00000000", -- 4475 - 0x117b  :    0 - 0x0
    "00000000", -- 4476 - 0x117c  :    0 - 0x0
    "00000000", -- 4477 - 0x117d  :    0 - 0x0
    "00000000", -- 4478 - 0x117e  :    0 - 0x0
    "00000000", -- 4479 - 0x117f  :    0 - 0x0
    "01111100", -- 4480 - 0x1180  :  124 - 0x7c
    "11000110", -- 4481 - 0x1181  :  198 - 0xc6
    "11000110", -- 4482 - 0x1182  :  198 - 0xc6
    "11000110", -- 4483 - 0x1183  :  198 - 0xc6
    "11000110", -- 4484 - 0x1184  :  198 - 0xc6
    "11000110", -- 4485 - 0x1185  :  198 - 0xc6
    "01111100", -- 4486 - 0x1186  :  124 - 0x7c
    "00000000", -- 4487 - 0x1187  :    0 - 0x0
    "00000000", -- 4488 - 0x1188  :    0 - 0x0
    "00000000", -- 4489 - 0x1189  :    0 - 0x0
    "00000000", -- 4490 - 0x118a  :    0 - 0x0
    "00000000", -- 4491 - 0x118b  :    0 - 0x0
    "00000000", -- 4492 - 0x118c  :    0 - 0x0
    "00000000", -- 4493 - 0x118d  :    0 - 0x0
    "00000000", -- 4494 - 0x118e  :    0 - 0x0
    "00000000", -- 4495 - 0x118f  :    0 - 0x0
    "11111100", -- 4496 - 0x1190  :  252 - 0xfc
    "11000110", -- 4497 - 0x1191  :  198 - 0xc6
    "11000110", -- 4498 - 0x1192  :  198 - 0xc6
    "11000110", -- 4499 - 0x1193  :  198 - 0xc6
    "11111100", -- 4500 - 0x1194  :  252 - 0xfc
    "11000000", -- 4501 - 0x1195  :  192 - 0xc0
    "11000000", -- 4502 - 0x1196  :  192 - 0xc0
    "00000000", -- 4503 - 0x1197  :    0 - 0x0
    "00000000", -- 4504 - 0x1198  :    0 - 0x0
    "00000000", -- 4505 - 0x1199  :    0 - 0x0
    "00000000", -- 4506 - 0x119a  :    0 - 0x0
    "00000000", -- 4507 - 0x119b  :    0 - 0x0
    "00000000", -- 4508 - 0x119c  :    0 - 0x0
    "00000000", -- 4509 - 0x119d  :    0 - 0x0
    "00000000", -- 4510 - 0x119e  :    0 - 0x0
    "00000000", -- 4511 - 0x119f  :    0 - 0x0
    "01111100", -- 4512 - 0x11a0  :  124 - 0x7c
    "11000110", -- 4513 - 0x11a1  :  198 - 0xc6
    "11000110", -- 4514 - 0x11a2  :  198 - 0xc6
    "11000110", -- 4515 - 0x11a3  :  198 - 0xc6
    "11011110", -- 4516 - 0x11a4  :  222 - 0xde
    "11001100", -- 4517 - 0x11a5  :  204 - 0xcc
    "01111010", -- 4518 - 0x11a6  :  122 - 0x7a
    "00000000", -- 4519 - 0x11a7  :    0 - 0x0
    "00000000", -- 4520 - 0x11a8  :    0 - 0x0
    "00000000", -- 4521 - 0x11a9  :    0 - 0x0
    "00000000", -- 4522 - 0x11aa  :    0 - 0x0
    "00000000", -- 4523 - 0x11ab  :    0 - 0x0
    "00000000", -- 4524 - 0x11ac  :    0 - 0x0
    "00000000", -- 4525 - 0x11ad  :    0 - 0x0
    "00000000", -- 4526 - 0x11ae  :    0 - 0x0
    "00000000", -- 4527 - 0x11af  :    0 - 0x0
    "11111100", -- 4528 - 0x11b0  :  252 - 0xfc
    "11000110", -- 4529 - 0x11b1  :  198 - 0xc6
    "11000110", -- 4530 - 0x11b2  :  198 - 0xc6
    "11001110", -- 4531 - 0x11b3  :  206 - 0xce
    "11111000", -- 4532 - 0x11b4  :  248 - 0xf8
    "11011100", -- 4533 - 0x11b5  :  220 - 0xdc
    "11001110", -- 4534 - 0x11b6  :  206 - 0xce
    "00000000", -- 4535 - 0x11b7  :    0 - 0x0
    "00000000", -- 4536 - 0x11b8  :    0 - 0x0
    "00000000", -- 4537 - 0x11b9  :    0 - 0x0
    "00000000", -- 4538 - 0x11ba  :    0 - 0x0
    "00000000", -- 4539 - 0x11bb  :    0 - 0x0
    "00000000", -- 4540 - 0x11bc  :    0 - 0x0
    "00000000", -- 4541 - 0x11bd  :    0 - 0x0
    "00000000", -- 4542 - 0x11be  :    0 - 0x0
    "00000000", -- 4543 - 0x11bf  :    0 - 0x0
    "01111000", -- 4544 - 0x11c0  :  120 - 0x78
    "11001100", -- 4545 - 0x11c1  :  204 - 0xcc
    "11000000", -- 4546 - 0x11c2  :  192 - 0xc0
    "01111100", -- 4547 - 0x11c3  :  124 - 0x7c
    "00000110", -- 4548 - 0x11c4  :    6 - 0x6
    "11000110", -- 4549 - 0x11c5  :  198 - 0xc6
    "01111100", -- 4550 - 0x11c6  :  124 - 0x7c
    "00000000", -- 4551 - 0x11c7  :    0 - 0x0
    "00000000", -- 4552 - 0x11c8  :    0 - 0x0
    "00000000", -- 4553 - 0x11c9  :    0 - 0x0
    "00000000", -- 4554 - 0x11ca  :    0 - 0x0
    "00000000", -- 4555 - 0x11cb  :    0 - 0x0
    "00000000", -- 4556 - 0x11cc  :    0 - 0x0
    "00000000", -- 4557 - 0x11cd  :    0 - 0x0
    "00000000", -- 4558 - 0x11ce  :    0 - 0x0
    "00000000", -- 4559 - 0x11cf  :    0 - 0x0
    "01111110", -- 4560 - 0x11d0  :  126 - 0x7e
    "00011000", -- 4561 - 0x11d1  :   24 - 0x18
    "00011000", -- 4562 - 0x11d2  :   24 - 0x18
    "00011000", -- 4563 - 0x11d3  :   24 - 0x18
    "00011000", -- 4564 - 0x11d4  :   24 - 0x18
    "00011000", -- 4565 - 0x11d5  :   24 - 0x18
    "00011000", -- 4566 - 0x11d6  :   24 - 0x18
    "00000000", -- 4567 - 0x11d7  :    0 - 0x0
    "00000000", -- 4568 - 0x11d8  :    0 - 0x0
    "00000000", -- 4569 - 0x11d9  :    0 - 0x0
    "00000000", -- 4570 - 0x11da  :    0 - 0x0
    "00000000", -- 4571 - 0x11db  :    0 - 0x0
    "00000000", -- 4572 - 0x11dc  :    0 - 0x0
    "00000000", -- 4573 - 0x11dd  :    0 - 0x0
    "00000000", -- 4574 - 0x11de  :    0 - 0x0
    "00000000", -- 4575 - 0x11df  :    0 - 0x0
    "11000110", -- 4576 - 0x11e0  :  198 - 0xc6
    "11000110", -- 4577 - 0x11e1  :  198 - 0xc6
    "11000110", -- 4578 - 0x11e2  :  198 - 0xc6
    "11000110", -- 4579 - 0x11e3  :  198 - 0xc6
    "11000110", -- 4580 - 0x11e4  :  198 - 0xc6
    "11000110", -- 4581 - 0x11e5  :  198 - 0xc6
    "01111100", -- 4582 - 0x11e6  :  124 - 0x7c
    "00000000", -- 4583 - 0x11e7  :    0 - 0x0
    "00000000", -- 4584 - 0x11e8  :    0 - 0x0
    "00000000", -- 4585 - 0x11e9  :    0 - 0x0
    "00000000", -- 4586 - 0x11ea  :    0 - 0x0
    "00000000", -- 4587 - 0x11eb  :    0 - 0x0
    "00000000", -- 4588 - 0x11ec  :    0 - 0x0
    "00000000", -- 4589 - 0x11ed  :    0 - 0x0
    "00000000", -- 4590 - 0x11ee  :    0 - 0x0
    "00000000", -- 4591 - 0x11ef  :    0 - 0x0
    "11000110", -- 4592 - 0x11f0  :  198 - 0xc6
    "11000110", -- 4593 - 0x11f1  :  198 - 0xc6
    "11000110", -- 4594 - 0x11f2  :  198 - 0xc6
    "11101110", -- 4595 - 0x11f3  :  238 - 0xee
    "01111100", -- 4596 - 0x11f4  :  124 - 0x7c
    "00111000", -- 4597 - 0x11f5  :   56 - 0x38
    "00010000", -- 4598 - 0x11f6  :   16 - 0x10
    "00000000", -- 4599 - 0x11f7  :    0 - 0x0
    "00000000", -- 4600 - 0x11f8  :    0 - 0x0
    "00000000", -- 4601 - 0x11f9  :    0 - 0x0
    "00000000", -- 4602 - 0x11fa  :    0 - 0x0
    "00000000", -- 4603 - 0x11fb  :    0 - 0x0
    "00000000", -- 4604 - 0x11fc  :    0 - 0x0
    "00000000", -- 4605 - 0x11fd  :    0 - 0x0
    "00000000", -- 4606 - 0x11fe  :    0 - 0x0
    "00000000", -- 4607 - 0x11ff  :    0 - 0x0
    "11000110", -- 4608 - 0x1200  :  198 - 0xc6
    "11000110", -- 4609 - 0x1201  :  198 - 0xc6
    "11010110", -- 4610 - 0x1202  :  214 - 0xd6
    "11111110", -- 4611 - 0x1203  :  254 - 0xfe
    "11111110", -- 4612 - 0x1204  :  254 - 0xfe
    "11101110", -- 4613 - 0x1205  :  238 - 0xee
    "11000110", -- 4614 - 0x1206  :  198 - 0xc6
    "00000000", -- 4615 - 0x1207  :    0 - 0x0
    "00000000", -- 4616 - 0x1208  :    0 - 0x0
    "00000000", -- 4617 - 0x1209  :    0 - 0x0
    "00000000", -- 4618 - 0x120a  :    0 - 0x0
    "00000000", -- 4619 - 0x120b  :    0 - 0x0
    "00000000", -- 4620 - 0x120c  :    0 - 0x0
    "00000000", -- 4621 - 0x120d  :    0 - 0x0
    "00000000", -- 4622 - 0x120e  :    0 - 0x0
    "00000000", -- 4623 - 0x120f  :    0 - 0x0
    "11000110", -- 4624 - 0x1210  :  198 - 0xc6
    "11101110", -- 4625 - 0x1211  :  238 - 0xee
    "01111100", -- 4626 - 0x1212  :  124 - 0x7c
    "00111000", -- 4627 - 0x1213  :   56 - 0x38
    "01111100", -- 4628 - 0x1214  :  124 - 0x7c
    "11101110", -- 4629 - 0x1215  :  238 - 0xee
    "11000110", -- 4630 - 0x1216  :  198 - 0xc6
    "00000000", -- 4631 - 0x1217  :    0 - 0x0
    "00000000", -- 4632 - 0x1218  :    0 - 0x0
    "00000000", -- 4633 - 0x1219  :    0 - 0x0
    "00000000", -- 4634 - 0x121a  :    0 - 0x0
    "00000000", -- 4635 - 0x121b  :    0 - 0x0
    "00000000", -- 4636 - 0x121c  :    0 - 0x0
    "00000000", -- 4637 - 0x121d  :    0 - 0x0
    "00000000", -- 4638 - 0x121e  :    0 - 0x0
    "00000000", -- 4639 - 0x121f  :    0 - 0x0
    "01100110", -- 4640 - 0x1220  :  102 - 0x66
    "01100110", -- 4641 - 0x1221  :  102 - 0x66
    "01100110", -- 4642 - 0x1222  :  102 - 0x66
    "00111100", -- 4643 - 0x1223  :   60 - 0x3c
    "00011000", -- 4644 - 0x1224  :   24 - 0x18
    "00011000", -- 4645 - 0x1225  :   24 - 0x18
    "00011000", -- 4646 - 0x1226  :   24 - 0x18
    "00000000", -- 4647 - 0x1227  :    0 - 0x0
    "00000000", -- 4648 - 0x1228  :    0 - 0x0
    "00000000", -- 4649 - 0x1229  :    0 - 0x0
    "00000000", -- 4650 - 0x122a  :    0 - 0x0
    "00000000", -- 4651 - 0x122b  :    0 - 0x0
    "00000000", -- 4652 - 0x122c  :    0 - 0x0
    "00000000", -- 4653 - 0x122d  :    0 - 0x0
    "00000000", -- 4654 - 0x122e  :    0 - 0x0
    "00000000", -- 4655 - 0x122f  :    0 - 0x0
    "11111110", -- 4656 - 0x1230  :  254 - 0xfe
    "00001110", -- 4657 - 0x1231  :   14 - 0xe
    "00011100", -- 4658 - 0x1232  :   28 - 0x1c
    "00111000", -- 4659 - 0x1233  :   56 - 0x38
    "01110000", -- 4660 - 0x1234  :  112 - 0x70
    "11100000", -- 4661 - 0x1235  :  224 - 0xe0
    "11111110", -- 4662 - 0x1236  :  254 - 0xfe
    "00000000", -- 4663 - 0x1237  :    0 - 0x0
    "00000000", -- 4664 - 0x1238  :    0 - 0x0
    "00000000", -- 4665 - 0x1239  :    0 - 0x0
    "00000000", -- 4666 - 0x123a  :    0 - 0x0
    "00000000", -- 4667 - 0x123b  :    0 - 0x0
    "00000000", -- 4668 - 0x123c  :    0 - 0x0
    "00000000", -- 4669 - 0x123d  :    0 - 0x0
    "00000000", -- 4670 - 0x123e  :    0 - 0x0
    "00000000", -- 4671 - 0x123f  :    0 - 0x0
    "00000000", -- 4672 - 0x1240  :    0 - 0x0
    "00000000", -- 4673 - 0x1241  :    0 - 0x0
    "00000000", -- 4674 - 0x1242  :    0 - 0x0
    "00000000", -- 4675 - 0x1243  :    0 - 0x0
    "00000000", -- 4676 - 0x1244  :    0 - 0x0
    "00000000", -- 4677 - 0x1245  :    0 - 0x0
    "00000000", -- 4678 - 0x1246  :    0 - 0x0
    "00000000", -- 4679 - 0x1247  :    0 - 0x0
    "00000000", -- 4680 - 0x1248  :    0 - 0x0
    "00000000", -- 4681 - 0x1249  :    0 - 0x0
    "00000000", -- 4682 - 0x124a  :    0 - 0x0
    "00000000", -- 4683 - 0x124b  :    0 - 0x0
    "00000000", -- 4684 - 0x124c  :    0 - 0x0
    "00000000", -- 4685 - 0x124d  :    0 - 0x0
    "00000000", -- 4686 - 0x124e  :    0 - 0x0
    "00000000", -- 4687 - 0x124f  :    0 - 0x0
    "11111111", -- 4688 - 0x1250  :  255 - 0xff
    "11111111", -- 4689 - 0x1251  :  255 - 0xff
    "11111111", -- 4690 - 0x1252  :  255 - 0xff
    "11111111", -- 4691 - 0x1253  :  255 - 0xff
    "11111111", -- 4692 - 0x1254  :  255 - 0xff
    "11111111", -- 4693 - 0x1255  :  255 - 0xff
    "11111111", -- 4694 - 0x1256  :  255 - 0xff
    "11111111", -- 4695 - 0x1257  :  255 - 0xff
    "00000000", -- 4696 - 0x1258  :    0 - 0x0
    "00000000", -- 4697 - 0x1259  :    0 - 0x0
    "00000000", -- 4698 - 0x125a  :    0 - 0x0
    "00000000", -- 4699 - 0x125b  :    0 - 0x0
    "00000000", -- 4700 - 0x125c  :    0 - 0x0
    "00000000", -- 4701 - 0x125d  :    0 - 0x0
    "00000000", -- 4702 - 0x125e  :    0 - 0x0
    "00000000", -- 4703 - 0x125f  :    0 - 0x0
    "00000000", -- 4704 - 0x1260  :    0 - 0x0
    "00000000", -- 4705 - 0x1261  :    0 - 0x0
    "00000000", -- 4706 - 0x1262  :    0 - 0x0
    "00000000", -- 4707 - 0x1263  :    0 - 0x0
    "00000000", -- 4708 - 0x1264  :    0 - 0x0
    "00000000", -- 4709 - 0x1265  :    0 - 0x0
    "00000000", -- 4710 - 0x1266  :    0 - 0x0
    "00000000", -- 4711 - 0x1267  :    0 - 0x0
    "11111111", -- 4712 - 0x1268  :  255 - 0xff
    "11111111", -- 4713 - 0x1269  :  255 - 0xff
    "11111111", -- 4714 - 0x126a  :  255 - 0xff
    "11111111", -- 4715 - 0x126b  :  255 - 0xff
    "11111111", -- 4716 - 0x126c  :  255 - 0xff
    "11111111", -- 4717 - 0x126d  :  255 - 0xff
    "11111111", -- 4718 - 0x126e  :  255 - 0xff
    "11111111", -- 4719 - 0x126f  :  255 - 0xff
    "11111111", -- 4720 - 0x1270  :  255 - 0xff
    "11111111", -- 4721 - 0x1271  :  255 - 0xff
    "11111111", -- 4722 - 0x1272  :  255 - 0xff
    "11111111", -- 4723 - 0x1273  :  255 - 0xff
    "11111111", -- 4724 - 0x1274  :  255 - 0xff
    "11111111", -- 4725 - 0x1275  :  255 - 0xff
    "11111111", -- 4726 - 0x1276  :  255 - 0xff
    "11111111", -- 4727 - 0x1277  :  255 - 0xff
    "11111111", -- 4728 - 0x1278  :  255 - 0xff
    "11111111", -- 4729 - 0x1279  :  255 - 0xff
    "11111111", -- 4730 - 0x127a  :  255 - 0xff
    "11111111", -- 4731 - 0x127b  :  255 - 0xff
    "11111111", -- 4732 - 0x127c  :  255 - 0xff
    "11111111", -- 4733 - 0x127d  :  255 - 0xff
    "11111111", -- 4734 - 0x127e  :  255 - 0xff
    "11111111", -- 4735 - 0x127f  :  255 - 0xff
    "00000000", -- 4736 - 0x1280  :    0 - 0x0
    "00000000", -- 4737 - 0x1281  :    0 - 0x0
    "00000000", -- 4738 - 0x1282  :    0 - 0x0
    "01111110", -- 4739 - 0x1283  :  126 - 0x7e
    "01111110", -- 4740 - 0x1284  :  126 - 0x7e
    "00000000", -- 4741 - 0x1285  :    0 - 0x0
    "00000000", -- 4742 - 0x1286  :    0 - 0x0
    "00000000", -- 4743 - 0x1287  :    0 - 0x0
    "00000000", -- 4744 - 0x1288  :    0 - 0x0
    "00000000", -- 4745 - 0x1289  :    0 - 0x0
    "00000000", -- 4746 - 0x128a  :    0 - 0x0
    "00000000", -- 4747 - 0x128b  :    0 - 0x0
    "00000000", -- 4748 - 0x128c  :    0 - 0x0
    "00000000", -- 4749 - 0x128d  :    0 - 0x0
    "00000000", -- 4750 - 0x128e  :    0 - 0x0
    "00000000", -- 4751 - 0x128f  :    0 - 0x0
    "00000000", -- 4752 - 0x1290  :    0 - 0x0
    "00000000", -- 4753 - 0x1291  :    0 - 0x0
    "01000100", -- 4754 - 0x1292  :   68 - 0x44
    "00101000", -- 4755 - 0x1293  :   40 - 0x28
    "00010000", -- 4756 - 0x1294  :   16 - 0x10
    "00101000", -- 4757 - 0x1295  :   40 - 0x28
    "01000100", -- 4758 - 0x1296  :   68 - 0x44
    "00000000", -- 4759 - 0x1297  :    0 - 0x0
    "00000000", -- 4760 - 0x1298  :    0 - 0x0
    "00000000", -- 4761 - 0x1299  :    0 - 0x0
    "00000000", -- 4762 - 0x129a  :    0 - 0x0
    "00000000", -- 4763 - 0x129b  :    0 - 0x0
    "00000000", -- 4764 - 0x129c  :    0 - 0x0
    "00000000", -- 4765 - 0x129d  :    0 - 0x0
    "00000000", -- 4766 - 0x129e  :    0 - 0x0
    "00000000", -- 4767 - 0x129f  :    0 - 0x0
    "11111111", -- 4768 - 0x12a0  :  255 - 0xff
    "11111111", -- 4769 - 0x12a1  :  255 - 0xff
    "11111111", -- 4770 - 0x12a2  :  255 - 0xff
    "11111111", -- 4771 - 0x12a3  :  255 - 0xff
    "11111111", -- 4772 - 0x12a4  :  255 - 0xff
    "11111111", -- 4773 - 0x12a5  :  255 - 0xff
    "11111111", -- 4774 - 0x12a6  :  255 - 0xff
    "11111111", -- 4775 - 0x12a7  :  255 - 0xff
    "01111111", -- 4776 - 0x12a8  :  127 - 0x7f
    "01111111", -- 4777 - 0x12a9  :  127 - 0x7f
    "01111111", -- 4778 - 0x12aa  :  127 - 0x7f
    "01111111", -- 4779 - 0x12ab  :  127 - 0x7f
    "01111111", -- 4780 - 0x12ac  :  127 - 0x7f
    "01111111", -- 4781 - 0x12ad  :  127 - 0x7f
    "01111111", -- 4782 - 0x12ae  :  127 - 0x7f
    "01111111", -- 4783 - 0x12af  :  127 - 0x7f
    "00011000", -- 4784 - 0x12b0  :   24 - 0x18
    "00111100", -- 4785 - 0x12b1  :   60 - 0x3c
    "00111100", -- 4786 - 0x12b2  :   60 - 0x3c
    "00111100", -- 4787 - 0x12b3  :   60 - 0x3c
    "00011000", -- 4788 - 0x12b4  :   24 - 0x18
    "00011000", -- 4789 - 0x12b5  :   24 - 0x18
    "00000000", -- 4790 - 0x12b6  :    0 - 0x0
    "00011000", -- 4791 - 0x12b7  :   24 - 0x18
    "00000000", -- 4792 - 0x12b8  :    0 - 0x0
    "00000000", -- 4793 - 0x12b9  :    0 - 0x0
    "00000000", -- 4794 - 0x12ba  :    0 - 0x0
    "00000000", -- 4795 - 0x12bb  :    0 - 0x0
    "00000000", -- 4796 - 0x12bc  :    0 - 0x0
    "00000000", -- 4797 - 0x12bd  :    0 - 0x0
    "00000000", -- 4798 - 0x12be  :    0 - 0x0
    "00000000", -- 4799 - 0x12bf  :    0 - 0x0
    "11111111", -- 4800 - 0x12c0  :  255 - 0xff
    "01111111", -- 4801 - 0x12c1  :  127 - 0x7f
    "01111111", -- 4802 - 0x12c2  :  127 - 0x7f
    "01111111", -- 4803 - 0x12c3  :  127 - 0x7f
    "01111111", -- 4804 - 0x12c4  :  127 - 0x7f
    "11111111", -- 4805 - 0x12c5  :  255 - 0xff
    "11100011", -- 4806 - 0x12c6  :  227 - 0xe3
    "11000001", -- 4807 - 0x12c7  :  193 - 0xc1
    "11111111", -- 4808 - 0x12c8  :  255 - 0xff
    "10000000", -- 4809 - 0x12c9  :  128 - 0x80
    "10000000", -- 4810 - 0x12ca  :  128 - 0x80
    "10000000", -- 4811 - 0x12cb  :  128 - 0x80
    "10000000", -- 4812 - 0x12cc  :  128 - 0x80
    "00000000", -- 4813 - 0x12cd  :    0 - 0x0
    "00011100", -- 4814 - 0x12ce  :   28 - 0x1c
    "00111110", -- 4815 - 0x12cf  :   62 - 0x3e
    "10000000", -- 4816 - 0x12d0  :  128 - 0x80
    "10000000", -- 4817 - 0x12d1  :  128 - 0x80
    "10000000", -- 4818 - 0x12d2  :  128 - 0x80
    "11000001", -- 4819 - 0x12d3  :  193 - 0xc1
    "11100011", -- 4820 - 0x12d4  :  227 - 0xe3
    "11111111", -- 4821 - 0x12d5  :  255 - 0xff
    "11111111", -- 4822 - 0x12d6  :  255 - 0xff
    "11111111", -- 4823 - 0x12d7  :  255 - 0xff
    "01111111", -- 4824 - 0x12d8  :  127 - 0x7f
    "01111111", -- 4825 - 0x12d9  :  127 - 0x7f
    "01111111", -- 4826 - 0x12da  :  127 - 0x7f
    "00111110", -- 4827 - 0x12db  :   62 - 0x3e
    "00011100", -- 4828 - 0x12dc  :   28 - 0x1c
    "00000000", -- 4829 - 0x12dd  :    0 - 0x0
    "00000000", -- 4830 - 0x12de  :    0 - 0x0
    "11111111", -- 4831 - 0x12df  :  255 - 0xff
    "00111000", -- 4832 - 0x12e0  :   56 - 0x38
    "01111100", -- 4833 - 0x12e1  :  124 - 0x7c
    "01111100", -- 4834 - 0x12e2  :  124 - 0x7c
    "01111100", -- 4835 - 0x12e3  :  124 - 0x7c
    "01111100", -- 4836 - 0x12e4  :  124 - 0x7c
    "01111100", -- 4837 - 0x12e5  :  124 - 0x7c
    "00111000", -- 4838 - 0x12e6  :   56 - 0x38
    "00000000", -- 4839 - 0x12e7  :    0 - 0x0
    "00001000", -- 4840 - 0x12e8  :    8 - 0x8
    "00000100", -- 4841 - 0x12e9  :    4 - 0x4
    "00000100", -- 4842 - 0x12ea  :    4 - 0x4
    "00000100", -- 4843 - 0x12eb  :    4 - 0x4
    "00000100", -- 4844 - 0x12ec  :    4 - 0x4
    "00000100", -- 4845 - 0x12ed  :    4 - 0x4
    "00001000", -- 4846 - 0x12ee  :    8 - 0x8
    "00000000", -- 4847 - 0x12ef  :    0 - 0x0
    "00000011", -- 4848 - 0x12f0  :    3 - 0x3
    "00000110", -- 4849 - 0x12f1  :    6 - 0x6
    "00001100", -- 4850 - 0x12f2  :   12 - 0xc
    "00001100", -- 4851 - 0x12f3  :   12 - 0xc
    "00001000", -- 4852 - 0x12f4  :    8 - 0x8
    "00001000", -- 4853 - 0x12f5  :    8 - 0x8
    "00000100", -- 4854 - 0x12f6  :    4 - 0x4
    "00000011", -- 4855 - 0x12f7  :    3 - 0x3
    "00000011", -- 4856 - 0x12f8  :    3 - 0x3
    "00000101", -- 4857 - 0x12f9  :    5 - 0x5
    "00001011", -- 4858 - 0x12fa  :   11 - 0xb
    "00001011", -- 4859 - 0x12fb  :   11 - 0xb
    "00001111", -- 4860 - 0x12fc  :   15 - 0xf
    "00001111", -- 4861 - 0x12fd  :   15 - 0xf
    "00000111", -- 4862 - 0x12fe  :    7 - 0x7
    "00000011", -- 4863 - 0x12ff  :    3 - 0x3
    "00000001", -- 4864 - 0x1300  :    1 - 0x1
    "00000010", -- 4865 - 0x1301  :    2 - 0x2
    "00000100", -- 4866 - 0x1302  :    4 - 0x4
    "00001000", -- 4867 - 0x1303  :    8 - 0x8
    "00010000", -- 4868 - 0x1304  :   16 - 0x10
    "00100000", -- 4869 - 0x1305  :   32 - 0x20
    "01000000", -- 4870 - 0x1306  :   64 - 0x40
    "10000000", -- 4871 - 0x1307  :  128 - 0x80
    "00000001", -- 4872 - 0x1308  :    1 - 0x1
    "00000011", -- 4873 - 0x1309  :    3 - 0x3
    "00000111", -- 4874 - 0x130a  :    7 - 0x7
    "00001111", -- 4875 - 0x130b  :   15 - 0xf
    "00011111", -- 4876 - 0x130c  :   31 - 0x1f
    "00111111", -- 4877 - 0x130d  :   63 - 0x3f
    "01111111", -- 4878 - 0x130e  :  127 - 0x7f
    "11111111", -- 4879 - 0x130f  :  255 - 0xff
    "00000000", -- 4880 - 0x1310  :    0 - 0x0
    "00000000", -- 4881 - 0x1311  :    0 - 0x0
    "00000000", -- 4882 - 0x1312  :    0 - 0x0
    "00000000", -- 4883 - 0x1313  :    0 - 0x0
    "00000000", -- 4884 - 0x1314  :    0 - 0x0
    "00000111", -- 4885 - 0x1315  :    7 - 0x7
    "00111000", -- 4886 - 0x1316  :   56 - 0x38
    "11000000", -- 4887 - 0x1317  :  192 - 0xc0
    "00000000", -- 4888 - 0x1318  :    0 - 0x0
    "00000000", -- 4889 - 0x1319  :    0 - 0x0
    "00000000", -- 4890 - 0x131a  :    0 - 0x0
    "00000000", -- 4891 - 0x131b  :    0 - 0x0
    "00000000", -- 4892 - 0x131c  :    0 - 0x0
    "00000111", -- 4893 - 0x131d  :    7 - 0x7
    "00111111", -- 4894 - 0x131e  :   63 - 0x3f
    "11111111", -- 4895 - 0x131f  :  255 - 0xff
    "00000000", -- 4896 - 0x1320  :    0 - 0x0
    "00000000", -- 4897 - 0x1321  :    0 - 0x0
    "00000000", -- 4898 - 0x1322  :    0 - 0x0
    "00000000", -- 4899 - 0x1323  :    0 - 0x0
    "00000000", -- 4900 - 0x1324  :    0 - 0x0
    "11100000", -- 4901 - 0x1325  :  224 - 0xe0
    "00011100", -- 4902 - 0x1326  :   28 - 0x1c
    "00000011", -- 4903 - 0x1327  :    3 - 0x3
    "00000000", -- 4904 - 0x1328  :    0 - 0x0
    "00000000", -- 4905 - 0x1329  :    0 - 0x0
    "00000000", -- 4906 - 0x132a  :    0 - 0x0
    "00000000", -- 4907 - 0x132b  :    0 - 0x0
    "00000000", -- 4908 - 0x132c  :    0 - 0x0
    "11100000", -- 4909 - 0x132d  :  224 - 0xe0
    "11111100", -- 4910 - 0x132e  :  252 - 0xfc
    "11111111", -- 4911 - 0x132f  :  255 - 0xff
    "10000000", -- 4912 - 0x1330  :  128 - 0x80
    "01000000", -- 4913 - 0x1331  :   64 - 0x40
    "00100000", -- 4914 - 0x1332  :   32 - 0x20
    "00010000", -- 4915 - 0x1333  :   16 - 0x10
    "00001000", -- 4916 - 0x1334  :    8 - 0x8
    "00000100", -- 4917 - 0x1335  :    4 - 0x4
    "00000010", -- 4918 - 0x1336  :    2 - 0x2
    "00000001", -- 4919 - 0x1337  :    1 - 0x1
    "10000000", -- 4920 - 0x1338  :  128 - 0x80
    "11000000", -- 4921 - 0x1339  :  192 - 0xc0
    "11100000", -- 4922 - 0x133a  :  224 - 0xe0
    "11110000", -- 4923 - 0x133b  :  240 - 0xf0
    "11111000", -- 4924 - 0x133c  :  248 - 0xf8
    "11111100", -- 4925 - 0x133d  :  252 - 0xfc
    "11111110", -- 4926 - 0x133e  :  254 - 0xfe
    "11111111", -- 4927 - 0x133f  :  255 - 0xff
    "00000100", -- 4928 - 0x1340  :    4 - 0x4
    "00001110", -- 4929 - 0x1341  :   14 - 0xe
    "00001110", -- 4930 - 0x1342  :   14 - 0xe
    "00001110", -- 4931 - 0x1343  :   14 - 0xe
    "01101110", -- 4932 - 0x1344  :  110 - 0x6e
    "01100100", -- 4933 - 0x1345  :  100 - 0x64
    "01100000", -- 4934 - 0x1346  :   96 - 0x60
    "01100000", -- 4935 - 0x1347  :   96 - 0x60
    "11111111", -- 4936 - 0x1348  :  255 - 0xff
    "11111111", -- 4937 - 0x1349  :  255 - 0xff
    "11111111", -- 4938 - 0x134a  :  255 - 0xff
    "11111111", -- 4939 - 0x134b  :  255 - 0xff
    "11111111", -- 4940 - 0x134c  :  255 - 0xff
    "11111111", -- 4941 - 0x134d  :  255 - 0xff
    "11111111", -- 4942 - 0x134e  :  255 - 0xff
    "11111111", -- 4943 - 0x134f  :  255 - 0xff
    "00000111", -- 4944 - 0x1350  :    7 - 0x7
    "00001111", -- 4945 - 0x1351  :   15 - 0xf
    "00011111", -- 4946 - 0x1352  :   31 - 0x1f
    "00011111", -- 4947 - 0x1353  :   31 - 0x1f
    "01111111", -- 4948 - 0x1354  :  127 - 0x7f
    "11111111", -- 4949 - 0x1355  :  255 - 0xff
    "11111111", -- 4950 - 0x1356  :  255 - 0xff
    "01111111", -- 4951 - 0x1357  :  127 - 0x7f
    "00000111", -- 4952 - 0x1358  :    7 - 0x7
    "00001000", -- 4953 - 0x1359  :    8 - 0x8
    "00010000", -- 4954 - 0x135a  :   16 - 0x10
    "00000000", -- 4955 - 0x135b  :    0 - 0x0
    "01100000", -- 4956 - 0x135c  :   96 - 0x60
    "10000000", -- 4957 - 0x135d  :  128 - 0x80
    "10000000", -- 4958 - 0x135e  :  128 - 0x80
    "01000000", -- 4959 - 0x135f  :   64 - 0x40
    "00000011", -- 4960 - 0x1360  :    3 - 0x3
    "00000111", -- 4961 - 0x1361  :    7 - 0x7
    "00011111", -- 4962 - 0x1362  :   31 - 0x1f
    "00111111", -- 4963 - 0x1363  :   63 - 0x3f
    "00111111", -- 4964 - 0x1364  :   63 - 0x3f
    "00111111", -- 4965 - 0x1365  :   63 - 0x3f
    "01111001", -- 4966 - 0x1366  :  121 - 0x79
    "11110111", -- 4967 - 0x1367  :  247 - 0xf7
    "00000011", -- 4968 - 0x1368  :    3 - 0x3
    "00000100", -- 4969 - 0x1369  :    4 - 0x4
    "00011000", -- 4970 - 0x136a  :   24 - 0x18
    "00100000", -- 4971 - 0x136b  :   32 - 0x20
    "00100000", -- 4972 - 0x136c  :   32 - 0x20
    "00100000", -- 4973 - 0x136d  :   32 - 0x20
    "01000110", -- 4974 - 0x136e  :   70 - 0x46
    "10001000", -- 4975 - 0x136f  :  136 - 0x88
    "11000000", -- 4976 - 0x1370  :  192 - 0xc0
    "11100000", -- 4977 - 0x1371  :  224 - 0xe0
    "11110000", -- 4978 - 0x1372  :  240 - 0xf0
    "11110100", -- 4979 - 0x1373  :  244 - 0xf4
    "11111110", -- 4980 - 0x1374  :  254 - 0xfe
    "10111111", -- 4981 - 0x1375  :  191 - 0xbf
    "11011111", -- 4982 - 0x1376  :  223 - 0xdf
    "11111111", -- 4983 - 0x1377  :  255 - 0xff
    "11000000", -- 4984 - 0x1378  :  192 - 0xc0
    "00100000", -- 4985 - 0x1379  :   32 - 0x20
    "00010000", -- 4986 - 0x137a  :   16 - 0x10
    "00010100", -- 4987 - 0x137b  :   20 - 0x14
    "00001010", -- 4988 - 0x137c  :   10 - 0xa
    "01000001", -- 4989 - 0x137d  :   65 - 0x41
    "00100001", -- 4990 - 0x137e  :   33 - 0x21
    "00000001", -- 4991 - 0x137f  :    1 - 0x1
    "10010000", -- 4992 - 0x1380  :  144 - 0x90
    "10111000", -- 4993 - 0x1381  :  184 - 0xb8
    "11111000", -- 4994 - 0x1382  :  248 - 0xf8
    "11111010", -- 4995 - 0x1383  :  250 - 0xfa
    "11111111", -- 4996 - 0x1384  :  255 - 0xff
    "11111111", -- 4997 - 0x1385  :  255 - 0xff
    "11111111", -- 4998 - 0x1386  :  255 - 0xff
    "11111110", -- 4999 - 0x1387  :  254 - 0xfe
    "10010000", -- 5000 - 0x1388  :  144 - 0x90
    "10101000", -- 5001 - 0x1389  :  168 - 0xa8
    "01001000", -- 5002 - 0x138a  :   72 - 0x48
    "00001010", -- 5003 - 0x138b  :   10 - 0xa
    "00000101", -- 5004 - 0x138c  :    5 - 0x5
    "00000001", -- 5005 - 0x138d  :    1 - 0x1
    "00000001", -- 5006 - 0x138e  :    1 - 0x1
    "00000010", -- 5007 - 0x138f  :    2 - 0x2
    "00111011", -- 5008 - 0x1390  :   59 - 0x3b
    "00011101", -- 5009 - 0x1391  :   29 - 0x1d
    "00001110", -- 5010 - 0x1392  :   14 - 0xe
    "00001111", -- 5011 - 0x1393  :   15 - 0xf
    "00000111", -- 5012 - 0x1394  :    7 - 0x7
    "00000000", -- 5013 - 0x1395  :    0 - 0x0
    "00000000", -- 5014 - 0x1396  :    0 - 0x0
    "00000000", -- 5015 - 0x1397  :    0 - 0x0
    "00100100", -- 5016 - 0x1398  :   36 - 0x24
    "00010010", -- 5017 - 0x1399  :   18 - 0x12
    "00001001", -- 5018 - 0x139a  :    9 - 0x9
    "00001000", -- 5019 - 0x139b  :    8 - 0x8
    "00000111", -- 5020 - 0x139c  :    7 - 0x7
    "00000000", -- 5021 - 0x139d  :    0 - 0x0
    "00000000", -- 5022 - 0x139e  :    0 - 0x0
    "00000000", -- 5023 - 0x139f  :    0 - 0x0
    "11111111", -- 5024 - 0x13a0  :  255 - 0xff
    "10111111", -- 5025 - 0x13a1  :  191 - 0xbf
    "00011100", -- 5026 - 0x13a2  :   28 - 0x1c
    "11000000", -- 5027 - 0x13a3  :  192 - 0xc0
    "11110011", -- 5028 - 0x13a4  :  243 - 0xf3
    "11111111", -- 5029 - 0x13a5  :  255 - 0xff
    "01111110", -- 5030 - 0x13a6  :  126 - 0x7e
    "00011100", -- 5031 - 0x13a7  :   28 - 0x1c
    "00000000", -- 5032 - 0x13a8  :    0 - 0x0
    "01000000", -- 5033 - 0x13a9  :   64 - 0x40
    "11100011", -- 5034 - 0x13aa  :  227 - 0xe3
    "00111111", -- 5035 - 0x13ab  :   63 - 0x3f
    "00001100", -- 5036 - 0x13ac  :   12 - 0xc
    "10000001", -- 5037 - 0x13ad  :  129 - 0x81
    "01100010", -- 5038 - 0x13ae  :   98 - 0x62
    "00011100", -- 5039 - 0x13af  :   28 - 0x1c
    "10111111", -- 5040 - 0x13b0  :  191 - 0xbf
    "01111111", -- 5041 - 0x13b1  :  127 - 0x7f
    "00111101", -- 5042 - 0x13b2  :   61 - 0x3d
    "10000011", -- 5043 - 0x13b3  :  131 - 0x83
    "11000111", -- 5044 - 0x13b4  :  199 - 0xc7
    "11111111", -- 5045 - 0x13b5  :  255 - 0xff
    "11111111", -- 5046 - 0x13b6  :  255 - 0xff
    "00111100", -- 5047 - 0x13b7  :   60 - 0x3c
    "01000000", -- 5048 - 0x13b8  :   64 - 0x40
    "10000000", -- 5049 - 0x13b9  :  128 - 0x80
    "11000010", -- 5050 - 0x13ba  :  194 - 0xc2
    "01111100", -- 5051 - 0x13bb  :  124 - 0x7c
    "00111000", -- 5052 - 0x13bc  :   56 - 0x38
    "00000000", -- 5053 - 0x13bd  :    0 - 0x0
    "11000011", -- 5054 - 0x13be  :  195 - 0xc3
    "00111100", -- 5055 - 0x13bf  :   60 - 0x3c
    "11111100", -- 5056 - 0x13c0  :  252 - 0xfc
    "11111110", -- 5057 - 0x13c1  :  254 - 0xfe
    "11111111", -- 5058 - 0x13c2  :  255 - 0xff
    "11111110", -- 5059 - 0x13c3  :  254 - 0xfe
    "11111110", -- 5060 - 0x13c4  :  254 - 0xfe
    "11111000", -- 5061 - 0x13c5  :  248 - 0xf8
    "01100000", -- 5062 - 0x13c6  :   96 - 0x60
    "00000000", -- 5063 - 0x13c7  :    0 - 0x0
    "00000100", -- 5064 - 0x13c8  :    4 - 0x4
    "00000010", -- 5065 - 0x13c9  :    2 - 0x2
    "00000001", -- 5066 - 0x13ca  :    1 - 0x1
    "00000000", -- 5067 - 0x13cb  :    0 - 0x0
    "00000110", -- 5068 - 0x13cc  :    6 - 0x6
    "10011000", -- 5069 - 0x13cd  :  152 - 0x98
    "01100000", -- 5070 - 0x13ce  :   96 - 0x60
    "00000000", -- 5071 - 0x13cf  :    0 - 0x0
    "11000000", -- 5072 - 0x13d0  :  192 - 0xc0
    "00100000", -- 5073 - 0x13d1  :   32 - 0x20
    "00010000", -- 5074 - 0x13d2  :   16 - 0x10
    "00010000", -- 5075 - 0x13d3  :   16 - 0x10
    "00010000", -- 5076 - 0x13d4  :   16 - 0x10
    "00010000", -- 5077 - 0x13d5  :   16 - 0x10
    "00100000", -- 5078 - 0x13d6  :   32 - 0x20
    "11000000", -- 5079 - 0x13d7  :  192 - 0xc0
    "11000000", -- 5080 - 0x13d8  :  192 - 0xc0
    "11100000", -- 5081 - 0x13d9  :  224 - 0xe0
    "11110000", -- 5082 - 0x13da  :  240 - 0xf0
    "11110000", -- 5083 - 0x13db  :  240 - 0xf0
    "11110000", -- 5084 - 0x13dc  :  240 - 0xf0
    "11110000", -- 5085 - 0x13dd  :  240 - 0xf0
    "11100000", -- 5086 - 0x13de  :  224 - 0xe0
    "11000000", -- 5087 - 0x13df  :  192 - 0xc0
    "00000000", -- 5088 - 0x13e0  :    0 - 0x0
    "00000000", -- 5089 - 0x13e1  :    0 - 0x0
    "00000000", -- 5090 - 0x13e2  :    0 - 0x0
    "00000000", -- 5091 - 0x13e3  :    0 - 0x0
    "00111111", -- 5092 - 0x13e4  :   63 - 0x3f
    "01111111", -- 5093 - 0x13e5  :  127 - 0x7f
    "11100000", -- 5094 - 0x13e6  :  224 - 0xe0
    "11000000", -- 5095 - 0x13e7  :  192 - 0xc0
    "00000000", -- 5096 - 0x13e8  :    0 - 0x0
    "00000000", -- 5097 - 0x13e9  :    0 - 0x0
    "00000000", -- 5098 - 0x13ea  :    0 - 0x0
    "00000000", -- 5099 - 0x13eb  :    0 - 0x0
    "00000000", -- 5100 - 0x13ec  :    0 - 0x0
    "00000000", -- 5101 - 0x13ed  :    0 - 0x0
    "00011100", -- 5102 - 0x13ee  :   28 - 0x1c
    "00111110", -- 5103 - 0x13ef  :   62 - 0x3e
    "10001000", -- 5104 - 0x13f0  :  136 - 0x88
    "10011100", -- 5105 - 0x13f1  :  156 - 0x9c
    "10001000", -- 5106 - 0x13f2  :  136 - 0x88
    "10000000", -- 5107 - 0x13f3  :  128 - 0x80
    "10000000", -- 5108 - 0x13f4  :  128 - 0x80
    "10000000", -- 5109 - 0x13f5  :  128 - 0x80
    "10000000", -- 5110 - 0x13f6  :  128 - 0x80
    "10000000", -- 5111 - 0x13f7  :  128 - 0x80
    "01111111", -- 5112 - 0x13f8  :  127 - 0x7f
    "01111111", -- 5113 - 0x13f9  :  127 - 0x7f
    "01111111", -- 5114 - 0x13fa  :  127 - 0x7f
    "00111110", -- 5115 - 0x13fb  :   62 - 0x3e
    "00011100", -- 5116 - 0x13fc  :   28 - 0x1c
    "00000000", -- 5117 - 0x13fd  :    0 - 0x0
    "00000000", -- 5118 - 0x13fe  :    0 - 0x0
    "00000000", -- 5119 - 0x13ff  :    0 - 0x0
    "11111110", -- 5120 - 0x1400  :  254 - 0xfe
    "11111110", -- 5121 - 0x1401  :  254 - 0xfe
    "11111110", -- 5122 - 0x1402  :  254 - 0xfe
    "11111110", -- 5123 - 0x1403  :  254 - 0xfe
    "11111110", -- 5124 - 0x1404  :  254 - 0xfe
    "11111110", -- 5125 - 0x1405  :  254 - 0xfe
    "11111110", -- 5126 - 0x1406  :  254 - 0xfe
    "11111110", -- 5127 - 0x1407  :  254 - 0xfe
    "11111111", -- 5128 - 0x1408  :  255 - 0xff
    "11111111", -- 5129 - 0x1409  :  255 - 0xff
    "11111111", -- 5130 - 0x140a  :  255 - 0xff
    "11111111", -- 5131 - 0x140b  :  255 - 0xff
    "11111111", -- 5132 - 0x140c  :  255 - 0xff
    "11111111", -- 5133 - 0x140d  :  255 - 0xff
    "11111111", -- 5134 - 0x140e  :  255 - 0xff
    "11111111", -- 5135 - 0x140f  :  255 - 0xff
    "00001000", -- 5136 - 0x1410  :    8 - 0x8
    "00010100", -- 5137 - 0x1411  :   20 - 0x14
    "00100100", -- 5138 - 0x1412  :   36 - 0x24
    "11000100", -- 5139 - 0x1413  :  196 - 0xc4
    "00000011", -- 5140 - 0x1414  :    3 - 0x3
    "01000000", -- 5141 - 0x1415  :   64 - 0x40
    "10100001", -- 5142 - 0x1416  :  161 - 0xa1
    "00100110", -- 5143 - 0x1417  :   38 - 0x26
    "00000000", -- 5144 - 0x1418  :    0 - 0x0
    "00001000", -- 5145 - 0x1419  :    8 - 0x8
    "00011000", -- 5146 - 0x141a  :   24 - 0x18
    "00111000", -- 5147 - 0x141b  :   56 - 0x38
    "11111100", -- 5148 - 0x141c  :  252 - 0xfc
    "10111111", -- 5149 - 0x141d  :  191 - 0xbf
    "01011110", -- 5150 - 0x141e  :   94 - 0x5e
    "11011001", -- 5151 - 0x141f  :  217 - 0xd9
    "11111111", -- 5152 - 0x1420  :  255 - 0xff
    "11111111", -- 5153 - 0x1421  :  255 - 0xff
    "11111111", -- 5154 - 0x1422  :  255 - 0xff
    "11111111", -- 5155 - 0x1423  :  255 - 0xff
    "01111111", -- 5156 - 0x1424  :  127 - 0x7f
    "01111111", -- 5157 - 0x1425  :  127 - 0x7f
    "01111111", -- 5158 - 0x1426  :  127 - 0x7f
    "01111111", -- 5159 - 0x1427  :  127 - 0x7f
    "10000001", -- 5160 - 0x1428  :  129 - 0x81
    "10000001", -- 5161 - 0x1429  :  129 - 0x81
    "10000001", -- 5162 - 0x142a  :  129 - 0x81
    "10000001", -- 5163 - 0x142b  :  129 - 0x81
    "10000001", -- 5164 - 0x142c  :  129 - 0x81
    "10000001", -- 5165 - 0x142d  :  129 - 0x81
    "10000001", -- 5166 - 0x142e  :  129 - 0x81
    "10000001", -- 5167 - 0x142f  :  129 - 0x81
    "11111111", -- 5168 - 0x1430  :  255 - 0xff
    "11111111", -- 5169 - 0x1431  :  255 - 0xff
    "11111111", -- 5170 - 0x1432  :  255 - 0xff
    "11111111", -- 5171 - 0x1433  :  255 - 0xff
    "11111111", -- 5172 - 0x1434  :  255 - 0xff
    "11111111", -- 5173 - 0x1435  :  255 - 0xff
    "11111111", -- 5174 - 0x1436  :  255 - 0xff
    "11111111", -- 5175 - 0x1437  :  255 - 0xff
    "00000001", -- 5176 - 0x1438  :    1 - 0x1
    "00000001", -- 5177 - 0x1439  :    1 - 0x1
    "00000001", -- 5178 - 0x143a  :    1 - 0x1
    "00000001", -- 5179 - 0x143b  :    1 - 0x1
    "00000001", -- 5180 - 0x143c  :    1 - 0x1
    "00000001", -- 5181 - 0x143d  :    1 - 0x1
    "00000001", -- 5182 - 0x143e  :    1 - 0x1
    "00000001", -- 5183 - 0x143f  :    1 - 0x1
    "01111111", -- 5184 - 0x1440  :  127 - 0x7f
    "10000000", -- 5185 - 0x1441  :  128 - 0x80
    "10000000", -- 5186 - 0x1442  :  128 - 0x80
    "10011000", -- 5187 - 0x1443  :  152 - 0x98
    "10011100", -- 5188 - 0x1444  :  156 - 0x9c
    "10001100", -- 5189 - 0x1445  :  140 - 0x8c
    "10000000", -- 5190 - 0x1446  :  128 - 0x80
    "10000000", -- 5191 - 0x1447  :  128 - 0x80
    "00000000", -- 5192 - 0x1448  :    0 - 0x0
    "01111111", -- 5193 - 0x1449  :  127 - 0x7f
    "01111111", -- 5194 - 0x144a  :  127 - 0x7f
    "01100111", -- 5195 - 0x144b  :  103 - 0x67
    "01100111", -- 5196 - 0x144c  :  103 - 0x67
    "01111111", -- 5197 - 0x144d  :  127 - 0x7f
    "01111111", -- 5198 - 0x144e  :  127 - 0x7f
    "01111111", -- 5199 - 0x144f  :  127 - 0x7f
    "11111111", -- 5200 - 0x1450  :  255 - 0xff
    "00000001", -- 5201 - 0x1451  :    1 - 0x1
    "00000001", -- 5202 - 0x1452  :    1 - 0x1
    "11111111", -- 5203 - 0x1453  :  255 - 0xff
    "00010000", -- 5204 - 0x1454  :   16 - 0x10
    "00010000", -- 5205 - 0x1455  :   16 - 0x10
    "00010000", -- 5206 - 0x1456  :   16 - 0x10
    "11111111", -- 5207 - 0x1457  :  255 - 0xff
    "00000000", -- 5208 - 0x1458  :    0 - 0x0
    "11111111", -- 5209 - 0x1459  :  255 - 0xff
    "11111111", -- 5210 - 0x145a  :  255 - 0xff
    "11111111", -- 5211 - 0x145b  :  255 - 0xff
    "11111111", -- 5212 - 0x145c  :  255 - 0xff
    "11111111", -- 5213 - 0x145d  :  255 - 0xff
    "11111111", -- 5214 - 0x145e  :  255 - 0xff
    "11111111", -- 5215 - 0x145f  :  255 - 0xff
    "10000000", -- 5216 - 0x1460  :  128 - 0x80
    "10000000", -- 5217 - 0x1461  :  128 - 0x80
    "10000000", -- 5218 - 0x1462  :  128 - 0x80
    "10000000", -- 5219 - 0x1463  :  128 - 0x80
    "10000000", -- 5220 - 0x1464  :  128 - 0x80
    "10000000", -- 5221 - 0x1465  :  128 - 0x80
    "10000000", -- 5222 - 0x1466  :  128 - 0x80
    "10000000", -- 5223 - 0x1467  :  128 - 0x80
    "01111111", -- 5224 - 0x1468  :  127 - 0x7f
    "01111111", -- 5225 - 0x1469  :  127 - 0x7f
    "01111111", -- 5226 - 0x146a  :  127 - 0x7f
    "01111111", -- 5227 - 0x146b  :  127 - 0x7f
    "01111111", -- 5228 - 0x146c  :  127 - 0x7f
    "01111111", -- 5229 - 0x146d  :  127 - 0x7f
    "01111111", -- 5230 - 0x146e  :  127 - 0x7f
    "01111111", -- 5231 - 0x146f  :  127 - 0x7f
    "00000001", -- 5232 - 0x1470  :    1 - 0x1
    "00000001", -- 5233 - 0x1471  :    1 - 0x1
    "00000001", -- 5234 - 0x1472  :    1 - 0x1
    "11111111", -- 5235 - 0x1473  :  255 - 0xff
    "00010000", -- 5236 - 0x1474  :   16 - 0x10
    "00010000", -- 5237 - 0x1475  :   16 - 0x10
    "00010000", -- 5238 - 0x1476  :   16 - 0x10
    "11111111", -- 5239 - 0x1477  :  255 - 0xff
    "11111111", -- 5240 - 0x1478  :  255 - 0xff
    "11111111", -- 5241 - 0x1479  :  255 - 0xff
    "11111111", -- 5242 - 0x147a  :  255 - 0xff
    "11111111", -- 5243 - 0x147b  :  255 - 0xff
    "11111111", -- 5244 - 0x147c  :  255 - 0xff
    "11111111", -- 5245 - 0x147d  :  255 - 0xff
    "11111111", -- 5246 - 0x147e  :  255 - 0xff
    "11111111", -- 5247 - 0x147f  :  255 - 0xff
    "11111111", -- 5248 - 0x1480  :  255 - 0xff
    "00000000", -- 5249 - 0x1481  :    0 - 0x0
    "00000000", -- 5250 - 0x1482  :    0 - 0x0
    "00000000", -- 5251 - 0x1483  :    0 - 0x0
    "00000000", -- 5252 - 0x1484  :    0 - 0x0
    "00000000", -- 5253 - 0x1485  :    0 - 0x0
    "00000000", -- 5254 - 0x1486  :    0 - 0x0
    "00000000", -- 5255 - 0x1487  :    0 - 0x0
    "00000000", -- 5256 - 0x1488  :    0 - 0x0
    "11111111", -- 5257 - 0x1489  :  255 - 0xff
    "11111111", -- 5258 - 0x148a  :  255 - 0xff
    "11111111", -- 5259 - 0x148b  :  255 - 0xff
    "11111111", -- 5260 - 0x148c  :  255 - 0xff
    "11111111", -- 5261 - 0x148d  :  255 - 0xff
    "11111111", -- 5262 - 0x148e  :  255 - 0xff
    "11111111", -- 5263 - 0x148f  :  255 - 0xff
    "11111110", -- 5264 - 0x1490  :  254 - 0xfe
    "00000001", -- 5265 - 0x1491  :    1 - 0x1
    "00000001", -- 5266 - 0x1492  :    1 - 0x1
    "00011001", -- 5267 - 0x1493  :   25 - 0x19
    "00011101", -- 5268 - 0x1494  :   29 - 0x1d
    "00001101", -- 5269 - 0x1495  :   13 - 0xd
    "00000001", -- 5270 - 0x1496  :    1 - 0x1
    "00000001", -- 5271 - 0x1497  :    1 - 0x1
    "00000000", -- 5272 - 0x1498  :    0 - 0x0
    "11111111", -- 5273 - 0x1499  :  255 - 0xff
    "11111111", -- 5274 - 0x149a  :  255 - 0xff
    "11100111", -- 5275 - 0x149b  :  231 - 0xe7
    "11100111", -- 5276 - 0x149c  :  231 - 0xe7
    "11111111", -- 5277 - 0x149d  :  255 - 0xff
    "11111111", -- 5278 - 0x149e  :  255 - 0xff
    "11111111", -- 5279 - 0x149f  :  255 - 0xff
    "00000001", -- 5280 - 0x14a0  :    1 - 0x1
    "00000001", -- 5281 - 0x14a1  :    1 - 0x1
    "00000001", -- 5282 - 0x14a2  :    1 - 0x1
    "00000001", -- 5283 - 0x14a3  :    1 - 0x1
    "00000001", -- 5284 - 0x14a4  :    1 - 0x1
    "00000001", -- 5285 - 0x14a5  :    1 - 0x1
    "00000001", -- 5286 - 0x14a6  :    1 - 0x1
    "00000001", -- 5287 - 0x14a7  :    1 - 0x1
    "11111111", -- 5288 - 0x14a8  :  255 - 0xff
    "11111111", -- 5289 - 0x14a9  :  255 - 0xff
    "11111111", -- 5290 - 0x14aa  :  255 - 0xff
    "11111111", -- 5291 - 0x14ab  :  255 - 0xff
    "11111111", -- 5292 - 0x14ac  :  255 - 0xff
    "11111111", -- 5293 - 0x14ad  :  255 - 0xff
    "11111111", -- 5294 - 0x14ae  :  255 - 0xff
    "11111111", -- 5295 - 0x14af  :  255 - 0xff
    "00111111", -- 5296 - 0x14b0  :   63 - 0x3f
    "01111111", -- 5297 - 0x14b1  :  127 - 0x7f
    "01111111", -- 5298 - 0x14b2  :  127 - 0x7f
    "11111111", -- 5299 - 0x14b3  :  255 - 0xff
    "11111111", -- 5300 - 0x14b4  :  255 - 0xff
    "11111111", -- 5301 - 0x14b5  :  255 - 0xff
    "11111111", -- 5302 - 0x14b6  :  255 - 0xff
    "11111111", -- 5303 - 0x14b7  :  255 - 0xff
    "00111111", -- 5304 - 0x14b8  :   63 - 0x3f
    "01100000", -- 5305 - 0x14b9  :   96 - 0x60
    "01000000", -- 5306 - 0x14ba  :   64 - 0x40
    "11000000", -- 5307 - 0x14bb  :  192 - 0xc0
    "10000000", -- 5308 - 0x14bc  :  128 - 0x80
    "10000000", -- 5309 - 0x14bd  :  128 - 0x80
    "10000000", -- 5310 - 0x14be  :  128 - 0x80
    "10000000", -- 5311 - 0x14bf  :  128 - 0x80
    "11111111", -- 5312 - 0x14c0  :  255 - 0xff
    "11111111", -- 5313 - 0x14c1  :  255 - 0xff
    "11111111", -- 5314 - 0x14c2  :  255 - 0xff
    "11111111", -- 5315 - 0x14c3  :  255 - 0xff
    "11111111", -- 5316 - 0x14c4  :  255 - 0xff
    "11111111", -- 5317 - 0x14c5  :  255 - 0xff
    "01111110", -- 5318 - 0x14c6  :  126 - 0x7e
    "00111100", -- 5319 - 0x14c7  :   60 - 0x3c
    "10000000", -- 5320 - 0x14c8  :  128 - 0x80
    "10000000", -- 5321 - 0x14c9  :  128 - 0x80
    "10000000", -- 5322 - 0x14ca  :  128 - 0x80
    "10000000", -- 5323 - 0x14cb  :  128 - 0x80
    "10000000", -- 5324 - 0x14cc  :  128 - 0x80
    "10000001", -- 5325 - 0x14cd  :  129 - 0x81
    "01000010", -- 5326 - 0x14ce  :   66 - 0x42
    "00111100", -- 5327 - 0x14cf  :   60 - 0x3c
    "11111111", -- 5328 - 0x14d0  :  255 - 0xff
    "11111111", -- 5329 - 0x14d1  :  255 - 0xff
    "11111111", -- 5330 - 0x14d2  :  255 - 0xff
    "11111111", -- 5331 - 0x14d3  :  255 - 0xff
    "11111111", -- 5332 - 0x14d4  :  255 - 0xff
    "11111111", -- 5333 - 0x14d5  :  255 - 0xff
    "11111111", -- 5334 - 0x14d6  :  255 - 0xff
    "11111111", -- 5335 - 0x14d7  :  255 - 0xff
    "11111111", -- 5336 - 0x14d8  :  255 - 0xff
    "00000000", -- 5337 - 0x14d9  :    0 - 0x0
    "00000000", -- 5338 - 0x14da  :    0 - 0x0
    "00000000", -- 5339 - 0x14db  :    0 - 0x0
    "00000000", -- 5340 - 0x14dc  :    0 - 0x0
    "00000000", -- 5341 - 0x14dd  :    0 - 0x0
    "00000000", -- 5342 - 0x14de  :    0 - 0x0
    "00000000", -- 5343 - 0x14df  :    0 - 0x0
    "11111111", -- 5344 - 0x14e0  :  255 - 0xff
    "11111111", -- 5345 - 0x14e1  :  255 - 0xff
    "11111111", -- 5346 - 0x14e2  :  255 - 0xff
    "11111111", -- 5347 - 0x14e3  :  255 - 0xff
    "11111111", -- 5348 - 0x14e4  :  255 - 0xff
    "11111111", -- 5349 - 0x14e5  :  255 - 0xff
    "11111110", -- 5350 - 0x14e6  :  254 - 0xfe
    "01111100", -- 5351 - 0x14e7  :  124 - 0x7c
    "00000000", -- 5352 - 0x14e8  :    0 - 0x0
    "00000000", -- 5353 - 0x14e9  :    0 - 0x0
    "00000000", -- 5354 - 0x14ea  :    0 - 0x0
    "00000000", -- 5355 - 0x14eb  :    0 - 0x0
    "00000000", -- 5356 - 0x14ec  :    0 - 0x0
    "00000001", -- 5357 - 0x14ed  :    1 - 0x1
    "10000010", -- 5358 - 0x14ee  :  130 - 0x82
    "01111100", -- 5359 - 0x14ef  :  124 - 0x7c
    "11111111", -- 5360 - 0x14f0  :  255 - 0xff
    "11111111", -- 5361 - 0x14f1  :  255 - 0xff
    "11111111", -- 5362 - 0x14f2  :  255 - 0xff
    "11111111", -- 5363 - 0x14f3  :  255 - 0xff
    "11111111", -- 5364 - 0x14f4  :  255 - 0xff
    "11111111", -- 5365 - 0x14f5  :  255 - 0xff
    "11111110", -- 5366 - 0x14f6  :  254 - 0xfe
    "01111100", -- 5367 - 0x14f7  :  124 - 0x7c
    "00000000", -- 5368 - 0x14f8  :    0 - 0x0
    "00000000", -- 5369 - 0x14f9  :    0 - 0x0
    "00000000", -- 5370 - 0x14fa  :    0 - 0x0
    "00000000", -- 5371 - 0x14fb  :    0 - 0x0
    "00000000", -- 5372 - 0x14fc  :    0 - 0x0
    "00000001", -- 5373 - 0x14fd  :    1 - 0x1
    "10000011", -- 5374 - 0x14fe  :  131 - 0x83
    "11111111", -- 5375 - 0x14ff  :  255 - 0xff
    "11111000", -- 5376 - 0x1500  :  248 - 0xf8
    "11111100", -- 5377 - 0x1501  :  252 - 0xfc
    "11111110", -- 5378 - 0x1502  :  254 - 0xfe
    "11111110", -- 5379 - 0x1503  :  254 - 0xfe
    "11111111", -- 5380 - 0x1504  :  255 - 0xff
    "11111111", -- 5381 - 0x1505  :  255 - 0xff
    "11111111", -- 5382 - 0x1506  :  255 - 0xff
    "11111111", -- 5383 - 0x1507  :  255 - 0xff
    "11111000", -- 5384 - 0x1508  :  248 - 0xf8
    "00000100", -- 5385 - 0x1509  :    4 - 0x4
    "00000010", -- 5386 - 0x150a  :    2 - 0x2
    "00000010", -- 5387 - 0x150b  :    2 - 0x2
    "00000001", -- 5388 - 0x150c  :    1 - 0x1
    "00000001", -- 5389 - 0x150d  :    1 - 0x1
    "00000001", -- 5390 - 0x150e  :    1 - 0x1
    "00000001", -- 5391 - 0x150f  :    1 - 0x1
    "11111111", -- 5392 - 0x1510  :  255 - 0xff
    "11111111", -- 5393 - 0x1511  :  255 - 0xff
    "11111111", -- 5394 - 0x1512  :  255 - 0xff
    "11111111", -- 5395 - 0x1513  :  255 - 0xff
    "11111111", -- 5396 - 0x1514  :  255 - 0xff
    "11111111", -- 5397 - 0x1515  :  255 - 0xff
    "01111110", -- 5398 - 0x1516  :  126 - 0x7e
    "00111100", -- 5399 - 0x1517  :   60 - 0x3c
    "00000001", -- 5400 - 0x1518  :    1 - 0x1
    "00000001", -- 5401 - 0x1519  :    1 - 0x1
    "00000001", -- 5402 - 0x151a  :    1 - 0x1
    "00000001", -- 5403 - 0x151b  :    1 - 0x1
    "00000001", -- 5404 - 0x151c  :    1 - 0x1
    "10000001", -- 5405 - 0x151d  :  129 - 0x81
    "01000010", -- 5406 - 0x151e  :   66 - 0x42
    "00111100", -- 5407 - 0x151f  :   60 - 0x3c
    "00000000", -- 5408 - 0x1520  :    0 - 0x0
    "00001000", -- 5409 - 0x1521  :    8 - 0x8
    "00001000", -- 5410 - 0x1522  :    8 - 0x8
    "00001000", -- 5411 - 0x1523  :    8 - 0x8
    "00010000", -- 5412 - 0x1524  :   16 - 0x10
    "00010000", -- 5413 - 0x1525  :   16 - 0x10
    "00010000", -- 5414 - 0x1526  :   16 - 0x10
    "00000000", -- 5415 - 0x1527  :    0 - 0x0
    "11111111", -- 5416 - 0x1528  :  255 - 0xff
    "11111111", -- 5417 - 0x1529  :  255 - 0xff
    "11111111", -- 5418 - 0x152a  :  255 - 0xff
    "11111111", -- 5419 - 0x152b  :  255 - 0xff
    "11111111", -- 5420 - 0x152c  :  255 - 0xff
    "11111111", -- 5421 - 0x152d  :  255 - 0xff
    "11111111", -- 5422 - 0x152e  :  255 - 0xff
    "11111111", -- 5423 - 0x152f  :  255 - 0xff
    "00000000", -- 5424 - 0x1530  :    0 - 0x0
    "01111111", -- 5425 - 0x1531  :  127 - 0x7f
    "01111111", -- 5426 - 0x1532  :  127 - 0x7f
    "01111000", -- 5427 - 0x1533  :  120 - 0x78
    "01110011", -- 5428 - 0x1534  :  115 - 0x73
    "01110011", -- 5429 - 0x1535  :  115 - 0x73
    "01110011", -- 5430 - 0x1536  :  115 - 0x73
    "01111111", -- 5431 - 0x1537  :  127 - 0x7f
    "01111111", -- 5432 - 0x1538  :  127 - 0x7f
    "10000000", -- 5433 - 0x1539  :  128 - 0x80
    "10100000", -- 5434 - 0x153a  :  160 - 0xa0
    "10000111", -- 5435 - 0x153b  :  135 - 0x87
    "10001111", -- 5436 - 0x153c  :  143 - 0x8f
    "10001110", -- 5437 - 0x153d  :  142 - 0x8e
    "10001110", -- 5438 - 0x153e  :  142 - 0x8e
    "10000110", -- 5439 - 0x153f  :  134 - 0x86
    "00000000", -- 5440 - 0x1540  :    0 - 0x0
    "11111111", -- 5441 - 0x1541  :  255 - 0xff
    "11111111", -- 5442 - 0x1542  :  255 - 0xff
    "00111111", -- 5443 - 0x1543  :   63 - 0x3f
    "10011111", -- 5444 - 0x1544  :  159 - 0x9f
    "10011111", -- 5445 - 0x1545  :  159 - 0x9f
    "10011111", -- 5446 - 0x1546  :  159 - 0x9f
    "00011111", -- 5447 - 0x1547  :   31 - 0x1f
    "11111110", -- 5448 - 0x1548  :  254 - 0xfe
    "00000001", -- 5449 - 0x1549  :    1 - 0x1
    "00000101", -- 5450 - 0x154a  :    5 - 0x5
    "11000001", -- 5451 - 0x154b  :  193 - 0xc1
    "11100001", -- 5452 - 0x154c  :  225 - 0xe1
    "01110001", -- 5453 - 0x154d  :  113 - 0x71
    "01110001", -- 5454 - 0x154e  :  113 - 0x71
    "11110001", -- 5455 - 0x154f  :  241 - 0xf1
    "01111110", -- 5456 - 0x1550  :  126 - 0x7e
    "01111110", -- 5457 - 0x1551  :  126 - 0x7e
    "01111111", -- 5458 - 0x1552  :  127 - 0x7f
    "01111110", -- 5459 - 0x1553  :  126 - 0x7e
    "01111110", -- 5460 - 0x1554  :  126 - 0x7e
    "01111111", -- 5461 - 0x1555  :  127 - 0x7f
    "01111111", -- 5462 - 0x1556  :  127 - 0x7f
    "11111111", -- 5463 - 0x1557  :  255 - 0xff
    "10000001", -- 5464 - 0x1558  :  129 - 0x81
    "10000001", -- 5465 - 0x1559  :  129 - 0x81
    "10000000", -- 5466 - 0x155a  :  128 - 0x80
    "10000001", -- 5467 - 0x155b  :  129 - 0x81
    "10000001", -- 5468 - 0x155c  :  129 - 0x81
    "10100000", -- 5469 - 0x155d  :  160 - 0xa0
    "10000000", -- 5470 - 0x155e  :  128 - 0x80
    "11111111", -- 5471 - 0x155f  :  255 - 0xff
    "01111111", -- 5472 - 0x1560  :  127 - 0x7f
    "01111111", -- 5473 - 0x1561  :  127 - 0x7f
    "11111111", -- 5474 - 0x1562  :  255 - 0xff
    "01111111", -- 5475 - 0x1563  :  127 - 0x7f
    "01111111", -- 5476 - 0x1564  :  127 - 0x7f
    "11111111", -- 5477 - 0x1565  :  255 - 0xff
    "11111111", -- 5478 - 0x1566  :  255 - 0xff
    "11111111", -- 5479 - 0x1567  :  255 - 0xff
    "11110001", -- 5480 - 0x1568  :  241 - 0xf1
    "11000001", -- 5481 - 0x1569  :  193 - 0xc1
    "11000001", -- 5482 - 0x156a  :  193 - 0xc1
    "10000001", -- 5483 - 0x156b  :  129 - 0x81
    "11000001", -- 5484 - 0x156c  :  193 - 0xc1
    "11000101", -- 5485 - 0x156d  :  197 - 0xc5
    "00000001", -- 5486 - 0x156e  :    1 - 0x1
    "11111111", -- 5487 - 0x156f  :  255 - 0xff
    "01111111", -- 5488 - 0x1570  :  127 - 0x7f
    "10000000", -- 5489 - 0x1571  :  128 - 0x80
    "10100000", -- 5490 - 0x1572  :  160 - 0xa0
    "10000000", -- 5491 - 0x1573  :  128 - 0x80
    "10000000", -- 5492 - 0x1574  :  128 - 0x80
    "10000000", -- 5493 - 0x1575  :  128 - 0x80
    "10000000", -- 5494 - 0x1576  :  128 - 0x80
    "10000000", -- 5495 - 0x1577  :  128 - 0x80
    "01111111", -- 5496 - 0x1578  :  127 - 0x7f
    "11111111", -- 5497 - 0x1579  :  255 - 0xff
    "11111111", -- 5498 - 0x157a  :  255 - 0xff
    "11111111", -- 5499 - 0x157b  :  255 - 0xff
    "11111111", -- 5500 - 0x157c  :  255 - 0xff
    "11111111", -- 5501 - 0x157d  :  255 - 0xff
    "11111111", -- 5502 - 0x157e  :  255 - 0xff
    "11111111", -- 5503 - 0x157f  :  255 - 0xff
    "11111110", -- 5504 - 0x1580  :  254 - 0xfe
    "00000001", -- 5505 - 0x1581  :    1 - 0x1
    "00000101", -- 5506 - 0x1582  :    5 - 0x5
    "00000001", -- 5507 - 0x1583  :    1 - 0x1
    "00000001", -- 5508 - 0x1584  :    1 - 0x1
    "00000001", -- 5509 - 0x1585  :    1 - 0x1
    "00000001", -- 5510 - 0x1586  :    1 - 0x1
    "00000001", -- 5511 - 0x1587  :    1 - 0x1
    "11111110", -- 5512 - 0x1588  :  254 - 0xfe
    "11111111", -- 5513 - 0x1589  :  255 - 0xff
    "11111111", -- 5514 - 0x158a  :  255 - 0xff
    "11111111", -- 5515 - 0x158b  :  255 - 0xff
    "11111111", -- 5516 - 0x158c  :  255 - 0xff
    "11111111", -- 5517 - 0x158d  :  255 - 0xff
    "11111111", -- 5518 - 0x158e  :  255 - 0xff
    "11111111", -- 5519 - 0x158f  :  255 - 0xff
    "10000000", -- 5520 - 0x1590  :  128 - 0x80
    "10000000", -- 5521 - 0x1591  :  128 - 0x80
    "10000000", -- 5522 - 0x1592  :  128 - 0x80
    "10000000", -- 5523 - 0x1593  :  128 - 0x80
    "10000000", -- 5524 - 0x1594  :  128 - 0x80
    "10100000", -- 5525 - 0x1595  :  160 - 0xa0
    "10000000", -- 5526 - 0x1596  :  128 - 0x80
    "01111111", -- 5527 - 0x1597  :  127 - 0x7f
    "11111111", -- 5528 - 0x1598  :  255 - 0xff
    "11111111", -- 5529 - 0x1599  :  255 - 0xff
    "11111111", -- 5530 - 0x159a  :  255 - 0xff
    "11111111", -- 5531 - 0x159b  :  255 - 0xff
    "11111111", -- 5532 - 0x159c  :  255 - 0xff
    "11111111", -- 5533 - 0x159d  :  255 - 0xff
    "11111111", -- 5534 - 0x159e  :  255 - 0xff
    "01111111", -- 5535 - 0x159f  :  127 - 0x7f
    "00000001", -- 5536 - 0x15a0  :    1 - 0x1
    "00000001", -- 5537 - 0x15a1  :    1 - 0x1
    "00000001", -- 5538 - 0x15a2  :    1 - 0x1
    "00000001", -- 5539 - 0x15a3  :    1 - 0x1
    "00000001", -- 5540 - 0x15a4  :    1 - 0x1
    "00000101", -- 5541 - 0x15a5  :    5 - 0x5
    "00000001", -- 5542 - 0x15a6  :    1 - 0x1
    "11111110", -- 5543 - 0x15a7  :  254 - 0xfe
    "11111111", -- 5544 - 0x15a8  :  255 - 0xff
    "11111111", -- 5545 - 0x15a9  :  255 - 0xff
    "11111111", -- 5546 - 0x15aa  :  255 - 0xff
    "11111111", -- 5547 - 0x15ab  :  255 - 0xff
    "11111111", -- 5548 - 0x15ac  :  255 - 0xff
    "11111111", -- 5549 - 0x15ad  :  255 - 0xff
    "11111111", -- 5550 - 0x15ae  :  255 - 0xff
    "11111110", -- 5551 - 0x15af  :  254 - 0xfe
    "00000000", -- 5552 - 0x15b0  :    0 - 0x0
    "00000000", -- 5553 - 0x15b1  :    0 - 0x0
    "00000000", -- 5554 - 0x15b2  :    0 - 0x0
    "00000000", -- 5555 - 0x15b3  :    0 - 0x0
    "11111100", -- 5556 - 0x15b4  :  252 - 0xfc
    "11111110", -- 5557 - 0x15b5  :  254 - 0xfe
    "00000111", -- 5558 - 0x15b6  :    7 - 0x7
    "00000011", -- 5559 - 0x15b7  :    3 - 0x3
    "00000000", -- 5560 - 0x15b8  :    0 - 0x0
    "00000000", -- 5561 - 0x15b9  :    0 - 0x0
    "00000000", -- 5562 - 0x15ba  :    0 - 0x0
    "00000000", -- 5563 - 0x15bb  :    0 - 0x0
    "00000000", -- 5564 - 0x15bc  :    0 - 0x0
    "00000000", -- 5565 - 0x15bd  :    0 - 0x0
    "00111000", -- 5566 - 0x15be  :   56 - 0x38
    "01111100", -- 5567 - 0x15bf  :  124 - 0x7c
    "00010001", -- 5568 - 0x15c0  :   17 - 0x11
    "00111001", -- 5569 - 0x15c1  :   57 - 0x39
    "00010001", -- 5570 - 0x15c2  :   17 - 0x11
    "00000001", -- 5571 - 0x15c3  :    1 - 0x1
    "00000001", -- 5572 - 0x15c4  :    1 - 0x1
    "00000001", -- 5573 - 0x15c5  :    1 - 0x1
    "00000001", -- 5574 - 0x15c6  :    1 - 0x1
    "00000001", -- 5575 - 0x15c7  :    1 - 0x1
    "11111110", -- 5576 - 0x15c8  :  254 - 0xfe
    "11111110", -- 5577 - 0x15c9  :  254 - 0xfe
    "11111110", -- 5578 - 0x15ca  :  254 - 0xfe
    "01111100", -- 5579 - 0x15cb  :  124 - 0x7c
    "00111000", -- 5580 - 0x15cc  :   56 - 0x38
    "00000000", -- 5581 - 0x15cd  :    0 - 0x0
    "00000000", -- 5582 - 0x15ce  :    0 - 0x0
    "00000000", -- 5583 - 0x15cf  :    0 - 0x0
    "11101111", -- 5584 - 0x15d0  :  239 - 0xef
    "00101000", -- 5585 - 0x15d1  :   40 - 0x28
    "00101000", -- 5586 - 0x15d2  :   40 - 0x28
    "00101000", -- 5587 - 0x15d3  :   40 - 0x28
    "00101000", -- 5588 - 0x15d4  :   40 - 0x28
    "00101000", -- 5589 - 0x15d5  :   40 - 0x28
    "11101111", -- 5590 - 0x15d6  :  239 - 0xef
    "00000000", -- 5591 - 0x15d7  :    0 - 0x0
    "00100000", -- 5592 - 0x15d8  :   32 - 0x20
    "11100111", -- 5593 - 0x15d9  :  231 - 0xe7
    "11100111", -- 5594 - 0x15da  :  231 - 0xe7
    "11100111", -- 5595 - 0x15db  :  231 - 0xe7
    "11100111", -- 5596 - 0x15dc  :  231 - 0xe7
    "11100111", -- 5597 - 0x15dd  :  231 - 0xe7
    "11101111", -- 5598 - 0x15de  :  239 - 0xef
    "00000000", -- 5599 - 0x15df  :    0 - 0x0
    "11111110", -- 5600 - 0x15e0  :  254 - 0xfe
    "10000010", -- 5601 - 0x15e1  :  130 - 0x82
    "10000010", -- 5602 - 0x15e2  :  130 - 0x82
    "10000010", -- 5603 - 0x15e3  :  130 - 0x82
    "10000010", -- 5604 - 0x15e4  :  130 - 0x82
    "10000010", -- 5605 - 0x15e5  :  130 - 0x82
    "11111110", -- 5606 - 0x15e6  :  254 - 0xfe
    "00000000", -- 5607 - 0x15e7  :    0 - 0x0
    "00000010", -- 5608 - 0x15e8  :    2 - 0x2
    "01111110", -- 5609 - 0x15e9  :  126 - 0x7e
    "01111110", -- 5610 - 0x15ea  :  126 - 0x7e
    "01111110", -- 5611 - 0x15eb  :  126 - 0x7e
    "01111110", -- 5612 - 0x15ec  :  126 - 0x7e
    "01111110", -- 5613 - 0x15ed  :  126 - 0x7e
    "11111110", -- 5614 - 0x15ee  :  254 - 0xfe
    "00000000", -- 5615 - 0x15ef  :    0 - 0x0
    "10000000", -- 5616 - 0x15f0  :  128 - 0x80
    "10000000", -- 5617 - 0x15f1  :  128 - 0x80
    "10000000", -- 5618 - 0x15f2  :  128 - 0x80
    "10011000", -- 5619 - 0x15f3  :  152 - 0x98
    "10011100", -- 5620 - 0x15f4  :  156 - 0x9c
    "10001100", -- 5621 - 0x15f5  :  140 - 0x8c
    "10000000", -- 5622 - 0x15f6  :  128 - 0x80
    "01111111", -- 5623 - 0x15f7  :  127 - 0x7f
    "01111111", -- 5624 - 0x15f8  :  127 - 0x7f
    "01111111", -- 5625 - 0x15f9  :  127 - 0x7f
    "01111111", -- 5626 - 0x15fa  :  127 - 0x7f
    "01100111", -- 5627 - 0x15fb  :  103 - 0x67
    "01100111", -- 5628 - 0x15fc  :  103 - 0x67
    "01111111", -- 5629 - 0x15fd  :  127 - 0x7f
    "01111111", -- 5630 - 0x15fe  :  127 - 0x7f
    "01111111", -- 5631 - 0x15ff  :  127 - 0x7f
    "11111111", -- 5632 - 0x1600  :  255 - 0xff
    "11111111", -- 5633 - 0x1601  :  255 - 0xff
    "10000011", -- 5634 - 0x1602  :  131 - 0x83
    "11110011", -- 5635 - 0x1603  :  243 - 0xf3
    "11110011", -- 5636 - 0x1604  :  243 - 0xf3
    "11110011", -- 5637 - 0x1605  :  243 - 0xf3
    "11110011", -- 5638 - 0x1606  :  243 - 0xf3
    "11110011", -- 5639 - 0x1607  :  243 - 0xf3
    "11111111", -- 5640 - 0x1608  :  255 - 0xff
    "10000000", -- 5641 - 0x1609  :  128 - 0x80
    "11111100", -- 5642 - 0x160a  :  252 - 0xfc
    "10001100", -- 5643 - 0x160b  :  140 - 0x8c
    "10001100", -- 5644 - 0x160c  :  140 - 0x8c
    "10001100", -- 5645 - 0x160d  :  140 - 0x8c
    "10001100", -- 5646 - 0x160e  :  140 - 0x8c
    "10001100", -- 5647 - 0x160f  :  140 - 0x8c
    "11111111", -- 5648 - 0x1610  :  255 - 0xff
    "11111111", -- 5649 - 0x1611  :  255 - 0xff
    "11110000", -- 5650 - 0x1612  :  240 - 0xf0
    "11110110", -- 5651 - 0x1613  :  246 - 0xf6
    "11110110", -- 5652 - 0x1614  :  246 - 0xf6
    "11110110", -- 5653 - 0x1615  :  246 - 0xf6
    "11110110", -- 5654 - 0x1616  :  246 - 0xf6
    "11110110", -- 5655 - 0x1617  :  246 - 0xf6
    "11111111", -- 5656 - 0x1618  :  255 - 0xff
    "00000000", -- 5657 - 0x1619  :    0 - 0x0
    "00001111", -- 5658 - 0x161a  :   15 - 0xf
    "00001001", -- 5659 - 0x161b  :    9 - 0x9
    "00001001", -- 5660 - 0x161c  :    9 - 0x9
    "00001001", -- 5661 - 0x161d  :    9 - 0x9
    "00001001", -- 5662 - 0x161e  :    9 - 0x9
    "00001001", -- 5663 - 0x161f  :    9 - 0x9
    "11111111", -- 5664 - 0x1620  :  255 - 0xff
    "11111111", -- 5665 - 0x1621  :  255 - 0xff
    "00000000", -- 5666 - 0x1622  :    0 - 0x0
    "00000000", -- 5667 - 0x1623  :    0 - 0x0
    "00000000", -- 5668 - 0x1624  :    0 - 0x0
    "00000000", -- 5669 - 0x1625  :    0 - 0x0
    "00000000", -- 5670 - 0x1626  :    0 - 0x0
    "00000000", -- 5671 - 0x1627  :    0 - 0x0
    "11111111", -- 5672 - 0x1628  :  255 - 0xff
    "00000000", -- 5673 - 0x1629  :    0 - 0x0
    "11111111", -- 5674 - 0x162a  :  255 - 0xff
    "11111111", -- 5675 - 0x162b  :  255 - 0xff
    "11111111", -- 5676 - 0x162c  :  255 - 0xff
    "11111111", -- 5677 - 0x162d  :  255 - 0xff
    "11111111", -- 5678 - 0x162e  :  255 - 0xff
    "11111111", -- 5679 - 0x162f  :  255 - 0xff
    "11111111", -- 5680 - 0x1630  :  255 - 0xff
    "11111111", -- 5681 - 0x1631  :  255 - 0xff
    "00000001", -- 5682 - 0x1632  :    1 - 0x1
    "01010111", -- 5683 - 0x1633  :   87 - 0x57
    "00101111", -- 5684 - 0x1634  :   47 - 0x2f
    "01010111", -- 5685 - 0x1635  :   87 - 0x57
    "00101111", -- 5686 - 0x1636  :   47 - 0x2f
    "01010111", -- 5687 - 0x1637  :   87 - 0x57
    "11111111", -- 5688 - 0x1638  :  255 - 0xff
    "00000001", -- 5689 - 0x1639  :    1 - 0x1
    "11111111", -- 5690 - 0x163a  :  255 - 0xff
    "10101001", -- 5691 - 0x163b  :  169 - 0xa9
    "11010001", -- 5692 - 0x163c  :  209 - 0xd1
    "10101001", -- 5693 - 0x163d  :  169 - 0xa9
    "11010001", -- 5694 - 0x163e  :  209 - 0xd1
    "10101001", -- 5695 - 0x163f  :  169 - 0xa9
    "11110011", -- 5696 - 0x1640  :  243 - 0xf3
    "11110011", -- 5697 - 0x1641  :  243 - 0xf3
    "11110011", -- 5698 - 0x1642  :  243 - 0xf3
    "11110011", -- 5699 - 0x1643  :  243 - 0xf3
    "11110011", -- 5700 - 0x1644  :  243 - 0xf3
    "11110011", -- 5701 - 0x1645  :  243 - 0xf3
    "11111111", -- 5702 - 0x1646  :  255 - 0xff
    "00111111", -- 5703 - 0x1647  :   63 - 0x3f
    "10001100", -- 5704 - 0x1648  :  140 - 0x8c
    "10001100", -- 5705 - 0x1649  :  140 - 0x8c
    "10001100", -- 5706 - 0x164a  :  140 - 0x8c
    "10001100", -- 5707 - 0x164b  :  140 - 0x8c
    "10001100", -- 5708 - 0x164c  :  140 - 0x8c
    "10001100", -- 5709 - 0x164d  :  140 - 0x8c
    "11111111", -- 5710 - 0x164e  :  255 - 0xff
    "00111111", -- 5711 - 0x164f  :   63 - 0x3f
    "11110110", -- 5712 - 0x1650  :  246 - 0xf6
    "11110110", -- 5713 - 0x1651  :  246 - 0xf6
    "11110110", -- 5714 - 0x1652  :  246 - 0xf6
    "11110110", -- 5715 - 0x1653  :  246 - 0xf6
    "11110110", -- 5716 - 0x1654  :  246 - 0xf6
    "11110110", -- 5717 - 0x1655  :  246 - 0xf6
    "11111111", -- 5718 - 0x1656  :  255 - 0xff
    "11111111", -- 5719 - 0x1657  :  255 - 0xff
    "00001001", -- 5720 - 0x1658  :    9 - 0x9
    "00001001", -- 5721 - 0x1659  :    9 - 0x9
    "00001001", -- 5722 - 0x165a  :    9 - 0x9
    "00001001", -- 5723 - 0x165b  :    9 - 0x9
    "00001001", -- 5724 - 0x165c  :    9 - 0x9
    "00001001", -- 5725 - 0x165d  :    9 - 0x9
    "11111111", -- 5726 - 0x165e  :  255 - 0xff
    "11111111", -- 5727 - 0x165f  :  255 - 0xff
    "00000000", -- 5728 - 0x1660  :    0 - 0x0
    "00000000", -- 5729 - 0x1661  :    0 - 0x0
    "00000000", -- 5730 - 0x1662  :    0 - 0x0
    "00000000", -- 5731 - 0x1663  :    0 - 0x0
    "00000000", -- 5732 - 0x1664  :    0 - 0x0
    "00000000", -- 5733 - 0x1665  :    0 - 0x0
    "11111111", -- 5734 - 0x1666  :  255 - 0xff
    "11111111", -- 5735 - 0x1667  :  255 - 0xff
    "11111111", -- 5736 - 0x1668  :  255 - 0xff
    "11111111", -- 5737 - 0x1669  :  255 - 0xff
    "11111111", -- 5738 - 0x166a  :  255 - 0xff
    "11111111", -- 5739 - 0x166b  :  255 - 0xff
    "11111111", -- 5740 - 0x166c  :  255 - 0xff
    "11111111", -- 5741 - 0x166d  :  255 - 0xff
    "11111111", -- 5742 - 0x166e  :  255 - 0xff
    "11111111", -- 5743 - 0x166f  :  255 - 0xff
    "00101111", -- 5744 - 0x1670  :   47 - 0x2f
    "01010111", -- 5745 - 0x1671  :   87 - 0x57
    "00101111", -- 5746 - 0x1672  :   47 - 0x2f
    "01010111", -- 5747 - 0x1673  :   87 - 0x57
    "00101111", -- 5748 - 0x1674  :   47 - 0x2f
    "01010111", -- 5749 - 0x1675  :   87 - 0x57
    "11111111", -- 5750 - 0x1676  :  255 - 0xff
    "11111100", -- 5751 - 0x1677  :  252 - 0xfc
    "11010001", -- 5752 - 0x1678  :  209 - 0xd1
    "10101001", -- 5753 - 0x1679  :  169 - 0xa9
    "11010001", -- 5754 - 0x167a  :  209 - 0xd1
    "10101001", -- 5755 - 0x167b  :  169 - 0xa9
    "11010001", -- 5756 - 0x167c  :  209 - 0xd1
    "10101001", -- 5757 - 0x167d  :  169 - 0xa9
    "11111111", -- 5758 - 0x167e  :  255 - 0xff
    "11111100", -- 5759 - 0x167f  :  252 - 0xfc
    "00111100", -- 5760 - 0x1680  :   60 - 0x3c
    "00111100", -- 5761 - 0x1681  :   60 - 0x3c
    "00111100", -- 5762 - 0x1682  :   60 - 0x3c
    "00111100", -- 5763 - 0x1683  :   60 - 0x3c
    "00111100", -- 5764 - 0x1684  :   60 - 0x3c
    "00111100", -- 5765 - 0x1685  :   60 - 0x3c
    "00111100", -- 5766 - 0x1686  :   60 - 0x3c
    "00111100", -- 5767 - 0x1687  :   60 - 0x3c
    "00100011", -- 5768 - 0x1688  :   35 - 0x23
    "00100011", -- 5769 - 0x1689  :   35 - 0x23
    "00100011", -- 5770 - 0x168a  :   35 - 0x23
    "00100011", -- 5771 - 0x168b  :   35 - 0x23
    "00100011", -- 5772 - 0x168c  :   35 - 0x23
    "00100011", -- 5773 - 0x168d  :   35 - 0x23
    "00100011", -- 5774 - 0x168e  :   35 - 0x23
    "00100011", -- 5775 - 0x168f  :   35 - 0x23
    "11111011", -- 5776 - 0x1690  :  251 - 0xfb
    "11111011", -- 5777 - 0x1691  :  251 - 0xfb
    "11111011", -- 5778 - 0x1692  :  251 - 0xfb
    "11111011", -- 5779 - 0x1693  :  251 - 0xfb
    "11111011", -- 5780 - 0x1694  :  251 - 0xfb
    "11111011", -- 5781 - 0x1695  :  251 - 0xfb
    "11111011", -- 5782 - 0x1696  :  251 - 0xfb
    "11111011", -- 5783 - 0x1697  :  251 - 0xfb
    "00000100", -- 5784 - 0x1698  :    4 - 0x4
    "00000100", -- 5785 - 0x1699  :    4 - 0x4
    "00000100", -- 5786 - 0x169a  :    4 - 0x4
    "00000100", -- 5787 - 0x169b  :    4 - 0x4
    "00000100", -- 5788 - 0x169c  :    4 - 0x4
    "00000100", -- 5789 - 0x169d  :    4 - 0x4
    "00000100", -- 5790 - 0x169e  :    4 - 0x4
    "00000100", -- 5791 - 0x169f  :    4 - 0x4
    "10111100", -- 5792 - 0x16a0  :  188 - 0xbc
    "01011100", -- 5793 - 0x16a1  :   92 - 0x5c
    "10111100", -- 5794 - 0x16a2  :  188 - 0xbc
    "01011100", -- 5795 - 0x16a3  :   92 - 0x5c
    "10111100", -- 5796 - 0x16a4  :  188 - 0xbc
    "01011100", -- 5797 - 0x16a5  :   92 - 0x5c
    "10111100", -- 5798 - 0x16a6  :  188 - 0xbc
    "01011100", -- 5799 - 0x16a7  :   92 - 0x5c
    "01000100", -- 5800 - 0x16a8  :   68 - 0x44
    "10100100", -- 5801 - 0x16a9  :  164 - 0xa4
    "01000100", -- 5802 - 0x16aa  :   68 - 0x44
    "10100100", -- 5803 - 0x16ab  :  164 - 0xa4
    "01000100", -- 5804 - 0x16ac  :   68 - 0x44
    "10100100", -- 5805 - 0x16ad  :  164 - 0xa4
    "01000100", -- 5806 - 0x16ae  :   68 - 0x44
    "10100100", -- 5807 - 0x16af  :  164 - 0xa4
    "00011111", -- 5808 - 0x16b0  :   31 - 0x1f
    "00100000", -- 5809 - 0x16b1  :   32 - 0x20
    "01000000", -- 5810 - 0x16b2  :   64 - 0x40
    "01000000", -- 5811 - 0x16b3  :   64 - 0x40
    "10000000", -- 5812 - 0x16b4  :  128 - 0x80
    "10000000", -- 5813 - 0x16b5  :  128 - 0x80
    "10000000", -- 5814 - 0x16b6  :  128 - 0x80
    "10000001", -- 5815 - 0x16b7  :  129 - 0x81
    "00011111", -- 5816 - 0x16b8  :   31 - 0x1f
    "00111111", -- 5817 - 0x16b9  :   63 - 0x3f
    "01111111", -- 5818 - 0x16ba  :  127 - 0x7f
    "01111111", -- 5819 - 0x16bb  :  127 - 0x7f
    "11111111", -- 5820 - 0x16bc  :  255 - 0xff
    "11111111", -- 5821 - 0x16bd  :  255 - 0xff
    "11111111", -- 5822 - 0x16be  :  255 - 0xff
    "11111110", -- 5823 - 0x16bf  :  254 - 0xfe
    "11111111", -- 5824 - 0x16c0  :  255 - 0xff
    "10000000", -- 5825 - 0x16c1  :  128 - 0x80
    "10000000", -- 5826 - 0x16c2  :  128 - 0x80
    "11000000", -- 5827 - 0x16c3  :  192 - 0xc0
    "11111111", -- 5828 - 0x16c4  :  255 - 0xff
    "11111111", -- 5829 - 0x16c5  :  255 - 0xff
    "11111110", -- 5830 - 0x16c6  :  254 - 0xfe
    "11111110", -- 5831 - 0x16c7  :  254 - 0xfe
    "11111111", -- 5832 - 0x16c8  :  255 - 0xff
    "01111111", -- 5833 - 0x16c9  :  127 - 0x7f
    "01111111", -- 5834 - 0x16ca  :  127 - 0x7f
    "00111111", -- 5835 - 0x16cb  :   63 - 0x3f
    "00000000", -- 5836 - 0x16cc  :    0 - 0x0
    "00000000", -- 5837 - 0x16cd  :    0 - 0x0
    "00000001", -- 5838 - 0x16ce  :    1 - 0x1
    "00000001", -- 5839 - 0x16cf  :    1 - 0x1
    "11111111", -- 5840 - 0x16d0  :  255 - 0xff
    "01111111", -- 5841 - 0x16d1  :  127 - 0x7f
    "01111111", -- 5842 - 0x16d2  :  127 - 0x7f
    "11111111", -- 5843 - 0x16d3  :  255 - 0xff
    "11111111", -- 5844 - 0x16d4  :  255 - 0xff
    "00000111", -- 5845 - 0x16d5  :    7 - 0x7
    "00000011", -- 5846 - 0x16d6  :    3 - 0x3
    "00000011", -- 5847 - 0x16d7  :    3 - 0x3
    "11111111", -- 5848 - 0x16d8  :  255 - 0xff
    "10000000", -- 5849 - 0x16d9  :  128 - 0x80
    "10000000", -- 5850 - 0x16da  :  128 - 0x80
    "00000000", -- 5851 - 0x16db  :    0 - 0x0
    "00000000", -- 5852 - 0x16dc  :    0 - 0x0
    "11111000", -- 5853 - 0x16dd  :  248 - 0xf8
    "11111100", -- 5854 - 0x16de  :  252 - 0xfc
    "11111100", -- 5855 - 0x16df  :  252 - 0xfc
    "11111111", -- 5856 - 0x16e0  :  255 - 0xff
    "00000000", -- 5857 - 0x16e1  :    0 - 0x0
    "00000000", -- 5858 - 0x16e2  :    0 - 0x0
    "00000000", -- 5859 - 0x16e3  :    0 - 0x0
    "00000000", -- 5860 - 0x16e4  :    0 - 0x0
    "10000001", -- 5861 - 0x16e5  :  129 - 0x81
    "11000011", -- 5862 - 0x16e6  :  195 - 0xc3
    "11111111", -- 5863 - 0x16e7  :  255 - 0xff
    "11111111", -- 5864 - 0x16e8  :  255 - 0xff
    "11111111", -- 5865 - 0x16e9  :  255 - 0xff
    "11111111", -- 5866 - 0x16ea  :  255 - 0xff
    "11111111", -- 5867 - 0x16eb  :  255 - 0xff
    "11111111", -- 5868 - 0x16ec  :  255 - 0xff
    "01111110", -- 5869 - 0x16ed  :  126 - 0x7e
    "00111100", -- 5870 - 0x16ee  :   60 - 0x3c
    "00000000", -- 5871 - 0x16ef  :    0 - 0x0
    "11111000", -- 5872 - 0x16f0  :  248 - 0xf8
    "11111100", -- 5873 - 0x16f1  :  252 - 0xfc
    "11111110", -- 5874 - 0x16f2  :  254 - 0xfe
    "11111110", -- 5875 - 0x16f3  :  254 - 0xfe
    "11100011", -- 5876 - 0x16f4  :  227 - 0xe3
    "11000001", -- 5877 - 0x16f5  :  193 - 0xc1
    "10000001", -- 5878 - 0x16f6  :  129 - 0x81
    "10000001", -- 5879 - 0x16f7  :  129 - 0x81
    "11111000", -- 5880 - 0x16f8  :  248 - 0xf8
    "00000100", -- 5881 - 0x16f9  :    4 - 0x4
    "00000010", -- 5882 - 0x16fa  :    2 - 0x2
    "00000010", -- 5883 - 0x16fb  :    2 - 0x2
    "00011101", -- 5884 - 0x16fc  :   29 - 0x1d
    "00111111", -- 5885 - 0x16fd  :   63 - 0x3f
    "01111111", -- 5886 - 0x16fe  :  127 - 0x7f
    "01111111", -- 5887 - 0x16ff  :  127 - 0x7f
    "10000011", -- 5888 - 0x1700  :  131 - 0x83
    "11111111", -- 5889 - 0x1701  :  255 - 0xff
    "11111111", -- 5890 - 0x1702  :  255 - 0xff
    "11111111", -- 5891 - 0x1703  :  255 - 0xff
    "11111111", -- 5892 - 0x1704  :  255 - 0xff
    "11111111", -- 5893 - 0x1705  :  255 - 0xff
    "01111111", -- 5894 - 0x1706  :  127 - 0x7f
    "00011111", -- 5895 - 0x1707  :   31 - 0x1f
    "11111100", -- 5896 - 0x1708  :  252 - 0xfc
    "10000000", -- 5897 - 0x1709  :  128 - 0x80
    "10000000", -- 5898 - 0x170a  :  128 - 0x80
    "10000000", -- 5899 - 0x170b  :  128 - 0x80
    "10000000", -- 5900 - 0x170c  :  128 - 0x80
    "10000000", -- 5901 - 0x170d  :  128 - 0x80
    "01100000", -- 5902 - 0x170e  :   96 - 0x60
    "00011111", -- 5903 - 0x170f  :   31 - 0x1f
    "11111100", -- 5904 - 0x1710  :  252 - 0xfc
    "11111100", -- 5905 - 0x1711  :  252 - 0xfc
    "11111100", -- 5906 - 0x1712  :  252 - 0xfc
    "11111100", -- 5907 - 0x1713  :  252 - 0xfc
    "11111110", -- 5908 - 0x1714  :  254 - 0xfe
    "11111110", -- 5909 - 0x1715  :  254 - 0xfe
    "11111111", -- 5910 - 0x1716  :  255 - 0xff
    "11111111", -- 5911 - 0x1717  :  255 - 0xff
    "00000011", -- 5912 - 0x1718  :    3 - 0x3
    "00000011", -- 5913 - 0x1719  :    3 - 0x3
    "00000011", -- 5914 - 0x171a  :    3 - 0x3
    "00000011", -- 5915 - 0x171b  :    3 - 0x3
    "00000001", -- 5916 - 0x171c  :    1 - 0x1
    "00000001", -- 5917 - 0x171d  :    1 - 0x1
    "00000000", -- 5918 - 0x171e  :    0 - 0x0
    "11111111", -- 5919 - 0x171f  :  255 - 0xff
    "00000001", -- 5920 - 0x1720  :    1 - 0x1
    "00000001", -- 5921 - 0x1721  :    1 - 0x1
    "00000001", -- 5922 - 0x1722  :    1 - 0x1
    "00000001", -- 5923 - 0x1723  :    1 - 0x1
    "00000011", -- 5924 - 0x1724  :    3 - 0x3
    "00000011", -- 5925 - 0x1725  :    3 - 0x3
    "00000111", -- 5926 - 0x1726  :    7 - 0x7
    "11111111", -- 5927 - 0x1727  :  255 - 0xff
    "11111110", -- 5928 - 0x1728  :  254 - 0xfe
    "11111110", -- 5929 - 0x1729  :  254 - 0xfe
    "11111110", -- 5930 - 0x172a  :  254 - 0xfe
    "11111110", -- 5931 - 0x172b  :  254 - 0xfe
    "11111100", -- 5932 - 0x172c  :  252 - 0xfc
    "11111100", -- 5933 - 0x172d  :  252 - 0xfc
    "11111000", -- 5934 - 0x172e  :  248 - 0xf8
    "11111111", -- 5935 - 0x172f  :  255 - 0xff
    "11111111", -- 5936 - 0x1730  :  255 - 0xff
    "11111111", -- 5937 - 0x1731  :  255 - 0xff
    "11111111", -- 5938 - 0x1732  :  255 - 0xff
    "11111111", -- 5939 - 0x1733  :  255 - 0xff
    "11111111", -- 5940 - 0x1734  :  255 - 0xff
    "11111111", -- 5941 - 0x1735  :  255 - 0xff
    "11111111", -- 5942 - 0x1736  :  255 - 0xff
    "11111111", -- 5943 - 0x1737  :  255 - 0xff
    "00000000", -- 5944 - 0x1738  :    0 - 0x0
    "00000000", -- 5945 - 0x1739  :    0 - 0x0
    "00000000", -- 5946 - 0x173a  :    0 - 0x0
    "00000000", -- 5947 - 0x173b  :    0 - 0x0
    "00000000", -- 5948 - 0x173c  :    0 - 0x0
    "00000000", -- 5949 - 0x173d  :    0 - 0x0
    "00000000", -- 5950 - 0x173e  :    0 - 0x0
    "11111111", -- 5951 - 0x173f  :  255 - 0xff
    "10000001", -- 5952 - 0x1740  :  129 - 0x81
    "11000001", -- 5953 - 0x1741  :  193 - 0xc1
    "11100011", -- 5954 - 0x1742  :  227 - 0xe3
    "11111111", -- 5955 - 0x1743  :  255 - 0xff
    "11111111", -- 5956 - 0x1744  :  255 - 0xff
    "11111111", -- 5957 - 0x1745  :  255 - 0xff
    "11111111", -- 5958 - 0x1746  :  255 - 0xff
    "11111110", -- 5959 - 0x1747  :  254 - 0xfe
    "01111111", -- 5960 - 0x1748  :  127 - 0x7f
    "00111111", -- 5961 - 0x1749  :   63 - 0x3f
    "00011101", -- 5962 - 0x174a  :   29 - 0x1d
    "00000001", -- 5963 - 0x174b  :    1 - 0x1
    "00000001", -- 5964 - 0x174c  :    1 - 0x1
    "00000001", -- 5965 - 0x174d  :    1 - 0x1
    "00000011", -- 5966 - 0x174e  :    3 - 0x3
    "11111110", -- 5967 - 0x174f  :  254 - 0xfe
    "11111111", -- 5968 - 0x1750  :  255 - 0xff
    "11111111", -- 5969 - 0x1751  :  255 - 0xff
    "11111111", -- 5970 - 0x1752  :  255 - 0xff
    "11111111", -- 5971 - 0x1753  :  255 - 0xff
    "11111111", -- 5972 - 0x1754  :  255 - 0xff
    "11111011", -- 5973 - 0x1755  :  251 - 0xfb
    "10110101", -- 5974 - 0x1756  :  181 - 0xb5
    "11001110", -- 5975 - 0x1757  :  206 - 0xce
    "10000000", -- 5976 - 0x1758  :  128 - 0x80
    "10000000", -- 5977 - 0x1759  :  128 - 0x80
    "10000000", -- 5978 - 0x175a  :  128 - 0x80
    "10000000", -- 5979 - 0x175b  :  128 - 0x80
    "10000000", -- 5980 - 0x175c  :  128 - 0x80
    "10000100", -- 5981 - 0x175d  :  132 - 0x84
    "11001010", -- 5982 - 0x175e  :  202 - 0xca
    "10110001", -- 5983 - 0x175f  :  177 - 0xb1
    "11111111", -- 5984 - 0x1760  :  255 - 0xff
    "11111111", -- 5985 - 0x1761  :  255 - 0xff
    "11111111", -- 5986 - 0x1762  :  255 - 0xff
    "11111111", -- 5987 - 0x1763  :  255 - 0xff
    "11111111", -- 5988 - 0x1764  :  255 - 0xff
    "11011111", -- 5989 - 0x1765  :  223 - 0xdf
    "10101101", -- 5990 - 0x1766  :  173 - 0xad
    "01110011", -- 5991 - 0x1767  :  115 - 0x73
    "00000001", -- 5992 - 0x1768  :    1 - 0x1
    "00000001", -- 5993 - 0x1769  :    1 - 0x1
    "00000001", -- 5994 - 0x176a  :    1 - 0x1
    "00000001", -- 5995 - 0x176b  :    1 - 0x1
    "00000001", -- 5996 - 0x176c  :    1 - 0x1
    "00100001", -- 5997 - 0x176d  :   33 - 0x21
    "01010011", -- 5998 - 0x176e  :   83 - 0x53
    "10001101", -- 5999 - 0x176f  :  141 - 0x8d
    "01110111", -- 6000 - 0x1770  :  119 - 0x77
    "01110111", -- 6001 - 0x1771  :  119 - 0x77
    "01110111", -- 6002 - 0x1772  :  119 - 0x77
    "01110111", -- 6003 - 0x1773  :  119 - 0x77
    "01110111", -- 6004 - 0x1774  :  119 - 0x77
    "01110111", -- 6005 - 0x1775  :  119 - 0x77
    "01110111", -- 6006 - 0x1776  :  119 - 0x77
    "01110111", -- 6007 - 0x1777  :  119 - 0x77
    "00000000", -- 6008 - 0x1778  :    0 - 0x0
    "00000000", -- 6009 - 0x1779  :    0 - 0x0
    "00000000", -- 6010 - 0x177a  :    0 - 0x0
    "00000000", -- 6011 - 0x177b  :    0 - 0x0
    "01110111", -- 6012 - 0x177c  :  119 - 0x77
    "11111111", -- 6013 - 0x177d  :  255 - 0xff
    "11111111", -- 6014 - 0x177e  :  255 - 0xff
    "11111111", -- 6015 - 0x177f  :  255 - 0xff
    "00000000", -- 6016 - 0x1780  :    0 - 0x0
    "00000000", -- 6017 - 0x1781  :    0 - 0x0
    "00000000", -- 6018 - 0x1782  :    0 - 0x0
    "00000000", -- 6019 - 0x1783  :    0 - 0x0
    "00000000", -- 6020 - 0x1784  :    0 - 0x0
    "00000000", -- 6021 - 0x1785  :    0 - 0x0
    "00000000", -- 6022 - 0x1786  :    0 - 0x0
    "11111111", -- 6023 - 0x1787  :  255 - 0xff
    "11111111", -- 6024 - 0x1788  :  255 - 0xff
    "11111111", -- 6025 - 0x1789  :  255 - 0xff
    "11111111", -- 6026 - 0x178a  :  255 - 0xff
    "11111111", -- 6027 - 0x178b  :  255 - 0xff
    "11111111", -- 6028 - 0x178c  :  255 - 0xff
    "11111111", -- 6029 - 0x178d  :  255 - 0xff
    "11111111", -- 6030 - 0x178e  :  255 - 0xff
    "11111111", -- 6031 - 0x178f  :  255 - 0xff
    "01110111", -- 6032 - 0x1790  :  119 - 0x77
    "01110111", -- 6033 - 0x1791  :  119 - 0x77
    "01110111", -- 6034 - 0x1792  :  119 - 0x77
    "01110111", -- 6035 - 0x1793  :  119 - 0x77
    "00000000", -- 6036 - 0x1794  :    0 - 0x0
    "00000000", -- 6037 - 0x1795  :    0 - 0x0
    "00000000", -- 6038 - 0x1796  :    0 - 0x0
    "00000000", -- 6039 - 0x1797  :    0 - 0x0
    "11111111", -- 6040 - 0x1798  :  255 - 0xff
    "11111111", -- 6041 - 0x1799  :  255 - 0xff
    "11111111", -- 6042 - 0x179a  :  255 - 0xff
    "01110111", -- 6043 - 0x179b  :  119 - 0x77
    "01110111", -- 6044 - 0x179c  :  119 - 0x77
    "01110111", -- 6045 - 0x179d  :  119 - 0x77
    "01110111", -- 6046 - 0x179e  :  119 - 0x77
    "01110111", -- 6047 - 0x179f  :  119 - 0x77
    "00000001", -- 6048 - 0x17a0  :    1 - 0x1
    "00000001", -- 6049 - 0x17a1  :    1 - 0x1
    "00000001", -- 6050 - 0x17a2  :    1 - 0x1
    "00011001", -- 6051 - 0x17a3  :   25 - 0x19
    "00011101", -- 6052 - 0x17a4  :   29 - 0x1d
    "00001101", -- 6053 - 0x17a5  :   13 - 0xd
    "00000001", -- 6054 - 0x17a6  :    1 - 0x1
    "11111110", -- 6055 - 0x17a7  :  254 - 0xfe
    "11111111", -- 6056 - 0x17a8  :  255 - 0xff
    "11111111", -- 6057 - 0x17a9  :  255 - 0xff
    "11111111", -- 6058 - 0x17aa  :  255 - 0xff
    "11100111", -- 6059 - 0x17ab  :  231 - 0xe7
    "11100111", -- 6060 - 0x17ac  :  231 - 0xe7
    "11111111", -- 6061 - 0x17ad  :  255 - 0xff
    "11111111", -- 6062 - 0x17ae  :  255 - 0xff
    "11111110", -- 6063 - 0x17af  :  254 - 0xfe
    "00100000", -- 6064 - 0x17b0  :   32 - 0x20
    "01111000", -- 6065 - 0x17b1  :  120 - 0x78
    "01111111", -- 6066 - 0x17b2  :  127 - 0x7f
    "11111110", -- 6067 - 0x17b3  :  254 - 0xfe
    "11111110", -- 6068 - 0x17b4  :  254 - 0xfe
    "11111110", -- 6069 - 0x17b5  :  254 - 0xfe
    "11111110", -- 6070 - 0x17b6  :  254 - 0xfe
    "11111110", -- 6071 - 0x17b7  :  254 - 0xfe
    "00000000", -- 6072 - 0x17b8  :    0 - 0x0
    "00100001", -- 6073 - 0x17b9  :   33 - 0x21
    "00100001", -- 6074 - 0x17ba  :   33 - 0x21
    "01000001", -- 6075 - 0x17bb  :   65 - 0x41
    "01000001", -- 6076 - 0x17bc  :   65 - 0x41
    "01000001", -- 6077 - 0x17bd  :   65 - 0x41
    "01000001", -- 6078 - 0x17be  :   65 - 0x41
    "01000001", -- 6079 - 0x17bf  :   65 - 0x41
    "00000100", -- 6080 - 0x17c0  :    4 - 0x4
    "10011010", -- 6081 - 0x17c1  :  154 - 0x9a
    "11111010", -- 6082 - 0x17c2  :  250 - 0xfa
    "11111101", -- 6083 - 0x17c3  :  253 - 0xfd
    "11111101", -- 6084 - 0x17c4  :  253 - 0xfd
    "11111101", -- 6085 - 0x17c5  :  253 - 0xfd
    "11111101", -- 6086 - 0x17c6  :  253 - 0xfd
    "11111101", -- 6087 - 0x17c7  :  253 - 0xfd
    "00000000", -- 6088 - 0x17c8  :    0 - 0x0
    "10000000", -- 6089 - 0x17c9  :  128 - 0x80
    "10000000", -- 6090 - 0x17ca  :  128 - 0x80
    "10000000", -- 6091 - 0x17cb  :  128 - 0x80
    "10000000", -- 6092 - 0x17cc  :  128 - 0x80
    "10000000", -- 6093 - 0x17cd  :  128 - 0x80
    "10000000", -- 6094 - 0x17ce  :  128 - 0x80
    "10000000", -- 6095 - 0x17cf  :  128 - 0x80
    "01111110", -- 6096 - 0x17d0  :  126 - 0x7e
    "00111000", -- 6097 - 0x17d1  :   56 - 0x38
    "00100001", -- 6098 - 0x17d2  :   33 - 0x21
    "00000000", -- 6099 - 0x17d3  :    0 - 0x0
    "00000001", -- 6100 - 0x17d4  :    1 - 0x1
    "00000000", -- 6101 - 0x17d5  :    0 - 0x0
    "00000001", -- 6102 - 0x17d6  :    1 - 0x1
    "00000000", -- 6103 - 0x17d7  :    0 - 0x0
    "00100001", -- 6104 - 0x17d8  :   33 - 0x21
    "00100001", -- 6105 - 0x17d9  :   33 - 0x21
    "00000001", -- 6106 - 0x17da  :    1 - 0x1
    "00000001", -- 6107 - 0x17db  :    1 - 0x1
    "00000001", -- 6108 - 0x17dc  :    1 - 0x1
    "00000001", -- 6109 - 0x17dd  :    1 - 0x1
    "00000001", -- 6110 - 0x17de  :    1 - 0x1
    "00000001", -- 6111 - 0x17df  :    1 - 0x1
    "11111010", -- 6112 - 0x17e0  :  250 - 0xfa
    "10001010", -- 6113 - 0x17e1  :  138 - 0x8a
    "10000100", -- 6114 - 0x17e2  :  132 - 0x84
    "10000000", -- 6115 - 0x17e3  :  128 - 0x80
    "10000000", -- 6116 - 0x17e4  :  128 - 0x80
    "10000000", -- 6117 - 0x17e5  :  128 - 0x80
    "10000000", -- 6118 - 0x17e6  :  128 - 0x80
    "10000000", -- 6119 - 0x17e7  :  128 - 0x80
    "10000000", -- 6120 - 0x17e8  :  128 - 0x80
    "10000000", -- 6121 - 0x17e9  :  128 - 0x80
    "10000000", -- 6122 - 0x17ea  :  128 - 0x80
    "10000000", -- 6123 - 0x17eb  :  128 - 0x80
    "10000000", -- 6124 - 0x17ec  :  128 - 0x80
    "10000000", -- 6125 - 0x17ed  :  128 - 0x80
    "10000000", -- 6126 - 0x17ee  :  128 - 0x80
    "10000000", -- 6127 - 0x17ef  :  128 - 0x80
    "00000010", -- 6128 - 0x17f0  :    2 - 0x2
    "00000100", -- 6129 - 0x17f1  :    4 - 0x4
    "00000000", -- 6130 - 0x17f2  :    0 - 0x0
    "00010000", -- 6131 - 0x17f3  :   16 - 0x10
    "00000000", -- 6132 - 0x17f4  :    0 - 0x0
    "01000000", -- 6133 - 0x17f5  :   64 - 0x40
    "10000000", -- 6134 - 0x17f6  :  128 - 0x80
    "00000000", -- 6135 - 0x17f7  :    0 - 0x0
    "00000001", -- 6136 - 0x17f8  :    1 - 0x1
    "00000001", -- 6137 - 0x17f9  :    1 - 0x1
    "00000110", -- 6138 - 0x17fa  :    6 - 0x6
    "00001000", -- 6139 - 0x17fb  :    8 - 0x8
    "00011000", -- 6140 - 0x17fc  :   24 - 0x18
    "00100000", -- 6141 - 0x17fd  :   32 - 0x20
    "00100000", -- 6142 - 0x17fe  :   32 - 0x20
    "11000000", -- 6143 - 0x17ff  :  192 - 0xc0
    "00001011", -- 6144 - 0x1800  :   11 - 0xb
    "00001011", -- 6145 - 0x1801  :   11 - 0xb
    "00111011", -- 6146 - 0x1802  :   59 - 0x3b
    "00001011", -- 6147 - 0x1803  :   11 - 0xb
    "11111011", -- 6148 - 0x1804  :  251 - 0xfb
    "00001011", -- 6149 - 0x1805  :   11 - 0xb
    "00001011", -- 6150 - 0x1806  :   11 - 0xb
    "00001010", -- 6151 - 0x1807  :   10 - 0xa
    "00000100", -- 6152 - 0x1808  :    4 - 0x4
    "00000100", -- 6153 - 0x1809  :    4 - 0x4
    "11000100", -- 6154 - 0x180a  :  196 - 0xc4
    "11110100", -- 6155 - 0x180b  :  244 - 0xf4
    "11110100", -- 6156 - 0x180c  :  244 - 0xf4
    "00000100", -- 6157 - 0x180d  :    4 - 0x4
    "00000100", -- 6158 - 0x180e  :    4 - 0x4
    "00000101", -- 6159 - 0x180f  :    5 - 0x5
    "10010000", -- 6160 - 0x1810  :  144 - 0x90
    "00010000", -- 6161 - 0x1811  :   16 - 0x10
    "00011111", -- 6162 - 0x1812  :   31 - 0x1f
    "00010000", -- 6163 - 0x1813  :   16 - 0x10
    "00011111", -- 6164 - 0x1814  :   31 - 0x1f
    "00010000", -- 6165 - 0x1815  :   16 - 0x10
    "00010000", -- 6166 - 0x1816  :   16 - 0x10
    "10010000", -- 6167 - 0x1817  :  144 - 0x90
    "01110000", -- 6168 - 0x1818  :  112 - 0x70
    "11110000", -- 6169 - 0x1819  :  240 - 0xf0
    "11110000", -- 6170 - 0x181a  :  240 - 0xf0
    "11111111", -- 6171 - 0x181b  :  255 - 0xff
    "11111111", -- 6172 - 0x181c  :  255 - 0xff
    "11110000", -- 6173 - 0x181d  :  240 - 0xf0
    "11110000", -- 6174 - 0x181e  :  240 - 0xf0
    "01110000", -- 6175 - 0x181f  :  112 - 0x70
    "00111111", -- 6176 - 0x1820  :   63 - 0x3f
    "01111000", -- 6177 - 0x1821  :  120 - 0x78
    "11100111", -- 6178 - 0x1822  :  231 - 0xe7
    "11001111", -- 6179 - 0x1823  :  207 - 0xcf
    "01011000", -- 6180 - 0x1824  :   88 - 0x58
    "01011000", -- 6181 - 0x1825  :   88 - 0x58
    "01010000", -- 6182 - 0x1826  :   80 - 0x50
    "10010000", -- 6183 - 0x1827  :  144 - 0x90
    "11000000", -- 6184 - 0x1828  :  192 - 0xc0
    "10000111", -- 6185 - 0x1829  :  135 - 0x87
    "00011000", -- 6186 - 0x182a  :   24 - 0x18
    "10110000", -- 6187 - 0x182b  :  176 - 0xb0
    "11100111", -- 6188 - 0x182c  :  231 - 0xe7
    "11100111", -- 6189 - 0x182d  :  231 - 0xe7
    "11101111", -- 6190 - 0x182e  :  239 - 0xef
    "11101111", -- 6191 - 0x182f  :  239 - 0xef
    "10110000", -- 6192 - 0x1830  :  176 - 0xb0
    "11111100", -- 6193 - 0x1831  :  252 - 0xfc
    "11100010", -- 6194 - 0x1832  :  226 - 0xe2
    "11000001", -- 6195 - 0x1833  :  193 - 0xc1
    "11000001", -- 6196 - 0x1834  :  193 - 0xc1
    "10000011", -- 6197 - 0x1835  :  131 - 0x83
    "10001111", -- 6198 - 0x1836  :  143 - 0x8f
    "01111110", -- 6199 - 0x1837  :  126 - 0x7e
    "01101111", -- 6200 - 0x1838  :  111 - 0x6f
    "01000011", -- 6201 - 0x1839  :   67 - 0x43
    "01011101", -- 6202 - 0x183a  :   93 - 0x5d
    "00111111", -- 6203 - 0x183b  :   63 - 0x3f
    "00111111", -- 6204 - 0x183c  :   63 - 0x3f
    "01111111", -- 6205 - 0x183d  :  127 - 0x7f
    "01111111", -- 6206 - 0x183e  :  127 - 0x7f
    "11111111", -- 6207 - 0x183f  :  255 - 0xff
    "11111110", -- 6208 - 0x1840  :  254 - 0xfe
    "00000011", -- 6209 - 0x1841  :    3 - 0x3
    "00001111", -- 6210 - 0x1842  :   15 - 0xf
    "10010001", -- 6211 - 0x1843  :  145 - 0x91
    "01110000", -- 6212 - 0x1844  :  112 - 0x70
    "01100000", -- 6213 - 0x1845  :   96 - 0x60
    "00100000", -- 6214 - 0x1846  :   32 - 0x20
    "00110001", -- 6215 - 0x1847  :   49 - 0x31
    "00000011", -- 6216 - 0x1848  :    3 - 0x3
    "11111111", -- 6217 - 0x1849  :  255 - 0xff
    "11110001", -- 6218 - 0x184a  :  241 - 0xf1
    "01101110", -- 6219 - 0x184b  :  110 - 0x6e
    "11001111", -- 6220 - 0x184c  :  207 - 0xcf
    "11011111", -- 6221 - 0x184d  :  223 - 0xdf
    "11111111", -- 6222 - 0x184e  :  255 - 0xff
    "11111111", -- 6223 - 0x184f  :  255 - 0xff
    "00111111", -- 6224 - 0x1850  :   63 - 0x3f
    "00111111", -- 6225 - 0x1851  :   63 - 0x3f
    "00011101", -- 6226 - 0x1852  :   29 - 0x1d
    "00111001", -- 6227 - 0x1853  :   57 - 0x39
    "01111011", -- 6228 - 0x1854  :  123 - 0x7b
    "11110011", -- 6229 - 0x1855  :  243 - 0xf3
    "10000110", -- 6230 - 0x1856  :  134 - 0x86
    "11111110", -- 6231 - 0x1857  :  254 - 0xfe
    "11111101", -- 6232 - 0x1858  :  253 - 0xfd
    "11111011", -- 6233 - 0x1859  :  251 - 0xfb
    "11111011", -- 6234 - 0x185a  :  251 - 0xfb
    "11110111", -- 6235 - 0x185b  :  247 - 0xf7
    "11110111", -- 6236 - 0x185c  :  247 - 0xf7
    "00001111", -- 6237 - 0x185d  :   15 - 0xf
    "01111111", -- 6238 - 0x185e  :  127 - 0x7f
    "11111111", -- 6239 - 0x185f  :  255 - 0xff
    "11111111", -- 6240 - 0x1860  :  255 - 0xff
    "11111111", -- 6241 - 0x1861  :  255 - 0xff
    "11111111", -- 6242 - 0x1862  :  255 - 0xff
    "11111111", -- 6243 - 0x1863  :  255 - 0xff
    "11111111", -- 6244 - 0x1864  :  255 - 0xff
    "10000000", -- 6245 - 0x1865  :  128 - 0x80
    "10000000", -- 6246 - 0x1866  :  128 - 0x80
    "11111111", -- 6247 - 0x1867  :  255 - 0xff
    "11111111", -- 6248 - 0x1868  :  255 - 0xff
    "10000000", -- 6249 - 0x1869  :  128 - 0x80
    "10000000", -- 6250 - 0x186a  :  128 - 0x80
    "10000000", -- 6251 - 0x186b  :  128 - 0x80
    "10000000", -- 6252 - 0x186c  :  128 - 0x80
    "11111111", -- 6253 - 0x186d  :  255 - 0xff
    "11111111", -- 6254 - 0x186e  :  255 - 0xff
    "10000000", -- 6255 - 0x186f  :  128 - 0x80
    "11111110", -- 6256 - 0x1870  :  254 - 0xfe
    "11111111", -- 6257 - 0x1871  :  255 - 0xff
    "11111111", -- 6258 - 0x1872  :  255 - 0xff
    "11111111", -- 6259 - 0x1873  :  255 - 0xff
    "11111111", -- 6260 - 0x1874  :  255 - 0xff
    "00000011", -- 6261 - 0x1875  :    3 - 0x3
    "00000011", -- 6262 - 0x1876  :    3 - 0x3
    "11111111", -- 6263 - 0x1877  :  255 - 0xff
    "11111110", -- 6264 - 0x1878  :  254 - 0xfe
    "00000011", -- 6265 - 0x1879  :    3 - 0x3
    "00000011", -- 6266 - 0x187a  :    3 - 0x3
    "00000011", -- 6267 - 0x187b  :    3 - 0x3
    "00000011", -- 6268 - 0x187c  :    3 - 0x3
    "11111111", -- 6269 - 0x187d  :  255 - 0xff
    "11111111", -- 6270 - 0x187e  :  255 - 0xff
    "00000011", -- 6271 - 0x187f  :    3 - 0x3
    "00000000", -- 6272 - 0x1880  :    0 - 0x0
    "11111111", -- 6273 - 0x1881  :  255 - 0xff
    "11111111", -- 6274 - 0x1882  :  255 - 0xff
    "11111111", -- 6275 - 0x1883  :  255 - 0xff
    "11111111", -- 6276 - 0x1884  :  255 - 0xff
    "11111111", -- 6277 - 0x1885  :  255 - 0xff
    "00000000", -- 6278 - 0x1886  :    0 - 0x0
    "00000000", -- 6279 - 0x1887  :    0 - 0x0
    "00000000", -- 6280 - 0x1888  :    0 - 0x0
    "11111111", -- 6281 - 0x1889  :  255 - 0xff
    "00000000", -- 6282 - 0x188a  :    0 - 0x0
    "00000000", -- 6283 - 0x188b  :    0 - 0x0
    "00000000", -- 6284 - 0x188c  :    0 - 0x0
    "00000000", -- 6285 - 0x188d  :    0 - 0x0
    "11111111", -- 6286 - 0x188e  :  255 - 0xff
    "11111111", -- 6287 - 0x188f  :  255 - 0xff
    "00111100", -- 6288 - 0x1890  :   60 - 0x3c
    "11111100", -- 6289 - 0x1891  :  252 - 0xfc
    "11111100", -- 6290 - 0x1892  :  252 - 0xfc
    "11111100", -- 6291 - 0x1893  :  252 - 0xfc
    "11111100", -- 6292 - 0x1894  :  252 - 0xfc
    "11111100", -- 6293 - 0x1895  :  252 - 0xfc
    "00000100", -- 6294 - 0x1896  :    4 - 0x4
    "00000100", -- 6295 - 0x1897  :    4 - 0x4
    "00100011", -- 6296 - 0x1898  :   35 - 0x23
    "11110011", -- 6297 - 0x1899  :  243 - 0xf3
    "00001011", -- 6298 - 0x189a  :   11 - 0xb
    "00001011", -- 6299 - 0x189b  :   11 - 0xb
    "00001011", -- 6300 - 0x189c  :   11 - 0xb
    "00000111", -- 6301 - 0x189d  :    7 - 0x7
    "11111111", -- 6302 - 0x189e  :  255 - 0xff
    "11111111", -- 6303 - 0x189f  :  255 - 0xff
    "11111111", -- 6304 - 0x18a0  :  255 - 0xff
    "11111111", -- 6305 - 0x18a1  :  255 - 0xff
    "11111111", -- 6306 - 0x18a2  :  255 - 0xff
    "11111111", -- 6307 - 0x18a3  :  255 - 0xff
    "10000000", -- 6308 - 0x18a4  :  128 - 0x80
    "11111111", -- 6309 - 0x18a5  :  255 - 0xff
    "11111111", -- 6310 - 0x18a6  :  255 - 0xff
    "11111111", -- 6311 - 0x18a7  :  255 - 0xff
    "10000000", -- 6312 - 0x18a8  :  128 - 0x80
    "10000000", -- 6313 - 0x18a9  :  128 - 0x80
    "10000000", -- 6314 - 0x18aa  :  128 - 0x80
    "10000000", -- 6315 - 0x18ab  :  128 - 0x80
    "11111111", -- 6316 - 0x18ac  :  255 - 0xff
    "10000000", -- 6317 - 0x18ad  :  128 - 0x80
    "10000000", -- 6318 - 0x18ae  :  128 - 0x80
    "10000000", -- 6319 - 0x18af  :  128 - 0x80
    "11111111", -- 6320 - 0x18b0  :  255 - 0xff
    "11111111", -- 6321 - 0x18b1  :  255 - 0xff
    "11111111", -- 6322 - 0x18b2  :  255 - 0xff
    "11111111", -- 6323 - 0x18b3  :  255 - 0xff
    "00000011", -- 6324 - 0x18b4  :    3 - 0x3
    "11111111", -- 6325 - 0x18b5  :  255 - 0xff
    "11111111", -- 6326 - 0x18b6  :  255 - 0xff
    "11111111", -- 6327 - 0x18b7  :  255 - 0xff
    "00000011", -- 6328 - 0x18b8  :    3 - 0x3
    "00000011", -- 6329 - 0x18b9  :    3 - 0x3
    "00000011", -- 6330 - 0x18ba  :    3 - 0x3
    "00000011", -- 6331 - 0x18bb  :    3 - 0x3
    "11111111", -- 6332 - 0x18bc  :  255 - 0xff
    "00000011", -- 6333 - 0x18bd  :    3 - 0x3
    "00000011", -- 6334 - 0x18be  :    3 - 0x3
    "00000011", -- 6335 - 0x18bf  :    3 - 0x3
    "11111111", -- 6336 - 0x18c0  :  255 - 0xff
    "11111111", -- 6337 - 0x18c1  :  255 - 0xff
    "11111111", -- 6338 - 0x18c2  :  255 - 0xff
    "11111111", -- 6339 - 0x18c3  :  255 - 0xff
    "11111111", -- 6340 - 0x18c4  :  255 - 0xff
    "00000000", -- 6341 - 0x18c5  :    0 - 0x0
    "11111111", -- 6342 - 0x18c6  :  255 - 0xff
    "11111111", -- 6343 - 0x18c7  :  255 - 0xff
    "00000000", -- 6344 - 0x18c8  :    0 - 0x0
    "00000000", -- 6345 - 0x18c9  :    0 - 0x0
    "00000000", -- 6346 - 0x18ca  :    0 - 0x0
    "00000000", -- 6347 - 0x18cb  :    0 - 0x0
    "00000000", -- 6348 - 0x18cc  :    0 - 0x0
    "11111111", -- 6349 - 0x18cd  :  255 - 0xff
    "00000000", -- 6350 - 0x18ce  :    0 - 0x0
    "00000000", -- 6351 - 0x18cf  :    0 - 0x0
    "11111100", -- 6352 - 0x18d0  :  252 - 0xfc
    "11111100", -- 6353 - 0x18d1  :  252 - 0xfc
    "11111110", -- 6354 - 0x18d2  :  254 - 0xfe
    "11111110", -- 6355 - 0x18d3  :  254 - 0xfe
    "11111110", -- 6356 - 0x18d4  :  254 - 0xfe
    "00000010", -- 6357 - 0x18d5  :    2 - 0x2
    "11111110", -- 6358 - 0x18d6  :  254 - 0xfe
    "11111110", -- 6359 - 0x18d7  :  254 - 0xfe
    "00000111", -- 6360 - 0x18d8  :    7 - 0x7
    "00000111", -- 6361 - 0x18d9  :    7 - 0x7
    "00000011", -- 6362 - 0x18da  :    3 - 0x3
    "00000011", -- 6363 - 0x18db  :    3 - 0x3
    "00000011", -- 6364 - 0x18dc  :    3 - 0x3
    "11111111", -- 6365 - 0x18dd  :  255 - 0xff
    "00000011", -- 6366 - 0x18de  :    3 - 0x3
    "00000011", -- 6367 - 0x18df  :    3 - 0x3
    "11111111", -- 6368 - 0x18e0  :  255 - 0xff
    "10000000", -- 6369 - 0x18e1  :  128 - 0x80
    "10000000", -- 6370 - 0x18e2  :  128 - 0x80
    "10000000", -- 6371 - 0x18e3  :  128 - 0x80
    "10000000", -- 6372 - 0x18e4  :  128 - 0x80
    "10000000", -- 6373 - 0x18e5  :  128 - 0x80
    "10000000", -- 6374 - 0x18e6  :  128 - 0x80
    "10000000", -- 6375 - 0x18e7  :  128 - 0x80
    "10000000", -- 6376 - 0x18e8  :  128 - 0x80
    "11111111", -- 6377 - 0x18e9  :  255 - 0xff
    "11111111", -- 6378 - 0x18ea  :  255 - 0xff
    "11111111", -- 6379 - 0x18eb  :  255 - 0xff
    "11111111", -- 6380 - 0x18ec  :  255 - 0xff
    "11111111", -- 6381 - 0x18ed  :  255 - 0xff
    "11111111", -- 6382 - 0x18ee  :  255 - 0xff
    "11111111", -- 6383 - 0x18ef  :  255 - 0xff
    "11111111", -- 6384 - 0x18f0  :  255 - 0xff
    "00000011", -- 6385 - 0x18f1  :    3 - 0x3
    "00000011", -- 6386 - 0x18f2  :    3 - 0x3
    "00000011", -- 6387 - 0x18f3  :    3 - 0x3
    "00000011", -- 6388 - 0x18f4  :    3 - 0x3
    "00000011", -- 6389 - 0x18f5  :    3 - 0x3
    "00000011", -- 6390 - 0x18f6  :    3 - 0x3
    "00000011", -- 6391 - 0x18f7  :    3 - 0x3
    "00000011", -- 6392 - 0x18f8  :    3 - 0x3
    "11111111", -- 6393 - 0x18f9  :  255 - 0xff
    "11111111", -- 6394 - 0x18fa  :  255 - 0xff
    "11111111", -- 6395 - 0x18fb  :  255 - 0xff
    "11111111", -- 6396 - 0x18fc  :  255 - 0xff
    "11111111", -- 6397 - 0x18fd  :  255 - 0xff
    "11111111", -- 6398 - 0x18fe  :  255 - 0xff
    "11111111", -- 6399 - 0x18ff  :  255 - 0xff
    "00000010", -- 6400 - 0x1900  :    2 - 0x2
    "00000010", -- 6401 - 0x1901  :    2 - 0x2
    "00000010", -- 6402 - 0x1902  :    2 - 0x2
    "00000010", -- 6403 - 0x1903  :    2 - 0x2
    "00000010", -- 6404 - 0x1904  :    2 - 0x2
    "00000010", -- 6405 - 0x1905  :    2 - 0x2
    "00000100", -- 6406 - 0x1906  :    4 - 0x4
    "00000100", -- 6407 - 0x1907  :    4 - 0x4
    "11111111", -- 6408 - 0x1908  :  255 - 0xff
    "11111111", -- 6409 - 0x1909  :  255 - 0xff
    "11111111", -- 6410 - 0x190a  :  255 - 0xff
    "11111111", -- 6411 - 0x190b  :  255 - 0xff
    "11111111", -- 6412 - 0x190c  :  255 - 0xff
    "11111111", -- 6413 - 0x190d  :  255 - 0xff
    "11111111", -- 6414 - 0x190e  :  255 - 0xff
    "11111111", -- 6415 - 0x190f  :  255 - 0xff
    "10000000", -- 6416 - 0x1910  :  128 - 0x80
    "10000000", -- 6417 - 0x1911  :  128 - 0x80
    "10101010", -- 6418 - 0x1912  :  170 - 0xaa
    "11010101", -- 6419 - 0x1913  :  213 - 0xd5
    "10101010", -- 6420 - 0x1914  :  170 - 0xaa
    "11111111", -- 6421 - 0x1915  :  255 - 0xff
    "11111111", -- 6422 - 0x1916  :  255 - 0xff
    "11111111", -- 6423 - 0x1917  :  255 - 0xff
    "11111111", -- 6424 - 0x1918  :  255 - 0xff
    "11111111", -- 6425 - 0x1919  :  255 - 0xff
    "11010101", -- 6426 - 0x191a  :  213 - 0xd5
    "10101010", -- 6427 - 0x191b  :  170 - 0xaa
    "11010101", -- 6428 - 0x191c  :  213 - 0xd5
    "10000000", -- 6429 - 0x191d  :  128 - 0x80
    "10000000", -- 6430 - 0x191e  :  128 - 0x80
    "11111111", -- 6431 - 0x191f  :  255 - 0xff
    "00000011", -- 6432 - 0x1920  :    3 - 0x3
    "00000011", -- 6433 - 0x1921  :    3 - 0x3
    "10101011", -- 6434 - 0x1922  :  171 - 0xab
    "01010111", -- 6435 - 0x1923  :   87 - 0x57
    "10101011", -- 6436 - 0x1924  :  171 - 0xab
    "11111111", -- 6437 - 0x1925  :  255 - 0xff
    "11111111", -- 6438 - 0x1926  :  255 - 0xff
    "11111110", -- 6439 - 0x1927  :  254 - 0xfe
    "11111111", -- 6440 - 0x1928  :  255 - 0xff
    "11111111", -- 6441 - 0x1929  :  255 - 0xff
    "01010111", -- 6442 - 0x192a  :   87 - 0x57
    "10101011", -- 6443 - 0x192b  :  171 - 0xab
    "01010111", -- 6444 - 0x192c  :   87 - 0x57
    "00000011", -- 6445 - 0x192d  :    3 - 0x3
    "00000011", -- 6446 - 0x192e  :    3 - 0x3
    "11111110", -- 6447 - 0x192f  :  254 - 0xfe
    "00000000", -- 6448 - 0x1930  :    0 - 0x0
    "01010101", -- 6449 - 0x1931  :   85 - 0x55
    "10101010", -- 6450 - 0x1932  :  170 - 0xaa
    "01010101", -- 6451 - 0x1933  :   85 - 0x55
    "11111111", -- 6452 - 0x1934  :  255 - 0xff
    "11111111", -- 6453 - 0x1935  :  255 - 0xff
    "11111111", -- 6454 - 0x1936  :  255 - 0xff
    "00000000", -- 6455 - 0x1937  :    0 - 0x0
    "11111111", -- 6456 - 0x1938  :  255 - 0xff
    "10101010", -- 6457 - 0x1939  :  170 - 0xaa
    "01010101", -- 6458 - 0x193a  :   85 - 0x55
    "10101010", -- 6459 - 0x193b  :  170 - 0xaa
    "00000000", -- 6460 - 0x193c  :    0 - 0x0
    "00000000", -- 6461 - 0x193d  :    0 - 0x0
    "11111111", -- 6462 - 0x193e  :  255 - 0xff
    "00000000", -- 6463 - 0x193f  :    0 - 0x0
    "00000100", -- 6464 - 0x1940  :    4 - 0x4
    "01010100", -- 6465 - 0x1941  :   84 - 0x54
    "10101100", -- 6466 - 0x1942  :  172 - 0xac
    "01011100", -- 6467 - 0x1943  :   92 - 0x5c
    "11111100", -- 6468 - 0x1944  :  252 - 0xfc
    "11111100", -- 6469 - 0x1945  :  252 - 0xfc
    "11111100", -- 6470 - 0x1946  :  252 - 0xfc
    "00111100", -- 6471 - 0x1947  :   60 - 0x3c
    "11111111", -- 6472 - 0x1948  :  255 - 0xff
    "10101111", -- 6473 - 0x1949  :  175 - 0xaf
    "01010111", -- 6474 - 0x194a  :   87 - 0x57
    "10101011", -- 6475 - 0x194b  :  171 - 0xab
    "00001011", -- 6476 - 0x194c  :   11 - 0xb
    "00001011", -- 6477 - 0x194d  :   11 - 0xb
    "11110011", -- 6478 - 0x194e  :  243 - 0xf3
    "00100011", -- 6479 - 0x194f  :   35 - 0x23
    "00111111", -- 6480 - 0x1950  :   63 - 0x3f
    "00111111", -- 6481 - 0x1951  :   63 - 0x3f
    "00111111", -- 6482 - 0x1952  :   63 - 0x3f
    "00111111", -- 6483 - 0x1953  :   63 - 0x3f
    "00000000", -- 6484 - 0x1954  :    0 - 0x0
    "00000000", -- 6485 - 0x1955  :    0 - 0x0
    "00000000", -- 6486 - 0x1956  :    0 - 0x0
    "11111111", -- 6487 - 0x1957  :  255 - 0xff
    "11111111", -- 6488 - 0x1958  :  255 - 0xff
    "11111111", -- 6489 - 0x1959  :  255 - 0xff
    "11111111", -- 6490 - 0x195a  :  255 - 0xff
    "11111111", -- 6491 - 0x195b  :  255 - 0xff
    "11111111", -- 6492 - 0x195c  :  255 - 0xff
    "11111111", -- 6493 - 0x195d  :  255 - 0xff
    "11111111", -- 6494 - 0x195e  :  255 - 0xff
    "11111111", -- 6495 - 0x195f  :  255 - 0xff
    "01111110", -- 6496 - 0x1960  :  126 - 0x7e
    "01111100", -- 6497 - 0x1961  :  124 - 0x7c
    "01111100", -- 6498 - 0x1962  :  124 - 0x7c
    "01111000", -- 6499 - 0x1963  :  120 - 0x78
    "00000000", -- 6500 - 0x1964  :    0 - 0x0
    "00000000", -- 6501 - 0x1965  :    0 - 0x0
    "00000000", -- 6502 - 0x1966  :    0 - 0x0
    "11111111", -- 6503 - 0x1967  :  255 - 0xff
    "11111111", -- 6504 - 0x1968  :  255 - 0xff
    "11111111", -- 6505 - 0x1969  :  255 - 0xff
    "11111111", -- 6506 - 0x196a  :  255 - 0xff
    "11111111", -- 6507 - 0x196b  :  255 - 0xff
    "11111111", -- 6508 - 0x196c  :  255 - 0xff
    "11111111", -- 6509 - 0x196d  :  255 - 0xff
    "11111111", -- 6510 - 0x196e  :  255 - 0xff
    "11111111", -- 6511 - 0x196f  :  255 - 0xff
    "00011111", -- 6512 - 0x1970  :   31 - 0x1f
    "00001111", -- 6513 - 0x1971  :   15 - 0xf
    "00001111", -- 6514 - 0x1972  :   15 - 0xf
    "00000111", -- 6515 - 0x1973  :    7 - 0x7
    "00000000", -- 6516 - 0x1974  :    0 - 0x0
    "00000000", -- 6517 - 0x1975  :    0 - 0x0
    "00000000", -- 6518 - 0x1976  :    0 - 0x0
    "11111111", -- 6519 - 0x1977  :  255 - 0xff
    "11111111", -- 6520 - 0x1978  :  255 - 0xff
    "11111111", -- 6521 - 0x1979  :  255 - 0xff
    "11111111", -- 6522 - 0x197a  :  255 - 0xff
    "11111111", -- 6523 - 0x197b  :  255 - 0xff
    "11111111", -- 6524 - 0x197c  :  255 - 0xff
    "11111111", -- 6525 - 0x197d  :  255 - 0xff
    "11111111", -- 6526 - 0x197e  :  255 - 0xff
    "11111111", -- 6527 - 0x197f  :  255 - 0xff
    "11111110", -- 6528 - 0x1980  :  254 - 0xfe
    "11111100", -- 6529 - 0x1981  :  252 - 0xfc
    "11111100", -- 6530 - 0x1982  :  252 - 0xfc
    "11111000", -- 6531 - 0x1983  :  248 - 0xf8
    "00000000", -- 6532 - 0x1984  :    0 - 0x0
    "00000000", -- 6533 - 0x1985  :    0 - 0x0
    "00000000", -- 6534 - 0x1986  :    0 - 0x0
    "11111111", -- 6535 - 0x1987  :  255 - 0xff
    "11111111", -- 6536 - 0x1988  :  255 - 0xff
    "11111111", -- 6537 - 0x1989  :  255 - 0xff
    "11111111", -- 6538 - 0x198a  :  255 - 0xff
    "11111111", -- 6539 - 0x198b  :  255 - 0xff
    "11111111", -- 6540 - 0x198c  :  255 - 0xff
    "11111111", -- 6541 - 0x198d  :  255 - 0xff
    "11111111", -- 6542 - 0x198e  :  255 - 0xff
    "11111111", -- 6543 - 0x198f  :  255 - 0xff
    "00000000", -- 6544 - 0x1990  :    0 - 0x0
    "00000000", -- 6545 - 0x1991  :    0 - 0x0
    "00000000", -- 6546 - 0x1992  :    0 - 0x0
    "00000000", -- 6547 - 0x1993  :    0 - 0x0
    "11111111", -- 6548 - 0x1994  :  255 - 0xff
    "11111111", -- 6549 - 0x1995  :  255 - 0xff
    "00000000", -- 6550 - 0x1996  :    0 - 0x0
    "00000000", -- 6551 - 0x1997  :    0 - 0x0
    "00000000", -- 6552 - 0x1998  :    0 - 0x0
    "00000000", -- 6553 - 0x1999  :    0 - 0x0
    "00000000", -- 6554 - 0x199a  :    0 - 0x0
    "00000000", -- 6555 - 0x199b  :    0 - 0x0
    "00000000", -- 6556 - 0x199c  :    0 - 0x0
    "00000000", -- 6557 - 0x199d  :    0 - 0x0
    "00000000", -- 6558 - 0x199e  :    0 - 0x0
    "00000000", -- 6559 - 0x199f  :    0 - 0x0
    "00011000", -- 6560 - 0x19a0  :   24 - 0x18
    "00011000", -- 6561 - 0x19a1  :   24 - 0x18
    "00011000", -- 6562 - 0x19a2  :   24 - 0x18
    "00011000", -- 6563 - 0x19a3  :   24 - 0x18
    "00011000", -- 6564 - 0x19a4  :   24 - 0x18
    "00011000", -- 6565 - 0x19a5  :   24 - 0x18
    "00011000", -- 6566 - 0x19a6  :   24 - 0x18
    "00011000", -- 6567 - 0x19a7  :   24 - 0x18
    "00000000", -- 6568 - 0x19a8  :    0 - 0x0
    "00000000", -- 6569 - 0x19a9  :    0 - 0x0
    "00000000", -- 6570 - 0x19aa  :    0 - 0x0
    "00000000", -- 6571 - 0x19ab  :    0 - 0x0
    "00000000", -- 6572 - 0x19ac  :    0 - 0x0
    "00000000", -- 6573 - 0x19ad  :    0 - 0x0
    "00000000", -- 6574 - 0x19ae  :    0 - 0x0
    "00000000", -- 6575 - 0x19af  :    0 - 0x0
    "00000111", -- 6576 - 0x19b0  :    7 - 0x7
    "00011111", -- 6577 - 0x19b1  :   31 - 0x1f
    "00111111", -- 6578 - 0x19b2  :   63 - 0x3f
    "11111111", -- 6579 - 0x19b3  :  255 - 0xff
    "01111111", -- 6580 - 0x19b4  :  127 - 0x7f
    "01111111", -- 6581 - 0x19b5  :  127 - 0x7f
    "11111111", -- 6582 - 0x19b6  :  255 - 0xff
    "11111111", -- 6583 - 0x19b7  :  255 - 0xff
    "11111111", -- 6584 - 0x19b8  :  255 - 0xff
    "11111111", -- 6585 - 0x19b9  :  255 - 0xff
    "11111111", -- 6586 - 0x19ba  :  255 - 0xff
    "11111111", -- 6587 - 0x19bb  :  255 - 0xff
    "11111111", -- 6588 - 0x19bc  :  255 - 0xff
    "11111111", -- 6589 - 0x19bd  :  255 - 0xff
    "11111111", -- 6590 - 0x19be  :  255 - 0xff
    "11111111", -- 6591 - 0x19bf  :  255 - 0xff
    "11100001", -- 6592 - 0x19c0  :  225 - 0xe1
    "11111001", -- 6593 - 0x19c1  :  249 - 0xf9
    "11111101", -- 6594 - 0x19c2  :  253 - 0xfd
    "11111111", -- 6595 - 0x19c3  :  255 - 0xff
    "11111110", -- 6596 - 0x19c4  :  254 - 0xfe
    "11111110", -- 6597 - 0x19c5  :  254 - 0xfe
    "11111111", -- 6598 - 0x19c6  :  255 - 0xff
    "11111111", -- 6599 - 0x19c7  :  255 - 0xff
    "11111111", -- 6600 - 0x19c8  :  255 - 0xff
    "11111111", -- 6601 - 0x19c9  :  255 - 0xff
    "11111111", -- 6602 - 0x19ca  :  255 - 0xff
    "11111111", -- 6603 - 0x19cb  :  255 - 0xff
    "11111111", -- 6604 - 0x19cc  :  255 - 0xff
    "11111111", -- 6605 - 0x19cd  :  255 - 0xff
    "11111111", -- 6606 - 0x19ce  :  255 - 0xff
    "11111111", -- 6607 - 0x19cf  :  255 - 0xff
    "11110000", -- 6608 - 0x19d0  :  240 - 0xf0
    "00010000", -- 6609 - 0x19d1  :   16 - 0x10
    "00010000", -- 6610 - 0x19d2  :   16 - 0x10
    "00010000", -- 6611 - 0x19d3  :   16 - 0x10
    "00010000", -- 6612 - 0x19d4  :   16 - 0x10
    "00010000", -- 6613 - 0x19d5  :   16 - 0x10
    "00010000", -- 6614 - 0x19d6  :   16 - 0x10
    "11111111", -- 6615 - 0x19d7  :  255 - 0xff
    "00000000", -- 6616 - 0x19d8  :    0 - 0x0
    "11100000", -- 6617 - 0x19d9  :  224 - 0xe0
    "11100000", -- 6618 - 0x19da  :  224 - 0xe0
    "11100000", -- 6619 - 0x19db  :  224 - 0xe0
    "11100000", -- 6620 - 0x19dc  :  224 - 0xe0
    "11100000", -- 6621 - 0x19dd  :  224 - 0xe0
    "11100000", -- 6622 - 0x19de  :  224 - 0xe0
    "11100000", -- 6623 - 0x19df  :  224 - 0xe0
    "00011111", -- 6624 - 0x19e0  :   31 - 0x1f
    "00010000", -- 6625 - 0x19e1  :   16 - 0x10
    "00010000", -- 6626 - 0x19e2  :   16 - 0x10
    "00010000", -- 6627 - 0x19e3  :   16 - 0x10
    "00010000", -- 6628 - 0x19e4  :   16 - 0x10
    "00010000", -- 6629 - 0x19e5  :   16 - 0x10
    "00010000", -- 6630 - 0x19e6  :   16 - 0x10
    "11111111", -- 6631 - 0x19e7  :  255 - 0xff
    "00000000", -- 6632 - 0x19e8  :    0 - 0x0
    "00001111", -- 6633 - 0x19e9  :   15 - 0xf
    "00001111", -- 6634 - 0x19ea  :   15 - 0xf
    "00001111", -- 6635 - 0x19eb  :   15 - 0xf
    "00001111", -- 6636 - 0x19ec  :   15 - 0xf
    "00001111", -- 6637 - 0x19ed  :   15 - 0xf
    "00001111", -- 6638 - 0x19ee  :   15 - 0xf
    "00001111", -- 6639 - 0x19ef  :   15 - 0xf
    "10010010", -- 6640 - 0x19f0  :  146 - 0x92
    "10010010", -- 6641 - 0x19f1  :  146 - 0x92
    "10010010", -- 6642 - 0x19f2  :  146 - 0x92
    "11111110", -- 6643 - 0x19f3  :  254 - 0xfe
    "11111110", -- 6644 - 0x19f4  :  254 - 0xfe
    "00000000", -- 6645 - 0x19f5  :    0 - 0x0
    "00000000", -- 6646 - 0x19f6  :    0 - 0x0
    "00000000", -- 6647 - 0x19f7  :    0 - 0x0
    "01001000", -- 6648 - 0x19f8  :   72 - 0x48
    "01001000", -- 6649 - 0x19f9  :   72 - 0x48
    "01101100", -- 6650 - 0x19fa  :  108 - 0x6c
    "00000000", -- 6651 - 0x19fb  :    0 - 0x0
    "00000000", -- 6652 - 0x19fc  :    0 - 0x0
    "00000000", -- 6653 - 0x19fd  :    0 - 0x0
    "11111110", -- 6654 - 0x19fe  :  254 - 0xfe
    "00000000", -- 6655 - 0x19ff  :    0 - 0x0
    "00001010", -- 6656 - 0x1a00  :   10 - 0xa
    "00001010", -- 6657 - 0x1a01  :   10 - 0xa
    "00111010", -- 6658 - 0x1a02  :   58 - 0x3a
    "00001010", -- 6659 - 0x1a03  :   10 - 0xa
    "11111011", -- 6660 - 0x1a04  :  251 - 0xfb
    "00001011", -- 6661 - 0x1a05  :   11 - 0xb
    "00001011", -- 6662 - 0x1a06  :   11 - 0xb
    "00001011", -- 6663 - 0x1a07  :   11 - 0xb
    "00000101", -- 6664 - 0x1a08  :    5 - 0x5
    "00000101", -- 6665 - 0x1a09  :    5 - 0x5
    "11000101", -- 6666 - 0x1a0a  :  197 - 0xc5
    "11110101", -- 6667 - 0x1a0b  :  245 - 0xf5
    "11110100", -- 6668 - 0x1a0c  :  244 - 0xf4
    "00000100", -- 6669 - 0x1a0d  :    4 - 0x4
    "00000100", -- 6670 - 0x1a0e  :    4 - 0x4
    "00000100", -- 6671 - 0x1a0f  :    4 - 0x4
    "10010000", -- 6672 - 0x1a10  :  144 - 0x90
    "10010000", -- 6673 - 0x1a11  :  144 - 0x90
    "10011111", -- 6674 - 0x1a12  :  159 - 0x9f
    "10010000", -- 6675 - 0x1a13  :  144 - 0x90
    "10011111", -- 6676 - 0x1a14  :  159 - 0x9f
    "10010000", -- 6677 - 0x1a15  :  144 - 0x90
    "10010000", -- 6678 - 0x1a16  :  144 - 0x90
    "10010000", -- 6679 - 0x1a17  :  144 - 0x90
    "01110000", -- 6680 - 0x1a18  :  112 - 0x70
    "01110000", -- 6681 - 0x1a19  :  112 - 0x70
    "01110000", -- 6682 - 0x1a1a  :  112 - 0x70
    "01111111", -- 6683 - 0x1a1b  :  127 - 0x7f
    "01111111", -- 6684 - 0x1a1c  :  127 - 0x7f
    "01110000", -- 6685 - 0x1a1d  :  112 - 0x70
    "01110000", -- 6686 - 0x1a1e  :  112 - 0x70
    "01110000", -- 6687 - 0x1a1f  :  112 - 0x70
    "00000001", -- 6688 - 0x1a20  :    1 - 0x1
    "00000001", -- 6689 - 0x1a21  :    1 - 0x1
    "00000001", -- 6690 - 0x1a22  :    1 - 0x1
    "00000001", -- 6691 - 0x1a23  :    1 - 0x1
    "00000001", -- 6692 - 0x1a24  :    1 - 0x1
    "00000001", -- 6693 - 0x1a25  :    1 - 0x1
    "00000001", -- 6694 - 0x1a26  :    1 - 0x1
    "00000001", -- 6695 - 0x1a27  :    1 - 0x1
    "00000000", -- 6696 - 0x1a28  :    0 - 0x0
    "00000000", -- 6697 - 0x1a29  :    0 - 0x0
    "00000000", -- 6698 - 0x1a2a  :    0 - 0x0
    "00000000", -- 6699 - 0x1a2b  :    0 - 0x0
    "00000000", -- 6700 - 0x1a2c  :    0 - 0x0
    "00000000", -- 6701 - 0x1a2d  :    0 - 0x0
    "00000000", -- 6702 - 0x1a2e  :    0 - 0x0
    "00000000", -- 6703 - 0x1a2f  :    0 - 0x0
    "10000000", -- 6704 - 0x1a30  :  128 - 0x80
    "10000000", -- 6705 - 0x1a31  :  128 - 0x80
    "10000000", -- 6706 - 0x1a32  :  128 - 0x80
    "10000000", -- 6707 - 0x1a33  :  128 - 0x80
    "10000000", -- 6708 - 0x1a34  :  128 - 0x80
    "10000000", -- 6709 - 0x1a35  :  128 - 0x80
    "10000000", -- 6710 - 0x1a36  :  128 - 0x80
    "10000000", -- 6711 - 0x1a37  :  128 - 0x80
    "00000000", -- 6712 - 0x1a38  :    0 - 0x0
    "00000000", -- 6713 - 0x1a39  :    0 - 0x0
    "00000000", -- 6714 - 0x1a3a  :    0 - 0x0
    "00000000", -- 6715 - 0x1a3b  :    0 - 0x0
    "00000000", -- 6716 - 0x1a3c  :    0 - 0x0
    "00000000", -- 6717 - 0x1a3d  :    0 - 0x0
    "00000000", -- 6718 - 0x1a3e  :    0 - 0x0
    "00000000", -- 6719 - 0x1a3f  :    0 - 0x0
    "00001000", -- 6720 - 0x1a40  :    8 - 0x8
    "10001000", -- 6721 - 0x1a41  :  136 - 0x88
    "10010001", -- 6722 - 0x1a42  :  145 - 0x91
    "11010001", -- 6723 - 0x1a43  :  209 - 0xd1
    "01010011", -- 6724 - 0x1a44  :   83 - 0x53
    "01010011", -- 6725 - 0x1a45  :   83 - 0x53
    "01110011", -- 6726 - 0x1a46  :  115 - 0x73
    "00111111", -- 6727 - 0x1a47  :   63 - 0x3f
    "11111111", -- 6728 - 0x1a48  :  255 - 0xff
    "11111111", -- 6729 - 0x1a49  :  255 - 0xff
    "11111111", -- 6730 - 0x1a4a  :  255 - 0xff
    "11111111", -- 6731 - 0x1a4b  :  255 - 0xff
    "11111111", -- 6732 - 0x1a4c  :  255 - 0xff
    "11111110", -- 6733 - 0x1a4d  :  254 - 0xfe
    "10111110", -- 6734 - 0x1a4e  :  190 - 0xbe
    "11001110", -- 6735 - 0x1a4f  :  206 - 0xce
    "00000000", -- 6736 - 0x1a50  :    0 - 0x0
    "00000000", -- 6737 - 0x1a51  :    0 - 0x0
    "00000111", -- 6738 - 0x1a52  :    7 - 0x7
    "00001111", -- 6739 - 0x1a53  :   15 - 0xf
    "00001100", -- 6740 - 0x1a54  :   12 - 0xc
    "00011011", -- 6741 - 0x1a55  :   27 - 0x1b
    "00011011", -- 6742 - 0x1a56  :   27 - 0x1b
    "00011011", -- 6743 - 0x1a57  :   27 - 0x1b
    "00000000", -- 6744 - 0x1a58  :    0 - 0x0
    "00000000", -- 6745 - 0x1a59  :    0 - 0x0
    "00000000", -- 6746 - 0x1a5a  :    0 - 0x0
    "00000000", -- 6747 - 0x1a5b  :    0 - 0x0
    "00000011", -- 6748 - 0x1a5c  :    3 - 0x3
    "00000100", -- 6749 - 0x1a5d  :    4 - 0x4
    "00000100", -- 6750 - 0x1a5e  :    4 - 0x4
    "00000100", -- 6751 - 0x1a5f  :    4 - 0x4
    "00000000", -- 6752 - 0x1a60  :    0 - 0x0
    "00000000", -- 6753 - 0x1a61  :    0 - 0x0
    "11100000", -- 6754 - 0x1a62  :  224 - 0xe0
    "11110000", -- 6755 - 0x1a63  :  240 - 0xf0
    "11110000", -- 6756 - 0x1a64  :  240 - 0xf0
    "11111000", -- 6757 - 0x1a65  :  248 - 0xf8
    "11111000", -- 6758 - 0x1a66  :  248 - 0xf8
    "11111000", -- 6759 - 0x1a67  :  248 - 0xf8
    "00000000", -- 6760 - 0x1a68  :    0 - 0x0
    "00000000", -- 6761 - 0x1a69  :    0 - 0x0
    "01100000", -- 6762 - 0x1a6a  :   96 - 0x60
    "00110000", -- 6763 - 0x1a6b  :   48 - 0x30
    "00110000", -- 6764 - 0x1a6c  :   48 - 0x30
    "10011000", -- 6765 - 0x1a6d  :  152 - 0x98
    "10011000", -- 6766 - 0x1a6e  :  152 - 0x98
    "10011000", -- 6767 - 0x1a6f  :  152 - 0x98
    "00011011", -- 6768 - 0x1a70  :   27 - 0x1b
    "00011011", -- 6769 - 0x1a71  :   27 - 0x1b
    "00011011", -- 6770 - 0x1a72  :   27 - 0x1b
    "00011011", -- 6771 - 0x1a73  :   27 - 0x1b
    "00011011", -- 6772 - 0x1a74  :   27 - 0x1b
    "00001111", -- 6773 - 0x1a75  :   15 - 0xf
    "00001111", -- 6774 - 0x1a76  :   15 - 0xf
    "00000111", -- 6775 - 0x1a77  :    7 - 0x7
    "00000100", -- 6776 - 0x1a78  :    4 - 0x4
    "00000100", -- 6777 - 0x1a79  :    4 - 0x4
    "00000100", -- 6778 - 0x1a7a  :    4 - 0x4
    "00000100", -- 6779 - 0x1a7b  :    4 - 0x4
    "00000100", -- 6780 - 0x1a7c  :    4 - 0x4
    "00000011", -- 6781 - 0x1a7d  :    3 - 0x3
    "00000000", -- 6782 - 0x1a7e  :    0 - 0x0
    "00000000", -- 6783 - 0x1a7f  :    0 - 0x0
    "11111000", -- 6784 - 0x1a80  :  248 - 0xf8
    "11111000", -- 6785 - 0x1a81  :  248 - 0xf8
    "11111000", -- 6786 - 0x1a82  :  248 - 0xf8
    "11111000", -- 6787 - 0x1a83  :  248 - 0xf8
    "11111000", -- 6788 - 0x1a84  :  248 - 0xf8
    "11110000", -- 6789 - 0x1a85  :  240 - 0xf0
    "11110000", -- 6790 - 0x1a86  :  240 - 0xf0
    "11100000", -- 6791 - 0x1a87  :  224 - 0xe0
    "10011000", -- 6792 - 0x1a88  :  152 - 0x98
    "10011000", -- 6793 - 0x1a89  :  152 - 0x98
    "10011000", -- 6794 - 0x1a8a  :  152 - 0x98
    "10011000", -- 6795 - 0x1a8b  :  152 - 0x98
    "10011000", -- 6796 - 0x1a8c  :  152 - 0x98
    "00110000", -- 6797 - 0x1a8d  :   48 - 0x30
    "00110000", -- 6798 - 0x1a8e  :   48 - 0x30
    "01100000", -- 6799 - 0x1a8f  :   96 - 0x60
    "11110001", -- 6800 - 0x1a90  :  241 - 0xf1
    "00010001", -- 6801 - 0x1a91  :   17 - 0x11
    "00010001", -- 6802 - 0x1a92  :   17 - 0x11
    "00011111", -- 6803 - 0x1a93  :   31 - 0x1f
    "00010000", -- 6804 - 0x1a94  :   16 - 0x10
    "00010000", -- 6805 - 0x1a95  :   16 - 0x10
    "00010000", -- 6806 - 0x1a96  :   16 - 0x10
    "11111111", -- 6807 - 0x1a97  :  255 - 0xff
    "00001111", -- 6808 - 0x1a98  :   15 - 0xf
    "11101111", -- 6809 - 0x1a99  :  239 - 0xef
    "11101111", -- 6810 - 0x1a9a  :  239 - 0xef
    "11101111", -- 6811 - 0x1a9b  :  239 - 0xef
    "11101111", -- 6812 - 0x1a9c  :  239 - 0xef
    "11101111", -- 6813 - 0x1a9d  :  239 - 0xef
    "11101111", -- 6814 - 0x1a9e  :  239 - 0xef
    "11100000", -- 6815 - 0x1a9f  :  224 - 0xe0
    "00011111", -- 6816 - 0x1aa0  :   31 - 0x1f
    "00010000", -- 6817 - 0x1aa1  :   16 - 0x10
    "00010000", -- 6818 - 0x1aa2  :   16 - 0x10
    "11110000", -- 6819 - 0x1aa3  :  240 - 0xf0
    "00010000", -- 6820 - 0x1aa4  :   16 - 0x10
    "00010000", -- 6821 - 0x1aa5  :   16 - 0x10
    "00010000", -- 6822 - 0x1aa6  :   16 - 0x10
    "11111111", -- 6823 - 0x1aa7  :  255 - 0xff
    "11100000", -- 6824 - 0x1aa8  :  224 - 0xe0
    "11101111", -- 6825 - 0x1aa9  :  239 - 0xef
    "11101111", -- 6826 - 0x1aaa  :  239 - 0xef
    "11101111", -- 6827 - 0x1aab  :  239 - 0xef
    "11101111", -- 6828 - 0x1aac  :  239 - 0xef
    "11101111", -- 6829 - 0x1aad  :  239 - 0xef
    "11101111", -- 6830 - 0x1aae  :  239 - 0xef
    "00001111", -- 6831 - 0x1aaf  :   15 - 0xf
    "01111111", -- 6832 - 0x1ab0  :  127 - 0x7f
    "10111111", -- 6833 - 0x1ab1  :  191 - 0xbf
    "11011111", -- 6834 - 0x1ab2  :  223 - 0xdf
    "11101111", -- 6835 - 0x1ab3  :  239 - 0xef
    "11110000", -- 6836 - 0x1ab4  :  240 - 0xf0
    "11110000", -- 6837 - 0x1ab5  :  240 - 0xf0
    "11110000", -- 6838 - 0x1ab6  :  240 - 0xf0
    "11110000", -- 6839 - 0x1ab7  :  240 - 0xf0
    "10000000", -- 6840 - 0x1ab8  :  128 - 0x80
    "01000000", -- 6841 - 0x1ab9  :   64 - 0x40
    "00100000", -- 6842 - 0x1aba  :   32 - 0x20
    "00010000", -- 6843 - 0x1abb  :   16 - 0x10
    "00001111", -- 6844 - 0x1abc  :   15 - 0xf
    "00001111", -- 6845 - 0x1abd  :   15 - 0xf
    "00001111", -- 6846 - 0x1abe  :   15 - 0xf
    "00001111", -- 6847 - 0x1abf  :   15 - 0xf
    "11110000", -- 6848 - 0x1ac0  :  240 - 0xf0
    "11110000", -- 6849 - 0x1ac1  :  240 - 0xf0
    "11110000", -- 6850 - 0x1ac2  :  240 - 0xf0
    "11110000", -- 6851 - 0x1ac3  :  240 - 0xf0
    "11111111", -- 6852 - 0x1ac4  :  255 - 0xff
    "11111111", -- 6853 - 0x1ac5  :  255 - 0xff
    "11111111", -- 6854 - 0x1ac6  :  255 - 0xff
    "11111111", -- 6855 - 0x1ac7  :  255 - 0xff
    "00001111", -- 6856 - 0x1ac8  :   15 - 0xf
    "00001111", -- 6857 - 0x1ac9  :   15 - 0xf
    "00001111", -- 6858 - 0x1aca  :   15 - 0xf
    "00001111", -- 6859 - 0x1acb  :   15 - 0xf
    "00011111", -- 6860 - 0x1acc  :   31 - 0x1f
    "00111111", -- 6861 - 0x1acd  :   63 - 0x3f
    "01111111", -- 6862 - 0x1ace  :  127 - 0x7f
    "11111111", -- 6863 - 0x1acf  :  255 - 0xff
    "11111111", -- 6864 - 0x1ad0  :  255 - 0xff
    "11111111", -- 6865 - 0x1ad1  :  255 - 0xff
    "11111111", -- 6866 - 0x1ad2  :  255 - 0xff
    "11111111", -- 6867 - 0x1ad3  :  255 - 0xff
    "00001111", -- 6868 - 0x1ad4  :   15 - 0xf
    "00001111", -- 6869 - 0x1ad5  :   15 - 0xf
    "00001111", -- 6870 - 0x1ad6  :   15 - 0xf
    "00001111", -- 6871 - 0x1ad7  :   15 - 0xf
    "00000001", -- 6872 - 0x1ad8  :    1 - 0x1
    "00000011", -- 6873 - 0x1ad9  :    3 - 0x3
    "00000111", -- 6874 - 0x1ada  :    7 - 0x7
    "00001111", -- 6875 - 0x1adb  :   15 - 0xf
    "11111111", -- 6876 - 0x1adc  :  255 - 0xff
    "11111111", -- 6877 - 0x1add  :  255 - 0xff
    "11111111", -- 6878 - 0x1ade  :  255 - 0xff
    "11111111", -- 6879 - 0x1adf  :  255 - 0xff
    "00001111", -- 6880 - 0x1ae0  :   15 - 0xf
    "00001111", -- 6881 - 0x1ae1  :   15 - 0xf
    "00001111", -- 6882 - 0x1ae2  :   15 - 0xf
    "00001111", -- 6883 - 0x1ae3  :   15 - 0xf
    "11110111", -- 6884 - 0x1ae4  :  247 - 0xf7
    "11111011", -- 6885 - 0x1ae5  :  251 - 0xfb
    "11111101", -- 6886 - 0x1ae6  :  253 - 0xfd
    "11111110", -- 6887 - 0x1ae7  :  254 - 0xfe
    "11111111", -- 6888 - 0x1ae8  :  255 - 0xff
    "11111111", -- 6889 - 0x1ae9  :  255 - 0xff
    "11111111", -- 6890 - 0x1aea  :  255 - 0xff
    "11111111", -- 6891 - 0x1aeb  :  255 - 0xff
    "11111111", -- 6892 - 0x1aec  :  255 - 0xff
    "11111111", -- 6893 - 0x1aed  :  255 - 0xff
    "11111111", -- 6894 - 0x1aee  :  255 - 0xff
    "11111111", -- 6895 - 0x1aef  :  255 - 0xff
    "00000000", -- 6896 - 0x1af0  :    0 - 0x0
    "00000000", -- 6897 - 0x1af1  :    0 - 0x0
    "00000000", -- 6898 - 0x1af2  :    0 - 0x0
    "00000000", -- 6899 - 0x1af3  :    0 - 0x0
    "00000000", -- 6900 - 0x1af4  :    0 - 0x0
    "00000000", -- 6901 - 0x1af5  :    0 - 0x0
    "00011000", -- 6902 - 0x1af6  :   24 - 0x18
    "00011000", -- 6903 - 0x1af7  :   24 - 0x18
    "00000000", -- 6904 - 0x1af8  :    0 - 0x0
    "00000000", -- 6905 - 0x1af9  :    0 - 0x0
    "00000000", -- 6906 - 0x1afa  :    0 - 0x0
    "00000000", -- 6907 - 0x1afb  :    0 - 0x0
    "00000000", -- 6908 - 0x1afc  :    0 - 0x0
    "00000000", -- 6909 - 0x1afd  :    0 - 0x0
    "00000000", -- 6910 - 0x1afe  :    0 - 0x0
    "00000000", -- 6911 - 0x1aff  :    0 - 0x0
    "00011111", -- 6912 - 0x1b00  :   31 - 0x1f
    "00111111", -- 6913 - 0x1b01  :   63 - 0x3f
    "01111111", -- 6914 - 0x1b02  :  127 - 0x7f
    "01111111", -- 6915 - 0x1b03  :  127 - 0x7f
    "01111111", -- 6916 - 0x1b04  :  127 - 0x7f
    "11111111", -- 6917 - 0x1b05  :  255 - 0xff
    "11111111", -- 6918 - 0x1b06  :  255 - 0xff
    "11111111", -- 6919 - 0x1b07  :  255 - 0xff
    "00011111", -- 6920 - 0x1b08  :   31 - 0x1f
    "00100000", -- 6921 - 0x1b09  :   32 - 0x20
    "01000000", -- 6922 - 0x1b0a  :   64 - 0x40
    "01000000", -- 6923 - 0x1b0b  :   64 - 0x40
    "01000000", -- 6924 - 0x1b0c  :   64 - 0x40
    "10000000", -- 6925 - 0x1b0d  :  128 - 0x80
    "10000010", -- 6926 - 0x1b0e  :  130 - 0x82
    "10000010", -- 6927 - 0x1b0f  :  130 - 0x82
    "11111111", -- 6928 - 0x1b10  :  255 - 0xff
    "11111111", -- 6929 - 0x1b11  :  255 - 0xff
    "11111111", -- 6930 - 0x1b12  :  255 - 0xff
    "01111111", -- 6931 - 0x1b13  :  127 - 0x7f
    "01111111", -- 6932 - 0x1b14  :  127 - 0x7f
    "01111111", -- 6933 - 0x1b15  :  127 - 0x7f
    "00111111", -- 6934 - 0x1b16  :   63 - 0x3f
    "00011110", -- 6935 - 0x1b17  :   30 - 0x1e
    "10000010", -- 6936 - 0x1b18  :  130 - 0x82
    "10000000", -- 6937 - 0x1b19  :  128 - 0x80
    "10100000", -- 6938 - 0x1b1a  :  160 - 0xa0
    "01000100", -- 6939 - 0x1b1b  :   68 - 0x44
    "01000011", -- 6940 - 0x1b1c  :   67 - 0x43
    "01000000", -- 6941 - 0x1b1d  :   64 - 0x40
    "00100001", -- 6942 - 0x1b1e  :   33 - 0x21
    "00011110", -- 6943 - 0x1b1f  :   30 - 0x1e
    "11111000", -- 6944 - 0x1b20  :  248 - 0xf8
    "11111100", -- 6945 - 0x1b21  :  252 - 0xfc
    "11111110", -- 6946 - 0x1b22  :  254 - 0xfe
    "11111110", -- 6947 - 0x1b23  :  254 - 0xfe
    "11111110", -- 6948 - 0x1b24  :  254 - 0xfe
    "11111111", -- 6949 - 0x1b25  :  255 - 0xff
    "11111111", -- 6950 - 0x1b26  :  255 - 0xff
    "11111111", -- 6951 - 0x1b27  :  255 - 0xff
    "11111000", -- 6952 - 0x1b28  :  248 - 0xf8
    "00000100", -- 6953 - 0x1b29  :    4 - 0x4
    "00000010", -- 6954 - 0x1b2a  :    2 - 0x2
    "00000010", -- 6955 - 0x1b2b  :    2 - 0x2
    "00000010", -- 6956 - 0x1b2c  :    2 - 0x2
    "00000001", -- 6957 - 0x1b2d  :    1 - 0x1
    "01000001", -- 6958 - 0x1b2e  :   65 - 0x41
    "01000001", -- 6959 - 0x1b2f  :   65 - 0x41
    "11111111", -- 6960 - 0x1b30  :  255 - 0xff
    "11111111", -- 6961 - 0x1b31  :  255 - 0xff
    "11111111", -- 6962 - 0x1b32  :  255 - 0xff
    "11111110", -- 6963 - 0x1b33  :  254 - 0xfe
    "11111110", -- 6964 - 0x1b34  :  254 - 0xfe
    "11111110", -- 6965 - 0x1b35  :  254 - 0xfe
    "11111100", -- 6966 - 0x1b36  :  252 - 0xfc
    "01111000", -- 6967 - 0x1b37  :  120 - 0x78
    "01000001", -- 6968 - 0x1b38  :   65 - 0x41
    "00000001", -- 6969 - 0x1b39  :    1 - 0x1
    "00000101", -- 6970 - 0x1b3a  :    5 - 0x5
    "00100010", -- 6971 - 0x1b3b  :   34 - 0x22
    "11000010", -- 6972 - 0x1b3c  :  194 - 0xc2
    "00000010", -- 6973 - 0x1b3d  :    2 - 0x2
    "10000100", -- 6974 - 0x1b3e  :  132 - 0x84
    "01111000", -- 6975 - 0x1b3f  :  120 - 0x78
    "01111111", -- 6976 - 0x1b40  :  127 - 0x7f
    "10000000", -- 6977 - 0x1b41  :  128 - 0x80
    "10000000", -- 6978 - 0x1b42  :  128 - 0x80
    "10000000", -- 6979 - 0x1b43  :  128 - 0x80
    "10000000", -- 6980 - 0x1b44  :  128 - 0x80
    "10000000", -- 6981 - 0x1b45  :  128 - 0x80
    "10000000", -- 6982 - 0x1b46  :  128 - 0x80
    "10000000", -- 6983 - 0x1b47  :  128 - 0x80
    "10000000", -- 6984 - 0x1b48  :  128 - 0x80
    "01111111", -- 6985 - 0x1b49  :  127 - 0x7f
    "01111111", -- 6986 - 0x1b4a  :  127 - 0x7f
    "01111111", -- 6987 - 0x1b4b  :  127 - 0x7f
    "01111111", -- 6988 - 0x1b4c  :  127 - 0x7f
    "01111111", -- 6989 - 0x1b4d  :  127 - 0x7f
    "01111111", -- 6990 - 0x1b4e  :  127 - 0x7f
    "01111111", -- 6991 - 0x1b4f  :  127 - 0x7f
    "11011110", -- 6992 - 0x1b50  :  222 - 0xde
    "01100001", -- 6993 - 0x1b51  :   97 - 0x61
    "01100001", -- 6994 - 0x1b52  :   97 - 0x61
    "01100001", -- 6995 - 0x1b53  :   97 - 0x61
    "01110001", -- 6996 - 0x1b54  :  113 - 0x71
    "01011110", -- 6997 - 0x1b55  :   94 - 0x5e
    "01111111", -- 6998 - 0x1b56  :  127 - 0x7f
    "01100001", -- 6999 - 0x1b57  :   97 - 0x61
    "01100001", -- 7000 - 0x1b58  :   97 - 0x61
    "11011111", -- 7001 - 0x1b59  :  223 - 0xdf
    "11011111", -- 7002 - 0x1b5a  :  223 - 0xdf
    "11011111", -- 7003 - 0x1b5b  :  223 - 0xdf
    "11011111", -- 7004 - 0x1b5c  :  223 - 0xdf
    "11111111", -- 7005 - 0x1b5d  :  255 - 0xff
    "11000001", -- 7006 - 0x1b5e  :  193 - 0xc1
    "11011111", -- 7007 - 0x1b5f  :  223 - 0xdf
    "10000000", -- 7008 - 0x1b60  :  128 - 0x80
    "10000000", -- 7009 - 0x1b61  :  128 - 0x80
    "11000000", -- 7010 - 0x1b62  :  192 - 0xc0
    "11110000", -- 7011 - 0x1b63  :  240 - 0xf0
    "10111111", -- 7012 - 0x1b64  :  191 - 0xbf
    "10001111", -- 7013 - 0x1b65  :  143 - 0x8f
    "10000001", -- 7014 - 0x1b66  :  129 - 0x81
    "01111110", -- 7015 - 0x1b67  :  126 - 0x7e
    "01111111", -- 7016 - 0x1b68  :  127 - 0x7f
    "01111111", -- 7017 - 0x1b69  :  127 - 0x7f
    "11111111", -- 7018 - 0x1b6a  :  255 - 0xff
    "00111111", -- 7019 - 0x1b6b  :   63 - 0x3f
    "01001111", -- 7020 - 0x1b6c  :   79 - 0x4f
    "01110001", -- 7021 - 0x1b6d  :  113 - 0x71
    "01111111", -- 7022 - 0x1b6e  :  127 - 0x7f
    "11111111", -- 7023 - 0x1b6f  :  255 - 0xff
    "01100001", -- 7024 - 0x1b70  :   97 - 0x61
    "01100001", -- 7025 - 0x1b71  :   97 - 0x61
    "11000001", -- 7026 - 0x1b72  :  193 - 0xc1
    "11000001", -- 7027 - 0x1b73  :  193 - 0xc1
    "10000001", -- 7028 - 0x1b74  :  129 - 0x81
    "10000001", -- 7029 - 0x1b75  :  129 - 0x81
    "10000011", -- 7030 - 0x1b76  :  131 - 0x83
    "11111110", -- 7031 - 0x1b77  :  254 - 0xfe
    "11011111", -- 7032 - 0x1b78  :  223 - 0xdf
    "11011111", -- 7033 - 0x1b79  :  223 - 0xdf
    "10111111", -- 7034 - 0x1b7a  :  191 - 0xbf
    "10111111", -- 7035 - 0x1b7b  :  191 - 0xbf
    "01111111", -- 7036 - 0x1b7c  :  127 - 0x7f
    "01111111", -- 7037 - 0x1b7d  :  127 - 0x7f
    "01111111", -- 7038 - 0x1b7e  :  127 - 0x7f
    "01111111", -- 7039 - 0x1b7f  :  127 - 0x7f
    "00000000", -- 7040 - 0x1b80  :    0 - 0x0
    "00000000", -- 7041 - 0x1b81  :    0 - 0x0
    "00000011", -- 7042 - 0x1b82  :    3 - 0x3
    "00001111", -- 7043 - 0x1b83  :   15 - 0xf
    "00011111", -- 7044 - 0x1b84  :   31 - 0x1f
    "00111111", -- 7045 - 0x1b85  :   63 - 0x3f
    "01111111", -- 7046 - 0x1b86  :  127 - 0x7f
    "01111111", -- 7047 - 0x1b87  :  127 - 0x7f
    "00000000", -- 7048 - 0x1b88  :    0 - 0x0
    "00000000", -- 7049 - 0x1b89  :    0 - 0x0
    "00000011", -- 7050 - 0x1b8a  :    3 - 0x3
    "00001100", -- 7051 - 0x1b8b  :   12 - 0xc
    "00010000", -- 7052 - 0x1b8c  :   16 - 0x10
    "00100000", -- 7053 - 0x1b8d  :   32 - 0x20
    "01000000", -- 7054 - 0x1b8e  :   64 - 0x40
    "01000000", -- 7055 - 0x1b8f  :   64 - 0x40
    "00000000", -- 7056 - 0x1b90  :    0 - 0x0
    "00000000", -- 7057 - 0x1b91  :    0 - 0x0
    "11000000", -- 7058 - 0x1b92  :  192 - 0xc0
    "11110000", -- 7059 - 0x1b93  :  240 - 0xf0
    "11111000", -- 7060 - 0x1b94  :  248 - 0xf8
    "11111100", -- 7061 - 0x1b95  :  252 - 0xfc
    "11111110", -- 7062 - 0x1b96  :  254 - 0xfe
    "11111110", -- 7063 - 0x1b97  :  254 - 0xfe
    "00000000", -- 7064 - 0x1b98  :    0 - 0x0
    "00000000", -- 7065 - 0x1b99  :    0 - 0x0
    "11000000", -- 7066 - 0x1b9a  :  192 - 0xc0
    "00110000", -- 7067 - 0x1b9b  :   48 - 0x30
    "00001000", -- 7068 - 0x1b9c  :    8 - 0x8
    "00000100", -- 7069 - 0x1b9d  :    4 - 0x4
    "00000010", -- 7070 - 0x1b9e  :    2 - 0x2
    "00000010", -- 7071 - 0x1b9f  :    2 - 0x2
    "11111111", -- 7072 - 0x1ba0  :  255 - 0xff
    "11111111", -- 7073 - 0x1ba1  :  255 - 0xff
    "11111111", -- 7074 - 0x1ba2  :  255 - 0xff
    "11111111", -- 7075 - 0x1ba3  :  255 - 0xff
    "11111111", -- 7076 - 0x1ba4  :  255 - 0xff
    "11111111", -- 7077 - 0x1ba5  :  255 - 0xff
    "11111111", -- 7078 - 0x1ba6  :  255 - 0xff
    "11111111", -- 7079 - 0x1ba7  :  255 - 0xff
    "10000000", -- 7080 - 0x1ba8  :  128 - 0x80
    "10000000", -- 7081 - 0x1ba9  :  128 - 0x80
    "10000000", -- 7082 - 0x1baa  :  128 - 0x80
    "10000000", -- 7083 - 0x1bab  :  128 - 0x80
    "10000000", -- 7084 - 0x1bac  :  128 - 0x80
    "10000000", -- 7085 - 0x1bad  :  128 - 0x80
    "10000000", -- 7086 - 0x1bae  :  128 - 0x80
    "10000000", -- 7087 - 0x1baf  :  128 - 0x80
    "11111111", -- 7088 - 0x1bb0  :  255 - 0xff
    "11111111", -- 7089 - 0x1bb1  :  255 - 0xff
    "11111111", -- 7090 - 0x1bb2  :  255 - 0xff
    "11111111", -- 7091 - 0x1bb3  :  255 - 0xff
    "11111111", -- 7092 - 0x1bb4  :  255 - 0xff
    "11111111", -- 7093 - 0x1bb5  :  255 - 0xff
    "11111111", -- 7094 - 0x1bb6  :  255 - 0xff
    "11111111", -- 7095 - 0x1bb7  :  255 - 0xff
    "00000001", -- 7096 - 0x1bb8  :    1 - 0x1
    "00000001", -- 7097 - 0x1bb9  :    1 - 0x1
    "00000001", -- 7098 - 0x1bba  :    1 - 0x1
    "00000001", -- 7099 - 0x1bbb  :    1 - 0x1
    "00000001", -- 7100 - 0x1bbc  :    1 - 0x1
    "00000001", -- 7101 - 0x1bbd  :    1 - 0x1
    "00000001", -- 7102 - 0x1bbe  :    1 - 0x1
    "00000001", -- 7103 - 0x1bbf  :    1 - 0x1
    "01111111", -- 7104 - 0x1bc0  :  127 - 0x7f
    "01111111", -- 7105 - 0x1bc1  :  127 - 0x7f
    "01111111", -- 7106 - 0x1bc2  :  127 - 0x7f
    "00111111", -- 7107 - 0x1bc3  :   63 - 0x3f
    "00111111", -- 7108 - 0x1bc4  :   63 - 0x3f
    "00011111", -- 7109 - 0x1bc5  :   31 - 0x1f
    "00001111", -- 7110 - 0x1bc6  :   15 - 0xf
    "00000111", -- 7111 - 0x1bc7  :    7 - 0x7
    "01000000", -- 7112 - 0x1bc8  :   64 - 0x40
    "01000000", -- 7113 - 0x1bc9  :   64 - 0x40
    "01000000", -- 7114 - 0x1bca  :   64 - 0x40
    "00100000", -- 7115 - 0x1bcb  :   32 - 0x20
    "00110000", -- 7116 - 0x1bcc  :   48 - 0x30
    "00011100", -- 7117 - 0x1bcd  :   28 - 0x1c
    "00001111", -- 7118 - 0x1bce  :   15 - 0xf
    "00000111", -- 7119 - 0x1bcf  :    7 - 0x7
    "11111110", -- 7120 - 0x1bd0  :  254 - 0xfe
    "11111110", -- 7121 - 0x1bd1  :  254 - 0xfe
    "11111110", -- 7122 - 0x1bd2  :  254 - 0xfe
    "11111100", -- 7123 - 0x1bd3  :  252 - 0xfc
    "11111100", -- 7124 - 0x1bd4  :  252 - 0xfc
    "11111000", -- 7125 - 0x1bd5  :  248 - 0xf8
    "11110000", -- 7126 - 0x1bd6  :  240 - 0xf0
    "11110000", -- 7127 - 0x1bd7  :  240 - 0xf0
    "00000010", -- 7128 - 0x1bd8  :    2 - 0x2
    "00000010", -- 7129 - 0x1bd9  :    2 - 0x2
    "00000010", -- 7130 - 0x1bda  :    2 - 0x2
    "00000100", -- 7131 - 0x1bdb  :    4 - 0x4
    "00001100", -- 7132 - 0x1bdc  :   12 - 0xc
    "00111000", -- 7133 - 0x1bdd  :   56 - 0x38
    "11110000", -- 7134 - 0x1bde  :  240 - 0xf0
    "11110000", -- 7135 - 0x1bdf  :  240 - 0xf0
    "00001111", -- 7136 - 0x1be0  :   15 - 0xf
    "00001111", -- 7137 - 0x1be1  :   15 - 0xf
    "00001111", -- 7138 - 0x1be2  :   15 - 0xf
    "00001111", -- 7139 - 0x1be3  :   15 - 0xf
    "00001111", -- 7140 - 0x1be4  :   15 - 0xf
    "00001111", -- 7141 - 0x1be5  :   15 - 0xf
    "00000111", -- 7142 - 0x1be6  :    7 - 0x7
    "00001111", -- 7143 - 0x1be7  :   15 - 0xf
    "00001000", -- 7144 - 0x1be8  :    8 - 0x8
    "00001000", -- 7145 - 0x1be9  :    8 - 0x8
    "00001000", -- 7146 - 0x1bea  :    8 - 0x8
    "00001000", -- 7147 - 0x1beb  :    8 - 0x8
    "00001000", -- 7148 - 0x1bec  :    8 - 0x8
    "00001100", -- 7149 - 0x1bed  :   12 - 0xc
    "00000101", -- 7150 - 0x1bee  :    5 - 0x5
    "00001010", -- 7151 - 0x1bef  :   10 - 0xa
    "11110000", -- 7152 - 0x1bf0  :  240 - 0xf0
    "11110000", -- 7153 - 0x1bf1  :  240 - 0xf0
    "11110000", -- 7154 - 0x1bf2  :  240 - 0xf0
    "11110000", -- 7155 - 0x1bf3  :  240 - 0xf0
    "11110000", -- 7156 - 0x1bf4  :  240 - 0xf0
    "11110000", -- 7157 - 0x1bf5  :  240 - 0xf0
    "11100000", -- 7158 - 0x1bf6  :  224 - 0xe0
    "11110000", -- 7159 - 0x1bf7  :  240 - 0xf0
    "00010000", -- 7160 - 0x1bf8  :   16 - 0x10
    "01010000", -- 7161 - 0x1bf9  :   80 - 0x50
    "01010000", -- 7162 - 0x1bfa  :   80 - 0x50
    "01010000", -- 7163 - 0x1bfb  :   80 - 0x50
    "01010000", -- 7164 - 0x1bfc  :   80 - 0x50
    "00110000", -- 7165 - 0x1bfd  :   48 - 0x30
    "10100000", -- 7166 - 0x1bfe  :  160 - 0xa0
    "01010000", -- 7167 - 0x1bff  :   80 - 0x50
    "10000001", -- 7168 - 0x1c00  :  129 - 0x81
    "11000001", -- 7169 - 0x1c01  :  193 - 0xc1
    "10100011", -- 7170 - 0x1c02  :  163 - 0xa3
    "10100011", -- 7171 - 0x1c03  :  163 - 0xa3
    "10011101", -- 7172 - 0x1c04  :  157 - 0x9d
    "10000001", -- 7173 - 0x1c05  :  129 - 0x81
    "10000001", -- 7174 - 0x1c06  :  129 - 0x81
    "10000001", -- 7175 - 0x1c07  :  129 - 0x81
    "00000000", -- 7176 - 0x1c08  :    0 - 0x0
    "01000001", -- 7177 - 0x1c09  :   65 - 0x41
    "00100010", -- 7178 - 0x1c0a  :   34 - 0x22
    "00100010", -- 7179 - 0x1c0b  :   34 - 0x22
    "00011100", -- 7180 - 0x1c0c  :   28 - 0x1c
    "00000000", -- 7181 - 0x1c0d  :    0 - 0x0
    "00000000", -- 7182 - 0x1c0e  :    0 - 0x0
    "00000000", -- 7183 - 0x1c0f  :    0 - 0x0
    "11100011", -- 7184 - 0x1c10  :  227 - 0xe3
    "11110111", -- 7185 - 0x1c11  :  247 - 0xf7
    "11000001", -- 7186 - 0x1c12  :  193 - 0xc1
    "11000001", -- 7187 - 0x1c13  :  193 - 0xc1
    "11000001", -- 7188 - 0x1c14  :  193 - 0xc1
    "11000001", -- 7189 - 0x1c15  :  193 - 0xc1
    "11110111", -- 7190 - 0x1c16  :  247 - 0xf7
    "11100011", -- 7191 - 0x1c17  :  227 - 0xe3
    "11100011", -- 7192 - 0x1c18  :  227 - 0xe3
    "00010100", -- 7193 - 0x1c19  :   20 - 0x14
    "00111110", -- 7194 - 0x1c1a  :   62 - 0x3e
    "00111110", -- 7195 - 0x1c1b  :   62 - 0x3e
    "00111110", -- 7196 - 0x1c1c  :   62 - 0x3e
    "00111110", -- 7197 - 0x1c1d  :   62 - 0x3e
    "00010100", -- 7198 - 0x1c1e  :   20 - 0x14
    "11100011", -- 7199 - 0x1c1f  :  227 - 0xe3
    "00000000", -- 7200 - 0x1c20  :    0 - 0x0
    "00000000", -- 7201 - 0x1c21  :    0 - 0x0
    "00000111", -- 7202 - 0x1c22  :    7 - 0x7
    "00001111", -- 7203 - 0x1c23  :   15 - 0xf
    "00001100", -- 7204 - 0x1c24  :   12 - 0xc
    "00011011", -- 7205 - 0x1c25  :   27 - 0x1b
    "00011011", -- 7206 - 0x1c26  :   27 - 0x1b
    "00011011", -- 7207 - 0x1c27  :   27 - 0x1b
    "11111111", -- 7208 - 0x1c28  :  255 - 0xff
    "11111111", -- 7209 - 0x1c29  :  255 - 0xff
    "11111000", -- 7210 - 0x1c2a  :  248 - 0xf8
    "11110000", -- 7211 - 0x1c2b  :  240 - 0xf0
    "11110000", -- 7212 - 0x1c2c  :  240 - 0xf0
    "11100000", -- 7213 - 0x1c2d  :  224 - 0xe0
    "11100000", -- 7214 - 0x1c2e  :  224 - 0xe0
    "11100000", -- 7215 - 0x1c2f  :  224 - 0xe0
    "00000000", -- 7216 - 0x1c30  :    0 - 0x0
    "00000000", -- 7217 - 0x1c31  :    0 - 0x0
    "11100000", -- 7218 - 0x1c32  :  224 - 0xe0
    "11110000", -- 7219 - 0x1c33  :  240 - 0xf0
    "11110000", -- 7220 - 0x1c34  :  240 - 0xf0
    "11111000", -- 7221 - 0x1c35  :  248 - 0xf8
    "11111000", -- 7222 - 0x1c36  :  248 - 0xf8
    "11111000", -- 7223 - 0x1c37  :  248 - 0xf8
    "11111111", -- 7224 - 0x1c38  :  255 - 0xff
    "11111111", -- 7225 - 0x1c39  :  255 - 0xff
    "01111111", -- 7226 - 0x1c3a  :  127 - 0x7f
    "00111111", -- 7227 - 0x1c3b  :   63 - 0x3f
    "00111111", -- 7228 - 0x1c3c  :   63 - 0x3f
    "10011111", -- 7229 - 0x1c3d  :  159 - 0x9f
    "10011111", -- 7230 - 0x1c3e  :  159 - 0x9f
    "10011111", -- 7231 - 0x1c3f  :  159 - 0x9f
    "00011011", -- 7232 - 0x1c40  :   27 - 0x1b
    "00011011", -- 7233 - 0x1c41  :   27 - 0x1b
    "00011011", -- 7234 - 0x1c42  :   27 - 0x1b
    "00011011", -- 7235 - 0x1c43  :   27 - 0x1b
    "00011011", -- 7236 - 0x1c44  :   27 - 0x1b
    "00001111", -- 7237 - 0x1c45  :   15 - 0xf
    "00001111", -- 7238 - 0x1c46  :   15 - 0xf
    "00000111", -- 7239 - 0x1c47  :    7 - 0x7
    "11100000", -- 7240 - 0x1c48  :  224 - 0xe0
    "11100000", -- 7241 - 0x1c49  :  224 - 0xe0
    "11100000", -- 7242 - 0x1c4a  :  224 - 0xe0
    "11100000", -- 7243 - 0x1c4b  :  224 - 0xe0
    "11100000", -- 7244 - 0x1c4c  :  224 - 0xe0
    "11110011", -- 7245 - 0x1c4d  :  243 - 0xf3
    "11110000", -- 7246 - 0x1c4e  :  240 - 0xf0
    "11111000", -- 7247 - 0x1c4f  :  248 - 0xf8
    "11111000", -- 7248 - 0x1c50  :  248 - 0xf8
    "11111000", -- 7249 - 0x1c51  :  248 - 0xf8
    "11111000", -- 7250 - 0x1c52  :  248 - 0xf8
    "11111000", -- 7251 - 0x1c53  :  248 - 0xf8
    "11111000", -- 7252 - 0x1c54  :  248 - 0xf8
    "11110000", -- 7253 - 0x1c55  :  240 - 0xf0
    "11110000", -- 7254 - 0x1c56  :  240 - 0xf0
    "11100000", -- 7255 - 0x1c57  :  224 - 0xe0
    "10011111", -- 7256 - 0x1c58  :  159 - 0x9f
    "10011111", -- 7257 - 0x1c59  :  159 - 0x9f
    "10011111", -- 7258 - 0x1c5a  :  159 - 0x9f
    "10011111", -- 7259 - 0x1c5b  :  159 - 0x9f
    "10011111", -- 7260 - 0x1c5c  :  159 - 0x9f
    "00111111", -- 7261 - 0x1c5d  :   63 - 0x3f
    "00111111", -- 7262 - 0x1c5e  :   63 - 0x3f
    "01111111", -- 7263 - 0x1c5f  :  127 - 0x7f
    "11100000", -- 7264 - 0x1c60  :  224 - 0xe0
    "11111111", -- 7265 - 0x1c61  :  255 - 0xff
    "11111111", -- 7266 - 0x1c62  :  255 - 0xff
    "11111111", -- 7267 - 0x1c63  :  255 - 0xff
    "11111111", -- 7268 - 0x1c64  :  255 - 0xff
    "11111111", -- 7269 - 0x1c65  :  255 - 0xff
    "11111111", -- 7270 - 0x1c66  :  255 - 0xff
    "11111111", -- 7271 - 0x1c67  :  255 - 0xff
    "00000000", -- 7272 - 0x1c68  :    0 - 0x0
    "01110000", -- 7273 - 0x1c69  :  112 - 0x70
    "00011111", -- 7274 - 0x1c6a  :   31 - 0x1f
    "00010000", -- 7275 - 0x1c6b  :   16 - 0x10
    "01110000", -- 7276 - 0x1c6c  :  112 - 0x70
    "01111111", -- 7277 - 0x1c6d  :  127 - 0x7f
    "01111111", -- 7278 - 0x1c6e  :  127 - 0x7f
    "01111111", -- 7279 - 0x1c6f  :  127 - 0x7f
    "00000111", -- 7280 - 0x1c70  :    7 - 0x7
    "11111111", -- 7281 - 0x1c71  :  255 - 0xff
    "11111111", -- 7282 - 0x1c72  :  255 - 0xff
    "11111111", -- 7283 - 0x1c73  :  255 - 0xff
    "11111111", -- 7284 - 0x1c74  :  255 - 0xff
    "11111111", -- 7285 - 0x1c75  :  255 - 0xff
    "11111111", -- 7286 - 0x1c76  :  255 - 0xff
    "11111111", -- 7287 - 0x1c77  :  255 - 0xff
    "00000000", -- 7288 - 0x1c78  :    0 - 0x0
    "00000011", -- 7289 - 0x1c79  :    3 - 0x3
    "11111000", -- 7290 - 0x1c7a  :  248 - 0xf8
    "00000000", -- 7291 - 0x1c7b  :    0 - 0x0
    "00000011", -- 7292 - 0x1c7c  :    3 - 0x3
    "11111011", -- 7293 - 0x1c7d  :  251 - 0xfb
    "11111011", -- 7294 - 0x1c7e  :  251 - 0xfb
    "11111011", -- 7295 - 0x1c7f  :  251 - 0xfb
    "11111111", -- 7296 - 0x1c80  :  255 - 0xff
    "11111111", -- 7297 - 0x1c81  :  255 - 0xff
    "11111111", -- 7298 - 0x1c82  :  255 - 0xff
    "11111111", -- 7299 - 0x1c83  :  255 - 0xff
    "11111111", -- 7300 - 0x1c84  :  255 - 0xff
    "11111110", -- 7301 - 0x1c85  :  254 - 0xfe
    "11111111", -- 7302 - 0x1c86  :  255 - 0xff
    "11101111", -- 7303 - 0x1c87  :  239 - 0xef
    "01111100", -- 7304 - 0x1c88  :  124 - 0x7c
    "01111011", -- 7305 - 0x1c89  :  123 - 0x7b
    "01110110", -- 7306 - 0x1c8a  :  118 - 0x76
    "01110101", -- 7307 - 0x1c8b  :  117 - 0x75
    "01110101", -- 7308 - 0x1c8c  :  117 - 0x75
    "01110111", -- 7309 - 0x1c8d  :  119 - 0x77
    "00010111", -- 7310 - 0x1c8e  :   23 - 0x17
    "01100111", -- 7311 - 0x1c8f  :  103 - 0x67
    "11111111", -- 7312 - 0x1c90  :  255 - 0xff
    "11011111", -- 7313 - 0x1c91  :  223 - 0xdf
    "11101111", -- 7314 - 0x1c92  :  239 - 0xef
    "10101111", -- 7315 - 0x1c93  :  175 - 0xaf
    "10101111", -- 7316 - 0x1c94  :  175 - 0xaf
    "01101111", -- 7317 - 0x1c95  :  111 - 0x6f
    "11101111", -- 7318 - 0x1c96  :  239 - 0xef
    "11100111", -- 7319 - 0x1c97  :  231 - 0xe7
    "00111011", -- 7320 - 0x1c98  :   59 - 0x3b
    "11111011", -- 7321 - 0x1c99  :  251 - 0xfb
    "01111011", -- 7322 - 0x1c9a  :  123 - 0x7b
    "11111011", -- 7323 - 0x1c9b  :  251 - 0xfb
    "11111011", -- 7324 - 0x1c9c  :  251 - 0xfb
    "11110011", -- 7325 - 0x1c9d  :  243 - 0xf3
    "11111000", -- 7326 - 0x1c9e  :  248 - 0xf8
    "11110011", -- 7327 - 0x1c9f  :  243 - 0xf3
    "00011111", -- 7328 - 0x1ca0  :   31 - 0x1f
    "00011111", -- 7329 - 0x1ca1  :   31 - 0x1f
    "00111111", -- 7330 - 0x1ca2  :   63 - 0x3f
    "00111111", -- 7331 - 0x1ca3  :   63 - 0x3f
    "01110000", -- 7332 - 0x1ca4  :  112 - 0x70
    "01100011", -- 7333 - 0x1ca5  :   99 - 0x63
    "11100111", -- 7334 - 0x1ca6  :  231 - 0xe7
    "11100101", -- 7335 - 0x1ca7  :  229 - 0xe5
    "00001111", -- 7336 - 0x1ca8  :   15 - 0xf
    "00001111", -- 7337 - 0x1ca9  :   15 - 0xf
    "00011111", -- 7338 - 0x1caa  :   31 - 0x1f
    "00011111", -- 7339 - 0x1cab  :   31 - 0x1f
    "00111111", -- 7340 - 0x1cac  :   63 - 0x3f
    "00111100", -- 7341 - 0x1cad  :   60 - 0x3c
    "01111000", -- 7342 - 0x1cae  :  120 - 0x78
    "01111010", -- 7343 - 0x1caf  :  122 - 0x7a
    "11110000", -- 7344 - 0x1cb0  :  240 - 0xf0
    "11110000", -- 7345 - 0x1cb1  :  240 - 0xf0
    "11111000", -- 7346 - 0x1cb2  :  248 - 0xf8
    "11111000", -- 7347 - 0x1cb3  :  248 - 0xf8
    "00001100", -- 7348 - 0x1cb4  :   12 - 0xc
    "11000100", -- 7349 - 0x1cb5  :  196 - 0xc4
    "11100100", -- 7350 - 0x1cb6  :  228 - 0xe4
    "10100110", -- 7351 - 0x1cb7  :  166 - 0xa6
    "11111000", -- 7352 - 0x1cb8  :  248 - 0xf8
    "11111000", -- 7353 - 0x1cb9  :  248 - 0xf8
    "11111100", -- 7354 - 0x1cba  :  252 - 0xfc
    "11111100", -- 7355 - 0x1cbb  :  252 - 0xfc
    "11111110", -- 7356 - 0x1cbc  :  254 - 0xfe
    "00111110", -- 7357 - 0x1cbd  :   62 - 0x3e
    "00011110", -- 7358 - 0x1cbe  :   30 - 0x1e
    "01011111", -- 7359 - 0x1cbf  :   95 - 0x5f
    "11101001", -- 7360 - 0x1cc0  :  233 - 0xe9
    "11101001", -- 7361 - 0x1cc1  :  233 - 0xe9
    "11101001", -- 7362 - 0x1cc2  :  233 - 0xe9
    "11101111", -- 7363 - 0x1cc3  :  239 - 0xef
    "11100010", -- 7364 - 0x1cc4  :  226 - 0xe2
    "11100011", -- 7365 - 0x1cc5  :  227 - 0xe3
    "11110000", -- 7366 - 0x1cc6  :  240 - 0xf0
    "11111111", -- 7367 - 0x1cc7  :  255 - 0xff
    "01110110", -- 7368 - 0x1cc8  :  118 - 0x76
    "01110110", -- 7369 - 0x1cc9  :  118 - 0x76
    "01110110", -- 7370 - 0x1cca  :  118 - 0x76
    "01110000", -- 7371 - 0x1ccb  :  112 - 0x70
    "01111101", -- 7372 - 0x1ccc  :  125 - 0x7d
    "01111100", -- 7373 - 0x1ccd  :  124 - 0x7c
    "01111111", -- 7374 - 0x1cce  :  127 - 0x7f
    "01111111", -- 7375 - 0x1ccf  :  127 - 0x7f
    "10010110", -- 7376 - 0x1cd0  :  150 - 0x96
    "10010110", -- 7377 - 0x1cd1  :  150 - 0x96
    "10010110", -- 7378 - 0x1cd2  :  150 - 0x96
    "11110110", -- 7379 - 0x1cd3  :  246 - 0xf6
    "01000110", -- 7380 - 0x1cd4  :   70 - 0x46
    "11000110", -- 7381 - 0x1cd5  :  198 - 0xc6
    "00001110", -- 7382 - 0x1cd6  :   14 - 0xe
    "11111110", -- 7383 - 0x1cd7  :  254 - 0xfe
    "01101111", -- 7384 - 0x1cd8  :  111 - 0x6f
    "01101111", -- 7385 - 0x1cd9  :  111 - 0x6f
    "01101111", -- 7386 - 0x1cda  :  111 - 0x6f
    "00001111", -- 7387 - 0x1cdb  :   15 - 0xf
    "10111111", -- 7388 - 0x1cdc  :  191 - 0xbf
    "00111111", -- 7389 - 0x1cdd  :   63 - 0x3f
    "11111111", -- 7390 - 0x1cde  :  255 - 0xff
    "11111111", -- 7391 - 0x1cdf  :  255 - 0xff
    "00000000", -- 7392 - 0x1ce0  :    0 - 0x0
    "00000000", -- 7393 - 0x1ce1  :    0 - 0x0
    "00000000", -- 7394 - 0x1ce2  :    0 - 0x0
    "00000000", -- 7395 - 0x1ce3  :    0 - 0x0
    "00000000", -- 7396 - 0x1ce4  :    0 - 0x0
    "00000000", -- 7397 - 0x1ce5  :    0 - 0x0
    "01111110", -- 7398 - 0x1ce6  :  126 - 0x7e
    "00111100", -- 7399 - 0x1ce7  :   60 - 0x3c
    "00111100", -- 7400 - 0x1ce8  :   60 - 0x3c
    "01111110", -- 7401 - 0x1ce9  :  126 - 0x7e
    "01111110", -- 7402 - 0x1cea  :  126 - 0x7e
    "11111111", -- 7403 - 0x1ceb  :  255 - 0xff
    "11111111", -- 7404 - 0x1cec  :  255 - 0xff
    "11111111", -- 7405 - 0x1ced  :  255 - 0xff
    "01000010", -- 7406 - 0x1cee  :   66 - 0x42
    "00000000", -- 7407 - 0x1cef  :    0 - 0x0
    "00111100", -- 7408 - 0x1cf0  :   60 - 0x3c
    "01000010", -- 7409 - 0x1cf1  :   66 - 0x42
    "10011001", -- 7410 - 0x1cf2  :  153 - 0x99
    "10100001", -- 7411 - 0x1cf3  :  161 - 0xa1
    "10100001", -- 7412 - 0x1cf4  :  161 - 0xa1
    "10011001", -- 7413 - 0x1cf5  :  153 - 0x99
    "01000010", -- 7414 - 0x1cf6  :   66 - 0x42
    "00111100", -- 7415 - 0x1cf7  :   60 - 0x3c
    "00000000", -- 7416 - 0x1cf8  :    0 - 0x0
    "00000000", -- 7417 - 0x1cf9  :    0 - 0x0
    "00000000", -- 7418 - 0x1cfa  :    0 - 0x0
    "00000000", -- 7419 - 0x1cfb  :    0 - 0x0
    "00000000", -- 7420 - 0x1cfc  :    0 - 0x0
    "00000000", -- 7421 - 0x1cfd  :    0 - 0x0
    "00000000", -- 7422 - 0x1cfe  :    0 - 0x0
    "00000000", -- 7423 - 0x1cff  :    0 - 0x0
    "00001111", -- 7424 - 0x1d00  :   15 - 0xf
    "00011111", -- 7425 - 0x1d01  :   31 - 0x1f
    "00011111", -- 7426 - 0x1d02  :   31 - 0x1f
    "00111111", -- 7427 - 0x1d03  :   63 - 0x3f
    "00111111", -- 7428 - 0x1d04  :   63 - 0x3f
    "01111111", -- 7429 - 0x1d05  :  127 - 0x7f
    "01111111", -- 7430 - 0x1d06  :  127 - 0x7f
    "01111111", -- 7431 - 0x1d07  :  127 - 0x7f
    "11110000", -- 7432 - 0x1d08  :  240 - 0xf0
    "11100000", -- 7433 - 0x1d09  :  224 - 0xe0
    "11100000", -- 7434 - 0x1d0a  :  224 - 0xe0
    "11000000", -- 7435 - 0x1d0b  :  192 - 0xc0
    "11000000", -- 7436 - 0x1d0c  :  192 - 0xc0
    "10000000", -- 7437 - 0x1d0d  :  128 - 0x80
    "10000000", -- 7438 - 0x1d0e  :  128 - 0x80
    "10000000", -- 7439 - 0x1d0f  :  128 - 0x80
    "11110000", -- 7440 - 0x1d10  :  240 - 0xf0
    "11111000", -- 7441 - 0x1d11  :  248 - 0xf8
    "11111000", -- 7442 - 0x1d12  :  248 - 0xf8
    "11111100", -- 7443 - 0x1d13  :  252 - 0xfc
    "11111100", -- 7444 - 0x1d14  :  252 - 0xfc
    "11111110", -- 7445 - 0x1d15  :  254 - 0xfe
    "11111110", -- 7446 - 0x1d16  :  254 - 0xfe
    "11111110", -- 7447 - 0x1d17  :  254 - 0xfe
    "00001111", -- 7448 - 0x1d18  :   15 - 0xf
    "00000111", -- 7449 - 0x1d19  :    7 - 0x7
    "00000111", -- 7450 - 0x1d1a  :    7 - 0x7
    "00000011", -- 7451 - 0x1d1b  :    3 - 0x3
    "00000011", -- 7452 - 0x1d1c  :    3 - 0x3
    "00000001", -- 7453 - 0x1d1d  :    1 - 0x1
    "00000001", -- 7454 - 0x1d1e  :    1 - 0x1
    "00000001", -- 7455 - 0x1d1f  :    1 - 0x1
    "01111111", -- 7456 - 0x1d20  :  127 - 0x7f
    "01111111", -- 7457 - 0x1d21  :  127 - 0x7f
    "00111111", -- 7458 - 0x1d22  :   63 - 0x3f
    "00111111", -- 7459 - 0x1d23  :   63 - 0x3f
    "00111111", -- 7460 - 0x1d24  :   63 - 0x3f
    "00111111", -- 7461 - 0x1d25  :   63 - 0x3f
    "00011111", -- 7462 - 0x1d26  :   31 - 0x1f
    "00011111", -- 7463 - 0x1d27  :   31 - 0x1f
    "10000000", -- 7464 - 0x1d28  :  128 - 0x80
    "10000000", -- 7465 - 0x1d29  :  128 - 0x80
    "11000000", -- 7466 - 0x1d2a  :  192 - 0xc0
    "11000000", -- 7467 - 0x1d2b  :  192 - 0xc0
    "11100000", -- 7468 - 0x1d2c  :  224 - 0xe0
    "11111000", -- 7469 - 0x1d2d  :  248 - 0xf8
    "11111110", -- 7470 - 0x1d2e  :  254 - 0xfe
    "11111111", -- 7471 - 0x1d2f  :  255 - 0xff
    "11111110", -- 7472 - 0x1d30  :  254 - 0xfe
    "11111111", -- 7473 - 0x1d31  :  255 - 0xff
    "11111111", -- 7474 - 0x1d32  :  255 - 0xff
    "11111111", -- 7475 - 0x1d33  :  255 - 0xff
    "11111100", -- 7476 - 0x1d34  :  252 - 0xfc
    "11111100", -- 7477 - 0x1d35  :  252 - 0xfc
    "11111110", -- 7478 - 0x1d36  :  254 - 0xfe
    "11111110", -- 7479 - 0x1d37  :  254 - 0xfe
    "11111111", -- 7480 - 0x1d38  :  255 - 0xff
    "01111111", -- 7481 - 0x1d39  :  127 - 0x7f
    "00011111", -- 7482 - 0x1d3a  :   31 - 0x1f
    "00000111", -- 7483 - 0x1d3b  :    7 - 0x7
    "00000011", -- 7484 - 0x1d3c  :    3 - 0x3
    "00000011", -- 7485 - 0x1d3d  :    3 - 0x3
    "00000001", -- 7486 - 0x1d3e  :    1 - 0x1
    "10000001", -- 7487 - 0x1d3f  :  129 - 0x81
    "01111111", -- 7488 - 0x1d40  :  127 - 0x7f
    "01111111", -- 7489 - 0x1d41  :  127 - 0x7f
    "01111111", -- 7490 - 0x1d42  :  127 - 0x7f
    "00111111", -- 7491 - 0x1d43  :   63 - 0x3f
    "00111111", -- 7492 - 0x1d44  :   63 - 0x3f
    "00111111", -- 7493 - 0x1d45  :   63 - 0x3f
    "00111111", -- 7494 - 0x1d46  :   63 - 0x3f
    "00011111", -- 7495 - 0x1d47  :   31 - 0x1f
    "10000000", -- 7496 - 0x1d48  :  128 - 0x80
    "10000000", -- 7497 - 0x1d49  :  128 - 0x80
    "10000000", -- 7498 - 0x1d4a  :  128 - 0x80
    "11000000", -- 7499 - 0x1d4b  :  192 - 0xc0
    "11000000", -- 7500 - 0x1d4c  :  192 - 0xc0
    "11100000", -- 7501 - 0x1d4d  :  224 - 0xe0
    "11100000", -- 7502 - 0x1d4e  :  224 - 0xe0
    "11110000", -- 7503 - 0x1d4f  :  240 - 0xf0
    "11111110", -- 7504 - 0x1d50  :  254 - 0xfe
    "11111110", -- 7505 - 0x1d51  :  254 - 0xfe
    "11111111", -- 7506 - 0x1d52  :  255 - 0xff
    "11111111", -- 7507 - 0x1d53  :  255 - 0xff
    "11111111", -- 7508 - 0x1d54  :  255 - 0xff
    "11111111", -- 7509 - 0x1d55  :  255 - 0xff
    "11111111", -- 7510 - 0x1d56  :  255 - 0xff
    "11111110", -- 7511 - 0x1d57  :  254 - 0xfe
    "00000001", -- 7512 - 0x1d58  :    1 - 0x1
    "00000001", -- 7513 - 0x1d59  :    1 - 0x1
    "00000001", -- 7514 - 0x1d5a  :    1 - 0x1
    "00000011", -- 7515 - 0x1d5b  :    3 - 0x3
    "00000011", -- 7516 - 0x1d5c  :    3 - 0x3
    "00000111", -- 7517 - 0x1d5d  :    7 - 0x7
    "00000111", -- 7518 - 0x1d5e  :    7 - 0x7
    "00001111", -- 7519 - 0x1d5f  :   15 - 0xf
    "00011111", -- 7520 - 0x1d60  :   31 - 0x1f
    "00001111", -- 7521 - 0x1d61  :   15 - 0xf
    "00001111", -- 7522 - 0x1d62  :   15 - 0xf
    "00000111", -- 7523 - 0x1d63  :    7 - 0x7
    "00000000", -- 7524 - 0x1d64  :    0 - 0x0
    "00000000", -- 7525 - 0x1d65  :    0 - 0x0
    "00000000", -- 7526 - 0x1d66  :    0 - 0x0
    "00000000", -- 7527 - 0x1d67  :    0 - 0x0
    "11111111", -- 7528 - 0x1d68  :  255 - 0xff
    "11111111", -- 7529 - 0x1d69  :  255 - 0xff
    "11111111", -- 7530 - 0x1d6a  :  255 - 0xff
    "11111111", -- 7531 - 0x1d6b  :  255 - 0xff
    "11111111", -- 7532 - 0x1d6c  :  255 - 0xff
    "11111111", -- 7533 - 0x1d6d  :  255 - 0xff
    "11111111", -- 7534 - 0x1d6e  :  255 - 0xff
    "11111111", -- 7535 - 0x1d6f  :  255 - 0xff
    "11111110", -- 7536 - 0x1d70  :  254 - 0xfe
    "11111100", -- 7537 - 0x1d71  :  252 - 0xfc
    "11111100", -- 7538 - 0x1d72  :  252 - 0xfc
    "11111000", -- 7539 - 0x1d73  :  248 - 0xf8
    "00000000", -- 7540 - 0x1d74  :    0 - 0x0
    "00000000", -- 7541 - 0x1d75  :    0 - 0x0
    "00000000", -- 7542 - 0x1d76  :    0 - 0x0
    "00000000", -- 7543 - 0x1d77  :    0 - 0x0
    "11111111", -- 7544 - 0x1d78  :  255 - 0xff
    "11111111", -- 7545 - 0x1d79  :  255 - 0xff
    "11111111", -- 7546 - 0x1d7a  :  255 - 0xff
    "11111111", -- 7547 - 0x1d7b  :  255 - 0xff
    "11111111", -- 7548 - 0x1d7c  :  255 - 0xff
    "11111111", -- 7549 - 0x1d7d  :  255 - 0xff
    "11111111", -- 7550 - 0x1d7e  :  255 - 0xff
    "11111111", -- 7551 - 0x1d7f  :  255 - 0xff
    "01111110", -- 7552 - 0x1d80  :  126 - 0x7e
    "01111110", -- 7553 - 0x1d81  :  126 - 0x7e
    "01111110", -- 7554 - 0x1d82  :  126 - 0x7e
    "01111110", -- 7555 - 0x1d83  :  126 - 0x7e
    "01111111", -- 7556 - 0x1d84  :  127 - 0x7f
    "01111111", -- 7557 - 0x1d85  :  127 - 0x7f
    "01111111", -- 7558 - 0x1d86  :  127 - 0x7f
    "01111111", -- 7559 - 0x1d87  :  127 - 0x7f
    "10000001", -- 7560 - 0x1d88  :  129 - 0x81
    "10000001", -- 7561 - 0x1d89  :  129 - 0x81
    "10000001", -- 7562 - 0x1d8a  :  129 - 0x81
    "10000001", -- 7563 - 0x1d8b  :  129 - 0x81
    "10000001", -- 7564 - 0x1d8c  :  129 - 0x81
    "10000001", -- 7565 - 0x1d8d  :  129 - 0x81
    "10000001", -- 7566 - 0x1d8e  :  129 - 0x81
    "10000001", -- 7567 - 0x1d8f  :  129 - 0x81
    "11111111", -- 7568 - 0x1d90  :  255 - 0xff
    "11111111", -- 7569 - 0x1d91  :  255 - 0xff
    "11111111", -- 7570 - 0x1d92  :  255 - 0xff
    "11111111", -- 7571 - 0x1d93  :  255 - 0xff
    "11111111", -- 7572 - 0x1d94  :  255 - 0xff
    "11111111", -- 7573 - 0x1d95  :  255 - 0xff
    "11111111", -- 7574 - 0x1d96  :  255 - 0xff
    "11111110", -- 7575 - 0x1d97  :  254 - 0xfe
    "00000001", -- 7576 - 0x1d98  :    1 - 0x1
    "00000001", -- 7577 - 0x1d99  :    1 - 0x1
    "00000001", -- 7578 - 0x1d9a  :    1 - 0x1
    "00000011", -- 7579 - 0x1d9b  :    3 - 0x3
    "00000011", -- 7580 - 0x1d9c  :    3 - 0x3
    "00000111", -- 7581 - 0x1d9d  :    7 - 0x7
    "00000111", -- 7582 - 0x1d9e  :    7 - 0x7
    "00001111", -- 7583 - 0x1d9f  :   15 - 0xf
    "11111110", -- 7584 - 0x1da0  :  254 - 0xfe
    "11111110", -- 7585 - 0x1da1  :  254 - 0xfe
    "11111110", -- 7586 - 0x1da2  :  254 - 0xfe
    "11111110", -- 7587 - 0x1da3  :  254 - 0xfe
    "11111111", -- 7588 - 0x1da4  :  255 - 0xff
    "11111111", -- 7589 - 0x1da5  :  255 - 0xff
    "11111111", -- 7590 - 0x1da6  :  255 - 0xff
    "11111111", -- 7591 - 0x1da7  :  255 - 0xff
    "00000001", -- 7592 - 0x1da8  :    1 - 0x1
    "00000001", -- 7593 - 0x1da9  :    1 - 0x1
    "00000001", -- 7594 - 0x1daa  :    1 - 0x1
    "00000001", -- 7595 - 0x1dab  :    1 - 0x1
    "00000001", -- 7596 - 0x1dac  :    1 - 0x1
    "00000001", -- 7597 - 0x1dad  :    1 - 0x1
    "00000001", -- 7598 - 0x1dae  :    1 - 0x1
    "00000001", -- 7599 - 0x1daf  :    1 - 0x1
    "01111111", -- 7600 - 0x1db0  :  127 - 0x7f
    "01111111", -- 7601 - 0x1db1  :  127 - 0x7f
    "01111111", -- 7602 - 0x1db2  :  127 - 0x7f
    "01111111", -- 7603 - 0x1db3  :  127 - 0x7f
    "01111111", -- 7604 - 0x1db4  :  127 - 0x7f
    "01111111", -- 7605 - 0x1db5  :  127 - 0x7f
    "01111111", -- 7606 - 0x1db6  :  127 - 0x7f
    "01111111", -- 7607 - 0x1db7  :  127 - 0x7f
    "10000001", -- 7608 - 0x1db8  :  129 - 0x81
    "10000001", -- 7609 - 0x1db9  :  129 - 0x81
    "10000001", -- 7610 - 0x1dba  :  129 - 0x81
    "10000001", -- 7611 - 0x1dbb  :  129 - 0x81
    "10000001", -- 7612 - 0x1dbc  :  129 - 0x81
    "10000001", -- 7613 - 0x1dbd  :  129 - 0x81
    "10000001", -- 7614 - 0x1dbe  :  129 - 0x81
    "10000001", -- 7615 - 0x1dbf  :  129 - 0x81
    "11111111", -- 7616 - 0x1dc0  :  255 - 0xff
    "11111111", -- 7617 - 0x1dc1  :  255 - 0xff
    "11111111", -- 7618 - 0x1dc2  :  255 - 0xff
    "11111111", -- 7619 - 0x1dc3  :  255 - 0xff
    "11111100", -- 7620 - 0x1dc4  :  252 - 0xfc
    "11111110", -- 7621 - 0x1dc5  :  254 - 0xfe
    "11111110", -- 7622 - 0x1dc6  :  254 - 0xfe
    "01111110", -- 7623 - 0x1dc7  :  126 - 0x7e
    "11111111", -- 7624 - 0x1dc8  :  255 - 0xff
    "00000011", -- 7625 - 0x1dc9  :    3 - 0x3
    "00000011", -- 7626 - 0x1dca  :    3 - 0x3
    "00000011", -- 7627 - 0x1dcb  :    3 - 0x3
    "00000011", -- 7628 - 0x1dcc  :    3 - 0x3
    "00000011", -- 7629 - 0x1dcd  :    3 - 0x3
    "00000011", -- 7630 - 0x1dce  :    3 - 0x3
    "11111111", -- 7631 - 0x1dcf  :  255 - 0xff
    "11111111", -- 7632 - 0x1dd0  :  255 - 0xff
    "11111111", -- 7633 - 0x1dd1  :  255 - 0xff
    "11111111", -- 7634 - 0x1dd2  :  255 - 0xff
    "11111111", -- 7635 - 0x1dd3  :  255 - 0xff
    "00000000", -- 7636 - 0x1dd4  :    0 - 0x0
    "00000000", -- 7637 - 0x1dd5  :    0 - 0x0
    "00000000", -- 7638 - 0x1dd6  :    0 - 0x0
    "00000000", -- 7639 - 0x1dd7  :    0 - 0x0
    "11111111", -- 7640 - 0x1dd8  :  255 - 0xff
    "11111111", -- 7641 - 0x1dd9  :  255 - 0xff
    "11111111", -- 7642 - 0x1dda  :  255 - 0xff
    "11111111", -- 7643 - 0x1ddb  :  255 - 0xff
    "11111111", -- 7644 - 0x1ddc  :  255 - 0xff
    "11111111", -- 7645 - 0x1ddd  :  255 - 0xff
    "11111111", -- 7646 - 0x1dde  :  255 - 0xff
    "11111111", -- 7647 - 0x1ddf  :  255 - 0xff
    "01111111", -- 7648 - 0x1de0  :  127 - 0x7f
    "01111111", -- 7649 - 0x1de1  :  127 - 0x7f
    "01111111", -- 7650 - 0x1de2  :  127 - 0x7f
    "01111111", -- 7651 - 0x1de3  :  127 - 0x7f
    "01111111", -- 7652 - 0x1de4  :  127 - 0x7f
    "01111111", -- 7653 - 0x1de5  :  127 - 0x7f
    "01111111", -- 7654 - 0x1de6  :  127 - 0x7f
    "01111111", -- 7655 - 0x1de7  :  127 - 0x7f
    "10000000", -- 7656 - 0x1de8  :  128 - 0x80
    "10000000", -- 7657 - 0x1de9  :  128 - 0x80
    "10000000", -- 7658 - 0x1dea  :  128 - 0x80
    "10000000", -- 7659 - 0x1deb  :  128 - 0x80
    "10000000", -- 7660 - 0x1dec  :  128 - 0x80
    "10000000", -- 7661 - 0x1ded  :  128 - 0x80
    "10000000", -- 7662 - 0x1dee  :  128 - 0x80
    "10000000", -- 7663 - 0x1def  :  128 - 0x80
    "11111111", -- 7664 - 0x1df0  :  255 - 0xff
    "11111111", -- 7665 - 0x1df1  :  255 - 0xff
    "11111111", -- 7666 - 0x1df2  :  255 - 0xff
    "11111111", -- 7667 - 0x1df3  :  255 - 0xff
    "11111111", -- 7668 - 0x1df4  :  255 - 0xff
    "11111111", -- 7669 - 0x1df5  :  255 - 0xff
    "11111111", -- 7670 - 0x1df6  :  255 - 0xff
    "11111110", -- 7671 - 0x1df7  :  254 - 0xfe
    "00000001", -- 7672 - 0x1df8  :    1 - 0x1
    "00000001", -- 7673 - 0x1df9  :    1 - 0x1
    "00000001", -- 7674 - 0x1dfa  :    1 - 0x1
    "00000011", -- 7675 - 0x1dfb  :    3 - 0x3
    "00000111", -- 7676 - 0x1dfc  :    7 - 0x7
    "00000011", -- 7677 - 0x1dfd  :    3 - 0x3
    "00000001", -- 7678 - 0x1dfe  :    1 - 0x1
    "00000001", -- 7679 - 0x1dff  :    1 - 0x1
    "01111110", -- 7680 - 0x1e00  :  126 - 0x7e
    "01111110", -- 7681 - 0x1e01  :  126 - 0x7e
    "01111111", -- 7682 - 0x1e02  :  127 - 0x7f
    "01111111", -- 7683 - 0x1e03  :  127 - 0x7f
    "01111111", -- 7684 - 0x1e04  :  127 - 0x7f
    "01111111", -- 7685 - 0x1e05  :  127 - 0x7f
    "01111111", -- 7686 - 0x1e06  :  127 - 0x7f
    "01111111", -- 7687 - 0x1e07  :  127 - 0x7f
    "10000001", -- 7688 - 0x1e08  :  129 - 0x81
    "10000001", -- 7689 - 0x1e09  :  129 - 0x81
    "10000001", -- 7690 - 0x1e0a  :  129 - 0x81
    "10000001", -- 7691 - 0x1e0b  :  129 - 0x81
    "10000001", -- 7692 - 0x1e0c  :  129 - 0x81
    "10000001", -- 7693 - 0x1e0d  :  129 - 0x81
    "10000001", -- 7694 - 0x1e0e  :  129 - 0x81
    "10000001", -- 7695 - 0x1e0f  :  129 - 0x81
    "00111111", -- 7696 - 0x1e10  :   63 - 0x3f
    "00111111", -- 7697 - 0x1e11  :   63 - 0x3f
    "00111111", -- 7698 - 0x1e12  :   63 - 0x3f
    "00111111", -- 7699 - 0x1e13  :   63 - 0x3f
    "00000000", -- 7700 - 0x1e14  :    0 - 0x0
    "00000000", -- 7701 - 0x1e15  :    0 - 0x0
    "00000000", -- 7702 - 0x1e16  :    0 - 0x0
    "00000000", -- 7703 - 0x1e17  :    0 - 0x0
    "11111111", -- 7704 - 0x1e18  :  255 - 0xff
    "11111111", -- 7705 - 0x1e19  :  255 - 0xff
    "11111111", -- 7706 - 0x1e1a  :  255 - 0xff
    "11111111", -- 7707 - 0x1e1b  :  255 - 0xff
    "11111111", -- 7708 - 0x1e1c  :  255 - 0xff
    "11111111", -- 7709 - 0x1e1d  :  255 - 0xff
    "11111111", -- 7710 - 0x1e1e  :  255 - 0xff
    "11111111", -- 7711 - 0x1e1f  :  255 - 0xff
    "01111110", -- 7712 - 0x1e20  :  126 - 0x7e
    "01111100", -- 7713 - 0x1e21  :  124 - 0x7c
    "01111100", -- 7714 - 0x1e22  :  124 - 0x7c
    "01111000", -- 7715 - 0x1e23  :  120 - 0x78
    "00000000", -- 7716 - 0x1e24  :    0 - 0x0
    "00000000", -- 7717 - 0x1e25  :    0 - 0x0
    "00000000", -- 7718 - 0x1e26  :    0 - 0x0
    "00000000", -- 7719 - 0x1e27  :    0 - 0x0
    "11111111", -- 7720 - 0x1e28  :  255 - 0xff
    "11111111", -- 7721 - 0x1e29  :  255 - 0xff
    "11111111", -- 7722 - 0x1e2a  :  255 - 0xff
    "11111111", -- 7723 - 0x1e2b  :  255 - 0xff
    "11111111", -- 7724 - 0x1e2c  :  255 - 0xff
    "11111111", -- 7725 - 0x1e2d  :  255 - 0xff
    "11111111", -- 7726 - 0x1e2e  :  255 - 0xff
    "11111111", -- 7727 - 0x1e2f  :  255 - 0xff
    "11111110", -- 7728 - 0x1e30  :  254 - 0xfe
    "11111110", -- 7729 - 0x1e31  :  254 - 0xfe
    "11111111", -- 7730 - 0x1e32  :  255 - 0xff
    "11111111", -- 7731 - 0x1e33  :  255 - 0xff
    "01111111", -- 7732 - 0x1e34  :  127 - 0x7f
    "01111111", -- 7733 - 0x1e35  :  127 - 0x7f
    "01111111", -- 7734 - 0x1e36  :  127 - 0x7f
    "01111111", -- 7735 - 0x1e37  :  127 - 0x7f
    "10000001", -- 7736 - 0x1e38  :  129 - 0x81
    "10000001", -- 7737 - 0x1e39  :  129 - 0x81
    "10000001", -- 7738 - 0x1e3a  :  129 - 0x81
    "10000001", -- 7739 - 0x1e3b  :  129 - 0x81
    "10000001", -- 7740 - 0x1e3c  :  129 - 0x81
    "10000001", -- 7741 - 0x1e3d  :  129 - 0x81
    "10000001", -- 7742 - 0x1e3e  :  129 - 0x81
    "10000001", -- 7743 - 0x1e3f  :  129 - 0x81
    "01111111", -- 7744 - 0x1e40  :  127 - 0x7f
    "01111111", -- 7745 - 0x1e41  :  127 - 0x7f
    "00111111", -- 7746 - 0x1e42  :   63 - 0x3f
    "00111111", -- 7747 - 0x1e43  :   63 - 0x3f
    "00111111", -- 7748 - 0x1e44  :   63 - 0x3f
    "00111111", -- 7749 - 0x1e45  :   63 - 0x3f
    "00011111", -- 7750 - 0x1e46  :   31 - 0x1f
    "00011111", -- 7751 - 0x1e47  :   31 - 0x1f
    "10000000", -- 7752 - 0x1e48  :  128 - 0x80
    "10000000", -- 7753 - 0x1e49  :  128 - 0x80
    "11000000", -- 7754 - 0x1e4a  :  192 - 0xc0
    "11000000", -- 7755 - 0x1e4b  :  192 - 0xc0
    "11100000", -- 7756 - 0x1e4c  :  224 - 0xe0
    "11111000", -- 7757 - 0x1e4d  :  248 - 0xf8
    "11111110", -- 7758 - 0x1e4e  :  254 - 0xfe
    "11111111", -- 7759 - 0x1e4f  :  255 - 0xff
    "00111111", -- 7760 - 0x1e50  :   63 - 0x3f
    "10111111", -- 7761 - 0x1e51  :  191 - 0xbf
    "11111111", -- 7762 - 0x1e52  :  255 - 0xff
    "11111111", -- 7763 - 0x1e53  :  255 - 0xff
    "11111100", -- 7764 - 0x1e54  :  252 - 0xfc
    "11111100", -- 7765 - 0x1e55  :  252 - 0xfc
    "11111110", -- 7766 - 0x1e56  :  254 - 0xfe
    "11111110", -- 7767 - 0x1e57  :  254 - 0xfe
    "11111111", -- 7768 - 0x1e58  :  255 - 0xff
    "01111111", -- 7769 - 0x1e59  :  127 - 0x7f
    "00011111", -- 7770 - 0x1e5a  :   31 - 0x1f
    "00000111", -- 7771 - 0x1e5b  :    7 - 0x7
    "00000011", -- 7772 - 0x1e5c  :    3 - 0x3
    "00000011", -- 7773 - 0x1e5d  :    3 - 0x3
    "00000001", -- 7774 - 0x1e5e  :    1 - 0x1
    "10000001", -- 7775 - 0x1e5f  :  129 - 0x81
    "01111111", -- 7776 - 0x1e60  :  127 - 0x7f
    "01111111", -- 7777 - 0x1e61  :  127 - 0x7f
    "01111110", -- 7778 - 0x1e62  :  126 - 0x7e
    "01111110", -- 7779 - 0x1e63  :  126 - 0x7e
    "01111111", -- 7780 - 0x1e64  :  127 - 0x7f
    "01111111", -- 7781 - 0x1e65  :  127 - 0x7f
    "01111111", -- 7782 - 0x1e66  :  127 - 0x7f
    "01111111", -- 7783 - 0x1e67  :  127 - 0x7f
    "10000001", -- 7784 - 0x1e68  :  129 - 0x81
    "10000001", -- 7785 - 0x1e69  :  129 - 0x81
    "10000001", -- 7786 - 0x1e6a  :  129 - 0x81
    "10000001", -- 7787 - 0x1e6b  :  129 - 0x81
    "10000001", -- 7788 - 0x1e6c  :  129 - 0x81
    "10000001", -- 7789 - 0x1e6d  :  129 - 0x81
    "10000001", -- 7790 - 0x1e6e  :  129 - 0x81
    "10000001", -- 7791 - 0x1e6f  :  129 - 0x81
    "01111110", -- 7792 - 0x1e70  :  126 - 0x7e
    "01111110", -- 7793 - 0x1e71  :  126 - 0x7e
    "01111110", -- 7794 - 0x1e72  :  126 - 0x7e
    "01111110", -- 7795 - 0x1e73  :  126 - 0x7e
    "01111111", -- 7796 - 0x1e74  :  127 - 0x7f
    "01111111", -- 7797 - 0x1e75  :  127 - 0x7f
    "01111111", -- 7798 - 0x1e76  :  127 - 0x7f
    "01111111", -- 7799 - 0x1e77  :  127 - 0x7f
    "10000001", -- 7800 - 0x1e78  :  129 - 0x81
    "10000001", -- 7801 - 0x1e79  :  129 - 0x81
    "10000001", -- 7802 - 0x1e7a  :  129 - 0x81
    "10000001", -- 7803 - 0x1e7b  :  129 - 0x81
    "10000001", -- 7804 - 0x1e7c  :  129 - 0x81
    "10000001", -- 7805 - 0x1e7d  :  129 - 0x81
    "10000001", -- 7806 - 0x1e7e  :  129 - 0x81
    "10000001", -- 7807 - 0x1e7f  :  129 - 0x81
    "10000001", -- 7808 - 0x1e80  :  129 - 0x81
    "11000011", -- 7809 - 0x1e81  :  195 - 0xc3
    "11000011", -- 7810 - 0x1e82  :  195 - 0xc3
    "11100111", -- 7811 - 0x1e83  :  231 - 0xe7
    "11100111", -- 7812 - 0x1e84  :  231 - 0xe7
    "11111111", -- 7813 - 0x1e85  :  255 - 0xff
    "11111111", -- 7814 - 0x1e86  :  255 - 0xff
    "11111111", -- 7815 - 0x1e87  :  255 - 0xff
    "01111110", -- 7816 - 0x1e88  :  126 - 0x7e
    "00111100", -- 7817 - 0x1e89  :   60 - 0x3c
    "00111100", -- 7818 - 0x1e8a  :   60 - 0x3c
    "00011000", -- 7819 - 0x1e8b  :   24 - 0x18
    "00011000", -- 7820 - 0x1e8c  :   24 - 0x18
    "00000000", -- 7821 - 0x1e8d  :    0 - 0x0
    "00000000", -- 7822 - 0x1e8e  :    0 - 0x0
    "00000000", -- 7823 - 0x1e8f  :    0 - 0x0
    "00001111", -- 7824 - 0x1e90  :   15 - 0xf
    "01000011", -- 7825 - 0x1e91  :   67 - 0x43
    "01011011", -- 7826 - 0x1e92  :   91 - 0x5b
    "01010011", -- 7827 - 0x1e93  :   83 - 0x53
    "00110001", -- 7828 - 0x1e94  :   49 - 0x31
    "00011001", -- 7829 - 0x1e95  :   25 - 0x19
    "00001111", -- 7830 - 0x1e96  :   15 - 0xf
    "00000111", -- 7831 - 0x1e97  :    7 - 0x7
    "11110010", -- 7832 - 0x1e98  :  242 - 0xf2
    "11111110", -- 7833 - 0x1e99  :  254 - 0xfe
    "11111110", -- 7834 - 0x1e9a  :  254 - 0xfe
    "11111111", -- 7835 - 0x1e9b  :  255 - 0xff
    "11111111", -- 7836 - 0x1e9c  :  255 - 0xff
    "11101111", -- 7837 - 0x1e9d  :  239 - 0xef
    "11110111", -- 7838 - 0x1e9e  :  247 - 0xf7
    "11111000", -- 7839 - 0x1e9f  :  248 - 0xf8
    "11000001", -- 7840 - 0x1ea0  :  193 - 0xc1
    "11000011", -- 7841 - 0x1ea1  :  195 - 0xc3
    "11000110", -- 7842 - 0x1ea2  :  198 - 0xc6
    "10000100", -- 7843 - 0x1ea3  :  132 - 0x84
    "11111100", -- 7844 - 0x1ea4  :  252 - 0xfc
    "11111100", -- 7845 - 0x1ea5  :  252 - 0xfc
    "00001110", -- 7846 - 0x1ea6  :   14 - 0xe
    "00000010", -- 7847 - 0x1ea7  :    2 - 0x2
    "10111111", -- 7848 - 0x1ea8  :  191 - 0xbf
    "10111110", -- 7849 - 0x1ea9  :  190 - 0xbe
    "10111101", -- 7850 - 0x1eaa  :  189 - 0xbd
    "01111011", -- 7851 - 0x1eab  :  123 - 0x7b
    "01111011", -- 7852 - 0x1eac  :  123 - 0x7b
    "00000111", -- 7853 - 0x1ead  :    7 - 0x7
    "11110011", -- 7854 - 0x1eae  :  243 - 0xf3
    "11111101", -- 7855 - 0x1eaf  :  253 - 0xfd
    "00010000", -- 7856 - 0x1eb0  :   16 - 0x10
    "00100000", -- 7857 - 0x1eb1  :   32 - 0x20
    "00100010", -- 7858 - 0x1eb2  :   34 - 0x22
    "10111010", -- 7859 - 0x1eb3  :  186 - 0xba
    "11100110", -- 7860 - 0x1eb4  :  230 - 0xe6
    "11100001", -- 7861 - 0x1eb5  :  225 - 0xe1
    "11000000", -- 7862 - 0x1eb6  :  192 - 0xc0
    "11000000", -- 7863 - 0x1eb7  :  192 - 0xc0
    "11111111", -- 7864 - 0x1eb8  :  255 - 0xff
    "11111111", -- 7865 - 0x1eb9  :  255 - 0xff
    "11111111", -- 7866 - 0x1eba  :  255 - 0xff
    "01100111", -- 7867 - 0x1ebb  :  103 - 0x67
    "01011001", -- 7868 - 0x1ebc  :   89 - 0x59
    "10011110", -- 7869 - 0x1ebd  :  158 - 0x9e
    "10111111", -- 7870 - 0x1ebe  :  191 - 0xbf
    "10111111", -- 7871 - 0x1ebf  :  191 - 0xbf
    "00100000", -- 7872 - 0x1ec0  :   32 - 0x20
    "10100110", -- 7873 - 0x1ec1  :  166 - 0xa6
    "01010100", -- 7874 - 0x1ec2  :   84 - 0x54
    "00100110", -- 7875 - 0x1ec3  :   38 - 0x26
    "00100000", -- 7876 - 0x1ec4  :   32 - 0x20
    "11000110", -- 7877 - 0x1ec5  :  198 - 0xc6
    "01010100", -- 7878 - 0x1ec6  :   84 - 0x54
    "00100110", -- 7879 - 0x1ec7  :   38 - 0x26
    "00100000", -- 7880 - 0x1ec8  :   32 - 0x20
    "11100110", -- 7881 - 0x1ec9  :  230 - 0xe6
    "01010100", -- 7882 - 0x1eca  :   84 - 0x54
    "00100110", -- 7883 - 0x1ecb  :   38 - 0x26
    "00100001", -- 7884 - 0x1ecc  :   33 - 0x21
    "00000110", -- 7885 - 0x1ecd  :    6 - 0x6
    "01010100", -- 7886 - 0x1ece  :   84 - 0x54
    "00100110", -- 7887 - 0x1ecf  :   38 - 0x26
    "00100000", -- 7888 - 0x1ed0  :   32 - 0x20
    "10000101", -- 7889 - 0x1ed1  :  133 - 0x85
    "00000001", -- 7890 - 0x1ed2  :    1 - 0x1
    "01000100", -- 7891 - 0x1ed3  :   68 - 0x44
    "00100000", -- 7892 - 0x1ed4  :   32 - 0x20
    "10000110", -- 7893 - 0x1ed5  :  134 - 0x86
    "01010100", -- 7894 - 0x1ed6  :   84 - 0x54
    "01001000", -- 7895 - 0x1ed7  :   72 - 0x48
    "00100000", -- 7896 - 0x1ed8  :   32 - 0x20
    "10011010", -- 7897 - 0x1ed9  :  154 - 0x9a
    "00000001", -- 7898 - 0x1eda  :    1 - 0x1
    "01001001", -- 7899 - 0x1edb  :   73 - 0x49
    "00100000", -- 7900 - 0x1edc  :   32 - 0x20
    "10100101", -- 7901 - 0x1edd  :  165 - 0xa5
    "11001001", -- 7902 - 0x1ede  :  201 - 0xc9
    "01000110", -- 7903 - 0x1edf  :   70 - 0x46
    "00100000", -- 7904 - 0x1ee0  :   32 - 0x20
    "10111010", -- 7905 - 0x1ee1  :  186 - 0xba
    "11001001", -- 7906 - 0x1ee2  :  201 - 0xc9
    "01001010", -- 7907 - 0x1ee3  :   74 - 0x4a
    "00100000", -- 7908 - 0x1ee4  :   32 - 0x20
    "10100110", -- 7909 - 0x1ee5  :  166 - 0xa6
    "00001010", -- 7910 - 0x1ee6  :   10 - 0xa
    "11010000", -- 7911 - 0x1ee7  :  208 - 0xd0
    "11010001", -- 7912 - 0x1ee8  :  209 - 0xd1
    "11011000", -- 7913 - 0x1ee9  :  216 - 0xd8
    "11011000", -- 7914 - 0x1eea  :  216 - 0xd8
    "11011110", -- 7915 - 0x1eeb  :  222 - 0xde
    "11010001", -- 7916 - 0x1eec  :  209 - 0xd1
    "11010000", -- 7917 - 0x1eed  :  208 - 0xd0
    "11011010", -- 7918 - 0x1eee  :  218 - 0xda
    "11011110", -- 7919 - 0x1eef  :  222 - 0xde
    "11010001", -- 7920 - 0x1ef0  :  209 - 0xd1
    "00100000", -- 7921 - 0x1ef1  :   32 - 0x20
    "11000110", -- 7922 - 0x1ef2  :  198 - 0xc6
    "00001010", -- 7923 - 0x1ef3  :   10 - 0xa
    "11010010", -- 7924 - 0x1ef4  :  210 - 0xd2
    "11010011", -- 7925 - 0x1ef5  :  211 - 0xd3
    "11011011", -- 7926 - 0x1ef6  :  219 - 0xdb
    "11011011", -- 7927 - 0x1ef7  :  219 - 0xdb
    "11011011", -- 7928 - 0x1ef8  :  219 - 0xdb
    "11011001", -- 7929 - 0x1ef9  :  217 - 0xd9
    "11011011", -- 7930 - 0x1efa  :  219 - 0xdb
    "11011100", -- 7931 - 0x1efb  :  220 - 0xdc
    "11011011", -- 7932 - 0x1efc  :  219 - 0xdb
    "11011111", -- 7933 - 0x1efd  :  223 - 0xdf
    "00100000", -- 7934 - 0x1efe  :   32 - 0x20
    "11100110", -- 7935 - 0x1eff  :  230 - 0xe6
    "00001010", -- 7936 - 0x1f00  :   10 - 0xa
    "11010100", -- 7937 - 0x1f01  :  212 - 0xd4
    "11010101", -- 7938 - 0x1f02  :  213 - 0xd5
    "11010100", -- 7939 - 0x1f03  :  212 - 0xd4
    "11011001", -- 7940 - 0x1f04  :  217 - 0xd9
    "11011011", -- 7941 - 0x1f05  :  219 - 0xdb
    "11100010", -- 7942 - 0x1f06  :  226 - 0xe2
    "11010100", -- 7943 - 0x1f07  :  212 - 0xd4
    "11011010", -- 7944 - 0x1f08  :  218 - 0xda
    "11011011", -- 7945 - 0x1f09  :  219 - 0xdb
    "11100000", -- 7946 - 0x1f0a  :  224 - 0xe0
    "00100001", -- 7947 - 0x1f0b  :   33 - 0x21
    "00000110", -- 7948 - 0x1f0c  :    6 - 0x6
    "00001010", -- 7949 - 0x1f0d  :   10 - 0xa
    "11010110", -- 7950 - 0x1f0e  :  214 - 0xd6
    "11010111", -- 7951 - 0x1f0f  :  215 - 0xd7
    "11010110", -- 7952 - 0x1f10  :  214 - 0xd6
    "11010111", -- 7953 - 0x1f11  :  215 - 0xd7
    "11100001", -- 7954 - 0x1f12  :  225 - 0xe1
    "00100110", -- 7955 - 0x1f13  :   38 - 0x26
    "11010110", -- 7956 - 0x1f14  :  214 - 0xd6
    "11011101", -- 7957 - 0x1f15  :  221 - 0xdd
    "11100001", -- 7958 - 0x1f16  :  225 - 0xe1
    "11100001", -- 7959 - 0x1f17  :  225 - 0xe1
    "00100001", -- 7960 - 0x1f18  :   33 - 0x21
    "00100110", -- 7961 - 0x1f19  :   38 - 0x26
    "00010100", -- 7962 - 0x1f1a  :   20 - 0x14
    "11010000", -- 7963 - 0x1f1b  :  208 - 0xd0
    "11101000", -- 7964 - 0x1f1c  :  232 - 0xe8
    "11010001", -- 7965 - 0x1f1d  :  209 - 0xd1
    "11010000", -- 7966 - 0x1f1e  :  208 - 0xd0
    "11010001", -- 7967 - 0x1f1f  :  209 - 0xd1
    "11011110", -- 7968 - 0x1f20  :  222 - 0xde
    "11010001", -- 7969 - 0x1f21  :  209 - 0xd1
    "11011000", -- 7970 - 0x1f22  :  216 - 0xd8
    "11010000", -- 7971 - 0x1f23  :  208 - 0xd0
    "11010001", -- 7972 - 0x1f24  :  209 - 0xd1
    "00100110", -- 7973 - 0x1f25  :   38 - 0x26
    "11011110", -- 7974 - 0x1f26  :  222 - 0xde
    "11010001", -- 7975 - 0x1f27  :  209 - 0xd1
    "11011110", -- 7976 - 0x1f28  :  222 - 0xde
    "11010001", -- 7977 - 0x1f29  :  209 - 0xd1
    "11010000", -- 7978 - 0x1f2a  :  208 - 0xd0
    "11010001", -- 7979 - 0x1f2b  :  209 - 0xd1
    "11010000", -- 7980 - 0x1f2c  :  208 - 0xd0
    "11010001", -- 7981 - 0x1f2d  :  209 - 0xd1
    "00100110", -- 7982 - 0x1f2e  :   38 - 0x26
    "00100001", -- 7983 - 0x1f2f  :   33 - 0x21
    "01000110", -- 7984 - 0x1f30  :   70 - 0x46
    "00010100", -- 7985 - 0x1f31  :   20 - 0x14
    "11011011", -- 7986 - 0x1f32  :  219 - 0xdb
    "01000010", -- 7987 - 0x1f33  :   66 - 0x42
    "01000010", -- 7988 - 0x1f34  :   66 - 0x42
    "11011011", -- 7989 - 0x1f35  :  219 - 0xdb
    "01000010", -- 7990 - 0x1f36  :   66 - 0x42
    "11011011", -- 7991 - 0x1f37  :  219 - 0xdb
    "01000010", -- 7992 - 0x1f38  :   66 - 0x42
    "11011011", -- 7993 - 0x1f39  :  219 - 0xdb
    "11011011", -- 7994 - 0x1f3a  :  219 - 0xdb
    "01000010", -- 7995 - 0x1f3b  :   66 - 0x42
    "00100110", -- 7996 - 0x1f3c  :   38 - 0x26
    "11011011", -- 7997 - 0x1f3d  :  219 - 0xdb
    "01000010", -- 7998 - 0x1f3e  :   66 - 0x42
    "11011011", -- 7999 - 0x1f3f  :  219 - 0xdb
    "01000010", -- 8000 - 0x1f40  :   66 - 0x42
    "11011011", -- 8001 - 0x1f41  :  219 - 0xdb
    "01000010", -- 8002 - 0x1f42  :   66 - 0x42
    "11011011", -- 8003 - 0x1f43  :  219 - 0xdb
    "01000010", -- 8004 - 0x1f44  :   66 - 0x42
    "00100110", -- 8005 - 0x1f45  :   38 - 0x26
    "00100001", -- 8006 - 0x1f46  :   33 - 0x21
    "01100110", -- 8007 - 0x1f47  :  102 - 0x66
    "01000110", -- 8008 - 0x1f48  :   70 - 0x46
    "11011011", -- 8009 - 0x1f49  :  219 - 0xdb
    "00100001", -- 8010 - 0x1f4a  :   33 - 0x21
    "01101100", -- 8011 - 0x1f4b  :  108 - 0x6c
    "00001110", -- 8012 - 0x1f4c  :   14 - 0xe
    "11011111", -- 8013 - 0x1f4d  :  223 - 0xdf
    "11011011", -- 8014 - 0x1f4e  :  219 - 0xdb
    "11011011", -- 8015 - 0x1f4f  :  219 - 0xdb
    "11011011", -- 8016 - 0x1f50  :  219 - 0xdb
    "00100110", -- 8017 - 0x1f51  :   38 - 0x26
    "11011011", -- 8018 - 0x1f52  :  219 - 0xdb
    "11011111", -- 8019 - 0x1f53  :  223 - 0xdf
    "11011011", -- 8020 - 0x1f54  :  219 - 0xdb
    "11011111", -- 8021 - 0x1f55  :  223 - 0xdf
    "11011011", -- 8022 - 0x1f56  :  219 - 0xdb
    "11011011", -- 8023 - 0x1f57  :  219 - 0xdb
    "11100100", -- 8024 - 0x1f58  :  228 - 0xe4
    "11100101", -- 8025 - 0x1f59  :  229 - 0xe5
    "00100110", -- 8026 - 0x1f5a  :   38 - 0x26
    "00100001", -- 8027 - 0x1f5b  :   33 - 0x21
    "10000110", -- 8028 - 0x1f5c  :  134 - 0x86
    "00010100", -- 8029 - 0x1f5d  :   20 - 0x14
    "11011011", -- 8030 - 0x1f5e  :  219 - 0xdb
    "11011011", -- 8031 - 0x1f5f  :  219 - 0xdb
    "11011011", -- 8032 - 0x1f60  :  219 - 0xdb
    "11011110", -- 8033 - 0x1f61  :  222 - 0xde
    "01000011", -- 8034 - 0x1f62  :   67 - 0x43
    "11011011", -- 8035 - 0x1f63  :  219 - 0xdb
    "11100000", -- 8036 - 0x1f64  :  224 - 0xe0
    "11011011", -- 8037 - 0x1f65  :  219 - 0xdb
    "11011011", -- 8038 - 0x1f66  :  219 - 0xdb
    "11011011", -- 8039 - 0x1f67  :  219 - 0xdb
    "00100110", -- 8040 - 0x1f68  :   38 - 0x26
    "11011011", -- 8041 - 0x1f69  :  219 - 0xdb
    "11100011", -- 8042 - 0x1f6a  :  227 - 0xe3
    "11011011", -- 8043 - 0x1f6b  :  219 - 0xdb
    "11100000", -- 8044 - 0x1f6c  :  224 - 0xe0
    "11011011", -- 8045 - 0x1f6d  :  219 - 0xdb
    "11011011", -- 8046 - 0x1f6e  :  219 - 0xdb
    "11100110", -- 8047 - 0x1f6f  :  230 - 0xe6
    "11100011", -- 8048 - 0x1f70  :  227 - 0xe3
    "00100110", -- 8049 - 0x1f71  :   38 - 0x26
    "00100001", -- 8050 - 0x1f72  :   33 - 0x21
    "10100110", -- 8051 - 0x1f73  :  166 - 0xa6
    "00010100", -- 8052 - 0x1f74  :   20 - 0x14
    "11011011", -- 8053 - 0x1f75  :  219 - 0xdb
    "11011011", -- 8054 - 0x1f76  :  219 - 0xdb
    "11011011", -- 8055 - 0x1f77  :  219 - 0xdb
    "11011011", -- 8056 - 0x1f78  :  219 - 0xdb
    "01000010", -- 8057 - 0x1f79  :   66 - 0x42
    "11011011", -- 8058 - 0x1f7a  :  219 - 0xdb
    "11011011", -- 8059 - 0x1f7b  :  219 - 0xdb
    "11011011", -- 8060 - 0x1f7c  :  219 - 0xdb
    "11010100", -- 8061 - 0x1f7d  :  212 - 0xd4
    "11011001", -- 8062 - 0x1f7e  :  217 - 0xd9
    "00100110", -- 8063 - 0x1f7f  :   38 - 0x26
    "11011011", -- 8064 - 0x1f80  :  219 - 0xdb
    "11011001", -- 8065 - 0x1f81  :  217 - 0xd9
    "11011011", -- 8066 - 0x1f82  :  219 - 0xdb
    "11011011", -- 8067 - 0x1f83  :  219 - 0xdb
    "11010100", -- 8068 - 0x1f84  :  212 - 0xd4
    "11011001", -- 8069 - 0x1f85  :  217 - 0xd9
    "11010100", -- 8070 - 0x1f86  :  212 - 0xd4
    "11011001", -- 8071 - 0x1f87  :  217 - 0xd9
    "11100111", -- 8072 - 0x1f88  :  231 - 0xe7
    "00100001", -- 8073 - 0x1f89  :   33 - 0x21
    "11000101", -- 8074 - 0x1f8a  :  197 - 0xc5
    "00010110", -- 8075 - 0x1f8b  :   22 - 0x16
    "01011111", -- 8076 - 0x1f8c  :   95 - 0x5f
    "10010101", -- 8077 - 0x1f8d  :  149 - 0x95
    "10010101", -- 8078 - 0x1f8e  :  149 - 0x95
    "10010101", -- 8079 - 0x1f8f  :  149 - 0x95
    "10010101", -- 8080 - 0x1f90  :  149 - 0x95
    "10010101", -- 8081 - 0x1f91  :  149 - 0x95
    "10010101", -- 8082 - 0x1f92  :  149 - 0x95
    "10010101", -- 8083 - 0x1f93  :  149 - 0x95
    "10010101", -- 8084 - 0x1f94  :  149 - 0x95
    "10010111", -- 8085 - 0x1f95  :  151 - 0x97
    "10011000", -- 8086 - 0x1f96  :  152 - 0x98
    "01111000", -- 8087 - 0x1f97  :  120 - 0x78
    "10010101", -- 8088 - 0x1f98  :  149 - 0x95
    "10010110", -- 8089 - 0x1f99  :  150 - 0x96
    "10010101", -- 8090 - 0x1f9a  :  149 - 0x95
    "10010101", -- 8091 - 0x1f9b  :  149 - 0x95
    "10010111", -- 8092 - 0x1f9c  :  151 - 0x97
    "10011000", -- 8093 - 0x1f9d  :  152 - 0x98
    "10010111", -- 8094 - 0x1f9e  :  151 - 0x97
    "10011000", -- 8095 - 0x1f9f  :  152 - 0x98
    "10010101", -- 8096 - 0x1fa0  :  149 - 0x95
    "01111010", -- 8097 - 0x1fa1  :  122 - 0x7a
    "00100001", -- 8098 - 0x1fa2  :   33 - 0x21
    "11101101", -- 8099 - 0x1fa3  :  237 - 0xed
    "00001110", -- 8100 - 0x1fa4  :   14 - 0xe
    "11001111", -- 8101 - 0x1fa5  :  207 - 0xcf
    "00000001", -- 8102 - 0x1fa6  :    1 - 0x1
    "00001001", -- 8103 - 0x1fa7  :    9 - 0x9
    "00001000", -- 8104 - 0x1fa8  :    8 - 0x8
    "00000101", -- 8105 - 0x1fa9  :    5 - 0x5
    "00100100", -- 8106 - 0x1faa  :   36 - 0x24
    "00010111", -- 8107 - 0x1fab  :   23 - 0x17
    "00010010", -- 8108 - 0x1fac  :   18 - 0x12
    "00010111", -- 8109 - 0x1fad  :   23 - 0x17
    "00011101", -- 8110 - 0x1fae  :   29 - 0x1d
    "00001110", -- 8111 - 0x1faf  :   14 - 0xe
    "00010111", -- 8112 - 0x1fb0  :   23 - 0x17
    "00001101", -- 8113 - 0x1fb1  :   13 - 0xd
    "00011000", -- 8114 - 0x1fb2  :   24 - 0x18
    "00100010", -- 8115 - 0x1fb3  :   34 - 0x22
    "01001011", -- 8116 - 0x1fb4  :   75 - 0x4b
    "00001101", -- 8117 - 0x1fb5  :   13 - 0xd
    "00000001", -- 8118 - 0x1fb6  :    1 - 0x1
    "00100100", -- 8119 - 0x1fb7  :   36 - 0x24
    "00011001", -- 8120 - 0x1fb8  :   25 - 0x19
    "00010101", -- 8121 - 0x1fb9  :   21 - 0x15
    "00001010", -- 8122 - 0x1fba  :   10 - 0xa
    "00100010", -- 8123 - 0x1fbb  :   34 - 0x22
    "00001110", -- 8124 - 0x1fbc  :   14 - 0xe
    "00011011", -- 8125 - 0x1fbd  :   27 - 0x1b
    "00100100", -- 8126 - 0x1fbe  :   36 - 0x24
    "00010000", -- 8127 - 0x1fbf  :   16 - 0x10
    "00001010", -- 8128 - 0x1fc0  :   10 - 0xa
    "00010110", -- 8129 - 0x1fc1  :   22 - 0x16
    "00001110", -- 8130 - 0x1fc2  :   14 - 0xe
    "00100010", -- 8131 - 0x1fc3  :   34 - 0x22
    "10001011", -- 8132 - 0x1fc4  :  139 - 0x8b
    "00001101", -- 8133 - 0x1fc5  :   13 - 0xd
    "00000010", -- 8134 - 0x1fc6  :    2 - 0x2
    "00100100", -- 8135 - 0x1fc7  :   36 - 0x24
    "00011001", -- 8136 - 0x1fc8  :   25 - 0x19
    "00010101", -- 8137 - 0x1fc9  :   21 - 0x15
    "00001010", -- 8138 - 0x1fca  :   10 - 0xa
    "00100010", -- 8139 - 0x1fcb  :   34 - 0x22
    "00001110", -- 8140 - 0x1fcc  :   14 - 0xe
    "00011011", -- 8141 - 0x1fcd  :   27 - 0x1b
    "00100100", -- 8142 - 0x1fce  :   36 - 0x24
    "00010000", -- 8143 - 0x1fcf  :   16 - 0x10
    "00001010", -- 8144 - 0x1fd0  :   10 - 0xa
    "00010110", -- 8145 - 0x1fd1  :   22 - 0x16
    "00001110", -- 8146 - 0x1fd2  :   14 - 0xe
    "00100010", -- 8147 - 0x1fd3  :   34 - 0x22
    "11101100", -- 8148 - 0x1fd4  :  236 - 0xec
    "00000100", -- 8149 - 0x1fd5  :    4 - 0x4
    "00011101", -- 8150 - 0x1fd6  :   29 - 0x1d
    "00011000", -- 8151 - 0x1fd7  :   24 - 0x18
    "00011001", -- 8152 - 0x1fd8  :   25 - 0x19
    "00101000", -- 8153 - 0x1fd9  :   40 - 0x28
    "00100010", -- 8154 - 0x1fda  :   34 - 0x22
    "11110110", -- 8155 - 0x1fdb  :  246 - 0xf6
    "00000001", -- 8156 - 0x1fdc  :    1 - 0x1
    "00000000", -- 8157 - 0x1fdd  :    0 - 0x0
    "00100011", -- 8158 - 0x1fde  :   35 - 0x23
    "11001001", -- 8159 - 0x1fdf  :  201 - 0xc9
    "01010110", -- 8160 - 0x1fe0  :   86 - 0x56
    "01010101", -- 8161 - 0x1fe1  :   85 - 0x55
    "00100011", -- 8162 - 0x1fe2  :   35 - 0x23
    "11100010", -- 8163 - 0x1fe3  :  226 - 0xe2
    "00000100", -- 8164 - 0x1fe4  :    4 - 0x4
    "10011001", -- 8165 - 0x1fe5  :  153 - 0x99
    "10101010", -- 8166 - 0x1fe6  :  170 - 0xaa
    "10101010", -- 8167 - 0x1fe7  :  170 - 0xaa
    "10101010", -- 8168 - 0x1fe8  :  170 - 0xaa
    "00100011", -- 8169 - 0x1fe9  :   35 - 0x23
    "11101010", -- 8170 - 0x1fea  :  234 - 0xea
    "00000100", -- 8171 - 0x1feb  :    4 - 0x4
    "10011001", -- 8172 - 0x1fec  :  153 - 0x99
    "10101010", -- 8173 - 0x1fed  :  170 - 0xaa
    "10101010", -- 8174 - 0x1fee  :  170 - 0xaa
    "10101010", -- 8175 - 0x1fef  :  170 - 0xaa
    "00000000", -- 8176 - 0x1ff0  :    0 - 0x0
    "11111111", -- 8177 - 0x1ff1  :  255 - 0xff
    "11111111", -- 8178 - 0x1ff2  :  255 - 0xff
    "11111111", -- 8179 - 0x1ff3  :  255 - 0xff
    "11111111", -- 8180 - 0x1ff4  :  255 - 0xff
    "11111111", -- 8181 - 0x1ff5  :  255 - 0xff
    "11111111", -- 8182 - 0x1ff6  :  255 - 0xff
    "11111111", -- 8183 - 0x1ff7  :  255 - 0xff
    "11111111", -- 8184 - 0x1ff8  :  255 - 0xff
    "11111111", -- 8185 - 0x1ff9  :  255 - 0xff
    "11111111", -- 8186 - 0x1ffa  :  255 - 0xff
    "11111111", -- 8187 - 0x1ffb  :  255 - 0xff
    "11111111", -- 8188 - 0x1ffc  :  255 - 0xff
    "11111111", -- 8189 - 0x1ffd  :  255 - 0xff
    "11111111", -- 8190 - 0x1ffe  :  255 - 0xff
    "11111111" -- 8191 - 0x1fff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= nametable_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
