//-   Sprites Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: pacman_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_PACMAN_SPR
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table both color planes
      12'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout <= 8'b00000011; //    1 :   3 - 0x3
      12'h2: dout <= 8'b00001111; //    2 :  15 - 0xf
      12'h3: dout <= 8'b00011111; //    3 :  31 - 0x1f
      12'h4: dout <= 8'b00111111; //    4 :  63 - 0x3f
      12'h5: dout <= 8'b00111111; //    5 :  63 - 0x3f
      12'h6: dout <= 8'b01111111; //    6 : 127 - 0x7f
      12'h7: dout <= 8'b01111111; //    7 : 127 - 0x7f
      12'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- plane 1
      12'h9: dout <= 8'b00000000; //    9 :   0 - 0x0
      12'hA: dout <= 8'b00000000; //   10 :   0 - 0x0
      12'hB: dout <= 8'b00000000; //   11 :   0 - 0x0
      12'hC: dout <= 8'b00000000; //   12 :   0 - 0x0
      12'hD: dout <= 8'b00000000; //   13 :   0 - 0x0
      12'hE: dout <= 8'b00000000; //   14 :   0 - 0x0
      12'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      12'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x1
      12'h11: dout <= 8'b11000000; //   17 : 192 - 0xc0
      12'h12: dout <= 8'b11110000; //   18 : 240 - 0xf0
      12'h13: dout <= 8'b11111000; //   19 : 248 - 0xf8
      12'h14: dout <= 8'b11111000; //   20 : 248 - 0xf8
      12'h15: dout <= 8'b11111100; //   21 : 252 - 0xfc
      12'h16: dout <= 8'b11111100; //   22 : 252 - 0xfc
      12'h17: dout <= 8'b11111100; //   23 : 252 - 0xfc
      12'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- plane 1
      12'h19: dout <= 8'b00000000; //   25 :   0 - 0x0
      12'h1A: dout <= 8'b00000000; //   26 :   0 - 0x0
      12'h1B: dout <= 8'b00000000; //   27 :   0 - 0x0
      12'h1C: dout <= 8'b00000000; //   28 :   0 - 0x0
      12'h1D: dout <= 8'b00000000; //   29 :   0 - 0x0
      12'h1E: dout <= 8'b00000000; //   30 :   0 - 0x0
      12'h1F: dout <= 8'b00000000; //   31 :   0 - 0x0
      12'h20: dout <= 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x2
      12'h21: dout <= 8'b00000111; //   33 :   7 - 0x7
      12'h22: dout <= 8'b00011111; //   34 :  31 - 0x1f
      12'h23: dout <= 8'b00111111; //   35 :  63 - 0x3f
      12'h24: dout <= 8'b00111111; //   36 :  63 - 0x3f
      12'h25: dout <= 8'b00001111; //   37 :  15 - 0xf
      12'h26: dout <= 8'b00000011; //   38 :   3 - 0x3
      12'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout <= 8'b00000000; //   40 :   0 - 0x0 -- plane 1
      12'h29: dout <= 8'b00000000; //   41 :   0 - 0x0
      12'h2A: dout <= 8'b00000000; //   42 :   0 - 0x0
      12'h2B: dout <= 8'b00000000; //   43 :   0 - 0x0
      12'h2C: dout <= 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout <= 8'b00000000; //   45 :   0 - 0x0
      12'h2E: dout <= 8'b00000000; //   46 :   0 - 0x0
      12'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout <= 8'b00000000; //   48 :   0 - 0x0 -- Sprite 0x3
      12'h31: dout <= 8'b00000000; //   49 :   0 - 0x0
      12'h32: dout <= 8'b00000111; //   50 :   7 - 0x7
      12'h33: dout <= 8'b00011111; //   51 :  31 - 0x1f
      12'h34: dout <= 8'b00111111; //   52 :  63 - 0x3f
      12'h35: dout <= 8'b00111111; //   53 :  63 - 0x3f
      12'h36: dout <= 8'b01111111; //   54 : 127 - 0x7f
      12'h37: dout <= 8'b01111111; //   55 : 127 - 0x7f
      12'h38: dout <= 8'b00000000; //   56 :   0 - 0x0 -- plane 1
      12'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      12'h3A: dout <= 8'b00000000; //   58 :   0 - 0x0
      12'h3B: dout <= 8'b00000000; //   59 :   0 - 0x0
      12'h3C: dout <= 8'b00000000; //   60 :   0 - 0x0
      12'h3D: dout <= 8'b00000000; //   61 :   0 - 0x0
      12'h3E: dout <= 8'b00000000; //   62 :   0 - 0x0
      12'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout <= 8'b01111110; //   64 : 126 - 0x7e -- Sprite 0x4
      12'h41: dout <= 8'b01111110; //   65 : 126 - 0x7e
      12'h42: dout <= 8'b01111100; //   66 : 124 - 0x7c
      12'h43: dout <= 8'b00111100; //   67 :  60 - 0x3c
      12'h44: dout <= 8'b00111000; //   68 :  56 - 0x38
      12'h45: dout <= 8'b00011000; //   69 :  24 - 0x18
      12'h46: dout <= 8'b00000000; //   70 :   0 - 0x0
      12'h47: dout <= 8'b00000000; //   71 :   0 - 0x0
      12'h48: dout <= 8'b00000000; //   72 :   0 - 0x0 -- plane 1
      12'h49: dout <= 8'b00000000; //   73 :   0 - 0x0
      12'h4A: dout <= 8'b00000000; //   74 :   0 - 0x0
      12'h4B: dout <= 8'b00000000; //   75 :   0 - 0x0
      12'h4C: dout <= 8'b00000000; //   76 :   0 - 0x0
      12'h4D: dout <= 8'b00000000; //   77 :   0 - 0x0
      12'h4E: dout <= 8'b00000000; //   78 :   0 - 0x0
      12'h4F: dout <= 8'b00000000; //   79 :   0 - 0x0
      12'h50: dout <= 8'b00000000; //   80 :   0 - 0x0 -- Sprite 0x5
      12'h51: dout <= 8'b11000000; //   81 : 192 - 0xc0
      12'h52: dout <= 8'b11110000; //   82 : 240 - 0xf0
      12'h53: dout <= 8'b11111000; //   83 : 248 - 0xf8
      12'h54: dout <= 8'b11111000; //   84 : 248 - 0xf8
      12'h55: dout <= 8'b11111100; //   85 : 252 - 0xfc
      12'h56: dout <= 8'b01111100; //   86 : 124 - 0x7c
      12'h57: dout <= 8'b00111100; //   87 :  60 - 0x3c
      12'h58: dout <= 8'b00000000; //   88 :   0 - 0x0 -- plane 1
      12'h59: dout <= 8'b00000000; //   89 :   0 - 0x0
      12'h5A: dout <= 8'b00000000; //   90 :   0 - 0x0
      12'h5B: dout <= 8'b00000000; //   91 :   0 - 0x0
      12'h5C: dout <= 8'b00000000; //   92 :   0 - 0x0
      12'h5D: dout <= 8'b00000000; //   93 :   0 - 0x0
      12'h5E: dout <= 8'b00000000; //   94 :   0 - 0x0
      12'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0x6
      12'h61: dout <= 8'b00000111; //   97 :   7 - 0x7
      12'h62: dout <= 8'b00000111; //   98 :   7 - 0x7
      12'h63: dout <= 8'b00000011; //   99 :   3 - 0x3
      12'h64: dout <= 8'b00000001; //  100 :   1 - 0x1
      12'h65: dout <= 8'b00000000; //  101 :   0 - 0x0
      12'h66: dout <= 8'b00000000; //  102 :   0 - 0x0
      12'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      12'h68: dout <= 8'b00000000; //  104 :   0 - 0x0 -- plane 1
      12'h69: dout <= 8'b00000000; //  105 :   0 - 0x0
      12'h6A: dout <= 8'b00000000; //  106 :   0 - 0x0
      12'h6B: dout <= 8'b00000000; //  107 :   0 - 0x0
      12'h6C: dout <= 8'b00000000; //  108 :   0 - 0x0
      12'h6D: dout <= 8'b00000000; //  109 :   0 - 0x0
      12'h6E: dout <= 8'b00000000; //  110 :   0 - 0x0
      12'h6F: dout <= 8'b00000000; //  111 :   0 - 0x0
      12'h70: dout <= 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0x7
      12'h71: dout <= 8'b00000000; //  113 :   0 - 0x0
      12'h72: dout <= 8'b00000111; //  114 :   7 - 0x7
      12'h73: dout <= 8'b00011111; //  115 :  31 - 0x1f
      12'h74: dout <= 8'b00111111; //  116 :  63 - 0x3f
      12'h75: dout <= 8'b00111111; //  117 :  63 - 0x3f
      12'h76: dout <= 8'b01111110; //  118 : 126 - 0x7e
      12'h77: dout <= 8'b01111100; //  119 : 124 - 0x7c
      12'h78: dout <= 8'b00000000; //  120 :   0 - 0x0 -- plane 1
      12'h79: dout <= 8'b00000000; //  121 :   0 - 0x0
      12'h7A: dout <= 8'b00000000; //  122 :   0 - 0x0
      12'h7B: dout <= 8'b00000000; //  123 :   0 - 0x0
      12'h7C: dout <= 8'b00000000; //  124 :   0 - 0x0
      12'h7D: dout <= 8'b00000000; //  125 :   0 - 0x0
      12'h7E: dout <= 8'b00000000; //  126 :   0 - 0x0
      12'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout <= 8'b01111000; //  128 : 120 - 0x78 -- Sprite 0x8
      12'h81: dout <= 8'b01110000; //  129 : 112 - 0x70
      12'h82: dout <= 8'b01100000; //  130 :  96 - 0x60
      12'h83: dout <= 8'b00000000; //  131 :   0 - 0x0
      12'h84: dout <= 8'b00000000; //  132 :   0 - 0x0
      12'h85: dout <= 8'b00000000; //  133 :   0 - 0x0
      12'h86: dout <= 8'b00000000; //  134 :   0 - 0x0
      12'h87: dout <= 8'b00000000; //  135 :   0 - 0x0
      12'h88: dout <= 8'b00000000; //  136 :   0 - 0x0 -- plane 1
      12'h89: dout <= 8'b00000000; //  137 :   0 - 0x0
      12'h8A: dout <= 8'b00000000; //  138 :   0 - 0x0
      12'h8B: dout <= 8'b00000000; //  139 :   0 - 0x0
      12'h8C: dout <= 8'b00000000; //  140 :   0 - 0x0
      12'h8D: dout <= 8'b00000000; //  141 :   0 - 0x0
      12'h8E: dout <= 8'b00000000; //  142 :   0 - 0x0
      12'h8F: dout <= 8'b00000000; //  143 :   0 - 0x0
      12'h90: dout <= 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x9
      12'h91: dout <= 8'b00000000; //  145 :   0 - 0x0
      12'h92: dout <= 8'b00000000; //  146 :   0 - 0x0
      12'h93: dout <= 8'b00000000; //  147 :   0 - 0x0
      12'h94: dout <= 8'b00000000; //  148 :   0 - 0x0
      12'h95: dout <= 8'b01000000; //  149 :  64 - 0x40
      12'h96: dout <= 8'b11110000; //  150 : 240 - 0xf0
      12'h97: dout <= 8'b11111000; //  151 : 248 - 0xf8
      12'h98: dout <= 8'b00000000; //  152 :   0 - 0x0 -- plane 1
      12'h99: dout <= 8'b00000000; //  153 :   0 - 0x0
      12'h9A: dout <= 8'b00000000; //  154 :   0 - 0x0
      12'h9B: dout <= 8'b00000000; //  155 :   0 - 0x0
      12'h9C: dout <= 8'b00000000; //  156 :   0 - 0x0
      12'h9D: dout <= 8'b00000000; //  157 :   0 - 0x0
      12'h9E: dout <= 8'b00000000; //  158 :   0 - 0x0
      12'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      12'hA0: dout <= 8'b11111110; //  160 : 254 - 0xfe -- Sprite 0xa
      12'hA1: dout <= 8'b01111111; //  161 : 127 - 0x7f
      12'hA2: dout <= 8'b01111111; //  162 : 127 - 0x7f
      12'hA3: dout <= 8'b00111111; //  163 :  63 - 0x3f
      12'hA4: dout <= 8'b00001110; //  164 :  14 - 0xe
      12'hA5: dout <= 8'b00000000; //  165 :   0 - 0x0
      12'hA6: dout <= 8'b00000000; //  166 :   0 - 0x0
      12'hA7: dout <= 8'b00000000; //  167 :   0 - 0x0
      12'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0 -- plane 1
      12'hA9: dout <= 8'b00000000; //  169 :   0 - 0x0
      12'hAA: dout <= 8'b00000000; //  170 :   0 - 0x0
      12'hAB: dout <= 8'b00000000; //  171 :   0 - 0x0
      12'hAC: dout <= 8'b00000000; //  172 :   0 - 0x0
      12'hAD: dout <= 8'b00000000; //  173 :   0 - 0x0
      12'hAE: dout <= 8'b00000000; //  174 :   0 - 0x0
      12'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      12'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0xb
      12'hB1: dout <= 8'b00000000; //  177 :   0 - 0x0
      12'hB2: dout <= 8'b00000000; //  178 :   0 - 0x0
      12'hB3: dout <= 8'b00000000; //  179 :   0 - 0x0
      12'hB4: dout <= 8'b00000000; //  180 :   0 - 0x0
      12'hB5: dout <= 8'b00000000; //  181 :   0 - 0x0
      12'hB6: dout <= 8'b00000000; //  182 :   0 - 0x0
      12'hB7: dout <= 8'b11100000; //  183 : 224 - 0xe0
      12'hB8: dout <= 8'b00000000; //  184 :   0 - 0x0 -- plane 1
      12'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      12'hBA: dout <= 8'b00000000; //  186 :   0 - 0x0
      12'hBB: dout <= 8'b00000000; //  187 :   0 - 0x0
      12'hBC: dout <= 8'b00000000; //  188 :   0 - 0x0
      12'hBD: dout <= 8'b00000000; //  189 :   0 - 0x0
      12'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      12'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout <= 8'b11111100; //  192 : 252 - 0xfc -- Sprite 0xc
      12'hC1: dout <= 8'b11111111; //  193 : 255 - 0xff
      12'hC2: dout <= 8'b01111111; //  194 : 127 - 0x7f
      12'hC3: dout <= 8'b00111111; //  195 :  63 - 0x3f
      12'hC4: dout <= 8'b00001110; //  196 :  14 - 0xe
      12'hC5: dout <= 8'b00000000; //  197 :   0 - 0x0
      12'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      12'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      12'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0 -- plane 1
      12'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      12'hCA: dout <= 8'b00000000; //  202 :   0 - 0x0
      12'hCB: dout <= 8'b00000000; //  203 :   0 - 0x0
      12'hCC: dout <= 8'b00000000; //  204 :   0 - 0x0
      12'hCD: dout <= 8'b00000000; //  205 :   0 - 0x0
      12'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      12'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      12'hD0: dout <= 8'b11110000; //  208 : 240 - 0xf0 -- Sprite 0xd
      12'hD1: dout <= 8'b11111111; //  209 : 255 - 0xff
      12'hD2: dout <= 8'b11111111; //  210 : 255 - 0xff
      12'hD3: dout <= 8'b01111111; //  211 : 127 - 0x7f
      12'hD4: dout <= 8'b00011110; //  212 :  30 - 0x1e
      12'hD5: dout <= 8'b00000000; //  213 :   0 - 0x0
      12'hD6: dout <= 8'b00000000; //  214 :   0 - 0x0
      12'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      12'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- plane 1
      12'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      12'hDA: dout <= 8'b00000000; //  218 :   0 - 0x0
      12'hDB: dout <= 8'b00000000; //  219 :   0 - 0x0
      12'hDC: dout <= 8'b00000000; //  220 :   0 - 0x0
      12'hDD: dout <= 8'b00000000; //  221 :   0 - 0x0
      12'hDE: dout <= 8'b00000000; //  222 :   0 - 0x0
      12'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      12'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0xe
      12'hE1: dout <= 8'b00001111; //  225 :  15 - 0xf
      12'hE2: dout <= 8'b11111111; //  226 : 255 - 0xff
      12'hE3: dout <= 8'b11111111; //  227 : 255 - 0xff
      12'hE4: dout <= 8'b01111111; //  228 : 127 - 0x7f
      12'hE5: dout <= 8'b00011110; //  229 :  30 - 0x1e
      12'hE6: dout <= 8'b00000000; //  230 :   0 - 0x0
      12'hE7: dout <= 8'b00000000; //  231 :   0 - 0x0
      12'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0 -- plane 1
      12'hE9: dout <= 8'b00000000; //  233 :   0 - 0x0
      12'hEA: dout <= 8'b00000000; //  234 :   0 - 0x0
      12'hEB: dout <= 8'b00000000; //  235 :   0 - 0x0
      12'hEC: dout <= 8'b00000000; //  236 :   0 - 0x0
      12'hED: dout <= 8'b00000000; //  237 :   0 - 0x0
      12'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      12'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      12'hF0: dout <= 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0xf
      12'hF1: dout <= 8'b00000011; //  241 :   3 - 0x3
      12'hF2: dout <= 8'b00001111; //  242 :  15 - 0xf
      12'hF3: dout <= 8'b01111111; //  243 : 127 - 0x7f
      12'hF4: dout <= 8'b11111111; //  244 : 255 - 0xff
      12'hF5: dout <= 8'b01111110; //  245 : 126 - 0x7e
      12'hF6: dout <= 8'b00011100; //  246 :  28 - 0x1c
      12'hF7: dout <= 8'b00000000; //  247 :   0 - 0x0
      12'hF8: dout <= 8'b00000000; //  248 :   0 - 0x0 -- plane 1
      12'hF9: dout <= 8'b00000000; //  249 :   0 - 0x0
      12'hFA: dout <= 8'b00000000; //  250 :   0 - 0x0
      12'hFB: dout <= 8'b00000000; //  251 :   0 - 0x0
      12'hFC: dout <= 8'b00000000; //  252 :   0 - 0x0
      12'hFD: dout <= 8'b00000000; //  253 :   0 - 0x0
      12'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      12'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x10
      12'h101: dout <= 8'b00000001; //  257 :   1 - 0x1
      12'h102: dout <= 8'b00000011; //  258 :   3 - 0x3
      12'h103: dout <= 8'b00001111; //  259 :  15 - 0xf
      12'h104: dout <= 8'b00011111; //  260 :  31 - 0x1f
      12'h105: dout <= 8'b01111111; //  261 : 127 - 0x7f
      12'h106: dout <= 8'b01111110; //  262 : 126 - 0x7e
      12'h107: dout <= 8'b00111100; //  263 :  60 - 0x3c
      12'h108: dout <= 8'b00000000; //  264 :   0 - 0x0 -- plane 1
      12'h109: dout <= 8'b00000000; //  265 :   0 - 0x0
      12'h10A: dout <= 8'b00000000; //  266 :   0 - 0x0
      12'h10B: dout <= 8'b00000000; //  267 :   0 - 0x0
      12'h10C: dout <= 8'b00000000; //  268 :   0 - 0x0
      12'h10D: dout <= 8'b00000000; //  269 :   0 - 0x0
      12'h10E: dout <= 8'b00000000; //  270 :   0 - 0x0
      12'h10F: dout <= 8'b00000000; //  271 :   0 - 0x0
      12'h110: dout <= 8'b00000000; //  272 :   0 - 0x0 -- Sprite 0x11
      12'h111: dout <= 8'b00000001; //  273 :   1 - 0x1
      12'h112: dout <= 8'b00000011; //  274 :   3 - 0x3
      12'h113: dout <= 8'b00000111; //  275 :   7 - 0x7
      12'h114: dout <= 8'b00000111; //  276 :   7 - 0x7
      12'h115: dout <= 8'b00001111; //  277 :  15 - 0xf
      12'h116: dout <= 8'b00011111; //  278 :  31 - 0x1f
      12'h117: dout <= 8'b00001110; //  279 :  14 - 0xe
      12'h118: dout <= 8'b00000000; //  280 :   0 - 0x0 -- plane 1
      12'h119: dout <= 8'b00000000; //  281 :   0 - 0x0
      12'h11A: dout <= 8'b00000000; //  282 :   0 - 0x0
      12'h11B: dout <= 8'b00000000; //  283 :   0 - 0x0
      12'h11C: dout <= 8'b00000000; //  284 :   0 - 0x0
      12'h11D: dout <= 8'b00000000; //  285 :   0 - 0x0
      12'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      12'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      12'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x12
      12'h121: dout <= 8'b00000000; //  289 :   0 - 0x0
      12'h122: dout <= 8'b00000001; //  290 :   1 - 0x1
      12'h123: dout <= 8'b00000011; //  291 :   3 - 0x3
      12'h124: dout <= 8'b00000011; //  292 :   3 - 0x3
      12'h125: dout <= 8'b00000011; //  293 :   3 - 0x3
      12'h126: dout <= 8'b00000111; //  294 :   7 - 0x7
      12'h127: dout <= 8'b00000010; //  295 :   2 - 0x2
      12'h128: dout <= 8'b00000000; //  296 :   0 - 0x0 -- plane 1
      12'h129: dout <= 8'b00000000; //  297 :   0 - 0x0
      12'h12A: dout <= 8'b00000000; //  298 :   0 - 0x0
      12'h12B: dout <= 8'b00000000; //  299 :   0 - 0x0
      12'h12C: dout <= 8'b00000000; //  300 :   0 - 0x0
      12'h12D: dout <= 8'b00000000; //  301 :   0 - 0x0
      12'h12E: dout <= 8'b00000000; //  302 :   0 - 0x0
      12'h12F: dout <= 8'b00000000; //  303 :   0 - 0x0
      12'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x13
      12'h131: dout <= 8'b00000000; //  305 :   0 - 0x0
      12'h132: dout <= 8'b00000001; //  306 :   1 - 0x1
      12'h133: dout <= 8'b00000001; //  307 :   1 - 0x1
      12'h134: dout <= 8'b00000001; //  308 :   1 - 0x1
      12'h135: dout <= 8'b00000001; //  309 :   1 - 0x1
      12'h136: dout <= 8'b00000001; //  310 :   1 - 0x1
      12'h137: dout <= 8'b00000001; //  311 :   1 - 0x1
      12'h138: dout <= 8'b00000000; //  312 :   0 - 0x0 -- plane 1
      12'h139: dout <= 8'b00000000; //  313 :   0 - 0x0
      12'h13A: dout <= 8'b00000000; //  314 :   0 - 0x0
      12'h13B: dout <= 8'b00000000; //  315 :   0 - 0x0
      12'h13C: dout <= 8'b00000000; //  316 :   0 - 0x0
      12'h13D: dout <= 8'b00000000; //  317 :   0 - 0x0
      12'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x14
      12'h141: dout <= 8'b00000000; //  321 :   0 - 0x0
      12'h142: dout <= 8'b00000000; //  322 :   0 - 0x0
      12'h143: dout <= 8'b00000000; //  323 :   0 - 0x0
      12'h144: dout <= 8'b00000000; //  324 :   0 - 0x0
      12'h145: dout <= 8'b00000000; //  325 :   0 - 0x0
      12'h146: dout <= 8'b00000100; //  326 :   4 - 0x4
      12'h147: dout <= 8'b00000010; //  327 :   2 - 0x2
      12'h148: dout <= 8'b00000000; //  328 :   0 - 0x0 -- plane 1
      12'h149: dout <= 8'b00000000; //  329 :   0 - 0x0
      12'h14A: dout <= 8'b00000000; //  330 :   0 - 0x0
      12'h14B: dout <= 8'b00000000; //  331 :   0 - 0x0
      12'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      12'h14D: dout <= 8'b00000000; //  333 :   0 - 0x0
      12'h14E: dout <= 8'b00000000; //  334 :   0 - 0x0
      12'h14F: dout <= 8'b00000000; //  335 :   0 - 0x0
      12'h150: dout <= 8'b00000000; //  336 :   0 - 0x0 -- Sprite 0x15
      12'h151: dout <= 8'b00000000; //  337 :   0 - 0x0
      12'h152: dout <= 8'b00000000; //  338 :   0 - 0x0
      12'h153: dout <= 8'b00000000; //  339 :   0 - 0x0
      12'h154: dout <= 8'b00000000; //  340 :   0 - 0x0
      12'h155: dout <= 8'b00000000; //  341 :   0 - 0x0
      12'h156: dout <= 8'b00100000; //  342 :  32 - 0x20
      12'h157: dout <= 8'b01001000; //  343 :  72 - 0x48
      12'h158: dout <= 8'b00000000; //  344 :   0 - 0x0 -- plane 1
      12'h159: dout <= 8'b00000000; //  345 :   0 - 0x0
      12'h15A: dout <= 8'b00000000; //  346 :   0 - 0x0
      12'h15B: dout <= 8'b00000000; //  347 :   0 - 0x0
      12'h15C: dout <= 8'b00000000; //  348 :   0 - 0x0
      12'h15D: dout <= 8'b00000000; //  349 :   0 - 0x0
      12'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      12'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout <= 8'b00010000; //  352 :  16 - 0x10 -- Sprite 0x16
      12'h161: dout <= 8'b00001000; //  353 :   8 - 0x8
      12'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      12'h163: dout <= 8'b00110000; //  355 :  48 - 0x30
      12'h164: dout <= 8'b00000000; //  356 :   0 - 0x0
      12'h165: dout <= 8'b00001000; //  357 :   8 - 0x8
      12'h166: dout <= 8'b00010010; //  358 :  18 - 0x12
      12'h167: dout <= 8'b00000100; //  359 :   4 - 0x4
      12'h168: dout <= 8'b00000000; //  360 :   0 - 0x0 -- plane 1
      12'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      12'h16A: dout <= 8'b00000000; //  362 :   0 - 0x0
      12'h16B: dout <= 8'b00000000; //  363 :   0 - 0x0
      12'h16C: dout <= 8'b00000000; //  364 :   0 - 0x0
      12'h16D: dout <= 8'b00000000; //  365 :   0 - 0x0
      12'h16E: dout <= 8'b00000000; //  366 :   0 - 0x0
      12'h16F: dout <= 8'b00000000; //  367 :   0 - 0x0
      12'h170: dout <= 8'b00010000; //  368 :  16 - 0x10 -- Sprite 0x17
      12'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      12'h172: dout <= 8'b00001100; //  370 :  12 - 0xc
      12'h173: dout <= 8'b00000000; //  371 :   0 - 0x0
      12'h174: dout <= 8'b00010000; //  372 :  16 - 0x10
      12'h175: dout <= 8'b00001000; //  373 :   8 - 0x8
      12'h176: dout <= 8'b01000000; //  374 :  64 - 0x40
      12'h177: dout <= 8'b00100000; //  375 :  32 - 0x20
      12'h178: dout <= 8'b00000000; //  376 :   0 - 0x0 -- plane 1
      12'h179: dout <= 8'b00000000; //  377 :   0 - 0x0
      12'h17A: dout <= 8'b00000000; //  378 :   0 - 0x0
      12'h17B: dout <= 8'b00000000; //  379 :   0 - 0x0
      12'h17C: dout <= 8'b00000000; //  380 :   0 - 0x0
      12'h17D: dout <= 8'b00000000; //  381 :   0 - 0x0
      12'h17E: dout <= 8'b00000000; //  382 :   0 - 0x0
      12'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      12'h180: dout <= 8'b00000000; //  384 :   0 - 0x0 -- Sprite 0x18
      12'h181: dout <= 8'b00000000; //  385 :   0 - 0x0
      12'h182: dout <= 8'b00000011; //  386 :   3 - 0x3
      12'h183: dout <= 8'b00000011; //  387 :   3 - 0x3
      12'h184: dout <= 8'b00000001; //  388 :   1 - 0x1
      12'h185: dout <= 8'b00100001; //  389 :  33 - 0x21
      12'h186: dout <= 8'b00100001; //  390 :  33 - 0x21
      12'h187: dout <= 8'b01110011; //  391 : 115 - 0x73
      12'h188: dout <= 8'b00000000; //  392 :   0 - 0x0 -- plane 1
      12'h189: dout <= 8'b00000000; //  393 :   0 - 0x0
      12'h18A: dout <= 8'b00000011; //  394 :   3 - 0x3
      12'h18B: dout <= 8'b00000011; //  395 :   3 - 0x3
      12'h18C: dout <= 8'b00010011; //  396 :  19 - 0x13
      12'h18D: dout <= 8'b00111111; //  397 :  63 - 0x3f
      12'h18E: dout <= 8'b00111111; //  398 :  63 - 0x3f
      12'h18F: dout <= 8'b01111111; //  399 : 127 - 0x7f
      12'h190: dout <= 8'b01111111; //  400 : 127 - 0x7f -- Sprite 0x19
      12'h191: dout <= 8'b01111111; //  401 : 127 - 0x7f
      12'h192: dout <= 8'b01111111; //  402 : 127 - 0x7f
      12'h193: dout <= 8'b01111111; //  403 : 127 - 0x7f
      12'h194: dout <= 8'b01101110; //  404 : 110 - 0x6e
      12'h195: dout <= 8'b01000110; //  405 :  70 - 0x46
      12'h196: dout <= 8'b00000000; //  406 :   0 - 0x0
      12'h197: dout <= 8'b00000000; //  407 :   0 - 0x0
      12'h198: dout <= 8'b01111111; //  408 : 127 - 0x7f -- plane 1
      12'h199: dout <= 8'b01111111; //  409 : 127 - 0x7f
      12'h19A: dout <= 8'b01111111; //  410 : 127 - 0x7f
      12'h19B: dout <= 8'b01111111; //  411 : 127 - 0x7f
      12'h19C: dout <= 8'b01101110; //  412 : 110 - 0x6e
      12'h19D: dout <= 8'b01000110; //  413 :  70 - 0x46
      12'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      12'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout <= 8'b01111111; //  416 : 127 - 0x7f -- Sprite 0x1a
      12'h1A1: dout <= 8'b01111111; //  417 : 127 - 0x7f
      12'h1A2: dout <= 8'b01111111; //  418 : 127 - 0x7f
      12'h1A3: dout <= 8'b01111111; //  419 : 127 - 0x7f
      12'h1A4: dout <= 8'b01111011; //  420 : 123 - 0x7b
      12'h1A5: dout <= 8'b00110001; //  421 :  49 - 0x31
      12'h1A6: dout <= 8'b00000000; //  422 :   0 - 0x0
      12'h1A7: dout <= 8'b00000000; //  423 :   0 - 0x0
      12'h1A8: dout <= 8'b01111111; //  424 : 127 - 0x7f -- plane 1
      12'h1A9: dout <= 8'b01111111; //  425 : 127 - 0x7f
      12'h1AA: dout <= 8'b01111111; //  426 : 127 - 0x7f
      12'h1AB: dout <= 8'b01111111; //  427 : 127 - 0x7f
      12'h1AC: dout <= 8'b01111011; //  428 : 123 - 0x7b
      12'h1AD: dout <= 8'b00110001; //  429 :  49 - 0x31
      12'h1AE: dout <= 8'b00000000; //  430 :   0 - 0x0
      12'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      12'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x1b
      12'h1B1: dout <= 8'b00000011; //  433 :   3 - 0x3
      12'h1B2: dout <= 8'b00001111; //  434 :  15 - 0xf
      12'h1B3: dout <= 8'b00011111; //  435 :  31 - 0x1f
      12'h1B4: dout <= 8'b00100111; //  436 :  39 - 0x27
      12'h1B5: dout <= 8'b00000011; //  437 :   3 - 0x3
      12'h1B6: dout <= 8'b00000011; //  438 :   3 - 0x3
      12'h1B7: dout <= 8'b01000011; //  439 :  67 - 0x43
      12'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0 -- plane 1
      12'h1B9: dout <= 8'b00000011; //  441 :   3 - 0x3
      12'h1BA: dout <= 8'b00001111; //  442 :  15 - 0xf
      12'h1BB: dout <= 8'b00011111; //  443 :  31 - 0x1f
      12'h1BC: dout <= 8'b00111111; //  444 :  63 - 0x3f
      12'h1BD: dout <= 8'b00111111; //  445 :  63 - 0x3f
      12'h1BE: dout <= 8'b00001111; //  446 :  15 - 0xf
      12'h1BF: dout <= 8'b01001111; //  447 :  79 - 0x4f
      12'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x1c
      12'h1C1: dout <= 8'b11000000; //  449 : 192 - 0xc0
      12'h1C2: dout <= 8'b11110000; //  450 : 240 - 0xf0
      12'h1C3: dout <= 8'b11111000; //  451 : 248 - 0xf8
      12'h1C4: dout <= 8'b10011100; //  452 : 156 - 0x9c
      12'h1C5: dout <= 8'b00001100; //  453 :  12 - 0xc
      12'h1C6: dout <= 8'b00001100; //  454 :  12 - 0xc
      12'h1C7: dout <= 8'b00001110; //  455 :  14 - 0xe
      12'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0 -- plane 1
      12'h1C9: dout <= 8'b11000000; //  457 : 192 - 0xc0
      12'h1CA: dout <= 8'b11110000; //  458 : 240 - 0xf0
      12'h1CB: dout <= 8'b11111000; //  459 : 248 - 0xf8
      12'h1CC: dout <= 8'b11111100; //  460 : 252 - 0xfc
      12'h1CD: dout <= 8'b11111100; //  461 : 252 - 0xfc
      12'h1CE: dout <= 8'b00111100; //  462 :  60 - 0x3c
      12'h1CF: dout <= 8'b00111110; //  463 :  62 - 0x3e
      12'h1D0: dout <= 8'b01100111; //  464 : 103 - 0x67 -- Sprite 0x1d
      12'h1D1: dout <= 8'b01111111; //  465 : 127 - 0x7f
      12'h1D2: dout <= 8'b01111111; //  466 : 127 - 0x7f
      12'h1D3: dout <= 8'b01111111; //  467 : 127 - 0x7f
      12'h1D4: dout <= 8'b01101110; //  468 : 110 - 0x6e
      12'h1D5: dout <= 8'b01000110; //  469 :  70 - 0x46
      12'h1D6: dout <= 8'b00000000; //  470 :   0 - 0x0
      12'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      12'h1D8: dout <= 8'b01111111; //  472 : 127 - 0x7f -- plane 1
      12'h1D9: dout <= 8'b01111111; //  473 : 127 - 0x7f
      12'h1DA: dout <= 8'b01111111; //  474 : 127 - 0x7f
      12'h1DB: dout <= 8'b01111111; //  475 : 127 - 0x7f
      12'h1DC: dout <= 8'b01101110; //  476 : 110 - 0x6e
      12'h1DD: dout <= 8'b01000110; //  477 :  70 - 0x46
      12'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b01100111; //  480 : 103 - 0x67 -- Sprite 0x1e
      12'h1E1: dout <= 8'b01111111; //  481 : 127 - 0x7f
      12'h1E2: dout <= 8'b01111111; //  482 : 127 - 0x7f
      12'h1E3: dout <= 8'b01111111; //  483 : 127 - 0x7f
      12'h1E4: dout <= 8'b01111011; //  484 : 123 - 0x7b
      12'h1E5: dout <= 8'b00110001; //  485 :  49 - 0x31
      12'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      12'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout <= 8'b01111111; //  488 : 127 - 0x7f -- plane 1
      12'h1E9: dout <= 8'b01111111; //  489 : 127 - 0x7f
      12'h1EA: dout <= 8'b01111111; //  490 : 127 - 0x7f
      12'h1EB: dout <= 8'b01111111; //  491 : 127 - 0x7f
      12'h1EC: dout <= 8'b01111011; //  492 : 123 - 0x7b
      12'h1ED: dout <= 8'b00110001; //  493 :  49 - 0x31
      12'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      12'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout <= 8'b10011110; //  496 : 158 - 0x9e -- Sprite 0x1f
      12'h1F1: dout <= 8'b11111110; //  497 : 254 - 0xfe
      12'h1F2: dout <= 8'b11111110; //  498 : 254 - 0xfe
      12'h1F3: dout <= 8'b11111110; //  499 : 254 - 0xfe
      12'h1F4: dout <= 8'b01110110; //  500 : 118 - 0x76
      12'h1F5: dout <= 8'b01100010; //  501 :  98 - 0x62
      12'h1F6: dout <= 8'b00000000; //  502 :   0 - 0x0
      12'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      12'h1F8: dout <= 8'b11111110; //  504 : 254 - 0xfe -- plane 1
      12'h1F9: dout <= 8'b11111110; //  505 : 254 - 0xfe
      12'h1FA: dout <= 8'b11111110; //  506 : 254 - 0xfe
      12'h1FB: dout <= 8'b11111110; //  507 : 254 - 0xfe
      12'h1FC: dout <= 8'b01110110; //  508 : 118 - 0x76
      12'h1FD: dout <= 8'b01100010; //  509 :  98 - 0x62
      12'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout <= 8'b10011110; //  512 : 158 - 0x9e -- Sprite 0x20
      12'h201: dout <= 8'b11111110; //  513 : 254 - 0xfe
      12'h202: dout <= 8'b11111110; //  514 : 254 - 0xfe
      12'h203: dout <= 8'b11111110; //  515 : 254 - 0xfe
      12'h204: dout <= 8'b11011110; //  516 : 222 - 0xde
      12'h205: dout <= 8'b10001100; //  517 : 140 - 0x8c
      12'h206: dout <= 8'b00000000; //  518 :   0 - 0x0
      12'h207: dout <= 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout <= 8'b11111110; //  520 : 254 - 0xfe -- plane 1
      12'h209: dout <= 8'b11111110; //  521 : 254 - 0xfe
      12'h20A: dout <= 8'b11111110; //  522 : 254 - 0xfe
      12'h20B: dout <= 8'b11111110; //  523 : 254 - 0xfe
      12'h20C: dout <= 8'b11011110; //  524 : 222 - 0xde
      12'h20D: dout <= 8'b10001100; //  525 : 140 - 0x8c
      12'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      12'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout <= 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x21
      12'h211: dout <= 8'b00000011; //  529 :   3 - 0x3
      12'h212: dout <= 8'b00001111; //  530 :  15 - 0xf
      12'h213: dout <= 8'b00011111; //  531 :  31 - 0x1f
      12'h214: dout <= 8'b00111111; //  532 :  63 - 0x3f
      12'h215: dout <= 8'b00110011; //  533 :  51 - 0x33
      12'h216: dout <= 8'b00100001; //  534 :  33 - 0x21
      12'h217: dout <= 8'b01100001; //  535 :  97 - 0x61
      12'h218: dout <= 8'b00000000; //  536 :   0 - 0x0 -- plane 1
      12'h219: dout <= 8'b00000011; //  537 :   3 - 0x3
      12'h21A: dout <= 8'b00001111; //  538 :  15 - 0xf
      12'h21B: dout <= 8'b00011111; //  539 :  31 - 0x1f
      12'h21C: dout <= 8'b00111111; //  540 :  63 - 0x3f
      12'h21D: dout <= 8'b00111111; //  541 :  63 - 0x3f
      12'h21E: dout <= 8'b00111111; //  542 :  63 - 0x3f
      12'h21F: dout <= 8'b01111111; //  543 : 127 - 0x7f
      12'h220: dout <= 8'b01100001; //  544 :  97 - 0x61 -- Sprite 0x22
      12'h221: dout <= 8'b01110011; //  545 : 115 - 0x73
      12'h222: dout <= 8'b01111111; //  546 : 127 - 0x7f
      12'h223: dout <= 8'b01111111; //  547 : 127 - 0x7f
      12'h224: dout <= 8'b01101110; //  548 : 110 - 0x6e
      12'h225: dout <= 8'b01000110; //  549 :  70 - 0x46
      12'h226: dout <= 8'b00000000; //  550 :   0 - 0x0
      12'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      12'h228: dout <= 8'b01110011; //  552 : 115 - 0x73 -- plane 1
      12'h229: dout <= 8'b01110011; //  553 : 115 - 0x73
      12'h22A: dout <= 8'b01111111; //  554 : 127 - 0x7f
      12'h22B: dout <= 8'b01111111; //  555 : 127 - 0x7f
      12'h22C: dout <= 8'b01101110; //  556 : 110 - 0x6e
      12'h22D: dout <= 8'b01000110; //  557 :  70 - 0x46
      12'h22E: dout <= 8'b00000000; //  558 :   0 - 0x0
      12'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout <= 8'b01100001; //  560 :  97 - 0x61 -- Sprite 0x23
      12'h231: dout <= 8'b01110011; //  561 : 115 - 0x73
      12'h232: dout <= 8'b01111111; //  562 : 127 - 0x7f
      12'h233: dout <= 8'b01111111; //  563 : 127 - 0x7f
      12'h234: dout <= 8'b01110111; //  564 : 119 - 0x77
      12'h235: dout <= 8'b00100011; //  565 :  35 - 0x23
      12'h236: dout <= 8'b00000000; //  566 :   0 - 0x0
      12'h237: dout <= 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout <= 8'b01110011; //  568 : 115 - 0x73 -- plane 1
      12'h239: dout <= 8'b01110011; //  569 : 115 - 0x73
      12'h23A: dout <= 8'b01111111; //  570 : 127 - 0x7f
      12'h23B: dout <= 8'b01111111; //  571 : 127 - 0x7f
      12'h23C: dout <= 8'b01110111; //  572 : 119 - 0x77
      12'h23D: dout <= 8'b00100011; //  573 :  35 - 0x23
      12'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x24
      12'h241: dout <= 8'b00000011; //  577 :   3 - 0x3
      12'h242: dout <= 8'b00001111; //  578 :  15 - 0xf
      12'h243: dout <= 8'b00011111; //  579 :  31 - 0x1f
      12'h244: dout <= 8'b00111111; //  580 :  63 - 0x3f
      12'h245: dout <= 8'b00111111; //  581 :  63 - 0x3f
      12'h246: dout <= 8'b00111111; //  582 :  63 - 0x3f
      12'h247: dout <= 8'b01111111; //  583 : 127 - 0x7f
      12'h248: dout <= 8'b00000000; //  584 :   0 - 0x0 -- plane 1
      12'h249: dout <= 8'b00000000; //  585 :   0 - 0x0
      12'h24A: dout <= 8'b00000000; //  586 :   0 - 0x0
      12'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      12'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      12'h24D: dout <= 8'b00000110; //  589 :   6 - 0x6
      12'h24E: dout <= 8'b00000110; //  590 :   6 - 0x6
      12'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout <= 8'b01111111; //  592 : 127 - 0x7f -- Sprite 0x25
      12'h251: dout <= 8'b01111111; //  593 : 127 - 0x7f
      12'h252: dout <= 8'b01111111; //  594 : 127 - 0x7f
      12'h253: dout <= 8'b01111111; //  595 : 127 - 0x7f
      12'h254: dout <= 8'b01101110; //  596 : 110 - 0x6e
      12'h255: dout <= 8'b01000110; //  597 :  70 - 0x46
      12'h256: dout <= 8'b00000000; //  598 :   0 - 0x0
      12'h257: dout <= 8'b00000000; //  599 :   0 - 0x0
      12'h258: dout <= 8'b00000000; //  600 :   0 - 0x0 -- plane 1
      12'h259: dout <= 8'b00011001; //  601 :  25 - 0x19
      12'h25A: dout <= 8'b00100110; //  602 :  38 - 0x26
      12'h25B: dout <= 8'b00000000; //  603 :   0 - 0x0
      12'h25C: dout <= 8'b00000000; //  604 :   0 - 0x0
      12'h25D: dout <= 8'b00000000; //  605 :   0 - 0x0
      12'h25E: dout <= 8'b00000000; //  606 :   0 - 0x0
      12'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout <= 8'b01111111; //  608 : 127 - 0x7f -- Sprite 0x26
      12'h261: dout <= 8'b01111111; //  609 : 127 - 0x7f
      12'h262: dout <= 8'b01111111; //  610 : 127 - 0x7f
      12'h263: dout <= 8'b01111111; //  611 : 127 - 0x7f
      12'h264: dout <= 8'b01111011; //  612 : 123 - 0x7b
      12'h265: dout <= 8'b00110001; //  613 :  49 - 0x31
      12'h266: dout <= 8'b00000000; //  614 :   0 - 0x0
      12'h267: dout <= 8'b00000000; //  615 :   0 - 0x0
      12'h268: dout <= 8'b00000000; //  616 :   0 - 0x0 -- plane 1
      12'h269: dout <= 8'b00011001; //  617 :  25 - 0x19
      12'h26A: dout <= 8'b00100110; //  618 :  38 - 0x26
      12'h26B: dout <= 8'b00000000; //  619 :   0 - 0x0
      12'h26C: dout <= 8'b00000000; //  620 :   0 - 0x0
      12'h26D: dout <= 8'b00000000; //  621 :   0 - 0x0
      12'h26E: dout <= 8'b00000000; //  622 :   0 - 0x0
      12'h26F: dout <= 8'b00000000; //  623 :   0 - 0x0
      12'h270: dout <= 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x27
      12'h271: dout <= 8'b00000000; //  625 :   0 - 0x0
      12'h272: dout <= 8'b00000000; //  626 :   0 - 0x0
      12'h273: dout <= 8'b00000000; //  627 :   0 - 0x0
      12'h274: dout <= 8'b00000000; //  628 :   0 - 0x0
      12'h275: dout <= 8'b00000000; //  629 :   0 - 0x0
      12'h276: dout <= 8'b00000000; //  630 :   0 - 0x0
      12'h277: dout <= 8'b00000000; //  631 :   0 - 0x0
      12'h278: dout <= 8'b00000000; //  632 :   0 - 0x0 -- plane 1
      12'h279: dout <= 8'b00001100; //  633 :  12 - 0xc
      12'h27A: dout <= 8'b00010010; //  634 :  18 - 0x12
      12'h27B: dout <= 8'b00010010; //  635 :  18 - 0x12
      12'h27C: dout <= 8'b00011110; //  636 :  30 - 0x1e
      12'h27D: dout <= 8'b00001100; //  637 :  12 - 0xc
      12'h27E: dout <= 8'b00000000; //  638 :   0 - 0x0
      12'h27F: dout <= 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout <= 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x28
      12'h281: dout <= 8'b00000000; //  641 :   0 - 0x0
      12'h282: dout <= 8'b00000000; //  642 :   0 - 0x0
      12'h283: dout <= 8'b00000000; //  643 :   0 - 0x0
      12'h284: dout <= 8'b00000000; //  644 :   0 - 0x0
      12'h285: dout <= 8'b00000000; //  645 :   0 - 0x0
      12'h286: dout <= 8'b00000000; //  646 :   0 - 0x0
      12'h287: dout <= 8'b00000000; //  647 :   0 - 0x0
      12'h288: dout <= 8'b00000000; //  648 :   0 - 0x0 -- plane 1
      12'h289: dout <= 8'b00000000; //  649 :   0 - 0x0
      12'h28A: dout <= 8'b00000000; //  650 :   0 - 0x0
      12'h28B: dout <= 8'b00000000; //  651 :   0 - 0x0
      12'h28C: dout <= 8'b00000000; //  652 :   0 - 0x0
      12'h28D: dout <= 8'b00111000; //  653 :  56 - 0x38
      12'h28E: dout <= 8'b01001101; //  654 :  77 - 0x4d
      12'h28F: dout <= 8'b01001101; //  655 :  77 - 0x4d
      12'h290: dout <= 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x29
      12'h291: dout <= 8'b00000000; //  657 :   0 - 0x0
      12'h292: dout <= 8'b00000000; //  658 :   0 - 0x0
      12'h293: dout <= 8'b00000000; //  659 :   0 - 0x0
      12'h294: dout <= 8'b00000000; //  660 :   0 - 0x0
      12'h295: dout <= 8'b00000000; //  661 :   0 - 0x0
      12'h296: dout <= 8'b00000000; //  662 :   0 - 0x0
      12'h297: dout <= 8'b00000000; //  663 :   0 - 0x0
      12'h298: dout <= 8'b00000000; //  664 :   0 - 0x0 -- plane 1
      12'h299: dout <= 8'b00000000; //  665 :   0 - 0x0
      12'h29A: dout <= 8'b00000000; //  666 :   0 - 0x0
      12'h29B: dout <= 8'b00000000; //  667 :   0 - 0x0
      12'h29C: dout <= 8'b00000000; //  668 :   0 - 0x0
      12'h29D: dout <= 8'b11100000; //  669 : 224 - 0xe0
      12'h29E: dout <= 8'b00110000; //  670 :  48 - 0x30
      12'h29F: dout <= 8'b00110000; //  671 :  48 - 0x30
      12'h2A0: dout <= 8'b00000000; //  672 :   0 - 0x0 -- Sprite 0x2a
      12'h2A1: dout <= 8'b00000000; //  673 :   0 - 0x0
      12'h2A2: dout <= 8'b00000000; //  674 :   0 - 0x0
      12'h2A3: dout <= 8'b00000000; //  675 :   0 - 0x0
      12'h2A4: dout <= 8'b00000000; //  676 :   0 - 0x0
      12'h2A5: dout <= 8'b00000000; //  677 :   0 - 0x0
      12'h2A6: dout <= 8'b00000000; //  678 :   0 - 0x0
      12'h2A7: dout <= 8'b00000000; //  679 :   0 - 0x0
      12'h2A8: dout <= 8'b00111000; //  680 :  56 - 0x38 -- plane 1
      12'h2A9: dout <= 8'b00000000; //  681 :   0 - 0x0
      12'h2AA: dout <= 8'b00000000; //  682 :   0 - 0x0
      12'h2AB: dout <= 8'b00000000; //  683 :   0 - 0x0
      12'h2AC: dout <= 8'b00000000; //  684 :   0 - 0x0
      12'h2AD: dout <= 8'b00000000; //  685 :   0 - 0x0
      12'h2AE: dout <= 8'b00000000; //  686 :   0 - 0x0
      12'h2AF: dout <= 8'b00000000; //  687 :   0 - 0x0
      12'h2B0: dout <= 8'b00000000; //  688 :   0 - 0x0 -- Sprite 0x2b
      12'h2B1: dout <= 8'b00000000; //  689 :   0 - 0x0
      12'h2B2: dout <= 8'b00000000; //  690 :   0 - 0x0
      12'h2B3: dout <= 8'b00000000; //  691 :   0 - 0x0
      12'h2B4: dout <= 8'b00000000; //  692 :   0 - 0x0
      12'h2B5: dout <= 8'b00000000; //  693 :   0 - 0x0
      12'h2B6: dout <= 8'b00000000; //  694 :   0 - 0x0
      12'h2B7: dout <= 8'b00000000; //  695 :   0 - 0x0
      12'h2B8: dout <= 8'b11100000; //  696 : 224 - 0xe0 -- plane 1
      12'h2B9: dout <= 8'b00000000; //  697 :   0 - 0x0
      12'h2BA: dout <= 8'b00000000; //  698 :   0 - 0x0
      12'h2BB: dout <= 8'b00000000; //  699 :   0 - 0x0
      12'h2BC: dout <= 8'b00000000; //  700 :   0 - 0x0
      12'h2BD: dout <= 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout <= 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x2c
      12'h2C1: dout <= 8'b00000000; //  705 :   0 - 0x0
      12'h2C2: dout <= 8'b00000000; //  706 :   0 - 0x0
      12'h2C3: dout <= 8'b00000000; //  707 :   0 - 0x0
      12'h2C4: dout <= 8'b00000000; //  708 :   0 - 0x0
      12'h2C5: dout <= 8'b00000000; //  709 :   0 - 0x0
      12'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      12'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0 -- plane 1
      12'h2C9: dout <= 8'b00000000; //  713 :   0 - 0x0
      12'h2CA: dout <= 8'b00000000; //  714 :   0 - 0x0
      12'h2CB: dout <= 8'b00000000; //  715 :   0 - 0x0
      12'h2CC: dout <= 8'b00000000; //  716 :   0 - 0x0
      12'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      12'h2CE: dout <= 8'b00001100; //  718 :  12 - 0xc
      12'h2CF: dout <= 8'b00011110; //  719 :  30 - 0x1e
      12'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x2d
      12'h2D1: dout <= 8'b00000000; //  721 :   0 - 0x0
      12'h2D2: dout <= 8'b00000000; //  722 :   0 - 0x0
      12'h2D3: dout <= 8'b00000000; //  723 :   0 - 0x0
      12'h2D4: dout <= 8'b00000000; //  724 :   0 - 0x0
      12'h2D5: dout <= 8'b00000000; //  725 :   0 - 0x0
      12'h2D6: dout <= 8'b00000000; //  726 :   0 - 0x0
      12'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      12'h2D8: dout <= 8'b00010010; //  728 :  18 - 0x12 -- plane 1
      12'h2D9: dout <= 8'b00010010; //  729 :  18 - 0x12
      12'h2DA: dout <= 8'b00001100; //  730 :  12 - 0xc
      12'h2DB: dout <= 8'b00000000; //  731 :   0 - 0x0
      12'h2DC: dout <= 8'b00000000; //  732 :   0 - 0x0
      12'h2DD: dout <= 8'b00000000; //  733 :   0 - 0x0
      12'h2DE: dout <= 8'b00000000; //  734 :   0 - 0x0
      12'h2DF: dout <= 8'b00000000; //  735 :   0 - 0x0
      12'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x2e
      12'h2E1: dout <= 8'b00000000; //  737 :   0 - 0x0
      12'h2E2: dout <= 8'b00000000; //  738 :   0 - 0x0
      12'h2E3: dout <= 8'b00000000; //  739 :   0 - 0x0
      12'h2E4: dout <= 8'b00000000; //  740 :   0 - 0x0
      12'h2E5: dout <= 8'b00000000; //  741 :   0 - 0x0
      12'h2E6: dout <= 8'b00000000; //  742 :   0 - 0x0
      12'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0 -- plane 1
      12'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      12'h2EA: dout <= 8'b00000000; //  746 :   0 - 0x0
      12'h2EB: dout <= 8'b00010001; //  747 :  17 - 0x11
      12'h2EC: dout <= 8'b00110010; //  748 :  50 - 0x32
      12'h2ED: dout <= 8'b00010010; //  749 :  18 - 0x12
      12'h2EE: dout <= 8'b00010010; //  750 :  18 - 0x12
      12'h2EF: dout <= 8'b00010010; //  751 :  18 - 0x12
      12'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x2f
      12'h2F1: dout <= 8'b00000000; //  753 :   0 - 0x0
      12'h2F2: dout <= 8'b00000000; //  754 :   0 - 0x0
      12'h2F3: dout <= 8'b00000000; //  755 :   0 - 0x0
      12'h2F4: dout <= 8'b00000000; //  756 :   0 - 0x0
      12'h2F5: dout <= 8'b00000000; //  757 :   0 - 0x0
      12'h2F6: dout <= 8'b00000000; //  758 :   0 - 0x0
      12'h2F7: dout <= 8'b00000000; //  759 :   0 - 0x0
      12'h2F8: dout <= 8'b00000000; //  760 :   0 - 0x0 -- plane 1
      12'h2F9: dout <= 8'b00000000; //  761 :   0 - 0x0
      12'h2FA: dout <= 8'b00000000; //  762 :   0 - 0x0
      12'h2FB: dout <= 8'b10001100; //  763 : 140 - 0x8c
      12'h2FC: dout <= 8'b01010010; //  764 :  82 - 0x52
      12'h2FD: dout <= 8'b01010010; //  765 :  82 - 0x52
      12'h2FE: dout <= 8'b01010010; //  766 :  82 - 0x52
      12'h2FF: dout <= 8'b01010010; //  767 :  82 - 0x52
      12'h300: dout <= 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x30
      12'h301: dout <= 8'b00000000; //  769 :   0 - 0x0
      12'h302: dout <= 8'b00000000; //  770 :   0 - 0x0
      12'h303: dout <= 8'b00000000; //  771 :   0 - 0x0
      12'h304: dout <= 8'b00000000; //  772 :   0 - 0x0
      12'h305: dout <= 8'b00000000; //  773 :   0 - 0x0
      12'h306: dout <= 8'b00000000; //  774 :   0 - 0x0
      12'h307: dout <= 8'b00000000; //  775 :   0 - 0x0
      12'h308: dout <= 8'b00010010; //  776 :  18 - 0x12 -- plane 1
      12'h309: dout <= 8'b00111001; //  777 :  57 - 0x39
      12'h30A: dout <= 8'b00000000; //  778 :   0 - 0x0
      12'h30B: dout <= 8'b00000000; //  779 :   0 - 0x0
      12'h30C: dout <= 8'b00000000; //  780 :   0 - 0x0
      12'h30D: dout <= 8'b00000000; //  781 :   0 - 0x0
      12'h30E: dout <= 8'b00000000; //  782 :   0 - 0x0
      12'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      12'h310: dout <= 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x31
      12'h311: dout <= 8'b00000000; //  785 :   0 - 0x0
      12'h312: dout <= 8'b00000000; //  786 :   0 - 0x0
      12'h313: dout <= 8'b00000000; //  787 :   0 - 0x0
      12'h314: dout <= 8'b00000000; //  788 :   0 - 0x0
      12'h315: dout <= 8'b00000000; //  789 :   0 - 0x0
      12'h316: dout <= 8'b00000000; //  790 :   0 - 0x0
      12'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout <= 8'b01010010; //  792 :  82 - 0x52 -- plane 1
      12'h319: dout <= 8'b10001100; //  793 : 140 - 0x8c
      12'h31A: dout <= 8'b00000000; //  794 :   0 - 0x0
      12'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      12'h31C: dout <= 8'b00000000; //  796 :   0 - 0x0
      12'h31D: dout <= 8'b00000000; //  797 :   0 - 0x0
      12'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      12'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout <= 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x32
      12'h321: dout <= 8'b00000000; //  801 :   0 - 0x0
      12'h322: dout <= 8'b00000000; //  802 :   0 - 0x0
      12'h323: dout <= 8'b00000000; //  803 :   0 - 0x0
      12'h324: dout <= 8'b00000000; //  804 :   0 - 0x0
      12'h325: dout <= 8'b00000000; //  805 :   0 - 0x0
      12'h326: dout <= 8'b00000000; //  806 :   0 - 0x0
      12'h327: dout <= 8'b00000000; //  807 :   0 - 0x0
      12'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- plane 1
      12'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      12'h32B: dout <= 8'b01110001; //  811 : 113 - 0x71
      12'h32C: dout <= 8'b10001010; //  812 : 138 - 0x8a
      12'h32D: dout <= 8'b00001010; //  813 :  10 - 0xa
      12'h32E: dout <= 8'b00010010; //  814 :  18 - 0x12
      12'h32F: dout <= 8'b00100010; //  815 :  34 - 0x22
      12'h330: dout <= 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x33
      12'h331: dout <= 8'b00000000; //  817 :   0 - 0x0
      12'h332: dout <= 8'b00000000; //  818 :   0 - 0x0
      12'h333: dout <= 8'b00000000; //  819 :   0 - 0x0
      12'h334: dout <= 8'b00000000; //  820 :   0 - 0x0
      12'h335: dout <= 8'b00000000; //  821 :   0 - 0x0
      12'h336: dout <= 8'b00000000; //  822 :   0 - 0x0
      12'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      12'h338: dout <= 8'b01000010; //  824 :  66 - 0x42 -- plane 1
      12'h339: dout <= 8'b11111001; //  825 : 249 - 0xf9
      12'h33A: dout <= 8'b00000000; //  826 :   0 - 0x0
      12'h33B: dout <= 8'b00000000; //  827 :   0 - 0x0
      12'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      12'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      12'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x34
      12'h341: dout <= 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout <= 8'b00000000; //  834 :   0 - 0x0
      12'h343: dout <= 8'b00000000; //  835 :   0 - 0x0
      12'h344: dout <= 8'b00000000; //  836 :   0 - 0x0
      12'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      12'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout <= 8'b00000000; //  840 :   0 - 0x0 -- plane 1
      12'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout <= 8'b00000000; //  842 :   0 - 0x0
      12'h34B: dout <= 8'b00110001; //  843 :  49 - 0x31
      12'h34C: dout <= 8'b01001010; //  844 :  74 - 0x4a
      12'h34D: dout <= 8'b00001010; //  845 :  10 - 0xa
      12'h34E: dout <= 8'b00110010; //  846 :  50 - 0x32
      12'h34F: dout <= 8'b00001010; //  847 :  10 - 0xa
      12'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x35
      12'h351: dout <= 8'b00000000; //  849 :   0 - 0x0
      12'h352: dout <= 8'b00000000; //  850 :   0 - 0x0
      12'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      12'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      12'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout <= 8'b01001010; //  856 :  74 - 0x4a -- plane 1
      12'h359: dout <= 8'b00110001; //  857 :  49 - 0x31
      12'h35A: dout <= 8'b00000000; //  858 :   0 - 0x0
      12'h35B: dout <= 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout <= 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x36
      12'h361: dout <= 8'b00000000; //  865 :   0 - 0x0
      12'h362: dout <= 8'b00000000; //  866 :   0 - 0x0
      12'h363: dout <= 8'b00000000; //  867 :   0 - 0x0
      12'h364: dout <= 8'b00000000; //  868 :   0 - 0x0
      12'h365: dout <= 8'b00000000; //  869 :   0 - 0x0
      12'h366: dout <= 8'b00000000; //  870 :   0 - 0x0
      12'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      12'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- plane 1
      12'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout <= 8'b00010001; //  875 :  17 - 0x11
      12'h36C: dout <= 8'b00110010; //  876 :  50 - 0x32
      12'h36D: dout <= 8'b01010010; //  877 :  82 - 0x52
      12'h36E: dout <= 8'b10010010; //  878 : 146 - 0x92
      12'h36F: dout <= 8'b11111010; //  879 : 250 - 0xfa
      12'h370: dout <= 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x37
      12'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout <= 8'b00000000; //  882 :   0 - 0x0
      12'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      12'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      12'h375: dout <= 8'b00000000; //  885 :   0 - 0x0
      12'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout <= 8'b00010010; //  888 :  18 - 0x12 -- plane 1
      12'h379: dout <= 8'b00010001; //  889 :  17 - 0x11
      12'h37A: dout <= 8'b00000000; //  890 :   0 - 0x0
      12'h37B: dout <= 8'b00000000; //  891 :   0 - 0x0
      12'h37C: dout <= 8'b00000000; //  892 :   0 - 0x0
      12'h37D: dout <= 8'b00000000; //  893 :   0 - 0x0
      12'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x38
      12'h381: dout <= 8'b00000000; //  897 :   0 - 0x0
      12'h382: dout <= 8'b00000000; //  898 :   0 - 0x0
      12'h383: dout <= 8'b00000000; //  899 :   0 - 0x0
      12'h384: dout <= 8'b00000000; //  900 :   0 - 0x0
      12'h385: dout <= 8'b00000000; //  901 :   0 - 0x0
      12'h386: dout <= 8'b00000000; //  902 :   0 - 0x0
      12'h387: dout <= 8'b00000000; //  903 :   0 - 0x0
      12'h388: dout <= 8'b00000000; //  904 :   0 - 0x0 -- plane 1
      12'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      12'h38B: dout <= 8'b01110001; //  907 : 113 - 0x71
      12'h38C: dout <= 8'b01000010; //  908 :  66 - 0x42
      12'h38D: dout <= 8'b01000010; //  909 :  66 - 0x42
      12'h38E: dout <= 8'b01110010; //  910 : 114 - 0x72
      12'h38F: dout <= 8'b00001010; //  911 :  10 - 0xa
      12'h390: dout <= 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x39
      12'h391: dout <= 8'b00000000; //  913 :   0 - 0x0
      12'h392: dout <= 8'b00000000; //  914 :   0 - 0x0
      12'h393: dout <= 8'b00000000; //  915 :   0 - 0x0
      12'h394: dout <= 8'b00000000; //  916 :   0 - 0x0
      12'h395: dout <= 8'b00000000; //  917 :   0 - 0x0
      12'h396: dout <= 8'b00000000; //  918 :   0 - 0x0
      12'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout <= 8'b00001010; //  920 :  10 - 0xa -- plane 1
      12'h399: dout <= 8'b01110001; //  921 : 113 - 0x71
      12'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      12'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      12'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      12'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      12'h39E: dout <= 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x3a
      12'h3A1: dout <= 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout <= 8'b00000000; //  930 :   0 - 0x0
      12'h3A3: dout <= 8'b00000000; //  931 :   0 - 0x0
      12'h3A4: dout <= 8'b00000000; //  932 :   0 - 0x0
      12'h3A5: dout <= 8'b00000000; //  933 :   0 - 0x0
      12'h3A6: dout <= 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0 -- plane 1
      12'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout <= 8'b00000000; //  938 :   0 - 0x0
      12'h3AB: dout <= 8'b01110001; //  939 : 113 - 0x71
      12'h3AC: dout <= 8'b00001010; //  940 :  10 - 0xa
      12'h3AD: dout <= 8'b00010010; //  941 :  18 - 0x12
      12'h3AE: dout <= 8'b00010010; //  942 :  18 - 0x12
      12'h3AF: dout <= 8'b00100010; //  943 :  34 - 0x22
      12'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x3b
      12'h3B1: dout <= 8'b00000000; //  945 :   0 - 0x0
      12'h3B2: dout <= 8'b00000000; //  946 :   0 - 0x0
      12'h3B3: dout <= 8'b00000000; //  947 :   0 - 0x0
      12'h3B4: dout <= 8'b00000000; //  948 :   0 - 0x0
      12'h3B5: dout <= 8'b00000000; //  949 :   0 - 0x0
      12'h3B6: dout <= 8'b00000000; //  950 :   0 - 0x0
      12'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout <= 8'b00100010; //  952 :  34 - 0x22 -- plane 1
      12'h3B9: dout <= 8'b00100001; //  953 :  33 - 0x21
      12'h3BA: dout <= 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout <= 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout <= 8'b00000000; //  956 :   0 - 0x0
      12'h3BD: dout <= 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout <= 8'b00000000; //  958 :   0 - 0x0
      12'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x3c
      12'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      12'h3C4: dout <= 8'b00000000; //  964 :   0 - 0x0
      12'h3C5: dout <= 8'b00000000; //  965 :   0 - 0x0
      12'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- plane 1
      12'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout <= 8'b01110001; //  971 : 113 - 0x71
      12'h3CC: dout <= 8'b10001010; //  972 : 138 - 0x8a
      12'h3CD: dout <= 8'b10001010; //  973 : 138 - 0x8a
      12'h3CE: dout <= 8'b01110010; //  974 : 114 - 0x72
      12'h3CF: dout <= 8'b10001010; //  975 : 138 - 0x8a
      12'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x3d
      12'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      12'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      12'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout <= 8'b10001010; //  984 : 138 - 0x8a -- plane 1
      12'h3D9: dout <= 8'b01110001; //  985 : 113 - 0x71
      12'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      12'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x3e
      12'h3E1: dout <= 8'b00000000; //  993 :   0 - 0x0
      12'h3E2: dout <= 8'b00000000; //  994 :   0 - 0x0
      12'h3E3: dout <= 8'b00000000; //  995 :   0 - 0x0
      12'h3E4: dout <= 8'b00000000; //  996 :   0 - 0x0
      12'h3E5: dout <= 8'b00000000; //  997 :   0 - 0x0
      12'h3E6: dout <= 8'b00000000; //  998 :   0 - 0x0
      12'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      12'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0 -- plane 1
      12'h3E9: dout <= 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout <= 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout <= 8'b10011000; // 1003 : 152 - 0x98
      12'h3EC: dout <= 8'b10100101; // 1004 : 165 - 0xa5
      12'h3ED: dout <= 8'b10100101; // 1005 : 165 - 0xa5
      12'h3EE: dout <= 8'b10100101; // 1006 : 165 - 0xa5
      12'h3EF: dout <= 8'b10100101; // 1007 : 165 - 0xa5
      12'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x3f
      12'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout <= 8'b00000000; // 1012 :   0 - 0x0
      12'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0 -- plane 1
      12'h3F9: dout <= 8'b00000000; // 1017 :   0 - 0x0
      12'h3FA: dout <= 8'b00000000; // 1018 :   0 - 0x0
      12'h3FB: dout <= 8'b11000110; // 1019 : 198 - 0xc6
      12'h3FC: dout <= 8'b00101001; // 1020 :  41 - 0x29
      12'h3FD: dout <= 8'b00101001; // 1021 :  41 - 0x29
      12'h3FE: dout <= 8'b00101001; // 1022 :  41 - 0x29
      12'h3FF: dout <= 8'b00101001; // 1023 :  41 - 0x29
      12'h400: dout <= 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x40
      12'h401: dout <= 8'b00000000; // 1025 :   0 - 0x0
      12'h402: dout <= 8'b00000000; // 1026 :   0 - 0x0
      12'h403: dout <= 8'b00000000; // 1027 :   0 - 0x0
      12'h404: dout <= 8'b00000000; // 1028 :   0 - 0x0
      12'h405: dout <= 8'b00000000; // 1029 :   0 - 0x0
      12'h406: dout <= 8'b00000000; // 1030 :   0 - 0x0
      12'h407: dout <= 8'b00000000; // 1031 :   0 - 0x0
      12'h408: dout <= 8'b10100101; // 1032 : 165 - 0xa5 -- plane 1
      12'h409: dout <= 8'b10011000; // 1033 : 152 - 0x98
      12'h40A: dout <= 8'b00000000; // 1034 :   0 - 0x0
      12'h40B: dout <= 8'b00000000; // 1035 :   0 - 0x0
      12'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      12'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      12'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout <= 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x41
      12'h411: dout <= 8'b00000000; // 1041 :   0 - 0x0
      12'h412: dout <= 8'b00000000; // 1042 :   0 - 0x0
      12'h413: dout <= 8'b00000000; // 1043 :   0 - 0x0
      12'h414: dout <= 8'b00000000; // 1044 :   0 - 0x0
      12'h415: dout <= 8'b00000000; // 1045 :   0 - 0x0
      12'h416: dout <= 8'b00000000; // 1046 :   0 - 0x0
      12'h417: dout <= 8'b00000000; // 1047 :   0 - 0x0
      12'h418: dout <= 8'b00101001; // 1048 :  41 - 0x29 -- plane 1
      12'h419: dout <= 8'b11000110; // 1049 : 198 - 0xc6
      12'h41A: dout <= 8'b00000000; // 1050 :   0 - 0x0
      12'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      12'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout <= 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x42
      12'h421: dout <= 8'b00000000; // 1057 :   0 - 0x0
      12'h422: dout <= 8'b00000000; // 1058 :   0 - 0x0
      12'h423: dout <= 8'b00000000; // 1059 :   0 - 0x0
      12'h424: dout <= 8'b00000000; // 1060 :   0 - 0x0
      12'h425: dout <= 8'b00000000; // 1061 :   0 - 0x0
      12'h426: dout <= 8'b00000000; // 1062 :   0 - 0x0
      12'h427: dout <= 8'b00000000; // 1063 :   0 - 0x0
      12'h428: dout <= 8'b00000000; // 1064 :   0 - 0x0 -- plane 1
      12'h429: dout <= 8'b00000000; // 1065 :   0 - 0x0
      12'h42A: dout <= 8'b00000000; // 1066 :   0 - 0x0
      12'h42B: dout <= 8'b10011100; // 1067 : 156 - 0x9c
      12'h42C: dout <= 8'b10100001; // 1068 : 161 - 0xa1
      12'h42D: dout <= 8'b10100001; // 1069 : 161 - 0xa1
      12'h42E: dout <= 8'b10111101; // 1070 : 189 - 0xbd
      12'h42F: dout <= 8'b10100101; // 1071 : 165 - 0xa5
      12'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x43
      12'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      12'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      12'h433: dout <= 8'b00000000; // 1075 :   0 - 0x0
      12'h434: dout <= 8'b00000000; // 1076 :   0 - 0x0
      12'h435: dout <= 8'b00000000; // 1077 :   0 - 0x0
      12'h436: dout <= 8'b00000000; // 1078 :   0 - 0x0
      12'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout <= 8'b10100101; // 1080 : 165 - 0xa5 -- plane 1
      12'h439: dout <= 8'b10011000; // 1081 : 152 - 0x98
      12'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      12'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      12'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      12'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout <= 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x44
      12'h441: dout <= 8'b00000000; // 1089 :   0 - 0x0
      12'h442: dout <= 8'b00000000; // 1090 :   0 - 0x0
      12'h443: dout <= 8'b00000000; // 1091 :   0 - 0x0
      12'h444: dout <= 8'b00000000; // 1092 :   0 - 0x0
      12'h445: dout <= 8'b00000000; // 1093 :   0 - 0x0
      12'h446: dout <= 8'b00000000; // 1094 :   0 - 0x0
      12'h447: dout <= 8'b00000000; // 1095 :   0 - 0x0
      12'h448: dout <= 8'b00000000; // 1096 :   0 - 0x0 -- plane 1
      12'h449: dout <= 8'b00000000; // 1097 :   0 - 0x0
      12'h44A: dout <= 8'b00000000; // 1098 :   0 - 0x0
      12'h44B: dout <= 8'b01100010; // 1099 :  98 - 0x62
      12'h44C: dout <= 8'b10010101; // 1100 : 149 - 0x95
      12'h44D: dout <= 8'b00010101; // 1101 :  21 - 0x15
      12'h44E: dout <= 8'b00100101; // 1102 :  37 - 0x25
      12'h44F: dout <= 8'b01000101; // 1103 :  69 - 0x45
      12'h450: dout <= 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x45
      12'h451: dout <= 8'b00000000; // 1105 :   0 - 0x0
      12'h452: dout <= 8'b00000000; // 1106 :   0 - 0x0
      12'h453: dout <= 8'b00000000; // 1107 :   0 - 0x0
      12'h454: dout <= 8'b00000000; // 1108 :   0 - 0x0
      12'h455: dout <= 8'b00000000; // 1109 :   0 - 0x0
      12'h456: dout <= 8'b00000000; // 1110 :   0 - 0x0
      12'h457: dout <= 8'b00000000; // 1111 :   0 - 0x0
      12'h458: dout <= 8'b00000000; // 1112 :   0 - 0x0 -- plane 1
      12'h459: dout <= 8'b00000000; // 1113 :   0 - 0x0
      12'h45A: dout <= 8'b00000000; // 1114 :   0 - 0x0
      12'h45B: dout <= 8'b00100010; // 1115 :  34 - 0x22
      12'h45C: dout <= 8'b01010101; // 1116 :  85 - 0x55
      12'h45D: dout <= 8'b01010101; // 1117 :  85 - 0x55
      12'h45E: dout <= 8'b01010101; // 1118 :  85 - 0x55
      12'h45F: dout <= 8'b01010101; // 1119 :  85 - 0x55
      12'h460: dout <= 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x46
      12'h461: dout <= 8'b00000000; // 1121 :   0 - 0x0
      12'h462: dout <= 8'b00000000; // 1122 :   0 - 0x0
      12'h463: dout <= 8'b00000000; // 1123 :   0 - 0x0
      12'h464: dout <= 8'b00000000; // 1124 :   0 - 0x0
      12'h465: dout <= 8'b00000000; // 1125 :   0 - 0x0
      12'h466: dout <= 8'b00000000; // 1126 :   0 - 0x0
      12'h467: dout <= 8'b00000000; // 1127 :   0 - 0x0
      12'h468: dout <= 8'b10000101; // 1128 : 133 - 0x85 -- plane 1
      12'h469: dout <= 8'b11110010; // 1129 : 242 - 0xf2
      12'h46A: dout <= 8'b00000000; // 1130 :   0 - 0x0
      12'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      12'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      12'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      12'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      12'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      12'h470: dout <= 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x47
      12'h471: dout <= 8'b00000000; // 1137 :   0 - 0x0
      12'h472: dout <= 8'b00000000; // 1138 :   0 - 0x0
      12'h473: dout <= 8'b00000000; // 1139 :   0 - 0x0
      12'h474: dout <= 8'b00000000; // 1140 :   0 - 0x0
      12'h475: dout <= 8'b00000000; // 1141 :   0 - 0x0
      12'h476: dout <= 8'b00000000; // 1142 :   0 - 0x0
      12'h477: dout <= 8'b00000000; // 1143 :   0 - 0x0
      12'h478: dout <= 8'b01010101; // 1144 :  85 - 0x55 -- plane 1
      12'h479: dout <= 8'b00100010; // 1145 :  34 - 0x22
      12'h47A: dout <= 8'b00000000; // 1146 :   0 - 0x0
      12'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      12'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      12'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      12'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      12'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x48
      12'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      12'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      12'h483: dout <= 8'b00000000; // 1155 :   0 - 0x0
      12'h484: dout <= 8'b00000000; // 1156 :   0 - 0x0
      12'h485: dout <= 8'b00000000; // 1157 :   0 - 0x0
      12'h486: dout <= 8'b00000000; // 1158 :   0 - 0x0
      12'h487: dout <= 8'b00000000; // 1159 :   0 - 0x0
      12'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0 -- plane 1
      12'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      12'h48A: dout <= 8'b00000000; // 1162 :   0 - 0x0
      12'h48B: dout <= 8'b01100010; // 1163 :  98 - 0x62
      12'h48C: dout <= 8'b10010101; // 1164 : 149 - 0x95
      12'h48D: dout <= 8'b00010101; // 1165 :  21 - 0x15
      12'h48E: dout <= 8'b01100101; // 1166 : 101 - 0x65
      12'h48F: dout <= 8'b00010101; // 1167 :  21 - 0x15
      12'h490: dout <= 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x49
      12'h491: dout <= 8'b00000000; // 1169 :   0 - 0x0
      12'h492: dout <= 8'b00000000; // 1170 :   0 - 0x0
      12'h493: dout <= 8'b00000000; // 1171 :   0 - 0x0
      12'h494: dout <= 8'b00000000; // 1172 :   0 - 0x0
      12'h495: dout <= 8'b00000000; // 1173 :   0 - 0x0
      12'h496: dout <= 8'b00000000; // 1174 :   0 - 0x0
      12'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      12'h498: dout <= 8'b10010101; // 1176 : 149 - 0x95 -- plane 1
      12'h499: dout <= 8'b01100010; // 1177 :  98 - 0x62
      12'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      12'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      12'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      12'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      12'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      12'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      12'h4A0: dout <= 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x4a
      12'h4A1: dout <= 8'b00000000; // 1185 :   0 - 0x0
      12'h4A2: dout <= 8'b00000000; // 1186 :   0 - 0x0
      12'h4A3: dout <= 8'b00000000; // 1187 :   0 - 0x0
      12'h4A4: dout <= 8'b00000000; // 1188 :   0 - 0x0
      12'h4A5: dout <= 8'b00000000; // 1189 :   0 - 0x0
      12'h4A6: dout <= 8'b00000000; // 1190 :   0 - 0x0
      12'h4A7: dout <= 8'b00000000; // 1191 :   0 - 0x0
      12'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0 -- plane 1
      12'h4A9: dout <= 8'b00000000; // 1193 :   0 - 0x0
      12'h4AA: dout <= 8'b00000000; // 1194 :   0 - 0x0
      12'h4AB: dout <= 8'b11100010; // 1195 : 226 - 0xe2
      12'h4AC: dout <= 8'b10000101; // 1196 : 133 - 0x85
      12'h4AD: dout <= 8'b10000101; // 1197 : 133 - 0x85
      12'h4AE: dout <= 8'b11100101; // 1198 : 229 - 0xe5
      12'h4AF: dout <= 8'b00010101; // 1199 :  21 - 0x15
      12'h4B0: dout <= 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x4b
      12'h4B1: dout <= 8'b00000000; // 1201 :   0 - 0x0
      12'h4B2: dout <= 8'b00000000; // 1202 :   0 - 0x0
      12'h4B3: dout <= 8'b00000000; // 1203 :   0 - 0x0
      12'h4B4: dout <= 8'b00000000; // 1204 :   0 - 0x0
      12'h4B5: dout <= 8'b00000000; // 1205 :   0 - 0x0
      12'h4B6: dout <= 8'b00000000; // 1206 :   0 - 0x0
      12'h4B7: dout <= 8'b00000000; // 1207 :   0 - 0x0
      12'h4B8: dout <= 8'b00010101; // 1208 :  21 - 0x15 -- plane 1
      12'h4B9: dout <= 8'b11100010; // 1209 : 226 - 0xe2
      12'h4BA: dout <= 8'b00000000; // 1210 :   0 - 0x0
      12'h4BB: dout <= 8'b00000000; // 1211 :   0 - 0x0
      12'h4BC: dout <= 8'b00000000; // 1212 :   0 - 0x0
      12'h4BD: dout <= 8'b00000000; // 1213 :   0 - 0x0
      12'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      12'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      12'h4C0: dout <= 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x4c
      12'h4C1: dout <= 8'b00000000; // 1217 :   0 - 0x0
      12'h4C2: dout <= 8'b00000000; // 1218 :   0 - 0x0
      12'h4C3: dout <= 8'b00000000; // 1219 :   0 - 0x0
      12'h4C4: dout <= 8'b00000000; // 1220 :   0 - 0x0
      12'h4C5: dout <= 8'b00000000; // 1221 :   0 - 0x0
      12'h4C6: dout <= 8'b00000000; // 1222 :   0 - 0x0
      12'h4C7: dout <= 8'b00000000; // 1223 :   0 - 0x0
      12'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0 -- plane 1
      12'h4C9: dout <= 8'b00000000; // 1225 :   0 - 0x0
      12'h4CA: dout <= 8'b00000000; // 1226 :   0 - 0x0
      12'h4CB: dout <= 8'b00000000; // 1227 :   0 - 0x0
      12'h4CC: dout <= 8'b00000000; // 1228 :   0 - 0x0
      12'h4CD: dout <= 8'b00000000; // 1229 :   0 - 0x0
      12'h4CE: dout <= 8'b00000000; // 1230 :   0 - 0x0
      12'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      12'h4D0: dout <= 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x4d
      12'h4D1: dout <= 8'b00000000; // 1233 :   0 - 0x0
      12'h4D2: dout <= 8'b00000000; // 1234 :   0 - 0x0
      12'h4D3: dout <= 8'b00000001; // 1235 :   1 - 0x1
      12'h4D4: dout <= 8'b00000011; // 1236 :   3 - 0x3
      12'h4D5: dout <= 8'b00000111; // 1237 :   7 - 0x7
      12'h4D6: dout <= 8'b00001111; // 1238 :  15 - 0xf
      12'h4D7: dout <= 8'b00011111; // 1239 :  31 - 0x1f
      12'h4D8: dout <= 8'b00000000; // 1240 :   0 - 0x0 -- plane 1
      12'h4D9: dout <= 8'b00000000; // 1241 :   0 - 0x0
      12'h4DA: dout <= 8'b00000000; // 1242 :   0 - 0x0
      12'h4DB: dout <= 8'b00000000; // 1243 :   0 - 0x0
      12'h4DC: dout <= 8'b00000000; // 1244 :   0 - 0x0
      12'h4DD: dout <= 8'b00000000; // 1245 :   0 - 0x0
      12'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      12'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout <= 8'b00000000; // 1248 :   0 - 0x0 -- Sprite 0x4e
      12'h4E1: dout <= 8'b00001111; // 1249 :  15 - 0xf
      12'h4E2: dout <= 8'b01111111; // 1250 : 127 - 0x7f
      12'h4E3: dout <= 8'b11111111; // 1251 : 255 - 0xff
      12'h4E4: dout <= 8'b11111111; // 1252 : 255 - 0xff
      12'h4E5: dout <= 8'b11111111; // 1253 : 255 - 0xff
      12'h4E6: dout <= 8'b11111111; // 1254 : 255 - 0xff
      12'h4E7: dout <= 8'b11111111; // 1255 : 255 - 0xff
      12'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0 -- plane 1
      12'h4E9: dout <= 8'b00000000; // 1257 :   0 - 0x0
      12'h4EA: dout <= 8'b00000000; // 1258 :   0 - 0x0
      12'h4EB: dout <= 8'b00000000; // 1259 :   0 - 0x0
      12'h4EC: dout <= 8'b00000000; // 1260 :   0 - 0x0
      12'h4ED: dout <= 8'b00000000; // 1261 :   0 - 0x0
      12'h4EE: dout <= 8'b00000000; // 1262 :   0 - 0x0
      12'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout <= 8'b00011111; // 1264 :  31 - 0x1f -- Sprite 0x4f
      12'h4F1: dout <= 8'b00111111; // 1265 :  63 - 0x3f
      12'h4F2: dout <= 8'b00111111; // 1266 :  63 - 0x3f
      12'h4F3: dout <= 8'b00111111; // 1267 :  63 - 0x3f
      12'h4F4: dout <= 8'b01111111; // 1268 : 127 - 0x7f
      12'h4F5: dout <= 8'b01111111; // 1269 : 127 - 0x7f
      12'h4F6: dout <= 8'b01111111; // 1270 : 127 - 0x7f
      12'h4F7: dout <= 8'b01111111; // 1271 : 127 - 0x7f
      12'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0 -- plane 1
      12'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      12'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      12'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      12'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      12'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout <= 8'b11111111; // 1280 : 255 - 0xff -- Sprite 0x50
      12'h501: dout <= 8'b11111111; // 1281 : 255 - 0xff
      12'h502: dout <= 8'b11111111; // 1282 : 255 - 0xff
      12'h503: dout <= 8'b11111111; // 1283 : 255 - 0xff
      12'h504: dout <= 8'b11111111; // 1284 : 255 - 0xff
      12'h505: dout <= 8'b11111111; // 1285 : 255 - 0xff
      12'h506: dout <= 8'b11111111; // 1286 : 255 - 0xff
      12'h507: dout <= 8'b11111111; // 1287 : 255 - 0xff
      12'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0 -- plane 1
      12'h509: dout <= 8'b00000000; // 1289 :   0 - 0x0
      12'h50A: dout <= 8'b00000000; // 1290 :   0 - 0x0
      12'h50B: dout <= 8'b00000000; // 1291 :   0 - 0x0
      12'h50C: dout <= 8'b00000000; // 1292 :   0 - 0x0
      12'h50D: dout <= 8'b00000000; // 1293 :   0 - 0x0
      12'h50E: dout <= 8'b00000000; // 1294 :   0 - 0x0
      12'h50F: dout <= 8'b00000000; // 1295 :   0 - 0x0
      12'h510: dout <= 8'b11111111; // 1296 : 255 - 0xff -- Sprite 0x51
      12'h511: dout <= 8'b11111111; // 1297 : 255 - 0xff
      12'h512: dout <= 8'b11111111; // 1298 : 255 - 0xff
      12'h513: dout <= 8'b11111111; // 1299 : 255 - 0xff
      12'h514: dout <= 8'b11111111; // 1300 : 255 - 0xff
      12'h515: dout <= 8'b11111111; // 1301 : 255 - 0xff
      12'h516: dout <= 8'b11111111; // 1302 : 255 - 0xff
      12'h517: dout <= 8'b11111110; // 1303 : 254 - 0xfe
      12'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0 -- plane 1
      12'h519: dout <= 8'b00000000; // 1305 :   0 - 0x0
      12'h51A: dout <= 8'b00000000; // 1306 :   0 - 0x0
      12'h51B: dout <= 8'b00000000; // 1307 :   0 - 0x0
      12'h51C: dout <= 8'b00000000; // 1308 :   0 - 0x0
      12'h51D: dout <= 8'b00000000; // 1309 :   0 - 0x0
      12'h51E: dout <= 8'b00000000; // 1310 :   0 - 0x0
      12'h51F: dout <= 8'b00000000; // 1311 :   0 - 0x0
      12'h520: dout <= 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0x52
      12'h521: dout <= 8'b00000000; // 1313 :   0 - 0x0
      12'h522: dout <= 8'b00000000; // 1314 :   0 - 0x0
      12'h523: dout <= 8'b10000000; // 1315 : 128 - 0x80
      12'h524: dout <= 8'b11000000; // 1316 : 192 - 0xc0
      12'h525: dout <= 8'b11100000; // 1317 : 224 - 0xe0
      12'h526: dout <= 8'b11110000; // 1318 : 240 - 0xf0
      12'h527: dout <= 8'b11110000; // 1319 : 240 - 0xf0
      12'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0 -- plane 1
      12'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      12'h52A: dout <= 8'b00000000; // 1322 :   0 - 0x0
      12'h52B: dout <= 8'b00000000; // 1323 :   0 - 0x0
      12'h52C: dout <= 8'b00000000; // 1324 :   0 - 0x0
      12'h52D: dout <= 8'b00000000; // 1325 :   0 - 0x0
      12'h52E: dout <= 8'b00000000; // 1326 :   0 - 0x0
      12'h52F: dout <= 8'b00000000; // 1327 :   0 - 0x0
      12'h530: dout <= 8'b11111111; // 1328 : 255 - 0xff -- Sprite 0x53
      12'h531: dout <= 8'b11111111; // 1329 : 255 - 0xff
      12'h532: dout <= 8'b11111110; // 1330 : 254 - 0xfe
      12'h533: dout <= 8'b11111100; // 1331 : 252 - 0xfc
      12'h534: dout <= 8'b11110000; // 1332 : 240 - 0xf0
      12'h535: dout <= 8'b11100000; // 1333 : 224 - 0xe0
      12'h536: dout <= 8'b10000000; // 1334 : 128 - 0x80
      12'h537: dout <= 8'b00000000; // 1335 :   0 - 0x0
      12'h538: dout <= 8'b00000000; // 1336 :   0 - 0x0 -- plane 1
      12'h539: dout <= 8'b00000000; // 1337 :   0 - 0x0
      12'h53A: dout <= 8'b00000000; // 1338 :   0 - 0x0
      12'h53B: dout <= 8'b00000000; // 1339 :   0 - 0x0
      12'h53C: dout <= 8'b00000000; // 1340 :   0 - 0x0
      12'h53D: dout <= 8'b00000000; // 1341 :   0 - 0x0
      12'h53E: dout <= 8'b00000000; // 1342 :   0 - 0x0
      12'h53F: dout <= 8'b00000000; // 1343 :   0 - 0x0
      12'h540: dout <= 8'b11000000; // 1344 : 192 - 0xc0 -- Sprite 0x54
      12'h541: dout <= 8'b10000000; // 1345 : 128 - 0x80
      12'h542: dout <= 8'b00000000; // 1346 :   0 - 0x0
      12'h543: dout <= 8'b00000000; // 1347 :   0 - 0x0
      12'h544: dout <= 8'b00000000; // 1348 :   0 - 0x0
      12'h545: dout <= 8'b00000000; // 1349 :   0 - 0x0
      12'h546: dout <= 8'b00000000; // 1350 :   0 - 0x0
      12'h547: dout <= 8'b00000000; // 1351 :   0 - 0x0
      12'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0 -- plane 1
      12'h549: dout <= 8'b00000000; // 1353 :   0 - 0x0
      12'h54A: dout <= 8'b00000000; // 1354 :   0 - 0x0
      12'h54B: dout <= 8'b00000000; // 1355 :   0 - 0x0
      12'h54C: dout <= 8'b00000000; // 1356 :   0 - 0x0
      12'h54D: dout <= 8'b00000000; // 1357 :   0 - 0x0
      12'h54E: dout <= 8'b00000000; // 1358 :   0 - 0x0
      12'h54F: dout <= 8'b00000000; // 1359 :   0 - 0x0
      12'h550: dout <= 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0x55
      12'h551: dout <= 8'b11110000; // 1361 : 240 - 0xf0
      12'h552: dout <= 8'b11111110; // 1362 : 254 - 0xfe
      12'h553: dout <= 8'b11111110; // 1363 : 254 - 0xfe
      12'h554: dout <= 8'b11111110; // 1364 : 254 - 0xfe
      12'h555: dout <= 8'b11111100; // 1365 : 252 - 0xfc
      12'h556: dout <= 8'b11111000; // 1366 : 248 - 0xf8
      12'h557: dout <= 8'b11111000; // 1367 : 248 - 0xf8
      12'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0 -- plane 1
      12'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      12'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      12'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      12'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      12'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      12'h560: dout <= 8'b11110000; // 1376 : 240 - 0xf0 -- Sprite 0x56
      12'h561: dout <= 8'b11100000; // 1377 : 224 - 0xe0
      12'h562: dout <= 8'b11100000; // 1378 : 224 - 0xe0
      12'h563: dout <= 8'b11000000; // 1379 : 192 - 0xc0
      12'h564: dout <= 8'b10000000; // 1380 : 128 - 0x80
      12'h565: dout <= 8'b10000000; // 1381 : 128 - 0x80
      12'h566: dout <= 8'b00000000; // 1382 :   0 - 0x0
      12'h567: dout <= 8'b00000000; // 1383 :   0 - 0x0
      12'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0 -- plane 1
      12'h569: dout <= 8'b00000000; // 1385 :   0 - 0x0
      12'h56A: dout <= 8'b00000000; // 1386 :   0 - 0x0
      12'h56B: dout <= 8'b00000000; // 1387 :   0 - 0x0
      12'h56C: dout <= 8'b00000000; // 1388 :   0 - 0x0
      12'h56D: dout <= 8'b00000000; // 1389 :   0 - 0x0
      12'h56E: dout <= 8'b00000000; // 1390 :   0 - 0x0
      12'h56F: dout <= 8'b00000000; // 1391 :   0 - 0x0
      12'h570: dout <= 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0x57
      12'h571: dout <= 8'b00000000; // 1393 :   0 - 0x0
      12'h572: dout <= 8'b00000000; // 1394 :   0 - 0x0
      12'h573: dout <= 8'b00000000; // 1395 :   0 - 0x0
      12'h574: dout <= 8'b00000000; // 1396 :   0 - 0x0
      12'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      12'h576: dout <= 8'b00000000; // 1398 :   0 - 0x0
      12'h577: dout <= 8'b00000100; // 1399 :   4 - 0x4
      12'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0 -- plane 1
      12'h579: dout <= 8'b00000000; // 1401 :   0 - 0x0
      12'h57A: dout <= 8'b00000000; // 1402 :   0 - 0x0
      12'h57B: dout <= 8'b00000000; // 1403 :   0 - 0x0
      12'h57C: dout <= 8'b00000000; // 1404 :   0 - 0x0
      12'h57D: dout <= 8'b00000000; // 1405 :   0 - 0x0
      12'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      12'h57F: dout <= 8'b00000100; // 1407 :   4 - 0x4
      12'h580: dout <= 8'b00000110; // 1408 :   6 - 0x6 -- Sprite 0x58
      12'h581: dout <= 8'b00000110; // 1409 :   6 - 0x6
      12'h582: dout <= 8'b00000111; // 1410 :   7 - 0x7
      12'h583: dout <= 8'b00000111; // 1411 :   7 - 0x7
      12'h584: dout <= 8'b00000111; // 1412 :   7 - 0x7
      12'h585: dout <= 8'b00000111; // 1413 :   7 - 0x7
      12'h586: dout <= 8'b00000000; // 1414 :   0 - 0x0
      12'h587: dout <= 8'b00000000; // 1415 :   0 - 0x0
      12'h588: dout <= 8'b00000110; // 1416 :   6 - 0x6 -- plane 1
      12'h589: dout <= 8'b00000110; // 1417 :   6 - 0x6
      12'h58A: dout <= 8'b00000111; // 1418 :   7 - 0x7
      12'h58B: dout <= 8'b00000111; // 1419 :   7 - 0x7
      12'h58C: dout <= 8'b00000111; // 1420 :   7 - 0x7
      12'h58D: dout <= 8'b00000111; // 1421 :   7 - 0x7
      12'h58E: dout <= 8'b00000000; // 1422 :   0 - 0x0
      12'h58F: dout <= 8'b00000000; // 1423 :   0 - 0x0
      12'h590: dout <= 8'b00000000; // 1424 :   0 - 0x0 -- Sprite 0x59
      12'h591: dout <= 8'b00000000; // 1425 :   0 - 0x0
      12'h592: dout <= 8'b00000000; // 1426 :   0 - 0x0
      12'h593: dout <= 8'b00000000; // 1427 :   0 - 0x0
      12'h594: dout <= 8'b00000000; // 1428 :   0 - 0x0
      12'h595: dout <= 8'b00000000; // 1429 :   0 - 0x0
      12'h596: dout <= 8'b00000000; // 1430 :   0 - 0x0
      12'h597: dout <= 8'b00010000; // 1431 :  16 - 0x10
      12'h598: dout <= 8'b00000000; // 1432 :   0 - 0x0 -- plane 1
      12'h599: dout <= 8'b00000000; // 1433 :   0 - 0x0
      12'h59A: dout <= 8'b00000000; // 1434 :   0 - 0x0
      12'h59B: dout <= 8'b00000000; // 1435 :   0 - 0x0
      12'h59C: dout <= 8'b00000000; // 1436 :   0 - 0x0
      12'h59D: dout <= 8'b00000000; // 1437 :   0 - 0x0
      12'h59E: dout <= 8'b00000000; // 1438 :   0 - 0x0
      12'h59F: dout <= 8'b00010000; // 1439 :  16 - 0x10
      12'h5A0: dout <= 8'b00011100; // 1440 :  28 - 0x1c -- Sprite 0x5a
      12'h5A1: dout <= 8'b00011110; // 1441 :  30 - 0x1e
      12'h5A2: dout <= 8'b00011111; // 1442 :  31 - 0x1f
      12'h5A3: dout <= 8'b00011111; // 1443 :  31 - 0x1f
      12'h5A4: dout <= 8'b00011111; // 1444 :  31 - 0x1f
      12'h5A5: dout <= 8'b00011111; // 1445 :  31 - 0x1f
      12'h5A6: dout <= 8'b00000000; // 1446 :   0 - 0x0
      12'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      12'h5A8: dout <= 8'b00011100; // 1448 :  28 - 0x1c -- plane 1
      12'h5A9: dout <= 8'b00011110; // 1449 :  30 - 0x1e
      12'h5AA: dout <= 8'b00011111; // 1450 :  31 - 0x1f
      12'h5AB: dout <= 8'b00011111; // 1451 :  31 - 0x1f
      12'h5AC: dout <= 8'b00011111; // 1452 :  31 - 0x1f
      12'h5AD: dout <= 8'b00011111; // 1453 :  31 - 0x1f
      12'h5AE: dout <= 8'b00000000; // 1454 :   0 - 0x0
      12'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      12'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0x5b
      12'h5B1: dout <= 8'b00000000; // 1457 :   0 - 0x0
      12'h5B2: dout <= 8'b00000000; // 1458 :   0 - 0x0
      12'h5B3: dout <= 8'b00000000; // 1459 :   0 - 0x0
      12'h5B4: dout <= 8'b00000000; // 1460 :   0 - 0x0
      12'h5B5: dout <= 8'b00000000; // 1461 :   0 - 0x0
      12'h5B6: dout <= 8'b00000000; // 1462 :   0 - 0x0
      12'h5B7: dout <= 8'b11000000; // 1463 : 192 - 0xc0
      12'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0 -- plane 1
      12'h5B9: dout <= 8'b00000000; // 1465 :   0 - 0x0
      12'h5BA: dout <= 8'b00000000; // 1466 :   0 - 0x0
      12'h5BB: dout <= 8'b00000000; // 1467 :   0 - 0x0
      12'h5BC: dout <= 8'b00000000; // 1468 :   0 - 0x0
      12'h5BD: dout <= 8'b00000000; // 1469 :   0 - 0x0
      12'h5BE: dout <= 8'b00000000; // 1470 :   0 - 0x0
      12'h5BF: dout <= 8'b11000000; // 1471 : 192 - 0xc0
      12'h5C0: dout <= 8'b11110000; // 1472 : 240 - 0xf0 -- Sprite 0x5c
      12'h5C1: dout <= 8'b11111100; // 1473 : 252 - 0xfc
      12'h5C2: dout <= 8'b11111111; // 1474 : 255 - 0xff
      12'h5C3: dout <= 8'b11111111; // 1475 : 255 - 0xff
      12'h5C4: dout <= 8'b11111111; // 1476 : 255 - 0xff
      12'h5C5: dout <= 8'b11111111; // 1477 : 255 - 0xff
      12'h5C6: dout <= 8'b00000000; // 1478 :   0 - 0x0
      12'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout <= 8'b11110000; // 1480 : 240 - 0xf0 -- plane 1
      12'h5C9: dout <= 8'b11111100; // 1481 : 252 - 0xfc
      12'h5CA: dout <= 8'b11111111; // 1482 : 255 - 0xff
      12'h5CB: dout <= 8'b11111111; // 1483 : 255 - 0xff
      12'h5CC: dout <= 8'b11111111; // 1484 : 255 - 0xff
      12'h5CD: dout <= 8'b11111111; // 1485 : 255 - 0xff
      12'h5CE: dout <= 8'b00000000; // 1486 :   0 - 0x0
      12'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout <= 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0x5d
      12'h5D1: dout <= 8'b00000000; // 1489 :   0 - 0x0
      12'h5D2: dout <= 8'b00000001; // 1490 :   1 - 0x1
      12'h5D3: dout <= 8'b00000011; // 1491 :   3 - 0x3
      12'h5D4: dout <= 8'b00001111; // 1492 :  15 - 0xf
      12'h5D5: dout <= 8'b00001111; // 1493 :  15 - 0xf
      12'h5D6: dout <= 8'b00000000; // 1494 :   0 - 0x0
      12'h5D7: dout <= 8'b00000000; // 1495 :   0 - 0x0
      12'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0 -- plane 1
      12'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout <= 8'b00000001; // 1498 :   1 - 0x1
      12'h5DB: dout <= 8'b00000011; // 1499 :   3 - 0x3
      12'h5DC: dout <= 8'b00001111; // 1500 :  15 - 0xf
      12'h5DD: dout <= 8'b00001111; // 1501 :  15 - 0xf
      12'h5DE: dout <= 8'b00000000; // 1502 :   0 - 0x0
      12'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout <= 8'b11111100; // 1504 : 252 - 0xfc -- Sprite 0x5e
      12'h5E1: dout <= 8'b11111100; // 1505 : 252 - 0xfc
      12'h5E2: dout <= 8'b11111100; // 1506 : 252 - 0xfc
      12'h5E3: dout <= 8'b11111100; // 1507 : 252 - 0xfc
      12'h5E4: dout <= 8'b11111000; // 1508 : 248 - 0xf8
      12'h5E5: dout <= 8'b11111100; // 1509 : 252 - 0xfc
      12'h5E6: dout <= 8'b00111100; // 1510 :  60 - 0x3c
      12'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout <= 8'b11111000; // 1512 : 248 - 0xf8 -- plane 1
      12'h5E9: dout <= 8'b11110000; // 1513 : 240 - 0xf0
      12'h5EA: dout <= 8'b11100000; // 1514 : 224 - 0xe0
      12'h5EB: dout <= 8'b11110000; // 1515 : 240 - 0xf0
      12'h5EC: dout <= 8'b11100000; // 1516 : 224 - 0xe0
      12'h5ED: dout <= 8'b11000000; // 1517 : 192 - 0xc0
      12'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      12'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout <= 8'b00000100; // 1520 :   4 - 0x4 -- Sprite 0x5f
      12'h5F1: dout <= 8'b00001100; // 1521 :  12 - 0xc
      12'h5F2: dout <= 8'b00011100; // 1522 :  28 - 0x1c
      12'h5F3: dout <= 8'b00001100; // 1523 :  12 - 0xc
      12'h5F4: dout <= 8'b00011000; // 1524 :  24 - 0x18
      12'h5F5: dout <= 8'b00111100; // 1525 :  60 - 0x3c
      12'h5F6: dout <= 8'b00111100; // 1526 :  60 - 0x3c
      12'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      12'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- plane 1
      12'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      12'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      12'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      12'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      12'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      12'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0x60
      12'h601: dout <= 8'b00000011; // 1537 :   3 - 0x3
      12'h602: dout <= 8'b00001111; // 1538 :  15 - 0xf
      12'h603: dout <= 8'b00010011; // 1539 :  19 - 0x13
      12'h604: dout <= 8'b00100001; // 1540 :  33 - 0x21
      12'h605: dout <= 8'b00100001; // 1541 :  33 - 0x21
      12'h606: dout <= 8'b00100001; // 1542 :  33 - 0x21
      12'h607: dout <= 8'b01110011; // 1543 : 115 - 0x73
      12'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0 -- plane 1
      12'h609: dout <= 8'b00000011; // 1545 :   3 - 0x3
      12'h60A: dout <= 8'b00001111; // 1546 :  15 - 0xf
      12'h60B: dout <= 8'b00011111; // 1547 :  31 - 0x1f
      12'h60C: dout <= 8'b00111111; // 1548 :  63 - 0x3f
      12'h60D: dout <= 8'b00111111; // 1549 :  63 - 0x3f
      12'h60E: dout <= 8'b00111001; // 1550 :  57 - 0x39
      12'h60F: dout <= 8'b01111011; // 1551 : 123 - 0x7b
      12'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0x61
      12'h611: dout <= 8'b11000000; // 1553 : 192 - 0xc0
      12'h612: dout <= 8'b11110000; // 1554 : 240 - 0xf0
      12'h613: dout <= 8'b11001000; // 1555 : 200 - 0xc8
      12'h614: dout <= 8'b10000100; // 1556 : 132 - 0x84
      12'h615: dout <= 8'b10000100; // 1557 : 132 - 0x84
      12'h616: dout <= 8'b10000100; // 1558 : 132 - 0x84
      12'h617: dout <= 8'b11001110; // 1559 : 206 - 0xce
      12'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0 -- plane 1
      12'h619: dout <= 8'b11000000; // 1561 : 192 - 0xc0
      12'h61A: dout <= 8'b11110000; // 1562 : 240 - 0xf0
      12'h61B: dout <= 8'b11111000; // 1563 : 248 - 0xf8
      12'h61C: dout <= 8'b11111100; // 1564 : 252 - 0xfc
      12'h61D: dout <= 8'b11111100; // 1565 : 252 - 0xfc
      12'h61E: dout <= 8'b11100100; // 1566 : 228 - 0xe4
      12'h61F: dout <= 8'b11101110; // 1567 : 238 - 0xee
      12'h620: dout <= 8'b10010100; // 1568 : 148 - 0x94 -- Sprite 0x62
      12'h621: dout <= 8'b11101010; // 1569 : 234 - 0xea
      12'h622: dout <= 8'b11011110; // 1570 : 222 - 0xde
      12'h623: dout <= 8'b11101110; // 1571 : 238 - 0xee
      12'h624: dout <= 8'b11011110; // 1572 : 222 - 0xde
      12'h625: dout <= 8'b01100110; // 1573 : 102 - 0x66
      12'h626: dout <= 8'b01000010; // 1574 :  66 - 0x42
      12'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout <= 8'b11111110; // 1576 : 254 - 0xfe -- plane 1
      12'h629: dout <= 8'b11111110; // 1577 : 254 - 0xfe
      12'h62A: dout <= 8'b11111110; // 1578 : 254 - 0xfe
      12'h62B: dout <= 8'b11111110; // 1579 : 254 - 0xfe
      12'h62C: dout <= 8'b11111110; // 1580 : 254 - 0xfe
      12'h62D: dout <= 8'b01100110; // 1581 : 102 - 0x66
      12'h62E: dout <= 8'b01000010; // 1582 :  66 - 0x42
      12'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout <= 8'b10010100; // 1584 : 148 - 0x94 -- Sprite 0x63
      12'h631: dout <= 8'b11101010; // 1585 : 234 - 0xea
      12'h632: dout <= 8'b11011110; // 1586 : 222 - 0xde
      12'h633: dout <= 8'b11101110; // 1587 : 238 - 0xee
      12'h634: dout <= 8'b11011110; // 1588 : 222 - 0xde
      12'h635: dout <= 8'b11001110; // 1589 : 206 - 0xce
      12'h636: dout <= 8'b10001100; // 1590 : 140 - 0x8c
      12'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      12'h638: dout <= 8'b11111110; // 1592 : 254 - 0xfe -- plane 1
      12'h639: dout <= 8'b11111110; // 1593 : 254 - 0xfe
      12'h63A: dout <= 8'b11111110; // 1594 : 254 - 0xfe
      12'h63B: dout <= 8'b11111110; // 1595 : 254 - 0xfe
      12'h63C: dout <= 8'b11111110; // 1596 : 254 - 0xfe
      12'h63D: dout <= 8'b11011110; // 1597 : 222 - 0xde
      12'h63E: dout <= 8'b10001100; // 1598 : 140 - 0x8c
      12'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0x64
      12'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      12'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      12'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      12'h644: dout <= 8'b00000000; // 1604 :   0 - 0x0
      12'h645: dout <= 8'b00000000; // 1605 :   0 - 0x0
      12'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      12'h647: dout <= 8'b00000001; // 1607 :   1 - 0x1
      12'h648: dout <= 8'b00000000; // 1608 :   0 - 0x0 -- plane 1
      12'h649: dout <= 8'b00000000; // 1609 :   0 - 0x0
      12'h64A: dout <= 8'b00000000; // 1610 :   0 - 0x0
      12'h64B: dout <= 8'b00000000; // 1611 :   0 - 0x0
      12'h64C: dout <= 8'b00000000; // 1612 :   0 - 0x0
      12'h64D: dout <= 8'b00000000; // 1613 :   0 - 0x0
      12'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0x65
      12'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      12'h652: dout <= 8'b00000000; // 1618 :   0 - 0x0
      12'h653: dout <= 8'b00000000; // 1619 :   0 - 0x0
      12'h654: dout <= 8'b00000000; // 1620 :   0 - 0x0
      12'h655: dout <= 8'b00110110; // 1621 :  54 - 0x36
      12'h656: dout <= 8'b00110110; // 1622 :  54 - 0x36
      12'h657: dout <= 8'b10010000; // 1623 : 144 - 0x90
      12'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- plane 1
      12'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      12'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      12'h65C: dout <= 8'b01101100; // 1628 : 108 - 0x6c
      12'h65D: dout <= 8'b11111110; // 1629 : 254 - 0xfe
      12'h65E: dout <= 8'b11111110; // 1630 : 254 - 0xfe
      12'h65F: dout <= 8'b11111100; // 1631 : 252 - 0xfc
      12'h660: dout <= 8'b00000001; // 1632 :   1 - 0x1 -- Sprite 0x66
      12'h661: dout <= 8'b00000011; // 1633 :   3 - 0x3
      12'h662: dout <= 8'b00000111; // 1634 :   7 - 0x7
      12'h663: dout <= 8'b00000111; // 1635 :   7 - 0x7
      12'h664: dout <= 8'b00011111; // 1636 :  31 - 0x1f
      12'h665: dout <= 8'b00011111; // 1637 :  31 - 0x1f
      12'h666: dout <= 8'b00011100; // 1638 :  28 - 0x1c
      12'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      12'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- plane 1
      12'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout <= 8'b00000000; // 1643 :   0 - 0x0
      12'h66C: dout <= 8'b00000000; // 1644 :   0 - 0x0
      12'h66D: dout <= 8'b00000000; // 1645 :   0 - 0x0
      12'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      12'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      12'h670: dout <= 8'b11111000; // 1648 : 248 - 0xf8 -- Sprite 0x67
      12'h671: dout <= 8'b11111000; // 1649 : 248 - 0xf8
      12'h672: dout <= 8'b11111000; // 1650 : 248 - 0xf8
      12'h673: dout <= 8'b11111000; // 1651 : 248 - 0xf8
      12'h674: dout <= 8'b11111110; // 1652 : 254 - 0xfe
      12'h675: dout <= 8'b11111110; // 1653 : 254 - 0xfe
      12'h676: dout <= 8'b00001110; // 1654 :  14 - 0xe
      12'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      12'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- plane 1
      12'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      12'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      12'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      12'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout <= 8'b00000111; // 1664 :   7 - 0x7 -- Sprite 0x68
      12'h681: dout <= 8'b00001111; // 1665 :  15 - 0xf
      12'h682: dout <= 8'b00011111; // 1666 :  31 - 0x1f
      12'h683: dout <= 8'b00011111; // 1667 :  31 - 0x1f
      12'h684: dout <= 8'b00111111; // 1668 :  63 - 0x3f
      12'h685: dout <= 8'b00111111; // 1669 :  63 - 0x3f
      12'h686: dout <= 8'b00111000; // 1670 :  56 - 0x38
      12'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      12'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- plane 1
      12'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      12'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      12'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      12'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      12'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      12'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      12'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout <= 8'b11111000; // 1680 : 248 - 0xf8 -- Sprite 0x69
      12'h691: dout <= 8'b11110000; // 1681 : 240 - 0xf0
      12'h692: dout <= 8'b11110000; // 1682 : 240 - 0xf0
      12'h693: dout <= 8'b11100000; // 1683 : 224 - 0xe0
      12'h694: dout <= 8'b11111000; // 1684 : 248 - 0xf8
      12'h695: dout <= 8'b11111000; // 1685 : 248 - 0xf8
      12'h696: dout <= 8'b00111000; // 1686 :  56 - 0x38
      12'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      12'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0 -- plane 1
      12'h699: dout <= 8'b00000000; // 1689 :   0 - 0x0
      12'h69A: dout <= 8'b00000000; // 1690 :   0 - 0x0
      12'h69B: dout <= 8'b00000000; // 1691 :   0 - 0x0
      12'h69C: dout <= 8'b00000000; // 1692 :   0 - 0x0
      12'h69D: dout <= 8'b00000000; // 1693 :   0 - 0x0
      12'h69E: dout <= 8'b00000000; // 1694 :   0 - 0x0
      12'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      12'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0x6a
      12'h6A1: dout <= 8'b00011111; // 1697 :  31 - 0x1f
      12'h6A2: dout <= 8'b01111111; // 1698 : 127 - 0x7f
      12'h6A3: dout <= 8'b00111111; // 1699 :  63 - 0x3f
      12'h6A4: dout <= 8'b00001111; // 1700 :  15 - 0xf
      12'h6A5: dout <= 8'b00000111; // 1701 :   7 - 0x7
      12'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      12'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      12'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0 -- plane 1
      12'h6A9: dout <= 8'b00011111; // 1705 :  31 - 0x1f
      12'h6AA: dout <= 8'b01111111; // 1706 : 127 - 0x7f
      12'h6AB: dout <= 8'b00111111; // 1707 :  63 - 0x3f
      12'h6AC: dout <= 8'b00001111; // 1708 :  15 - 0xf
      12'h6AD: dout <= 8'b00000111; // 1709 :   7 - 0x7
      12'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      12'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0x6b
      12'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout <= 8'b11000000; // 1714 : 192 - 0xc0
      12'h6B3: dout <= 8'b11110000; // 1715 : 240 - 0xf0
      12'h6B4: dout <= 8'b11111000; // 1716 : 248 - 0xf8
      12'h6B5: dout <= 8'b11111000; // 1717 : 248 - 0xf8
      12'h6B6: dout <= 8'b11100000; // 1718 : 224 - 0xe0
      12'h6B7: dout <= 8'b00000000; // 1719 :   0 - 0x0
      12'h6B8: dout <= 8'b00000000; // 1720 :   0 - 0x0 -- plane 1
      12'h6B9: dout <= 8'b00000000; // 1721 :   0 - 0x0
      12'h6BA: dout <= 8'b11000000; // 1722 : 192 - 0xc0
      12'h6BB: dout <= 8'b11110000; // 1723 : 240 - 0xf0
      12'h6BC: dout <= 8'b11111000; // 1724 : 248 - 0xf8
      12'h6BD: dout <= 8'b11111000; // 1725 : 248 - 0xf8
      12'h6BE: dout <= 8'b11100000; // 1726 : 224 - 0xe0
      12'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout <= 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0x6c
      12'h6C1: dout <= 8'b00000000; // 1729 :   0 - 0x0
      12'h6C2: dout <= 8'b00000000; // 1730 :   0 - 0x0
      12'h6C3: dout <= 8'b00000000; // 1731 :   0 - 0x0
      12'h6C4: dout <= 8'b00000000; // 1732 :   0 - 0x0
      12'h6C5: dout <= 8'b00000000; // 1733 :   0 - 0x0
      12'h6C6: dout <= 8'b00000000; // 1734 :   0 - 0x0
      12'h6C7: dout <= 8'b00000000; // 1735 :   0 - 0x0
      12'h6C8: dout <= 8'b00000000; // 1736 :   0 - 0x0 -- plane 1
      12'h6C9: dout <= 8'b00000000; // 1737 :   0 - 0x0
      12'h6CA: dout <= 8'b00000000; // 1738 :   0 - 0x0
      12'h6CB: dout <= 8'b00000000; // 1739 :   0 - 0x0
      12'h6CC: dout <= 8'b00000000; // 1740 :   0 - 0x0
      12'h6CD: dout <= 8'b00000000; // 1741 :   0 - 0x0
      12'h6CE: dout <= 8'b00000000; // 1742 :   0 - 0x0
      12'h6CF: dout <= 8'b00000000; // 1743 :   0 - 0x0
      12'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0x6d
      12'h6D1: dout <= 8'b00000000; // 1745 :   0 - 0x0
      12'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      12'h6D3: dout <= 8'b00000000; // 1747 :   0 - 0x0
      12'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      12'h6D5: dout <= 8'b00000000; // 1749 :   0 - 0x0
      12'h6D6: dout <= 8'b00000000; // 1750 :   0 - 0x0
      12'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      12'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0 -- plane 1
      12'h6D9: dout <= 8'b00000000; // 1753 :   0 - 0x0
      12'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      12'h6DB: dout <= 8'b00000000; // 1755 :   0 - 0x0
      12'h6DC: dout <= 8'b00000000; // 1756 :   0 - 0x0
      12'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      12'h6DE: dout <= 8'b00000000; // 1758 :   0 - 0x0
      12'h6DF: dout <= 8'b00000000; // 1759 :   0 - 0x0
      12'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0x6e
      12'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      12'h6E5: dout <= 8'b00000000; // 1765 :   0 - 0x0
      12'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      12'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      12'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- plane 1
      12'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      12'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      12'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      12'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      12'h6ED: dout <= 8'b00000000; // 1773 :   0 - 0x0
      12'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      12'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      12'h6F0: dout <= 8'b00000000; // 1776 :   0 - 0x0 -- Sprite 0x6f
      12'h6F1: dout <= 8'b00000000; // 1777 :   0 - 0x0
      12'h6F2: dout <= 8'b00000000; // 1778 :   0 - 0x0
      12'h6F3: dout <= 8'b00000000; // 1779 :   0 - 0x0
      12'h6F4: dout <= 8'b00000000; // 1780 :   0 - 0x0
      12'h6F5: dout <= 8'b00000000; // 1781 :   0 - 0x0
      12'h6F6: dout <= 8'b00000000; // 1782 :   0 - 0x0
      12'h6F7: dout <= 8'b00000000; // 1783 :   0 - 0x0
      12'h6F8: dout <= 8'b00000000; // 1784 :   0 - 0x0 -- plane 1
      12'h6F9: dout <= 8'b00000000; // 1785 :   0 - 0x0
      12'h6FA: dout <= 8'b00000000; // 1786 :   0 - 0x0
      12'h6FB: dout <= 8'b00000000; // 1787 :   0 - 0x0
      12'h6FC: dout <= 8'b00000000; // 1788 :   0 - 0x0
      12'h6FD: dout <= 8'b00000000; // 1789 :   0 - 0x0
      12'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      12'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout <= 8'b11111111; // 1792 : 255 - 0xff -- Sprite 0x70
      12'h701: dout <= 8'b11111111; // 1793 : 255 - 0xff
      12'h702: dout <= 8'b11111111; // 1794 : 255 - 0xff
      12'h703: dout <= 8'b11111111; // 1795 : 255 - 0xff
      12'h704: dout <= 8'b11111111; // 1796 : 255 - 0xff
      12'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      12'h706: dout <= 8'b11111111; // 1798 : 255 - 0xff
      12'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      12'h708: dout <= 8'b11111111; // 1800 : 255 - 0xff -- plane 1
      12'h709: dout <= 8'b11111111; // 1801 : 255 - 0xff
      12'h70A: dout <= 8'b11111111; // 1802 : 255 - 0xff
      12'h70B: dout <= 8'b11111111; // 1803 : 255 - 0xff
      12'h70C: dout <= 8'b11111111; // 1804 : 255 - 0xff
      12'h70D: dout <= 8'b11111111; // 1805 : 255 - 0xff
      12'h70E: dout <= 8'b11111111; // 1806 : 255 - 0xff
      12'h70F: dout <= 8'b11111111; // 1807 : 255 - 0xff
      12'h710: dout <= 8'b11111111; // 1808 : 255 - 0xff -- Sprite 0x71
      12'h711: dout <= 8'b11111111; // 1809 : 255 - 0xff
      12'h712: dout <= 8'b11111111; // 1810 : 255 - 0xff
      12'h713: dout <= 8'b11111111; // 1811 : 255 - 0xff
      12'h714: dout <= 8'b11111111; // 1812 : 255 - 0xff
      12'h715: dout <= 8'b11111111; // 1813 : 255 - 0xff
      12'h716: dout <= 8'b11111111; // 1814 : 255 - 0xff
      12'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      12'h718: dout <= 8'b11111111; // 1816 : 255 - 0xff -- plane 1
      12'h719: dout <= 8'b11111111; // 1817 : 255 - 0xff
      12'h71A: dout <= 8'b11111111; // 1818 : 255 - 0xff
      12'h71B: dout <= 8'b11111111; // 1819 : 255 - 0xff
      12'h71C: dout <= 8'b11111111; // 1820 : 255 - 0xff
      12'h71D: dout <= 8'b11111111; // 1821 : 255 - 0xff
      12'h71E: dout <= 8'b11111111; // 1822 : 255 - 0xff
      12'h71F: dout <= 8'b11111111; // 1823 : 255 - 0xff
      12'h720: dout <= 8'b11111111; // 1824 : 255 - 0xff -- Sprite 0x72
      12'h721: dout <= 8'b11111111; // 1825 : 255 - 0xff
      12'h722: dout <= 8'b11111111; // 1826 : 255 - 0xff
      12'h723: dout <= 8'b11111111; // 1827 : 255 - 0xff
      12'h724: dout <= 8'b11111111; // 1828 : 255 - 0xff
      12'h725: dout <= 8'b11111111; // 1829 : 255 - 0xff
      12'h726: dout <= 8'b11111111; // 1830 : 255 - 0xff
      12'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      12'h728: dout <= 8'b11111111; // 1832 : 255 - 0xff -- plane 1
      12'h729: dout <= 8'b11111111; // 1833 : 255 - 0xff
      12'h72A: dout <= 8'b11111111; // 1834 : 255 - 0xff
      12'h72B: dout <= 8'b11111111; // 1835 : 255 - 0xff
      12'h72C: dout <= 8'b11111111; // 1836 : 255 - 0xff
      12'h72D: dout <= 8'b11111111; // 1837 : 255 - 0xff
      12'h72E: dout <= 8'b11111111; // 1838 : 255 - 0xff
      12'h72F: dout <= 8'b11111111; // 1839 : 255 - 0xff
      12'h730: dout <= 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0x73
      12'h731: dout <= 8'b11111111; // 1841 : 255 - 0xff
      12'h732: dout <= 8'b11111111; // 1842 : 255 - 0xff
      12'h733: dout <= 8'b11111111; // 1843 : 255 - 0xff
      12'h734: dout <= 8'b11111111; // 1844 : 255 - 0xff
      12'h735: dout <= 8'b11111111; // 1845 : 255 - 0xff
      12'h736: dout <= 8'b11111111; // 1846 : 255 - 0xff
      12'h737: dout <= 8'b11111111; // 1847 : 255 - 0xff
      12'h738: dout <= 8'b11111111; // 1848 : 255 - 0xff -- plane 1
      12'h739: dout <= 8'b11111111; // 1849 : 255 - 0xff
      12'h73A: dout <= 8'b11111111; // 1850 : 255 - 0xff
      12'h73B: dout <= 8'b11111111; // 1851 : 255 - 0xff
      12'h73C: dout <= 8'b11111111; // 1852 : 255 - 0xff
      12'h73D: dout <= 8'b11111111; // 1853 : 255 - 0xff
      12'h73E: dout <= 8'b11111111; // 1854 : 255 - 0xff
      12'h73F: dout <= 8'b11111111; // 1855 : 255 - 0xff
      12'h740: dout <= 8'b11111111; // 1856 : 255 - 0xff -- Sprite 0x74
      12'h741: dout <= 8'b11111111; // 1857 : 255 - 0xff
      12'h742: dout <= 8'b11111111; // 1858 : 255 - 0xff
      12'h743: dout <= 8'b11111111; // 1859 : 255 - 0xff
      12'h744: dout <= 8'b11111111; // 1860 : 255 - 0xff
      12'h745: dout <= 8'b11111111; // 1861 : 255 - 0xff
      12'h746: dout <= 8'b11111111; // 1862 : 255 - 0xff
      12'h747: dout <= 8'b11111111; // 1863 : 255 - 0xff
      12'h748: dout <= 8'b11111111; // 1864 : 255 - 0xff -- plane 1
      12'h749: dout <= 8'b11111111; // 1865 : 255 - 0xff
      12'h74A: dout <= 8'b11111111; // 1866 : 255 - 0xff
      12'h74B: dout <= 8'b11111111; // 1867 : 255 - 0xff
      12'h74C: dout <= 8'b11111111; // 1868 : 255 - 0xff
      12'h74D: dout <= 8'b11111111; // 1869 : 255 - 0xff
      12'h74E: dout <= 8'b11111111; // 1870 : 255 - 0xff
      12'h74F: dout <= 8'b11111111; // 1871 : 255 - 0xff
      12'h750: dout <= 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0x75
      12'h751: dout <= 8'b11111111; // 1873 : 255 - 0xff
      12'h752: dout <= 8'b11111111; // 1874 : 255 - 0xff
      12'h753: dout <= 8'b11111111; // 1875 : 255 - 0xff
      12'h754: dout <= 8'b11111111; // 1876 : 255 - 0xff
      12'h755: dout <= 8'b11111111; // 1877 : 255 - 0xff
      12'h756: dout <= 8'b11111111; // 1878 : 255 - 0xff
      12'h757: dout <= 8'b11111111; // 1879 : 255 - 0xff
      12'h758: dout <= 8'b11111111; // 1880 : 255 - 0xff -- plane 1
      12'h759: dout <= 8'b11111111; // 1881 : 255 - 0xff
      12'h75A: dout <= 8'b11111111; // 1882 : 255 - 0xff
      12'h75B: dout <= 8'b11111111; // 1883 : 255 - 0xff
      12'h75C: dout <= 8'b11111111; // 1884 : 255 - 0xff
      12'h75D: dout <= 8'b11111111; // 1885 : 255 - 0xff
      12'h75E: dout <= 8'b11111111; // 1886 : 255 - 0xff
      12'h75F: dout <= 8'b11111111; // 1887 : 255 - 0xff
      12'h760: dout <= 8'b11111111; // 1888 : 255 - 0xff -- Sprite 0x76
      12'h761: dout <= 8'b11111111; // 1889 : 255 - 0xff
      12'h762: dout <= 8'b11111111; // 1890 : 255 - 0xff
      12'h763: dout <= 8'b11111111; // 1891 : 255 - 0xff
      12'h764: dout <= 8'b11111111; // 1892 : 255 - 0xff
      12'h765: dout <= 8'b11111111; // 1893 : 255 - 0xff
      12'h766: dout <= 8'b11111111; // 1894 : 255 - 0xff
      12'h767: dout <= 8'b11111111; // 1895 : 255 - 0xff
      12'h768: dout <= 8'b11111111; // 1896 : 255 - 0xff -- plane 1
      12'h769: dout <= 8'b11111111; // 1897 : 255 - 0xff
      12'h76A: dout <= 8'b11111111; // 1898 : 255 - 0xff
      12'h76B: dout <= 8'b11111111; // 1899 : 255 - 0xff
      12'h76C: dout <= 8'b11111111; // 1900 : 255 - 0xff
      12'h76D: dout <= 8'b11111111; // 1901 : 255 - 0xff
      12'h76E: dout <= 8'b11111111; // 1902 : 255 - 0xff
      12'h76F: dout <= 8'b11111111; // 1903 : 255 - 0xff
      12'h770: dout <= 8'b11111111; // 1904 : 255 - 0xff -- Sprite 0x77
      12'h771: dout <= 8'b11111111; // 1905 : 255 - 0xff
      12'h772: dout <= 8'b11111111; // 1906 : 255 - 0xff
      12'h773: dout <= 8'b11111111; // 1907 : 255 - 0xff
      12'h774: dout <= 8'b11111111; // 1908 : 255 - 0xff
      12'h775: dout <= 8'b11111111; // 1909 : 255 - 0xff
      12'h776: dout <= 8'b11111111; // 1910 : 255 - 0xff
      12'h777: dout <= 8'b11111111; // 1911 : 255 - 0xff
      12'h778: dout <= 8'b11111111; // 1912 : 255 - 0xff -- plane 1
      12'h779: dout <= 8'b11111111; // 1913 : 255 - 0xff
      12'h77A: dout <= 8'b11111111; // 1914 : 255 - 0xff
      12'h77B: dout <= 8'b11111111; // 1915 : 255 - 0xff
      12'h77C: dout <= 8'b11111111; // 1916 : 255 - 0xff
      12'h77D: dout <= 8'b11111111; // 1917 : 255 - 0xff
      12'h77E: dout <= 8'b11111111; // 1918 : 255 - 0xff
      12'h77F: dout <= 8'b11111111; // 1919 : 255 - 0xff
      12'h780: dout <= 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0x78
      12'h781: dout <= 8'b11111111; // 1921 : 255 - 0xff
      12'h782: dout <= 8'b11111111; // 1922 : 255 - 0xff
      12'h783: dout <= 8'b11111111; // 1923 : 255 - 0xff
      12'h784: dout <= 8'b11111111; // 1924 : 255 - 0xff
      12'h785: dout <= 8'b11111111; // 1925 : 255 - 0xff
      12'h786: dout <= 8'b11111111; // 1926 : 255 - 0xff
      12'h787: dout <= 8'b11111111; // 1927 : 255 - 0xff
      12'h788: dout <= 8'b11111111; // 1928 : 255 - 0xff -- plane 1
      12'h789: dout <= 8'b11111111; // 1929 : 255 - 0xff
      12'h78A: dout <= 8'b11111111; // 1930 : 255 - 0xff
      12'h78B: dout <= 8'b11111111; // 1931 : 255 - 0xff
      12'h78C: dout <= 8'b11111111; // 1932 : 255 - 0xff
      12'h78D: dout <= 8'b11111111; // 1933 : 255 - 0xff
      12'h78E: dout <= 8'b11111111; // 1934 : 255 - 0xff
      12'h78F: dout <= 8'b11111111; // 1935 : 255 - 0xff
      12'h790: dout <= 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0x79
      12'h791: dout <= 8'b11111111; // 1937 : 255 - 0xff
      12'h792: dout <= 8'b11111111; // 1938 : 255 - 0xff
      12'h793: dout <= 8'b11111111; // 1939 : 255 - 0xff
      12'h794: dout <= 8'b11111111; // 1940 : 255 - 0xff
      12'h795: dout <= 8'b11111111; // 1941 : 255 - 0xff
      12'h796: dout <= 8'b11111111; // 1942 : 255 - 0xff
      12'h797: dout <= 8'b11111111; // 1943 : 255 - 0xff
      12'h798: dout <= 8'b11111111; // 1944 : 255 - 0xff -- plane 1
      12'h799: dout <= 8'b11111111; // 1945 : 255 - 0xff
      12'h79A: dout <= 8'b11111111; // 1946 : 255 - 0xff
      12'h79B: dout <= 8'b11111111; // 1947 : 255 - 0xff
      12'h79C: dout <= 8'b11111111; // 1948 : 255 - 0xff
      12'h79D: dout <= 8'b11111111; // 1949 : 255 - 0xff
      12'h79E: dout <= 8'b11111111; // 1950 : 255 - 0xff
      12'h79F: dout <= 8'b11111111; // 1951 : 255 - 0xff
      12'h7A0: dout <= 8'b11111111; // 1952 : 255 - 0xff -- Sprite 0x7a
      12'h7A1: dout <= 8'b11111111; // 1953 : 255 - 0xff
      12'h7A2: dout <= 8'b11111111; // 1954 : 255 - 0xff
      12'h7A3: dout <= 8'b11111111; // 1955 : 255 - 0xff
      12'h7A4: dout <= 8'b11111111; // 1956 : 255 - 0xff
      12'h7A5: dout <= 8'b11111111; // 1957 : 255 - 0xff
      12'h7A6: dout <= 8'b11111111; // 1958 : 255 - 0xff
      12'h7A7: dout <= 8'b11111111; // 1959 : 255 - 0xff
      12'h7A8: dout <= 8'b11111111; // 1960 : 255 - 0xff -- plane 1
      12'h7A9: dout <= 8'b11111111; // 1961 : 255 - 0xff
      12'h7AA: dout <= 8'b11111111; // 1962 : 255 - 0xff
      12'h7AB: dout <= 8'b11111111; // 1963 : 255 - 0xff
      12'h7AC: dout <= 8'b11111111; // 1964 : 255 - 0xff
      12'h7AD: dout <= 8'b11111111; // 1965 : 255 - 0xff
      12'h7AE: dout <= 8'b11111111; // 1966 : 255 - 0xff
      12'h7AF: dout <= 8'b11111111; // 1967 : 255 - 0xff
      12'h7B0: dout <= 8'b11111111; // 1968 : 255 - 0xff -- Sprite 0x7b
      12'h7B1: dout <= 8'b11111111; // 1969 : 255 - 0xff
      12'h7B2: dout <= 8'b11111111; // 1970 : 255 - 0xff
      12'h7B3: dout <= 8'b11111111; // 1971 : 255 - 0xff
      12'h7B4: dout <= 8'b11111111; // 1972 : 255 - 0xff
      12'h7B5: dout <= 8'b11111111; // 1973 : 255 - 0xff
      12'h7B6: dout <= 8'b11111111; // 1974 : 255 - 0xff
      12'h7B7: dout <= 8'b11111111; // 1975 : 255 - 0xff
      12'h7B8: dout <= 8'b11111111; // 1976 : 255 - 0xff -- plane 1
      12'h7B9: dout <= 8'b11111111; // 1977 : 255 - 0xff
      12'h7BA: dout <= 8'b11111111; // 1978 : 255 - 0xff
      12'h7BB: dout <= 8'b11111111; // 1979 : 255 - 0xff
      12'h7BC: dout <= 8'b11111111; // 1980 : 255 - 0xff
      12'h7BD: dout <= 8'b11111111; // 1981 : 255 - 0xff
      12'h7BE: dout <= 8'b11111111; // 1982 : 255 - 0xff
      12'h7BF: dout <= 8'b11111111; // 1983 : 255 - 0xff
      12'h7C0: dout <= 8'b11111111; // 1984 : 255 - 0xff -- Sprite 0x7c
      12'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      12'h7C2: dout <= 8'b11111111; // 1986 : 255 - 0xff
      12'h7C3: dout <= 8'b11111111; // 1987 : 255 - 0xff
      12'h7C4: dout <= 8'b11111111; // 1988 : 255 - 0xff
      12'h7C5: dout <= 8'b11111111; // 1989 : 255 - 0xff
      12'h7C6: dout <= 8'b11111111; // 1990 : 255 - 0xff
      12'h7C7: dout <= 8'b11111111; // 1991 : 255 - 0xff
      12'h7C8: dout <= 8'b11111111; // 1992 : 255 - 0xff -- plane 1
      12'h7C9: dout <= 8'b11111111; // 1993 : 255 - 0xff
      12'h7CA: dout <= 8'b11111111; // 1994 : 255 - 0xff
      12'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      12'h7CC: dout <= 8'b11111111; // 1996 : 255 - 0xff
      12'h7CD: dout <= 8'b11111111; // 1997 : 255 - 0xff
      12'h7CE: dout <= 8'b11111111; // 1998 : 255 - 0xff
      12'h7CF: dout <= 8'b11111111; // 1999 : 255 - 0xff
      12'h7D0: dout <= 8'b11111111; // 2000 : 255 - 0xff -- Sprite 0x7d
      12'h7D1: dout <= 8'b11111111; // 2001 : 255 - 0xff
      12'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      12'h7D3: dout <= 8'b11111111; // 2003 : 255 - 0xff
      12'h7D4: dout <= 8'b11111111; // 2004 : 255 - 0xff
      12'h7D5: dout <= 8'b11111111; // 2005 : 255 - 0xff
      12'h7D6: dout <= 8'b11111111; // 2006 : 255 - 0xff
      12'h7D7: dout <= 8'b11111111; // 2007 : 255 - 0xff
      12'h7D8: dout <= 8'b11111111; // 2008 : 255 - 0xff -- plane 1
      12'h7D9: dout <= 8'b11111111; // 2009 : 255 - 0xff
      12'h7DA: dout <= 8'b11111111; // 2010 : 255 - 0xff
      12'h7DB: dout <= 8'b11111111; // 2011 : 255 - 0xff
      12'h7DC: dout <= 8'b11111111; // 2012 : 255 - 0xff
      12'h7DD: dout <= 8'b11111111; // 2013 : 255 - 0xff
      12'h7DE: dout <= 8'b11111111; // 2014 : 255 - 0xff
      12'h7DF: dout <= 8'b11111111; // 2015 : 255 - 0xff
      12'h7E0: dout <= 8'b11111111; // 2016 : 255 - 0xff -- Sprite 0x7e
      12'h7E1: dout <= 8'b11111111; // 2017 : 255 - 0xff
      12'h7E2: dout <= 8'b11111111; // 2018 : 255 - 0xff
      12'h7E3: dout <= 8'b11111111; // 2019 : 255 - 0xff
      12'h7E4: dout <= 8'b11111111; // 2020 : 255 - 0xff
      12'h7E5: dout <= 8'b11111111; // 2021 : 255 - 0xff
      12'h7E6: dout <= 8'b11111111; // 2022 : 255 - 0xff
      12'h7E7: dout <= 8'b11111111; // 2023 : 255 - 0xff
      12'h7E8: dout <= 8'b11111111; // 2024 : 255 - 0xff -- plane 1
      12'h7E9: dout <= 8'b11111111; // 2025 : 255 - 0xff
      12'h7EA: dout <= 8'b11111111; // 2026 : 255 - 0xff
      12'h7EB: dout <= 8'b11111111; // 2027 : 255 - 0xff
      12'h7EC: dout <= 8'b11111111; // 2028 : 255 - 0xff
      12'h7ED: dout <= 8'b11111111; // 2029 : 255 - 0xff
      12'h7EE: dout <= 8'b11111111; // 2030 : 255 - 0xff
      12'h7EF: dout <= 8'b11111111; // 2031 : 255 - 0xff
      12'h7F0: dout <= 8'b11111111; // 2032 : 255 - 0xff -- Sprite 0x7f
      12'h7F1: dout <= 8'b11111111; // 2033 : 255 - 0xff
      12'h7F2: dout <= 8'b11111111; // 2034 : 255 - 0xff
      12'h7F3: dout <= 8'b11111111; // 2035 : 255 - 0xff
      12'h7F4: dout <= 8'b11111111; // 2036 : 255 - 0xff
      12'h7F5: dout <= 8'b11111111; // 2037 : 255 - 0xff
      12'h7F6: dout <= 8'b11111111; // 2038 : 255 - 0xff
      12'h7F7: dout <= 8'b11111111; // 2039 : 255 - 0xff
      12'h7F8: dout <= 8'b11111111; // 2040 : 255 - 0xff -- plane 1
      12'h7F9: dout <= 8'b11111111; // 2041 : 255 - 0xff
      12'h7FA: dout <= 8'b11111111; // 2042 : 255 - 0xff
      12'h7FB: dout <= 8'b11111111; // 2043 : 255 - 0xff
      12'h7FC: dout <= 8'b11111111; // 2044 : 255 - 0xff
      12'h7FD: dout <= 8'b11111111; // 2045 : 255 - 0xff
      12'h7FE: dout <= 8'b11111111; // 2046 : 255 - 0xff
      12'h7FF: dout <= 8'b11111111; // 2047 : 255 - 0xff
      12'h800: dout <= 8'b11111111; // 2048 : 255 - 0xff -- Sprite 0x80
      12'h801: dout <= 8'b11111111; // 2049 : 255 - 0xff
      12'h802: dout <= 8'b11111111; // 2050 : 255 - 0xff
      12'h803: dout <= 8'b11111111; // 2051 : 255 - 0xff
      12'h804: dout <= 8'b11111111; // 2052 : 255 - 0xff
      12'h805: dout <= 8'b11111111; // 2053 : 255 - 0xff
      12'h806: dout <= 8'b11111111; // 2054 : 255 - 0xff
      12'h807: dout <= 8'b11111111; // 2055 : 255 - 0xff
      12'h808: dout <= 8'b11111111; // 2056 : 255 - 0xff -- plane 1
      12'h809: dout <= 8'b11111111; // 2057 : 255 - 0xff
      12'h80A: dout <= 8'b11111111; // 2058 : 255 - 0xff
      12'h80B: dout <= 8'b11111111; // 2059 : 255 - 0xff
      12'h80C: dout <= 8'b11111111; // 2060 : 255 - 0xff
      12'h80D: dout <= 8'b11111111; // 2061 : 255 - 0xff
      12'h80E: dout <= 8'b11111111; // 2062 : 255 - 0xff
      12'h80F: dout <= 8'b11111111; // 2063 : 255 - 0xff
      12'h810: dout <= 8'b11111111; // 2064 : 255 - 0xff -- Sprite 0x81
      12'h811: dout <= 8'b11111111; // 2065 : 255 - 0xff
      12'h812: dout <= 8'b11111111; // 2066 : 255 - 0xff
      12'h813: dout <= 8'b11111111; // 2067 : 255 - 0xff
      12'h814: dout <= 8'b11111111; // 2068 : 255 - 0xff
      12'h815: dout <= 8'b11111111; // 2069 : 255 - 0xff
      12'h816: dout <= 8'b11111111; // 2070 : 255 - 0xff
      12'h817: dout <= 8'b11111111; // 2071 : 255 - 0xff
      12'h818: dout <= 8'b11111111; // 2072 : 255 - 0xff -- plane 1
      12'h819: dout <= 8'b11111111; // 2073 : 255 - 0xff
      12'h81A: dout <= 8'b11111111; // 2074 : 255 - 0xff
      12'h81B: dout <= 8'b11111111; // 2075 : 255 - 0xff
      12'h81C: dout <= 8'b11111111; // 2076 : 255 - 0xff
      12'h81D: dout <= 8'b11111111; // 2077 : 255 - 0xff
      12'h81E: dout <= 8'b11111111; // 2078 : 255 - 0xff
      12'h81F: dout <= 8'b11111111; // 2079 : 255 - 0xff
      12'h820: dout <= 8'b11111111; // 2080 : 255 - 0xff -- Sprite 0x82
      12'h821: dout <= 8'b11111111; // 2081 : 255 - 0xff
      12'h822: dout <= 8'b11111111; // 2082 : 255 - 0xff
      12'h823: dout <= 8'b11111111; // 2083 : 255 - 0xff
      12'h824: dout <= 8'b11111111; // 2084 : 255 - 0xff
      12'h825: dout <= 8'b11111111; // 2085 : 255 - 0xff
      12'h826: dout <= 8'b11111111; // 2086 : 255 - 0xff
      12'h827: dout <= 8'b11111111; // 2087 : 255 - 0xff
      12'h828: dout <= 8'b11111111; // 2088 : 255 - 0xff -- plane 1
      12'h829: dout <= 8'b11111111; // 2089 : 255 - 0xff
      12'h82A: dout <= 8'b11111111; // 2090 : 255 - 0xff
      12'h82B: dout <= 8'b11111111; // 2091 : 255 - 0xff
      12'h82C: dout <= 8'b11111111; // 2092 : 255 - 0xff
      12'h82D: dout <= 8'b11111111; // 2093 : 255 - 0xff
      12'h82E: dout <= 8'b11111111; // 2094 : 255 - 0xff
      12'h82F: dout <= 8'b11111111; // 2095 : 255 - 0xff
      12'h830: dout <= 8'b11111111; // 2096 : 255 - 0xff -- Sprite 0x83
      12'h831: dout <= 8'b11111111; // 2097 : 255 - 0xff
      12'h832: dout <= 8'b11111111; // 2098 : 255 - 0xff
      12'h833: dout <= 8'b11111111; // 2099 : 255 - 0xff
      12'h834: dout <= 8'b11111111; // 2100 : 255 - 0xff
      12'h835: dout <= 8'b11111111; // 2101 : 255 - 0xff
      12'h836: dout <= 8'b11111111; // 2102 : 255 - 0xff
      12'h837: dout <= 8'b11111111; // 2103 : 255 - 0xff
      12'h838: dout <= 8'b11111111; // 2104 : 255 - 0xff -- plane 1
      12'h839: dout <= 8'b11111111; // 2105 : 255 - 0xff
      12'h83A: dout <= 8'b11111111; // 2106 : 255 - 0xff
      12'h83B: dout <= 8'b11111111; // 2107 : 255 - 0xff
      12'h83C: dout <= 8'b11111111; // 2108 : 255 - 0xff
      12'h83D: dout <= 8'b11111111; // 2109 : 255 - 0xff
      12'h83E: dout <= 8'b11111111; // 2110 : 255 - 0xff
      12'h83F: dout <= 8'b11111111; // 2111 : 255 - 0xff
      12'h840: dout <= 8'b11111111; // 2112 : 255 - 0xff -- Sprite 0x84
      12'h841: dout <= 8'b11111111; // 2113 : 255 - 0xff
      12'h842: dout <= 8'b11111111; // 2114 : 255 - 0xff
      12'h843: dout <= 8'b11111111; // 2115 : 255 - 0xff
      12'h844: dout <= 8'b11111111; // 2116 : 255 - 0xff
      12'h845: dout <= 8'b11111111; // 2117 : 255 - 0xff
      12'h846: dout <= 8'b11111111; // 2118 : 255 - 0xff
      12'h847: dout <= 8'b11111111; // 2119 : 255 - 0xff
      12'h848: dout <= 8'b11111111; // 2120 : 255 - 0xff -- plane 1
      12'h849: dout <= 8'b11111111; // 2121 : 255 - 0xff
      12'h84A: dout <= 8'b11111111; // 2122 : 255 - 0xff
      12'h84B: dout <= 8'b11111111; // 2123 : 255 - 0xff
      12'h84C: dout <= 8'b11111111; // 2124 : 255 - 0xff
      12'h84D: dout <= 8'b11111111; // 2125 : 255 - 0xff
      12'h84E: dout <= 8'b11111111; // 2126 : 255 - 0xff
      12'h84F: dout <= 8'b11111111; // 2127 : 255 - 0xff
      12'h850: dout <= 8'b11111111; // 2128 : 255 - 0xff -- Sprite 0x85
      12'h851: dout <= 8'b11111111; // 2129 : 255 - 0xff
      12'h852: dout <= 8'b11111111; // 2130 : 255 - 0xff
      12'h853: dout <= 8'b11111111; // 2131 : 255 - 0xff
      12'h854: dout <= 8'b11111111; // 2132 : 255 - 0xff
      12'h855: dout <= 8'b11111111; // 2133 : 255 - 0xff
      12'h856: dout <= 8'b11111111; // 2134 : 255 - 0xff
      12'h857: dout <= 8'b11111111; // 2135 : 255 - 0xff
      12'h858: dout <= 8'b11111111; // 2136 : 255 - 0xff -- plane 1
      12'h859: dout <= 8'b11111111; // 2137 : 255 - 0xff
      12'h85A: dout <= 8'b11111111; // 2138 : 255 - 0xff
      12'h85B: dout <= 8'b11111111; // 2139 : 255 - 0xff
      12'h85C: dout <= 8'b11111111; // 2140 : 255 - 0xff
      12'h85D: dout <= 8'b11111111; // 2141 : 255 - 0xff
      12'h85E: dout <= 8'b11111111; // 2142 : 255 - 0xff
      12'h85F: dout <= 8'b11111111; // 2143 : 255 - 0xff
      12'h860: dout <= 8'b11111111; // 2144 : 255 - 0xff -- Sprite 0x86
      12'h861: dout <= 8'b11111111; // 2145 : 255 - 0xff
      12'h862: dout <= 8'b11111111; // 2146 : 255 - 0xff
      12'h863: dout <= 8'b11111111; // 2147 : 255 - 0xff
      12'h864: dout <= 8'b11111111; // 2148 : 255 - 0xff
      12'h865: dout <= 8'b11111111; // 2149 : 255 - 0xff
      12'h866: dout <= 8'b11111111; // 2150 : 255 - 0xff
      12'h867: dout <= 8'b11111111; // 2151 : 255 - 0xff
      12'h868: dout <= 8'b11111111; // 2152 : 255 - 0xff -- plane 1
      12'h869: dout <= 8'b11111111; // 2153 : 255 - 0xff
      12'h86A: dout <= 8'b11111111; // 2154 : 255 - 0xff
      12'h86B: dout <= 8'b11111111; // 2155 : 255 - 0xff
      12'h86C: dout <= 8'b11111111; // 2156 : 255 - 0xff
      12'h86D: dout <= 8'b11111111; // 2157 : 255 - 0xff
      12'h86E: dout <= 8'b11111111; // 2158 : 255 - 0xff
      12'h86F: dout <= 8'b11111111; // 2159 : 255 - 0xff
      12'h870: dout <= 8'b11111111; // 2160 : 255 - 0xff -- Sprite 0x87
      12'h871: dout <= 8'b11111111; // 2161 : 255 - 0xff
      12'h872: dout <= 8'b11111111; // 2162 : 255 - 0xff
      12'h873: dout <= 8'b11111111; // 2163 : 255 - 0xff
      12'h874: dout <= 8'b11111111; // 2164 : 255 - 0xff
      12'h875: dout <= 8'b11111111; // 2165 : 255 - 0xff
      12'h876: dout <= 8'b11111111; // 2166 : 255 - 0xff
      12'h877: dout <= 8'b11111111; // 2167 : 255 - 0xff
      12'h878: dout <= 8'b11111111; // 2168 : 255 - 0xff -- plane 1
      12'h879: dout <= 8'b11111111; // 2169 : 255 - 0xff
      12'h87A: dout <= 8'b11111111; // 2170 : 255 - 0xff
      12'h87B: dout <= 8'b11111111; // 2171 : 255 - 0xff
      12'h87C: dout <= 8'b11111111; // 2172 : 255 - 0xff
      12'h87D: dout <= 8'b11111111; // 2173 : 255 - 0xff
      12'h87E: dout <= 8'b11111111; // 2174 : 255 - 0xff
      12'h87F: dout <= 8'b11111111; // 2175 : 255 - 0xff
      12'h880: dout <= 8'b11111111; // 2176 : 255 - 0xff -- Sprite 0x88
      12'h881: dout <= 8'b11111111; // 2177 : 255 - 0xff
      12'h882: dout <= 8'b11111111; // 2178 : 255 - 0xff
      12'h883: dout <= 8'b11111111; // 2179 : 255 - 0xff
      12'h884: dout <= 8'b11111111; // 2180 : 255 - 0xff
      12'h885: dout <= 8'b11111111; // 2181 : 255 - 0xff
      12'h886: dout <= 8'b11111111; // 2182 : 255 - 0xff
      12'h887: dout <= 8'b11111111; // 2183 : 255 - 0xff
      12'h888: dout <= 8'b11111111; // 2184 : 255 - 0xff -- plane 1
      12'h889: dout <= 8'b11111111; // 2185 : 255 - 0xff
      12'h88A: dout <= 8'b11111111; // 2186 : 255 - 0xff
      12'h88B: dout <= 8'b11111111; // 2187 : 255 - 0xff
      12'h88C: dout <= 8'b11111111; // 2188 : 255 - 0xff
      12'h88D: dout <= 8'b11111111; // 2189 : 255 - 0xff
      12'h88E: dout <= 8'b11111111; // 2190 : 255 - 0xff
      12'h88F: dout <= 8'b11111111; // 2191 : 255 - 0xff
      12'h890: dout <= 8'b11111111; // 2192 : 255 - 0xff -- Sprite 0x89
      12'h891: dout <= 8'b11111111; // 2193 : 255 - 0xff
      12'h892: dout <= 8'b11111111; // 2194 : 255 - 0xff
      12'h893: dout <= 8'b11111111; // 2195 : 255 - 0xff
      12'h894: dout <= 8'b11111111; // 2196 : 255 - 0xff
      12'h895: dout <= 8'b11111111; // 2197 : 255 - 0xff
      12'h896: dout <= 8'b11111111; // 2198 : 255 - 0xff
      12'h897: dout <= 8'b11111111; // 2199 : 255 - 0xff
      12'h898: dout <= 8'b11111111; // 2200 : 255 - 0xff -- plane 1
      12'h899: dout <= 8'b11111111; // 2201 : 255 - 0xff
      12'h89A: dout <= 8'b11111111; // 2202 : 255 - 0xff
      12'h89B: dout <= 8'b11111111; // 2203 : 255 - 0xff
      12'h89C: dout <= 8'b11111111; // 2204 : 255 - 0xff
      12'h89D: dout <= 8'b11111111; // 2205 : 255 - 0xff
      12'h89E: dout <= 8'b11111111; // 2206 : 255 - 0xff
      12'h89F: dout <= 8'b11111111; // 2207 : 255 - 0xff
      12'h8A0: dout <= 8'b11111111; // 2208 : 255 - 0xff -- Sprite 0x8a
      12'h8A1: dout <= 8'b11111111; // 2209 : 255 - 0xff
      12'h8A2: dout <= 8'b11111111; // 2210 : 255 - 0xff
      12'h8A3: dout <= 8'b11111111; // 2211 : 255 - 0xff
      12'h8A4: dout <= 8'b11111111; // 2212 : 255 - 0xff
      12'h8A5: dout <= 8'b11111111; // 2213 : 255 - 0xff
      12'h8A6: dout <= 8'b11111111; // 2214 : 255 - 0xff
      12'h8A7: dout <= 8'b11111111; // 2215 : 255 - 0xff
      12'h8A8: dout <= 8'b11111111; // 2216 : 255 - 0xff -- plane 1
      12'h8A9: dout <= 8'b11111111; // 2217 : 255 - 0xff
      12'h8AA: dout <= 8'b11111111; // 2218 : 255 - 0xff
      12'h8AB: dout <= 8'b11111111; // 2219 : 255 - 0xff
      12'h8AC: dout <= 8'b11111111; // 2220 : 255 - 0xff
      12'h8AD: dout <= 8'b11111111; // 2221 : 255 - 0xff
      12'h8AE: dout <= 8'b11111111; // 2222 : 255 - 0xff
      12'h8AF: dout <= 8'b11111111; // 2223 : 255 - 0xff
      12'h8B0: dout <= 8'b11111111; // 2224 : 255 - 0xff -- Sprite 0x8b
      12'h8B1: dout <= 8'b11111111; // 2225 : 255 - 0xff
      12'h8B2: dout <= 8'b11111111; // 2226 : 255 - 0xff
      12'h8B3: dout <= 8'b11111111; // 2227 : 255 - 0xff
      12'h8B4: dout <= 8'b11111111; // 2228 : 255 - 0xff
      12'h8B5: dout <= 8'b11111111; // 2229 : 255 - 0xff
      12'h8B6: dout <= 8'b11111111; // 2230 : 255 - 0xff
      12'h8B7: dout <= 8'b11111111; // 2231 : 255 - 0xff
      12'h8B8: dout <= 8'b11111111; // 2232 : 255 - 0xff -- plane 1
      12'h8B9: dout <= 8'b11111111; // 2233 : 255 - 0xff
      12'h8BA: dout <= 8'b11111111; // 2234 : 255 - 0xff
      12'h8BB: dout <= 8'b11111111; // 2235 : 255 - 0xff
      12'h8BC: dout <= 8'b11111111; // 2236 : 255 - 0xff
      12'h8BD: dout <= 8'b11111111; // 2237 : 255 - 0xff
      12'h8BE: dout <= 8'b11111111; // 2238 : 255 - 0xff
      12'h8BF: dout <= 8'b11111111; // 2239 : 255 - 0xff
      12'h8C0: dout <= 8'b11111111; // 2240 : 255 - 0xff -- Sprite 0x8c
      12'h8C1: dout <= 8'b11111111; // 2241 : 255 - 0xff
      12'h8C2: dout <= 8'b11111111; // 2242 : 255 - 0xff
      12'h8C3: dout <= 8'b11111111; // 2243 : 255 - 0xff
      12'h8C4: dout <= 8'b11111111; // 2244 : 255 - 0xff
      12'h8C5: dout <= 8'b11111111; // 2245 : 255 - 0xff
      12'h8C6: dout <= 8'b11111111; // 2246 : 255 - 0xff
      12'h8C7: dout <= 8'b11111111; // 2247 : 255 - 0xff
      12'h8C8: dout <= 8'b11111111; // 2248 : 255 - 0xff -- plane 1
      12'h8C9: dout <= 8'b11111111; // 2249 : 255 - 0xff
      12'h8CA: dout <= 8'b11111111; // 2250 : 255 - 0xff
      12'h8CB: dout <= 8'b11111111; // 2251 : 255 - 0xff
      12'h8CC: dout <= 8'b11111111; // 2252 : 255 - 0xff
      12'h8CD: dout <= 8'b11111111; // 2253 : 255 - 0xff
      12'h8CE: dout <= 8'b11111111; // 2254 : 255 - 0xff
      12'h8CF: dout <= 8'b11111111; // 2255 : 255 - 0xff
      12'h8D0: dout <= 8'b11111111; // 2256 : 255 - 0xff -- Sprite 0x8d
      12'h8D1: dout <= 8'b11111111; // 2257 : 255 - 0xff
      12'h8D2: dout <= 8'b11111111; // 2258 : 255 - 0xff
      12'h8D3: dout <= 8'b11111111; // 2259 : 255 - 0xff
      12'h8D4: dout <= 8'b11111111; // 2260 : 255 - 0xff
      12'h8D5: dout <= 8'b11111111; // 2261 : 255 - 0xff
      12'h8D6: dout <= 8'b11111111; // 2262 : 255 - 0xff
      12'h8D7: dout <= 8'b11111111; // 2263 : 255 - 0xff
      12'h8D8: dout <= 8'b11111111; // 2264 : 255 - 0xff -- plane 1
      12'h8D9: dout <= 8'b11111111; // 2265 : 255 - 0xff
      12'h8DA: dout <= 8'b11111111; // 2266 : 255 - 0xff
      12'h8DB: dout <= 8'b11111111; // 2267 : 255 - 0xff
      12'h8DC: dout <= 8'b11111111; // 2268 : 255 - 0xff
      12'h8DD: dout <= 8'b11111111; // 2269 : 255 - 0xff
      12'h8DE: dout <= 8'b11111111; // 2270 : 255 - 0xff
      12'h8DF: dout <= 8'b11111111; // 2271 : 255 - 0xff
      12'h8E0: dout <= 8'b11111111; // 2272 : 255 - 0xff -- Sprite 0x8e
      12'h8E1: dout <= 8'b11111111; // 2273 : 255 - 0xff
      12'h8E2: dout <= 8'b11111111; // 2274 : 255 - 0xff
      12'h8E3: dout <= 8'b11111111; // 2275 : 255 - 0xff
      12'h8E4: dout <= 8'b11111111; // 2276 : 255 - 0xff
      12'h8E5: dout <= 8'b11111111; // 2277 : 255 - 0xff
      12'h8E6: dout <= 8'b11111111; // 2278 : 255 - 0xff
      12'h8E7: dout <= 8'b11111111; // 2279 : 255 - 0xff
      12'h8E8: dout <= 8'b11111111; // 2280 : 255 - 0xff -- plane 1
      12'h8E9: dout <= 8'b11111111; // 2281 : 255 - 0xff
      12'h8EA: dout <= 8'b11111111; // 2282 : 255 - 0xff
      12'h8EB: dout <= 8'b11111111; // 2283 : 255 - 0xff
      12'h8EC: dout <= 8'b11111111; // 2284 : 255 - 0xff
      12'h8ED: dout <= 8'b11111111; // 2285 : 255 - 0xff
      12'h8EE: dout <= 8'b11111111; // 2286 : 255 - 0xff
      12'h8EF: dout <= 8'b11111111; // 2287 : 255 - 0xff
      12'h8F0: dout <= 8'b11111111; // 2288 : 255 - 0xff -- Sprite 0x8f
      12'h8F1: dout <= 8'b11111111; // 2289 : 255 - 0xff
      12'h8F2: dout <= 8'b11111111; // 2290 : 255 - 0xff
      12'h8F3: dout <= 8'b11111111; // 2291 : 255 - 0xff
      12'h8F4: dout <= 8'b11111111; // 2292 : 255 - 0xff
      12'h8F5: dout <= 8'b11111111; // 2293 : 255 - 0xff
      12'h8F6: dout <= 8'b11111111; // 2294 : 255 - 0xff
      12'h8F7: dout <= 8'b11111111; // 2295 : 255 - 0xff
      12'h8F8: dout <= 8'b11111111; // 2296 : 255 - 0xff -- plane 1
      12'h8F9: dout <= 8'b11111111; // 2297 : 255 - 0xff
      12'h8FA: dout <= 8'b11111111; // 2298 : 255 - 0xff
      12'h8FB: dout <= 8'b11111111; // 2299 : 255 - 0xff
      12'h8FC: dout <= 8'b11111111; // 2300 : 255 - 0xff
      12'h8FD: dout <= 8'b11111111; // 2301 : 255 - 0xff
      12'h8FE: dout <= 8'b11111111; // 2302 : 255 - 0xff
      12'h8FF: dout <= 8'b11111111; // 2303 : 255 - 0xff
      12'h900: dout <= 8'b00000000; // 2304 :   0 - 0x0 -- Sprite 0x90
      12'h901: dout <= 8'b00000000; // 2305 :   0 - 0x0
      12'h902: dout <= 8'b00000000; // 2306 :   0 - 0x0
      12'h903: dout <= 8'b00000000; // 2307 :   0 - 0x0
      12'h904: dout <= 8'b00000000; // 2308 :   0 - 0x0
      12'h905: dout <= 8'b00000001; // 2309 :   1 - 0x1
      12'h906: dout <= 8'b00011110; // 2310 :  30 - 0x1e
      12'h907: dout <= 8'b00111011; // 2311 :  59 - 0x3b
      12'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0 -- plane 1
      12'h909: dout <= 8'b00000000; // 2313 :   0 - 0x0
      12'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout <= 8'b00000000; // 2315 :   0 - 0x0
      12'h90C: dout <= 8'b00000000; // 2316 :   0 - 0x0
      12'h90D: dout <= 8'b00000000; // 2317 :   0 - 0x0
      12'h90E: dout <= 8'b00000000; // 2318 :   0 - 0x0
      12'h90F: dout <= 8'b00000000; // 2319 :   0 - 0x0
      12'h910: dout <= 8'b00000000; // 2320 :   0 - 0x0 -- Sprite 0x91
      12'h911: dout <= 8'b00000000; // 2321 :   0 - 0x0
      12'h912: dout <= 8'b00001100; // 2322 :  12 - 0xc
      12'h913: dout <= 8'b00111100; // 2323 :  60 - 0x3c
      12'h914: dout <= 8'b11010000; // 2324 : 208 - 0xd0
      12'h915: dout <= 8'b00010000; // 2325 :  16 - 0x10
      12'h916: dout <= 8'b00100000; // 2326 :  32 - 0x20
      12'h917: dout <= 8'b01000000; // 2327 :  64 - 0x40
      12'h918: dout <= 8'b00000000; // 2328 :   0 - 0x0 -- plane 1
      12'h919: dout <= 8'b00000000; // 2329 :   0 - 0x0
      12'h91A: dout <= 8'b00000000; // 2330 :   0 - 0x0
      12'h91B: dout <= 8'b00000000; // 2331 :   0 - 0x0
      12'h91C: dout <= 8'b00000000; // 2332 :   0 - 0x0
      12'h91D: dout <= 8'b00000000; // 2333 :   0 - 0x0
      12'h91E: dout <= 8'b00000000; // 2334 :   0 - 0x0
      12'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout <= 8'b00111110; // 2336 :  62 - 0x3e -- Sprite 0x92
      12'h921: dout <= 8'b00101101; // 2337 :  45 - 0x2d
      12'h922: dout <= 8'b00110101; // 2338 :  53 - 0x35
      12'h923: dout <= 8'b00011101; // 2339 :  29 - 0x1d
      12'h924: dout <= 8'b00000001; // 2340 :   1 - 0x1
      12'h925: dout <= 8'b00000000; // 2341 :   0 - 0x0
      12'h926: dout <= 8'b00000000; // 2342 :   0 - 0x0
      12'h927: dout <= 8'b00000000; // 2343 :   0 - 0x0
      12'h928: dout <= 8'b00000000; // 2344 :   0 - 0x0 -- plane 1
      12'h929: dout <= 8'b00000000; // 2345 :   0 - 0x0
      12'h92A: dout <= 8'b00000000; // 2346 :   0 - 0x0
      12'h92B: dout <= 8'b00000000; // 2347 :   0 - 0x0
      12'h92C: dout <= 8'b00000000; // 2348 :   0 - 0x0
      12'h92D: dout <= 8'b00000000; // 2349 :   0 - 0x0
      12'h92E: dout <= 8'b00000000; // 2350 :   0 - 0x0
      12'h92F: dout <= 8'b00000000; // 2351 :   0 - 0x0
      12'h930: dout <= 8'b10110000; // 2352 : 176 - 0xb0 -- Sprite 0x93
      12'h931: dout <= 8'b10111000; // 2353 : 184 - 0xb8
      12'h932: dout <= 8'b11111000; // 2354 : 248 - 0xf8
      12'h933: dout <= 8'b01111000; // 2355 : 120 - 0x78
      12'h934: dout <= 8'b10011000; // 2356 : 152 - 0x98
      12'h935: dout <= 8'b11110000; // 2357 : 240 - 0xf0
      12'h936: dout <= 8'b00000000; // 2358 :   0 - 0x0
      12'h937: dout <= 8'b00000000; // 2359 :   0 - 0x0
      12'h938: dout <= 8'b00000000; // 2360 :   0 - 0x0 -- plane 1
      12'h939: dout <= 8'b00000000; // 2361 :   0 - 0x0
      12'h93A: dout <= 8'b00000000; // 2362 :   0 - 0x0
      12'h93B: dout <= 8'b00000000; // 2363 :   0 - 0x0
      12'h93C: dout <= 8'b00000000; // 2364 :   0 - 0x0
      12'h93D: dout <= 8'b00000000; // 2365 :   0 - 0x0
      12'h93E: dout <= 8'b00000000; // 2366 :   0 - 0x0
      12'h93F: dout <= 8'b00000000; // 2367 :   0 - 0x0
      12'h940: dout <= 8'b00000000; // 2368 :   0 - 0x0 -- Sprite 0x94
      12'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout <= 8'b00000111; // 2370 :   7 - 0x7
      12'h943: dout <= 8'b00000011; // 2371 :   3 - 0x3
      12'h944: dout <= 8'b00001101; // 2372 :  13 - 0xd
      12'h945: dout <= 8'b00011110; // 2373 :  30 - 0x1e
      12'h946: dout <= 8'b00010111; // 2374 :  23 - 0x17
      12'h947: dout <= 8'b00011101; // 2375 :  29 - 0x1d
      12'h948: dout <= 8'b00000000; // 2376 :   0 - 0x0 -- plane 1
      12'h949: dout <= 8'b00000000; // 2377 :   0 - 0x0
      12'h94A: dout <= 8'b00000000; // 2378 :   0 - 0x0
      12'h94B: dout <= 8'b00000000; // 2379 :   0 - 0x0
      12'h94C: dout <= 8'b00000000; // 2380 :   0 - 0x0
      12'h94D: dout <= 8'b00000000; // 2381 :   0 - 0x0
      12'h94E: dout <= 8'b00000000; // 2382 :   0 - 0x0
      12'h94F: dout <= 8'b00000000; // 2383 :   0 - 0x0
      12'h950: dout <= 8'b00000000; // 2384 :   0 - 0x0 -- Sprite 0x95
      12'h951: dout <= 8'b10000000; // 2385 : 128 - 0x80
      12'h952: dout <= 8'b01110000; // 2386 : 112 - 0x70
      12'h953: dout <= 8'b11100000; // 2387 : 224 - 0xe0
      12'h954: dout <= 8'b11011000; // 2388 : 216 - 0xd8
      12'h955: dout <= 8'b10111100; // 2389 : 188 - 0xbc
      12'h956: dout <= 8'b01110100; // 2390 : 116 - 0x74
      12'h957: dout <= 8'b11011100; // 2391 : 220 - 0xdc
      12'h958: dout <= 8'b00000000; // 2392 :   0 - 0x0 -- plane 1
      12'h959: dout <= 8'b00000000; // 2393 :   0 - 0x0
      12'h95A: dout <= 8'b00000000; // 2394 :   0 - 0x0
      12'h95B: dout <= 8'b00000000; // 2395 :   0 - 0x0
      12'h95C: dout <= 8'b00000000; // 2396 :   0 - 0x0
      12'h95D: dout <= 8'b00000000; // 2397 :   0 - 0x0
      12'h95E: dout <= 8'b00000000; // 2398 :   0 - 0x0
      12'h95F: dout <= 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout <= 8'b00011111; // 2400 :  31 - 0x1f -- Sprite 0x96
      12'h961: dout <= 8'b00001011; // 2401 :  11 - 0xb
      12'h962: dout <= 8'b00001111; // 2402 :  15 - 0xf
      12'h963: dout <= 8'b00000101; // 2403 :   5 - 0x5
      12'h964: dout <= 8'b00000011; // 2404 :   3 - 0x3
      12'h965: dout <= 8'b00000001; // 2405 :   1 - 0x1
      12'h966: dout <= 8'b00000000; // 2406 :   0 - 0x0
      12'h967: dout <= 8'b00000000; // 2407 :   0 - 0x0
      12'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0 -- plane 1
      12'h969: dout <= 8'b00000000; // 2409 :   0 - 0x0
      12'h96A: dout <= 8'b00000000; // 2410 :   0 - 0x0
      12'h96B: dout <= 8'b00000000; // 2411 :   0 - 0x0
      12'h96C: dout <= 8'b00000000; // 2412 :   0 - 0x0
      12'h96D: dout <= 8'b00000000; // 2413 :   0 - 0x0
      12'h96E: dout <= 8'b00000000; // 2414 :   0 - 0x0
      12'h96F: dout <= 8'b00000000; // 2415 :   0 - 0x0
      12'h970: dout <= 8'b11111100; // 2416 : 252 - 0xfc -- Sprite 0x97
      12'h971: dout <= 8'b01101000; // 2417 : 104 - 0x68
      12'h972: dout <= 8'b11111000; // 2418 : 248 - 0xf8
      12'h973: dout <= 8'b10110000; // 2419 : 176 - 0xb0
      12'h974: dout <= 8'b11100000; // 2420 : 224 - 0xe0
      12'h975: dout <= 8'b10000000; // 2421 : 128 - 0x80
      12'h976: dout <= 8'b00000000; // 2422 :   0 - 0x0
      12'h977: dout <= 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout <= 8'b00000000; // 2424 :   0 - 0x0 -- plane 1
      12'h979: dout <= 8'b00000000; // 2425 :   0 - 0x0
      12'h97A: dout <= 8'b00000000; // 2426 :   0 - 0x0
      12'h97B: dout <= 8'b00000000; // 2427 :   0 - 0x0
      12'h97C: dout <= 8'b00000000; // 2428 :   0 - 0x0
      12'h97D: dout <= 8'b00000000; // 2429 :   0 - 0x0
      12'h97E: dout <= 8'b00000000; // 2430 :   0 - 0x0
      12'h97F: dout <= 8'b00000000; // 2431 :   0 - 0x0
      12'h980: dout <= 8'b00000000; // 2432 :   0 - 0x0 -- Sprite 0x98
      12'h981: dout <= 8'b00000000; // 2433 :   0 - 0x0
      12'h982: dout <= 8'b00000000; // 2434 :   0 - 0x0
      12'h983: dout <= 8'b00000001; // 2435 :   1 - 0x1
      12'h984: dout <= 8'b00000001; // 2436 :   1 - 0x1
      12'h985: dout <= 8'b00001011; // 2437 :  11 - 0xb
      12'h986: dout <= 8'b00011100; // 2438 :  28 - 0x1c
      12'h987: dout <= 8'b00111111; // 2439 :  63 - 0x3f
      12'h988: dout <= 8'b00000000; // 2440 :   0 - 0x0 -- plane 1
      12'h989: dout <= 8'b00000000; // 2441 :   0 - 0x0
      12'h98A: dout <= 8'b00000000; // 2442 :   0 - 0x0
      12'h98B: dout <= 8'b00000000; // 2443 :   0 - 0x0
      12'h98C: dout <= 8'b00000000; // 2444 :   0 - 0x0
      12'h98D: dout <= 8'b00000000; // 2445 :   0 - 0x0
      12'h98E: dout <= 8'b00000000; // 2446 :   0 - 0x0
      12'h98F: dout <= 8'b00000000; // 2447 :   0 - 0x0
      12'h990: dout <= 8'b00000000; // 2448 :   0 - 0x0 -- Sprite 0x99
      12'h991: dout <= 8'b00000000; // 2449 :   0 - 0x0
      12'h992: dout <= 8'b00110000; // 2450 :  48 - 0x30
      12'h993: dout <= 8'b01111000; // 2451 : 120 - 0x78
      12'h994: dout <= 8'b10000000; // 2452 : 128 - 0x80
      12'h995: dout <= 8'b11110000; // 2453 : 240 - 0xf0
      12'h996: dout <= 8'b11111000; // 2454 : 248 - 0xf8
      12'h997: dout <= 8'b11111100; // 2455 : 252 - 0xfc
      12'h998: dout <= 8'b00000000; // 2456 :   0 - 0x0 -- plane 1
      12'h999: dout <= 8'b00000000; // 2457 :   0 - 0x0
      12'h99A: dout <= 8'b00000000; // 2458 :   0 - 0x0
      12'h99B: dout <= 8'b00000000; // 2459 :   0 - 0x0
      12'h99C: dout <= 8'b00000000; // 2460 :   0 - 0x0
      12'h99D: dout <= 8'b00000000; // 2461 :   0 - 0x0
      12'h99E: dout <= 8'b00000000; // 2462 :   0 - 0x0
      12'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout <= 8'b00111111; // 2464 :  63 - 0x3f -- Sprite 0x9a
      12'h9A1: dout <= 8'b00111111; // 2465 :  63 - 0x3f
      12'h9A2: dout <= 8'b00111111; // 2466 :  63 - 0x3f
      12'h9A3: dout <= 8'b00011111; // 2467 :  31 - 0x1f
      12'h9A4: dout <= 8'b00011111; // 2468 :  31 - 0x1f
      12'h9A5: dout <= 8'b00000111; // 2469 :   7 - 0x7
      12'h9A6: dout <= 8'b00000000; // 2470 :   0 - 0x0
      12'h9A7: dout <= 8'b00000000; // 2471 :   0 - 0x0
      12'h9A8: dout <= 8'b00000000; // 2472 :   0 - 0x0 -- plane 1
      12'h9A9: dout <= 8'b00000000; // 2473 :   0 - 0x0
      12'h9AA: dout <= 8'b00000000; // 2474 :   0 - 0x0
      12'h9AB: dout <= 8'b00000000; // 2475 :   0 - 0x0
      12'h9AC: dout <= 8'b00000000; // 2476 :   0 - 0x0
      12'h9AD: dout <= 8'b00000000; // 2477 :   0 - 0x0
      12'h9AE: dout <= 8'b00000000; // 2478 :   0 - 0x0
      12'h9AF: dout <= 8'b00000000; // 2479 :   0 - 0x0
      12'h9B0: dout <= 8'b11111100; // 2480 : 252 - 0xfc -- Sprite 0x9b
      12'h9B1: dout <= 8'b11101100; // 2481 : 236 - 0xec
      12'h9B2: dout <= 8'b11101100; // 2482 : 236 - 0xec
      12'h9B3: dout <= 8'b11011000; // 2483 : 216 - 0xd8
      12'h9B4: dout <= 8'b11111000; // 2484 : 248 - 0xf8
      12'h9B5: dout <= 8'b11100000; // 2485 : 224 - 0xe0
      12'h9B6: dout <= 8'b00000000; // 2486 :   0 - 0x0
      12'h9B7: dout <= 8'b00000000; // 2487 :   0 - 0x0
      12'h9B8: dout <= 8'b00000000; // 2488 :   0 - 0x0 -- plane 1
      12'h9B9: dout <= 8'b00000000; // 2489 :   0 - 0x0
      12'h9BA: dout <= 8'b00000000; // 2490 :   0 - 0x0
      12'h9BB: dout <= 8'b00000000; // 2491 :   0 - 0x0
      12'h9BC: dout <= 8'b00000000; // 2492 :   0 - 0x0
      12'h9BD: dout <= 8'b00000000; // 2493 :   0 - 0x0
      12'h9BE: dout <= 8'b00000000; // 2494 :   0 - 0x0
      12'h9BF: dout <= 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout <= 8'b00000000; // 2496 :   0 - 0x0 -- Sprite 0x9c
      12'h9C1: dout <= 8'b00000000; // 2497 :   0 - 0x0
      12'h9C2: dout <= 8'b00000001; // 2498 :   1 - 0x1
      12'h9C3: dout <= 8'b00011101; // 2499 :  29 - 0x1d
      12'h9C4: dout <= 8'b00111110; // 2500 :  62 - 0x3e
      12'h9C5: dout <= 8'b00111111; // 2501 :  63 - 0x3f
      12'h9C6: dout <= 8'b00111111; // 2502 :  63 - 0x3f
      12'h9C7: dout <= 8'b00111111; // 2503 :  63 - 0x3f
      12'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0 -- plane 1
      12'h9C9: dout <= 8'b00000000; // 2505 :   0 - 0x0
      12'h9CA: dout <= 8'b00000000; // 2506 :   0 - 0x0
      12'h9CB: dout <= 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout <= 8'b00000000; // 2508 :   0 - 0x0
      12'h9CD: dout <= 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout <= 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout <= 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout <= 8'b00000000; // 2512 :   0 - 0x0 -- Sprite 0x9d
      12'h9D1: dout <= 8'b10000000; // 2513 : 128 - 0x80
      12'h9D2: dout <= 8'b00000000; // 2514 :   0 - 0x0
      12'h9D3: dout <= 8'b01110000; // 2515 : 112 - 0x70
      12'h9D4: dout <= 8'b11111000; // 2516 : 248 - 0xf8
      12'h9D5: dout <= 8'b11111100; // 2517 : 252 - 0xfc
      12'h9D6: dout <= 8'b11111100; // 2518 : 252 - 0xfc
      12'h9D7: dout <= 8'b11111100; // 2519 : 252 - 0xfc
      12'h9D8: dout <= 8'b00000000; // 2520 :   0 - 0x0 -- plane 1
      12'h9D9: dout <= 8'b00000000; // 2521 :   0 - 0x0
      12'h9DA: dout <= 8'b00000000; // 2522 :   0 - 0x0
      12'h9DB: dout <= 8'b00000000; // 2523 :   0 - 0x0
      12'h9DC: dout <= 8'b00000000; // 2524 :   0 - 0x0
      12'h9DD: dout <= 8'b00000000; // 2525 :   0 - 0x0
      12'h9DE: dout <= 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout <= 8'b00111111; // 2528 :  63 - 0x3f -- Sprite 0x9e
      12'h9E1: dout <= 8'b00111111; // 2529 :  63 - 0x3f
      12'h9E2: dout <= 8'b00011111; // 2530 :  31 - 0x1f
      12'h9E3: dout <= 8'b00011111; // 2531 :  31 - 0x1f
      12'h9E4: dout <= 8'b00001111; // 2532 :  15 - 0xf
      12'h9E5: dout <= 8'b00000110; // 2533 :   6 - 0x6
      12'h9E6: dout <= 8'b00000000; // 2534 :   0 - 0x0
      12'h9E7: dout <= 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0 -- plane 1
      12'h9E9: dout <= 8'b00000000; // 2537 :   0 - 0x0
      12'h9EA: dout <= 8'b00000000; // 2538 :   0 - 0x0
      12'h9EB: dout <= 8'b00000000; // 2539 :   0 - 0x0
      12'h9EC: dout <= 8'b00000000; // 2540 :   0 - 0x0
      12'h9ED: dout <= 8'b00000000; // 2541 :   0 - 0x0
      12'h9EE: dout <= 8'b00000000; // 2542 :   0 - 0x0
      12'h9EF: dout <= 8'b00000000; // 2543 :   0 - 0x0
      12'h9F0: dout <= 8'b11101100; // 2544 : 236 - 0xec -- Sprite 0x9f
      12'h9F1: dout <= 8'b11101100; // 2545 : 236 - 0xec
      12'h9F2: dout <= 8'b11011000; // 2546 : 216 - 0xd8
      12'h9F3: dout <= 8'b11111000; // 2547 : 248 - 0xf8
      12'h9F4: dout <= 8'b11110000; // 2548 : 240 - 0xf0
      12'h9F5: dout <= 8'b11100000; // 2549 : 224 - 0xe0
      12'h9F6: dout <= 8'b00000000; // 2550 :   0 - 0x0
      12'h9F7: dout <= 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- plane 1
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout <= 8'b00000000; // 2560 :   0 - 0x0 -- Sprite 0xa0
      12'hA01: dout <= 8'b00000100; // 2561 :   4 - 0x4
      12'hA02: dout <= 8'b00000011; // 2562 :   3 - 0x3
      12'hA03: dout <= 8'b00000000; // 2563 :   0 - 0x0
      12'hA04: dout <= 8'b00000001; // 2564 :   1 - 0x1
      12'hA05: dout <= 8'b00000111; // 2565 :   7 - 0x7
      12'hA06: dout <= 8'b00001111; // 2566 :  15 - 0xf
      12'hA07: dout <= 8'b00001100; // 2567 :  12 - 0xc
      12'hA08: dout <= 8'b00000000; // 2568 :   0 - 0x0 -- plane 1
      12'hA09: dout <= 8'b00000000; // 2569 :   0 - 0x0
      12'hA0A: dout <= 8'b00000000; // 2570 :   0 - 0x0
      12'hA0B: dout <= 8'b00000000; // 2571 :   0 - 0x0
      12'hA0C: dout <= 8'b00000000; // 2572 :   0 - 0x0
      12'hA0D: dout <= 8'b00000000; // 2573 :   0 - 0x0
      12'hA0E: dout <= 8'b00000000; // 2574 :   0 - 0x0
      12'hA0F: dout <= 8'b00000000; // 2575 :   0 - 0x0
      12'hA10: dout <= 8'b00000000; // 2576 :   0 - 0x0 -- Sprite 0xa1
      12'hA11: dout <= 8'b00000000; // 2577 :   0 - 0x0
      12'hA12: dout <= 8'b11100000; // 2578 : 224 - 0xe0
      12'hA13: dout <= 8'b10000000; // 2579 : 128 - 0x80
      12'hA14: dout <= 8'b01000000; // 2580 :  64 - 0x40
      12'hA15: dout <= 8'b11110000; // 2581 : 240 - 0xf0
      12'hA16: dout <= 8'b10011000; // 2582 : 152 - 0x98
      12'hA17: dout <= 8'b11111000; // 2583 : 248 - 0xf8
      12'hA18: dout <= 8'b00000000; // 2584 :   0 - 0x0 -- plane 1
      12'hA19: dout <= 8'b00000000; // 2585 :   0 - 0x0
      12'hA1A: dout <= 8'b00000000; // 2586 :   0 - 0x0
      12'hA1B: dout <= 8'b00000000; // 2587 :   0 - 0x0
      12'hA1C: dout <= 8'b00000000; // 2588 :   0 - 0x0
      12'hA1D: dout <= 8'b00000000; // 2589 :   0 - 0x0
      12'hA1E: dout <= 8'b00000000; // 2590 :   0 - 0x0
      12'hA1F: dout <= 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout <= 8'b00011111; // 2592 :  31 - 0x1f -- Sprite 0xa2
      12'hA21: dout <= 8'b00010011; // 2593 :  19 - 0x13
      12'hA22: dout <= 8'b00011111; // 2594 :  31 - 0x1f
      12'hA23: dout <= 8'b00001111; // 2595 :  15 - 0xf
      12'hA24: dout <= 8'b00001001; // 2596 :   9 - 0x9
      12'hA25: dout <= 8'b00000111; // 2597 :   7 - 0x7
      12'hA26: dout <= 8'b00000001; // 2598 :   1 - 0x1
      12'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0 -- plane 1
      12'hA29: dout <= 8'b00000000; // 2601 :   0 - 0x0
      12'hA2A: dout <= 8'b00000000; // 2602 :   0 - 0x0
      12'hA2B: dout <= 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout <= 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout <= 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout <= 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout <= 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout <= 8'b11100100; // 2608 : 228 - 0xe4 -- Sprite 0xa3
      12'hA31: dout <= 8'b00111100; // 2609 :  60 - 0x3c
      12'hA32: dout <= 8'b11100100; // 2610 : 228 - 0xe4
      12'hA33: dout <= 8'b00111000; // 2611 :  56 - 0x38
      12'hA34: dout <= 8'b11111000; // 2612 : 248 - 0xf8
      12'hA35: dout <= 8'b11110000; // 2613 : 240 - 0xf0
      12'hA36: dout <= 8'b11000000; // 2614 : 192 - 0xc0
      12'hA37: dout <= 8'b00000000; // 2615 :   0 - 0x0
      12'hA38: dout <= 8'b00000000; // 2616 :   0 - 0x0 -- plane 1
      12'hA39: dout <= 8'b00000000; // 2617 :   0 - 0x0
      12'hA3A: dout <= 8'b00000000; // 2618 :   0 - 0x0
      12'hA3B: dout <= 8'b00000000; // 2619 :   0 - 0x0
      12'hA3C: dout <= 8'b00000000; // 2620 :   0 - 0x0
      12'hA3D: dout <= 8'b00000000; // 2621 :   0 - 0x0
      12'hA3E: dout <= 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout <= 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout <= 8'b00000000; // 2624 :   0 - 0x0 -- Sprite 0xa4
      12'hA41: dout <= 8'b00000000; // 2625 :   0 - 0x0
      12'hA42: dout <= 8'b00000000; // 2626 :   0 - 0x0
      12'hA43: dout <= 8'b00000000; // 2627 :   0 - 0x0
      12'hA44: dout <= 8'b00010001; // 2628 :  17 - 0x11
      12'hA45: dout <= 8'b00010011; // 2629 :  19 - 0x13
      12'hA46: dout <= 8'b00011111; // 2630 :  31 - 0x1f
      12'hA47: dout <= 8'b00011111; // 2631 :  31 - 0x1f
      12'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0 -- plane 1
      12'hA49: dout <= 8'b00000000; // 2633 :   0 - 0x0
      12'hA4A: dout <= 8'b00000000; // 2634 :   0 - 0x0
      12'hA4B: dout <= 8'b00000000; // 2635 :   0 - 0x0
      12'hA4C: dout <= 8'b00000000; // 2636 :   0 - 0x0
      12'hA4D: dout <= 8'b00000000; // 2637 :   0 - 0x0
      12'hA4E: dout <= 8'b00000000; // 2638 :   0 - 0x0
      12'hA4F: dout <= 8'b00000000; // 2639 :   0 - 0x0
      12'hA50: dout <= 8'b00000000; // 2640 :   0 - 0x0 -- Sprite 0xa5
      12'hA51: dout <= 8'b00000000; // 2641 :   0 - 0x0
      12'hA52: dout <= 8'b00000000; // 2642 :   0 - 0x0
      12'hA53: dout <= 8'b10000000; // 2643 : 128 - 0x80
      12'hA54: dout <= 8'b11000100; // 2644 : 196 - 0xc4
      12'hA55: dout <= 8'b11100100; // 2645 : 228 - 0xe4
      12'hA56: dout <= 8'b11111100; // 2646 : 252 - 0xfc
      12'hA57: dout <= 8'b11111100; // 2647 : 252 - 0xfc
      12'hA58: dout <= 8'b00000000; // 2648 :   0 - 0x0 -- plane 1
      12'hA59: dout <= 8'b00000000; // 2649 :   0 - 0x0
      12'hA5A: dout <= 8'b00000000; // 2650 :   0 - 0x0
      12'hA5B: dout <= 8'b00000000; // 2651 :   0 - 0x0
      12'hA5C: dout <= 8'b00000000; // 2652 :   0 - 0x0
      12'hA5D: dout <= 8'b00000000; // 2653 :   0 - 0x0
      12'hA5E: dout <= 8'b00000000; // 2654 :   0 - 0x0
      12'hA5F: dout <= 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout <= 8'b00011111; // 2656 :  31 - 0x1f -- Sprite 0xa6
      12'hA61: dout <= 8'b00001110; // 2657 :  14 - 0xe
      12'hA62: dout <= 8'b00000110; // 2658 :   6 - 0x6
      12'hA63: dout <= 8'b00000010; // 2659 :   2 - 0x2
      12'hA64: dout <= 8'b00000000; // 2660 :   0 - 0x0
      12'hA65: dout <= 8'b00000000; // 2661 :   0 - 0x0
      12'hA66: dout <= 8'b00000000; // 2662 :   0 - 0x0
      12'hA67: dout <= 8'b00000000; // 2663 :   0 - 0x0
      12'hA68: dout <= 8'b00000000; // 2664 :   0 - 0x0 -- plane 1
      12'hA69: dout <= 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout <= 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout <= 8'b00000000; // 2667 :   0 - 0x0
      12'hA6C: dout <= 8'b00000000; // 2668 :   0 - 0x0
      12'hA6D: dout <= 8'b00000000; // 2669 :   0 - 0x0
      12'hA6E: dout <= 8'b00000000; // 2670 :   0 - 0x0
      12'hA6F: dout <= 8'b00000000; // 2671 :   0 - 0x0
      12'hA70: dout <= 8'b11111100; // 2672 : 252 - 0xfc -- Sprite 0xa7
      12'hA71: dout <= 8'b10111000; // 2673 : 184 - 0xb8
      12'hA72: dout <= 8'b10110000; // 2674 : 176 - 0xb0
      12'hA73: dout <= 8'b10100000; // 2675 : 160 - 0xa0
      12'hA74: dout <= 8'b10000000; // 2676 : 128 - 0x80
      12'hA75: dout <= 8'b00000000; // 2677 :   0 - 0x0
      12'hA76: dout <= 8'b00000000; // 2678 :   0 - 0x0
      12'hA77: dout <= 8'b00000000; // 2679 :   0 - 0x0
      12'hA78: dout <= 8'b00000000; // 2680 :   0 - 0x0 -- plane 1
      12'hA79: dout <= 8'b00000000; // 2681 :   0 - 0x0
      12'hA7A: dout <= 8'b00000000; // 2682 :   0 - 0x0
      12'hA7B: dout <= 8'b00000000; // 2683 :   0 - 0x0
      12'hA7C: dout <= 8'b00000000; // 2684 :   0 - 0x0
      12'hA7D: dout <= 8'b00000000; // 2685 :   0 - 0x0
      12'hA7E: dout <= 8'b00000000; // 2686 :   0 - 0x0
      12'hA7F: dout <= 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout <= 8'b00000000; // 2688 :   0 - 0x0 -- Sprite 0xa8
      12'hA81: dout <= 8'b00000000; // 2689 :   0 - 0x0
      12'hA82: dout <= 8'b00000000; // 2690 :   0 - 0x0
      12'hA83: dout <= 8'b00000001; // 2691 :   1 - 0x1
      12'hA84: dout <= 8'b00000011; // 2692 :   3 - 0x3
      12'hA85: dout <= 8'b00000110; // 2693 :   6 - 0x6
      12'hA86: dout <= 8'b00000110; // 2694 :   6 - 0x6
      12'hA87: dout <= 8'b00001111; // 2695 :  15 - 0xf
      12'hA88: dout <= 8'b00000000; // 2696 :   0 - 0x0 -- plane 1
      12'hA89: dout <= 8'b00000000; // 2697 :   0 - 0x0
      12'hA8A: dout <= 8'b00000000; // 2698 :   0 - 0x0
      12'hA8B: dout <= 8'b00000000; // 2699 :   0 - 0x0
      12'hA8C: dout <= 8'b00000000; // 2700 :   0 - 0x0
      12'hA8D: dout <= 8'b00000000; // 2701 :   0 - 0x0
      12'hA8E: dout <= 8'b00000000; // 2702 :   0 - 0x0
      12'hA8F: dout <= 8'b00000000; // 2703 :   0 - 0x0
      12'hA90: dout <= 8'b00000000; // 2704 :   0 - 0x0 -- Sprite 0xa9
      12'hA91: dout <= 8'b00011000; // 2705 :  24 - 0x18
      12'hA92: dout <= 8'b11110100; // 2706 : 244 - 0xf4
      12'hA93: dout <= 8'b11111000; // 2707 : 248 - 0xf8
      12'hA94: dout <= 8'b00111000; // 2708 :  56 - 0x38
      12'hA95: dout <= 8'b01111100; // 2709 : 124 - 0x7c
      12'hA96: dout <= 8'b11111100; // 2710 : 252 - 0xfc
      12'hA97: dout <= 8'b11111100; // 2711 : 252 - 0xfc
      12'hA98: dout <= 8'b00000000; // 2712 :   0 - 0x0 -- plane 1
      12'hA99: dout <= 8'b00000000; // 2713 :   0 - 0x0
      12'hA9A: dout <= 8'b00000000; // 2714 :   0 - 0x0
      12'hA9B: dout <= 8'b00000000; // 2715 :   0 - 0x0
      12'hA9C: dout <= 8'b00000000; // 2716 :   0 - 0x0
      12'hA9D: dout <= 8'b00000000; // 2717 :   0 - 0x0
      12'hA9E: dout <= 8'b00000000; // 2718 :   0 - 0x0
      12'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout <= 8'b00001111; // 2720 :  15 - 0xf -- Sprite 0xaa
      12'hAA1: dout <= 8'b00011111; // 2721 :  31 - 0x1f
      12'hAA2: dout <= 8'b00110000; // 2722 :  48 - 0x30
      12'hAA3: dout <= 8'b00111000; // 2723 :  56 - 0x38
      12'hAA4: dout <= 8'b00011101; // 2724 :  29 - 0x1d
      12'hAA5: dout <= 8'b00000011; // 2725 :   3 - 0x3
      12'hAA6: dout <= 8'b00000011; // 2726 :   3 - 0x3
      12'hAA7: dout <= 8'b00000000; // 2727 :   0 - 0x0
      12'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0 -- plane 1
      12'hAA9: dout <= 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout <= 8'b00000000; // 2730 :   0 - 0x0
      12'hAAB: dout <= 8'b00000000; // 2731 :   0 - 0x0
      12'hAAC: dout <= 8'b00000000; // 2732 :   0 - 0x0
      12'hAAD: dout <= 8'b00000000; // 2733 :   0 - 0x0
      12'hAAE: dout <= 8'b00000000; // 2734 :   0 - 0x0
      12'hAAF: dout <= 8'b00000000; // 2735 :   0 - 0x0
      12'hAB0: dout <= 8'b11111100; // 2736 : 252 - 0xfc -- Sprite 0xab
      12'hAB1: dout <= 8'b11111100; // 2737 : 252 - 0xfc
      12'hAB2: dout <= 8'b01111100; // 2738 : 124 - 0x7c
      12'hAB3: dout <= 8'b10001110; // 2739 : 142 - 0x8e
      12'hAB4: dout <= 8'b10000110; // 2740 : 134 - 0x86
      12'hAB5: dout <= 8'b10011100; // 2741 : 156 - 0x9c
      12'hAB6: dout <= 8'b01111000; // 2742 : 120 - 0x78
      12'hAB7: dout <= 8'b00000000; // 2743 :   0 - 0x0
      12'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0 -- plane 1
      12'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout <= 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout <= 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout <= 8'b00000000; // 2752 :   0 - 0x0 -- Sprite 0xac
      12'hAC1: dout <= 8'b00000001; // 2753 :   1 - 0x1
      12'hAC2: dout <= 8'b00000110; // 2754 :   6 - 0x6
      12'hAC3: dout <= 8'b00000111; // 2755 :   7 - 0x7
      12'hAC4: dout <= 8'b00000111; // 2756 :   7 - 0x7
      12'hAC5: dout <= 8'b00000111; // 2757 :   7 - 0x7
      12'hAC6: dout <= 8'b00000001; // 2758 :   1 - 0x1
      12'hAC7: dout <= 8'b00000011; // 2759 :   3 - 0x3
      12'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0 -- plane 1
      12'hAC9: dout <= 8'b00000000; // 2761 :   0 - 0x0
      12'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout <= 8'b00000000; // 2763 :   0 - 0x0
      12'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      12'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout <= 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout <= 8'b00000000; // 2768 :   0 - 0x0 -- Sprite 0xad
      12'hAD1: dout <= 8'b11000000; // 2769 : 192 - 0xc0
      12'hAD2: dout <= 8'b00110000; // 2770 :  48 - 0x30
      12'hAD3: dout <= 8'b11110000; // 2771 : 240 - 0xf0
      12'hAD4: dout <= 8'b11110000; // 2772 : 240 - 0xf0
      12'hAD5: dout <= 8'b11110000; // 2773 : 240 - 0xf0
      12'hAD6: dout <= 8'b01000000; // 2774 :  64 - 0x40
      12'hAD7: dout <= 8'b01000000; // 2775 :  64 - 0x40
      12'hAD8: dout <= 8'b00000000; // 2776 :   0 - 0x0 -- plane 1
      12'hAD9: dout <= 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout <= 8'b00000000; // 2778 :   0 - 0x0
      12'hADB: dout <= 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout <= 8'b00000000; // 2780 :   0 - 0x0
      12'hADD: dout <= 8'b00000000; // 2781 :   0 - 0x0
      12'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      12'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout <= 8'b00000001; // 2784 :   1 - 0x1 -- Sprite 0xae
      12'hAE1: dout <= 8'b00000000; // 2785 :   0 - 0x0
      12'hAE2: dout <= 8'b00000001; // 2786 :   1 - 0x1
      12'hAE3: dout <= 8'b00000011; // 2787 :   3 - 0x3
      12'hAE4: dout <= 8'b00000001; // 2788 :   1 - 0x1
      12'hAE5: dout <= 8'b00000000; // 2789 :   0 - 0x0
      12'hAE6: dout <= 8'b00000000; // 2790 :   0 - 0x0
      12'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0 -- plane 1
      12'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout <= 8'b00000000; // 2794 :   0 - 0x0
      12'hAEB: dout <= 8'b00000000; // 2795 :   0 - 0x0
      12'hAEC: dout <= 8'b00000000; // 2796 :   0 - 0x0
      12'hAED: dout <= 8'b00000000; // 2797 :   0 - 0x0
      12'hAEE: dout <= 8'b00000000; // 2798 :   0 - 0x0
      12'hAEF: dout <= 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout <= 8'b01000000; // 2800 :  64 - 0x40 -- Sprite 0xaf
      12'hAF1: dout <= 8'b01000000; // 2801 :  64 - 0x40
      12'hAF2: dout <= 8'b01000000; // 2802 :  64 - 0x40
      12'hAF3: dout <= 8'b01000000; // 2803 :  64 - 0x40
      12'hAF4: dout <= 8'b01000000; // 2804 :  64 - 0x40
      12'hAF5: dout <= 8'b10000000; // 2805 : 128 - 0x80
      12'hAF6: dout <= 8'b00000000; // 2806 :   0 - 0x0
      12'hAF7: dout <= 8'b00000000; // 2807 :   0 - 0x0
      12'hAF8: dout <= 8'b00000000; // 2808 :   0 - 0x0 -- plane 1
      12'hAF9: dout <= 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout <= 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout <= 8'b00000000; // 2811 :   0 - 0x0
      12'hAFC: dout <= 8'b00000000; // 2812 :   0 - 0x0
      12'hAFD: dout <= 8'b00000000; // 2813 :   0 - 0x0
      12'hAFE: dout <= 8'b00000000; // 2814 :   0 - 0x0
      12'hAFF: dout <= 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout <= 8'b01111110; // 2816 : 126 - 0x7e -- Sprite 0xb0
      12'hB01: dout <= 8'b01100011; // 2817 :  99 - 0x63
      12'hB02: dout <= 8'b01100011; // 2818 :  99 - 0x63
      12'hB03: dout <= 8'b01100011; // 2819 :  99 - 0x63
      12'hB04: dout <= 8'b01111110; // 2820 : 126 - 0x7e
      12'hB05: dout <= 8'b01100000; // 2821 :  96 - 0x60
      12'hB06: dout <= 8'b01100000; // 2822 :  96 - 0x60
      12'hB07: dout <= 8'b00000000; // 2823 :   0 - 0x0
      12'hB08: dout <= 8'b01111110; // 2824 : 126 - 0x7e -- plane 1
      12'hB09: dout <= 8'b01100011; // 2825 :  99 - 0x63
      12'hB0A: dout <= 8'b01100011; // 2826 :  99 - 0x63
      12'hB0B: dout <= 8'b01100011; // 2827 :  99 - 0x63
      12'hB0C: dout <= 8'b01111110; // 2828 : 126 - 0x7e
      12'hB0D: dout <= 8'b01100000; // 2829 :  96 - 0x60
      12'hB0E: dout <= 8'b01100000; // 2830 :  96 - 0x60
      12'hB0F: dout <= 8'b00000000; // 2831 :   0 - 0x0
      12'hB10: dout <= 8'b01100000; // 2832 :  96 - 0x60 -- Sprite 0xb1
      12'hB11: dout <= 8'b01100000; // 2833 :  96 - 0x60
      12'hB12: dout <= 8'b01100000; // 2834 :  96 - 0x60
      12'hB13: dout <= 8'b01100000; // 2835 :  96 - 0x60
      12'hB14: dout <= 8'b01100000; // 2836 :  96 - 0x60
      12'hB15: dout <= 8'b01100000; // 2837 :  96 - 0x60
      12'hB16: dout <= 8'b01111111; // 2838 : 127 - 0x7f
      12'hB17: dout <= 8'b00000000; // 2839 :   0 - 0x0
      12'hB18: dout <= 8'b01100000; // 2840 :  96 - 0x60 -- plane 1
      12'hB19: dout <= 8'b01100000; // 2841 :  96 - 0x60
      12'hB1A: dout <= 8'b01100000; // 2842 :  96 - 0x60
      12'hB1B: dout <= 8'b01100000; // 2843 :  96 - 0x60
      12'hB1C: dout <= 8'b01100000; // 2844 :  96 - 0x60
      12'hB1D: dout <= 8'b01100000; // 2845 :  96 - 0x60
      12'hB1E: dout <= 8'b01111111; // 2846 : 127 - 0x7f
      12'hB1F: dout <= 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout <= 8'b00011100; // 2848 :  28 - 0x1c -- Sprite 0xb2
      12'hB21: dout <= 8'b00110110; // 2849 :  54 - 0x36
      12'hB22: dout <= 8'b01100011; // 2850 :  99 - 0x63
      12'hB23: dout <= 8'b01100011; // 2851 :  99 - 0x63
      12'hB24: dout <= 8'b01111111; // 2852 : 127 - 0x7f
      12'hB25: dout <= 8'b01100011; // 2853 :  99 - 0x63
      12'hB26: dout <= 8'b01100011; // 2854 :  99 - 0x63
      12'hB27: dout <= 8'b00000000; // 2855 :   0 - 0x0
      12'hB28: dout <= 8'b00011100; // 2856 :  28 - 0x1c -- plane 1
      12'hB29: dout <= 8'b00110110; // 2857 :  54 - 0x36
      12'hB2A: dout <= 8'b01100011; // 2858 :  99 - 0x63
      12'hB2B: dout <= 8'b01100011; // 2859 :  99 - 0x63
      12'hB2C: dout <= 8'b01111111; // 2860 : 127 - 0x7f
      12'hB2D: dout <= 8'b01100011; // 2861 :  99 - 0x63
      12'hB2E: dout <= 8'b01100011; // 2862 :  99 - 0x63
      12'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout <= 8'b00110011; // 2864 :  51 - 0x33 -- Sprite 0xb3
      12'hB31: dout <= 8'b00110011; // 2865 :  51 - 0x33
      12'hB32: dout <= 8'b00110011; // 2866 :  51 - 0x33
      12'hB33: dout <= 8'b00011110; // 2867 :  30 - 0x1e
      12'hB34: dout <= 8'b00001100; // 2868 :  12 - 0xc
      12'hB35: dout <= 8'b00001100; // 2869 :  12 - 0xc
      12'hB36: dout <= 8'b00001100; // 2870 :  12 - 0xc
      12'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      12'hB38: dout <= 8'b00110011; // 2872 :  51 - 0x33 -- plane 1
      12'hB39: dout <= 8'b00110011; // 2873 :  51 - 0x33
      12'hB3A: dout <= 8'b00110011; // 2874 :  51 - 0x33
      12'hB3B: dout <= 8'b00011110; // 2875 :  30 - 0x1e
      12'hB3C: dout <= 8'b00001100; // 2876 :  12 - 0xc
      12'hB3D: dout <= 8'b00001100; // 2877 :  12 - 0xc
      12'hB3E: dout <= 8'b00001100; // 2878 :  12 - 0xc
      12'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout <= 8'b01111111; // 2880 : 127 - 0x7f -- Sprite 0xb4
      12'hB41: dout <= 8'b01100000; // 2881 :  96 - 0x60
      12'hB42: dout <= 8'b01100000; // 2882 :  96 - 0x60
      12'hB43: dout <= 8'b01111110; // 2883 : 126 - 0x7e
      12'hB44: dout <= 8'b01100000; // 2884 :  96 - 0x60
      12'hB45: dout <= 8'b01100000; // 2885 :  96 - 0x60
      12'hB46: dout <= 8'b01111111; // 2886 : 127 - 0x7f
      12'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout <= 8'b01111111; // 2888 : 127 - 0x7f -- plane 1
      12'hB49: dout <= 8'b01100000; // 2889 :  96 - 0x60
      12'hB4A: dout <= 8'b01100000; // 2890 :  96 - 0x60
      12'hB4B: dout <= 8'b01111110; // 2891 : 126 - 0x7e
      12'hB4C: dout <= 8'b01100000; // 2892 :  96 - 0x60
      12'hB4D: dout <= 8'b01100000; // 2893 :  96 - 0x60
      12'hB4E: dout <= 8'b01111111; // 2894 : 127 - 0x7f
      12'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout <= 8'b01111110; // 2896 : 126 - 0x7e -- Sprite 0xb5
      12'hB51: dout <= 8'b01100011; // 2897 :  99 - 0x63
      12'hB52: dout <= 8'b01100011; // 2898 :  99 - 0x63
      12'hB53: dout <= 8'b01100111; // 2899 : 103 - 0x67
      12'hB54: dout <= 8'b01111100; // 2900 : 124 - 0x7c
      12'hB55: dout <= 8'b01101110; // 2901 : 110 - 0x6e
      12'hB56: dout <= 8'b01100111; // 2902 : 103 - 0x67
      12'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout <= 8'b01111110; // 2904 : 126 - 0x7e -- plane 1
      12'hB59: dout <= 8'b01100011; // 2905 :  99 - 0x63
      12'hB5A: dout <= 8'b01100011; // 2906 :  99 - 0x63
      12'hB5B: dout <= 8'b01100111; // 2907 : 103 - 0x67
      12'hB5C: dout <= 8'b01111100; // 2908 : 124 - 0x7c
      12'hB5D: dout <= 8'b01101110; // 2909 : 110 - 0x6e
      12'hB5E: dout <= 8'b01100111; // 2910 : 103 - 0x67
      12'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout <= 8'b00111110; // 2912 :  62 - 0x3e -- Sprite 0xb6
      12'hB61: dout <= 8'b01100011; // 2913 :  99 - 0x63
      12'hB62: dout <= 8'b01100011; // 2914 :  99 - 0x63
      12'hB63: dout <= 8'b01100011; // 2915 :  99 - 0x63
      12'hB64: dout <= 8'b01100011; // 2916 :  99 - 0x63
      12'hB65: dout <= 8'b01100011; // 2917 :  99 - 0x63
      12'hB66: dout <= 8'b00111110; // 2918 :  62 - 0x3e
      12'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout <= 8'b00111110; // 2920 :  62 - 0x3e -- plane 1
      12'hB69: dout <= 8'b01100011; // 2921 :  99 - 0x63
      12'hB6A: dout <= 8'b01100011; // 2922 :  99 - 0x63
      12'hB6B: dout <= 8'b01100011; // 2923 :  99 - 0x63
      12'hB6C: dout <= 8'b01100011; // 2924 :  99 - 0x63
      12'hB6D: dout <= 8'b01100011; // 2925 :  99 - 0x63
      12'hB6E: dout <= 8'b00111110; // 2926 :  62 - 0x3e
      12'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout <= 8'b01100011; // 2928 :  99 - 0x63 -- Sprite 0xb7
      12'hB71: dout <= 8'b01110011; // 2929 : 115 - 0x73
      12'hB72: dout <= 8'b01111011; // 2930 : 123 - 0x7b
      12'hB73: dout <= 8'b01111111; // 2931 : 127 - 0x7f
      12'hB74: dout <= 8'b01101111; // 2932 : 111 - 0x6f
      12'hB75: dout <= 8'b01100111; // 2933 : 103 - 0x67
      12'hB76: dout <= 8'b01100011; // 2934 :  99 - 0x63
      12'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout <= 8'b01100011; // 2936 :  99 - 0x63 -- plane 1
      12'hB79: dout <= 8'b01110011; // 2937 : 115 - 0x73
      12'hB7A: dout <= 8'b01111011; // 2938 : 123 - 0x7b
      12'hB7B: dout <= 8'b01111111; // 2939 : 127 - 0x7f
      12'hB7C: dout <= 8'b01101111; // 2940 : 111 - 0x6f
      12'hB7D: dout <= 8'b01100111; // 2941 : 103 - 0x67
      12'hB7E: dout <= 8'b01100011; // 2942 :  99 - 0x63
      12'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout <= 8'b00111111; // 2944 :  63 - 0x3f -- Sprite 0xb8
      12'hB81: dout <= 8'b00001100; // 2945 :  12 - 0xc
      12'hB82: dout <= 8'b00001100; // 2946 :  12 - 0xc
      12'hB83: dout <= 8'b00001100; // 2947 :  12 - 0xc
      12'hB84: dout <= 8'b00001100; // 2948 :  12 - 0xc
      12'hB85: dout <= 8'b00001100; // 2949 :  12 - 0xc
      12'hB86: dout <= 8'b00001100; // 2950 :  12 - 0xc
      12'hB87: dout <= 8'b00000000; // 2951 :   0 - 0x0
      12'hB88: dout <= 8'b00111111; // 2952 :  63 - 0x3f -- plane 1
      12'hB89: dout <= 8'b00001100; // 2953 :  12 - 0xc
      12'hB8A: dout <= 8'b00001100; // 2954 :  12 - 0xc
      12'hB8B: dout <= 8'b00001100; // 2955 :  12 - 0xc
      12'hB8C: dout <= 8'b00001100; // 2956 :  12 - 0xc
      12'hB8D: dout <= 8'b00001100; // 2957 :  12 - 0xc
      12'hB8E: dout <= 8'b00001100; // 2958 :  12 - 0xc
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b01100011; // 2960 :  99 - 0x63 -- Sprite 0xb9
      12'hB91: dout <= 8'b01100011; // 2961 :  99 - 0x63
      12'hB92: dout <= 8'b01101011; // 2962 : 107 - 0x6b
      12'hB93: dout <= 8'b01111111; // 2963 : 127 - 0x7f
      12'hB94: dout <= 8'b01111111; // 2964 : 127 - 0x7f
      12'hB95: dout <= 8'b01110111; // 2965 : 119 - 0x77
      12'hB96: dout <= 8'b01100011; // 2966 :  99 - 0x63
      12'hB97: dout <= 8'b00000000; // 2967 :   0 - 0x0
      12'hB98: dout <= 8'b01100011; // 2968 :  99 - 0x63 -- plane 1
      12'hB99: dout <= 8'b01100011; // 2969 :  99 - 0x63
      12'hB9A: dout <= 8'b01101011; // 2970 : 107 - 0x6b
      12'hB9B: dout <= 8'b01111111; // 2971 : 127 - 0x7f
      12'hB9C: dout <= 8'b01111111; // 2972 : 127 - 0x7f
      12'hB9D: dout <= 8'b01110111; // 2973 : 119 - 0x77
      12'hB9E: dout <= 8'b01100011; // 2974 :  99 - 0x63
      12'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout <= 8'b01111100; // 2976 : 124 - 0x7c -- Sprite 0xba
      12'hBA1: dout <= 8'b01100110; // 2977 : 102 - 0x66
      12'hBA2: dout <= 8'b01100011; // 2978 :  99 - 0x63
      12'hBA3: dout <= 8'b01100011; // 2979 :  99 - 0x63
      12'hBA4: dout <= 8'b01100011; // 2980 :  99 - 0x63
      12'hBA5: dout <= 8'b01100110; // 2981 : 102 - 0x66
      12'hBA6: dout <= 8'b01111100; // 2982 : 124 - 0x7c
      12'hBA7: dout <= 8'b00000000; // 2983 :   0 - 0x0
      12'hBA8: dout <= 8'b00000000; // 2984 :   0 - 0x0 -- plane 1
      12'hBA9: dout <= 8'b00000000; // 2985 :   0 - 0x0
      12'hBAA: dout <= 8'b00000000; // 2986 :   0 - 0x0
      12'hBAB: dout <= 8'b00000000; // 2987 :   0 - 0x0
      12'hBAC: dout <= 8'b00000000; // 2988 :   0 - 0x0
      12'hBAD: dout <= 8'b00000000; // 2989 :   0 - 0x0
      12'hBAE: dout <= 8'b00000000; // 2990 :   0 - 0x0
      12'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout <= 8'b00011100; // 2992 :  28 - 0x1c -- Sprite 0xbb
      12'hBB1: dout <= 8'b00011100; // 2993 :  28 - 0x1c
      12'hBB2: dout <= 8'b00011100; // 2994 :  28 - 0x1c
      12'hBB3: dout <= 8'b00011000; // 2995 :  24 - 0x18
      12'hBB4: dout <= 8'b00011000; // 2996 :  24 - 0x18
      12'hBB5: dout <= 8'b00000000; // 2997 :   0 - 0x0
      12'hBB6: dout <= 8'b00011000; // 2998 :  24 - 0x18
      12'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0 -- plane 1
      12'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      12'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      12'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      12'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      12'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b00011111; // 3008 :  31 - 0x1f -- Sprite 0xbc
      12'hBC1: dout <= 8'b00110000; // 3009 :  48 - 0x30
      12'hBC2: dout <= 8'b01100000; // 3010 :  96 - 0x60
      12'hBC3: dout <= 8'b01100111; // 3011 : 103 - 0x67
      12'hBC4: dout <= 8'b01100011; // 3012 :  99 - 0x63
      12'hBC5: dout <= 8'b00110011; // 3013 :  51 - 0x33
      12'hBC6: dout <= 8'b00011111; // 3014 :  31 - 0x1f
      12'hBC7: dout <= 8'b00000000; // 3015 :   0 - 0x0
      12'hBC8: dout <= 8'b00011111; // 3016 :  31 - 0x1f -- plane 1
      12'hBC9: dout <= 8'b00110000; // 3017 :  48 - 0x30
      12'hBCA: dout <= 8'b01100000; // 3018 :  96 - 0x60
      12'hBCB: dout <= 8'b01100111; // 3019 : 103 - 0x67
      12'hBCC: dout <= 8'b01100011; // 3020 :  99 - 0x63
      12'hBCD: dout <= 8'b00110011; // 3021 :  51 - 0x33
      12'hBCE: dout <= 8'b00011111; // 3022 :  31 - 0x1f
      12'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout <= 8'b01100011; // 3024 :  99 - 0x63 -- Sprite 0xbd
      12'hBD1: dout <= 8'b01110111; // 3025 : 119 - 0x77
      12'hBD2: dout <= 8'b01111111; // 3026 : 127 - 0x7f
      12'hBD3: dout <= 8'b01111111; // 3027 : 127 - 0x7f
      12'hBD4: dout <= 8'b01101011; // 3028 : 107 - 0x6b
      12'hBD5: dout <= 8'b01100011; // 3029 :  99 - 0x63
      12'hBD6: dout <= 8'b01100011; // 3030 :  99 - 0x63
      12'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout <= 8'b01100011; // 3032 :  99 - 0x63 -- plane 1
      12'hBD9: dout <= 8'b01110111; // 3033 : 119 - 0x77
      12'hBDA: dout <= 8'b01111111; // 3034 : 127 - 0x7f
      12'hBDB: dout <= 8'b01111111; // 3035 : 127 - 0x7f
      12'hBDC: dout <= 8'b01101011; // 3036 : 107 - 0x6b
      12'hBDD: dout <= 8'b01100011; // 3037 :  99 - 0x63
      12'hBDE: dout <= 8'b01100011; // 3038 :  99 - 0x63
      12'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout <= 8'b01100011; // 3040 :  99 - 0x63 -- Sprite 0xbe
      12'hBE1: dout <= 8'b01100011; // 3041 :  99 - 0x63
      12'hBE2: dout <= 8'b01100011; // 3042 :  99 - 0x63
      12'hBE3: dout <= 8'b01110111; // 3043 : 119 - 0x77
      12'hBE4: dout <= 8'b00111110; // 3044 :  62 - 0x3e
      12'hBE5: dout <= 8'b00011100; // 3045 :  28 - 0x1c
      12'hBE6: dout <= 8'b00001000; // 3046 :   8 - 0x8
      12'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      12'hBE8: dout <= 8'b01100011; // 3048 :  99 - 0x63 -- plane 1
      12'hBE9: dout <= 8'b01100011; // 3049 :  99 - 0x63
      12'hBEA: dout <= 8'b01100011; // 3050 :  99 - 0x63
      12'hBEB: dout <= 8'b01110111; // 3051 : 119 - 0x77
      12'hBEC: dout <= 8'b00111110; // 3052 :  62 - 0x3e
      12'hBED: dout <= 8'b00011100; // 3053 :  28 - 0x1c
      12'hBEE: dout <= 8'b00001000; // 3054 :   8 - 0x8
      12'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Sprite 0xbf
      12'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      12'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      12'hBF4: dout <= 8'b00000000; // 3060 :   0 - 0x0
      12'hBF5: dout <= 8'b00000000; // 3061 :   0 - 0x0
      12'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      12'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0 -- plane 1
      12'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      12'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      12'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      12'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout <= 8'b00011111; // 3072 :  31 - 0x1f -- Sprite 0xc0
      12'hC01: dout <= 8'b00110000; // 3073 :  48 - 0x30
      12'hC02: dout <= 8'b01100000; // 3074 :  96 - 0x60
      12'hC03: dout <= 8'b01100111; // 3075 : 103 - 0x67
      12'hC04: dout <= 8'b01100011; // 3076 :  99 - 0x63
      12'hC05: dout <= 8'b00110011; // 3077 :  51 - 0x33
      12'hC06: dout <= 8'b00011111; // 3078 :  31 - 0x1f
      12'hC07: dout <= 8'b00000000; // 3079 :   0 - 0x0
      12'hC08: dout <= 8'b00000000; // 3080 :   0 - 0x0 -- plane 1
      12'hC09: dout <= 8'b00000000; // 3081 :   0 - 0x0
      12'hC0A: dout <= 8'b00000000; // 3082 :   0 - 0x0
      12'hC0B: dout <= 8'b00000000; // 3083 :   0 - 0x0
      12'hC0C: dout <= 8'b00000000; // 3084 :   0 - 0x0
      12'hC0D: dout <= 8'b00000000; // 3085 :   0 - 0x0
      12'hC0E: dout <= 8'b00000000; // 3086 :   0 - 0x0
      12'hC0F: dout <= 8'b00000000; // 3087 :   0 - 0x0
      12'hC10: dout <= 8'b00011100; // 3088 :  28 - 0x1c -- Sprite 0xc1
      12'hC11: dout <= 8'b00110110; // 3089 :  54 - 0x36
      12'hC12: dout <= 8'b01100011; // 3090 :  99 - 0x63
      12'hC13: dout <= 8'b01100011; // 3091 :  99 - 0x63
      12'hC14: dout <= 8'b01111111; // 3092 : 127 - 0x7f
      12'hC15: dout <= 8'b01100011; // 3093 :  99 - 0x63
      12'hC16: dout <= 8'b01100011; // 3094 :  99 - 0x63
      12'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      12'hC18: dout <= 8'b00000000; // 3096 :   0 - 0x0 -- plane 1
      12'hC19: dout <= 8'b00000000; // 3097 :   0 - 0x0
      12'hC1A: dout <= 8'b00000000; // 3098 :   0 - 0x0
      12'hC1B: dout <= 8'b00000000; // 3099 :   0 - 0x0
      12'hC1C: dout <= 8'b00000000; // 3100 :   0 - 0x0
      12'hC1D: dout <= 8'b00000000; // 3101 :   0 - 0x0
      12'hC1E: dout <= 8'b00000000; // 3102 :   0 - 0x0
      12'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout <= 8'b01100011; // 3104 :  99 - 0x63 -- Sprite 0xc2
      12'hC21: dout <= 8'b01110111; // 3105 : 119 - 0x77
      12'hC22: dout <= 8'b01111111; // 3106 : 127 - 0x7f
      12'hC23: dout <= 8'b01111111; // 3107 : 127 - 0x7f
      12'hC24: dout <= 8'b01101011; // 3108 : 107 - 0x6b
      12'hC25: dout <= 8'b01100011; // 3109 :  99 - 0x63
      12'hC26: dout <= 8'b01100011; // 3110 :  99 - 0x63
      12'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      12'hC28: dout <= 8'b00000000; // 3112 :   0 - 0x0 -- plane 1
      12'hC29: dout <= 8'b00000000; // 3113 :   0 - 0x0
      12'hC2A: dout <= 8'b00000000; // 3114 :   0 - 0x0
      12'hC2B: dout <= 8'b00000000; // 3115 :   0 - 0x0
      12'hC2C: dout <= 8'b00000000; // 3116 :   0 - 0x0
      12'hC2D: dout <= 8'b00000000; // 3117 :   0 - 0x0
      12'hC2E: dout <= 8'b00000000; // 3118 :   0 - 0x0
      12'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      12'hC30: dout <= 8'b01111111; // 3120 : 127 - 0x7f -- Sprite 0xc3
      12'hC31: dout <= 8'b01100000; // 3121 :  96 - 0x60
      12'hC32: dout <= 8'b01100000; // 3122 :  96 - 0x60
      12'hC33: dout <= 8'b01111110; // 3123 : 126 - 0x7e
      12'hC34: dout <= 8'b01100000; // 3124 :  96 - 0x60
      12'hC35: dout <= 8'b01100000; // 3125 :  96 - 0x60
      12'hC36: dout <= 8'b01111111; // 3126 : 127 - 0x7f
      12'hC37: dout <= 8'b00000000; // 3127 :   0 - 0x0
      12'hC38: dout <= 8'b00000000; // 3128 :   0 - 0x0 -- plane 1
      12'hC39: dout <= 8'b00000000; // 3129 :   0 - 0x0
      12'hC3A: dout <= 8'b00000000; // 3130 :   0 - 0x0
      12'hC3B: dout <= 8'b00000000; // 3131 :   0 - 0x0
      12'hC3C: dout <= 8'b00000000; // 3132 :   0 - 0x0
      12'hC3D: dout <= 8'b00000000; // 3133 :   0 - 0x0
      12'hC3E: dout <= 8'b00000000; // 3134 :   0 - 0x0
      12'hC3F: dout <= 8'b00000000; // 3135 :   0 - 0x0
      12'hC40: dout <= 8'b00111110; // 3136 :  62 - 0x3e -- Sprite 0xc4
      12'hC41: dout <= 8'b01100011; // 3137 :  99 - 0x63
      12'hC42: dout <= 8'b01100011; // 3138 :  99 - 0x63
      12'hC43: dout <= 8'b01100011; // 3139 :  99 - 0x63
      12'hC44: dout <= 8'b01100011; // 3140 :  99 - 0x63
      12'hC45: dout <= 8'b01100011; // 3141 :  99 - 0x63
      12'hC46: dout <= 8'b00111110; // 3142 :  62 - 0x3e
      12'hC47: dout <= 8'b00000000; // 3143 :   0 - 0x0
      12'hC48: dout <= 8'b00000000; // 3144 :   0 - 0x0 -- plane 1
      12'hC49: dout <= 8'b00000000; // 3145 :   0 - 0x0
      12'hC4A: dout <= 8'b00000000; // 3146 :   0 - 0x0
      12'hC4B: dout <= 8'b00000000; // 3147 :   0 - 0x0
      12'hC4C: dout <= 8'b00000000; // 3148 :   0 - 0x0
      12'hC4D: dout <= 8'b00000000; // 3149 :   0 - 0x0
      12'hC4E: dout <= 8'b00000000; // 3150 :   0 - 0x0
      12'hC4F: dout <= 8'b00000000; // 3151 :   0 - 0x0
      12'hC50: dout <= 8'b01100011; // 3152 :  99 - 0x63 -- Sprite 0xc5
      12'hC51: dout <= 8'b01100011; // 3153 :  99 - 0x63
      12'hC52: dout <= 8'b01100011; // 3154 :  99 - 0x63
      12'hC53: dout <= 8'b01110111; // 3155 : 119 - 0x77
      12'hC54: dout <= 8'b00111110; // 3156 :  62 - 0x3e
      12'hC55: dout <= 8'b00011100; // 3157 :  28 - 0x1c
      12'hC56: dout <= 8'b00001000; // 3158 :   8 - 0x8
      12'hC57: dout <= 8'b00000000; // 3159 :   0 - 0x0
      12'hC58: dout <= 8'b00000000; // 3160 :   0 - 0x0 -- plane 1
      12'hC59: dout <= 8'b00000000; // 3161 :   0 - 0x0
      12'hC5A: dout <= 8'b00000000; // 3162 :   0 - 0x0
      12'hC5B: dout <= 8'b00000000; // 3163 :   0 - 0x0
      12'hC5C: dout <= 8'b00000000; // 3164 :   0 - 0x0
      12'hC5D: dout <= 8'b00000000; // 3165 :   0 - 0x0
      12'hC5E: dout <= 8'b00000000; // 3166 :   0 - 0x0
      12'hC5F: dout <= 8'b00000000; // 3167 :   0 - 0x0
      12'hC60: dout <= 8'b01111110; // 3168 : 126 - 0x7e -- Sprite 0xc6
      12'hC61: dout <= 8'b01100011; // 3169 :  99 - 0x63
      12'hC62: dout <= 8'b01100011; // 3170 :  99 - 0x63
      12'hC63: dout <= 8'b01100111; // 3171 : 103 - 0x67
      12'hC64: dout <= 8'b01111100; // 3172 : 124 - 0x7c
      12'hC65: dout <= 8'b01101110; // 3173 : 110 - 0x6e
      12'hC66: dout <= 8'b01100111; // 3174 : 103 - 0x67
      12'hC67: dout <= 8'b00000000; // 3175 :   0 - 0x0
      12'hC68: dout <= 8'b00000000; // 3176 :   0 - 0x0 -- plane 1
      12'hC69: dout <= 8'b00000000; // 3177 :   0 - 0x0
      12'hC6A: dout <= 8'b00000000; // 3178 :   0 - 0x0
      12'hC6B: dout <= 8'b00000000; // 3179 :   0 - 0x0
      12'hC6C: dout <= 8'b00000000; // 3180 :   0 - 0x0
      12'hC6D: dout <= 8'b00000000; // 3181 :   0 - 0x0
      12'hC6E: dout <= 8'b00000000; // 3182 :   0 - 0x0
      12'hC6F: dout <= 8'b00000000; // 3183 :   0 - 0x0
      12'hC70: dout <= 8'b00110011; // 3184 :  51 - 0x33 -- Sprite 0xc7
      12'hC71: dout <= 8'b00110011; // 3185 :  51 - 0x33
      12'hC72: dout <= 8'b00110011; // 3186 :  51 - 0x33
      12'hC73: dout <= 8'b00011110; // 3187 :  30 - 0x1e
      12'hC74: dout <= 8'b00001100; // 3188 :  12 - 0xc
      12'hC75: dout <= 8'b00001100; // 3189 :  12 - 0xc
      12'hC76: dout <= 8'b00001100; // 3190 :  12 - 0xc
      12'hC77: dout <= 8'b00000000; // 3191 :   0 - 0x0
      12'hC78: dout <= 8'b00000000; // 3192 :   0 - 0x0 -- plane 1
      12'hC79: dout <= 8'b00000000; // 3193 :   0 - 0x0
      12'hC7A: dout <= 8'b00000000; // 3194 :   0 - 0x0
      12'hC7B: dout <= 8'b00000000; // 3195 :   0 - 0x0
      12'hC7C: dout <= 8'b00000000; // 3196 :   0 - 0x0
      12'hC7D: dout <= 8'b00000000; // 3197 :   0 - 0x0
      12'hC7E: dout <= 8'b00000000; // 3198 :   0 - 0x0
      12'hC7F: dout <= 8'b00000000; // 3199 :   0 - 0x0
      12'hC80: dout <= 8'b00000000; // 3200 :   0 - 0x0 -- Sprite 0xc8
      12'hC81: dout <= 8'b00000000; // 3201 :   0 - 0x0
      12'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      12'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      12'hC84: dout <= 8'b00000000; // 3204 :   0 - 0x0
      12'hC85: dout <= 8'b00000000; // 3205 :   0 - 0x0
      12'hC86: dout <= 8'b00000000; // 3206 :   0 - 0x0
      12'hC87: dout <= 8'b00000000; // 3207 :   0 - 0x0
      12'hC88: dout <= 8'b00000000; // 3208 :   0 - 0x0 -- plane 1
      12'hC89: dout <= 8'b00000000; // 3209 :   0 - 0x0
      12'hC8A: dout <= 8'b00000000; // 3210 :   0 - 0x0
      12'hC8B: dout <= 8'b00000000; // 3211 :   0 - 0x0
      12'hC8C: dout <= 8'b00000000; // 3212 :   0 - 0x0
      12'hC8D: dout <= 8'b00000000; // 3213 :   0 - 0x0
      12'hC8E: dout <= 8'b00000000; // 3214 :   0 - 0x0
      12'hC8F: dout <= 8'b00000000; // 3215 :   0 - 0x0
      12'hC90: dout <= 8'b00000000; // 3216 :   0 - 0x0 -- Sprite 0xc9
      12'hC91: dout <= 8'b00000000; // 3217 :   0 - 0x0
      12'hC92: dout <= 8'b00000000; // 3218 :   0 - 0x0
      12'hC93: dout <= 8'b00000000; // 3219 :   0 - 0x0
      12'hC94: dout <= 8'b00000000; // 3220 :   0 - 0x0
      12'hC95: dout <= 8'b00000000; // 3221 :   0 - 0x0
      12'hC96: dout <= 8'b00000000; // 3222 :   0 - 0x0
      12'hC97: dout <= 8'b00000000; // 3223 :   0 - 0x0
      12'hC98: dout <= 8'b00000000; // 3224 :   0 - 0x0 -- plane 1
      12'hC99: dout <= 8'b00000000; // 3225 :   0 - 0x0
      12'hC9A: dout <= 8'b00000000; // 3226 :   0 - 0x0
      12'hC9B: dout <= 8'b00000000; // 3227 :   0 - 0x0
      12'hC9C: dout <= 8'b00000000; // 3228 :   0 - 0x0
      12'hC9D: dout <= 8'b00000000; // 3229 :   0 - 0x0
      12'hC9E: dout <= 8'b00000000; // 3230 :   0 - 0x0
      12'hC9F: dout <= 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout <= 8'b00000000; // 3232 :   0 - 0x0 -- Sprite 0xca
      12'hCA1: dout <= 8'b00000000; // 3233 :   0 - 0x0
      12'hCA2: dout <= 8'b00000000; // 3234 :   0 - 0x0
      12'hCA3: dout <= 8'b00000000; // 3235 :   0 - 0x0
      12'hCA4: dout <= 8'b00000000; // 3236 :   0 - 0x0
      12'hCA5: dout <= 8'b00000000; // 3237 :   0 - 0x0
      12'hCA6: dout <= 8'b00000000; // 3238 :   0 - 0x0
      12'hCA7: dout <= 8'b00000000; // 3239 :   0 - 0x0
      12'hCA8: dout <= 8'b00000000; // 3240 :   0 - 0x0 -- plane 1
      12'hCA9: dout <= 8'b00000000; // 3241 :   0 - 0x0
      12'hCAA: dout <= 8'b00000000; // 3242 :   0 - 0x0
      12'hCAB: dout <= 8'b00000000; // 3243 :   0 - 0x0
      12'hCAC: dout <= 8'b00000000; // 3244 :   0 - 0x0
      12'hCAD: dout <= 8'b00000000; // 3245 :   0 - 0x0
      12'hCAE: dout <= 8'b00000000; // 3246 :   0 - 0x0
      12'hCAF: dout <= 8'b00000000; // 3247 :   0 - 0x0
      12'hCB0: dout <= 8'b00000000; // 3248 :   0 - 0x0 -- Sprite 0xcb
      12'hCB1: dout <= 8'b00000000; // 3249 :   0 - 0x0
      12'hCB2: dout <= 8'b00000000; // 3250 :   0 - 0x0
      12'hCB3: dout <= 8'b00000000; // 3251 :   0 - 0x0
      12'hCB4: dout <= 8'b00000000; // 3252 :   0 - 0x0
      12'hCB5: dout <= 8'b00000000; // 3253 :   0 - 0x0
      12'hCB6: dout <= 8'b00000000; // 3254 :   0 - 0x0
      12'hCB7: dout <= 8'b00000000; // 3255 :   0 - 0x0
      12'hCB8: dout <= 8'b00000000; // 3256 :   0 - 0x0 -- plane 1
      12'hCB9: dout <= 8'b00000000; // 3257 :   0 - 0x0
      12'hCBA: dout <= 8'b00000000; // 3258 :   0 - 0x0
      12'hCBB: dout <= 8'b00000000; // 3259 :   0 - 0x0
      12'hCBC: dout <= 8'b00000000; // 3260 :   0 - 0x0
      12'hCBD: dout <= 8'b00000000; // 3261 :   0 - 0x0
      12'hCBE: dout <= 8'b00000000; // 3262 :   0 - 0x0
      12'hCBF: dout <= 8'b00000000; // 3263 :   0 - 0x0
      12'hCC0: dout <= 8'b00000000; // 3264 :   0 - 0x0 -- Sprite 0xcc
      12'hCC1: dout <= 8'b00000000; // 3265 :   0 - 0x0
      12'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      12'hCC3: dout <= 8'b00000000; // 3267 :   0 - 0x0
      12'hCC4: dout <= 8'b00000000; // 3268 :   0 - 0x0
      12'hCC5: dout <= 8'b00000000; // 3269 :   0 - 0x0
      12'hCC6: dout <= 8'b00000000; // 3270 :   0 - 0x0
      12'hCC7: dout <= 8'b00000000; // 3271 :   0 - 0x0
      12'hCC8: dout <= 8'b00000000; // 3272 :   0 - 0x0 -- plane 1
      12'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      12'hCCA: dout <= 8'b00000000; // 3274 :   0 - 0x0
      12'hCCB: dout <= 8'b00000000; // 3275 :   0 - 0x0
      12'hCCC: dout <= 8'b00000000; // 3276 :   0 - 0x0
      12'hCCD: dout <= 8'b00000000; // 3277 :   0 - 0x0
      12'hCCE: dout <= 8'b00000000; // 3278 :   0 - 0x0
      12'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout <= 8'b00000000; // 3280 :   0 - 0x0 -- Sprite 0xcd
      12'hCD1: dout <= 8'b00000000; // 3281 :   0 - 0x0
      12'hCD2: dout <= 8'b00000000; // 3282 :   0 - 0x0
      12'hCD3: dout <= 8'b00000000; // 3283 :   0 - 0x0
      12'hCD4: dout <= 8'b00000000; // 3284 :   0 - 0x0
      12'hCD5: dout <= 8'b00000000; // 3285 :   0 - 0x0
      12'hCD6: dout <= 8'b00000000; // 3286 :   0 - 0x0
      12'hCD7: dout <= 8'b00000000; // 3287 :   0 - 0x0
      12'hCD8: dout <= 8'b00000000; // 3288 :   0 - 0x0 -- plane 1
      12'hCD9: dout <= 8'b00000000; // 3289 :   0 - 0x0
      12'hCDA: dout <= 8'b00000000; // 3290 :   0 - 0x0
      12'hCDB: dout <= 8'b00000000; // 3291 :   0 - 0x0
      12'hCDC: dout <= 8'b00000000; // 3292 :   0 - 0x0
      12'hCDD: dout <= 8'b00000000; // 3293 :   0 - 0x0
      12'hCDE: dout <= 8'b00000000; // 3294 :   0 - 0x0
      12'hCDF: dout <= 8'b00000000; // 3295 :   0 - 0x0
      12'hCE0: dout <= 8'b00000000; // 3296 :   0 - 0x0 -- Sprite 0xce
      12'hCE1: dout <= 8'b00000000; // 3297 :   0 - 0x0
      12'hCE2: dout <= 8'b00000000; // 3298 :   0 - 0x0
      12'hCE3: dout <= 8'b00000000; // 3299 :   0 - 0x0
      12'hCE4: dout <= 8'b00000000; // 3300 :   0 - 0x0
      12'hCE5: dout <= 8'b00000000; // 3301 :   0 - 0x0
      12'hCE6: dout <= 8'b00000000; // 3302 :   0 - 0x0
      12'hCE7: dout <= 8'b00000000; // 3303 :   0 - 0x0
      12'hCE8: dout <= 8'b00000000; // 3304 :   0 - 0x0 -- plane 1
      12'hCE9: dout <= 8'b00000000; // 3305 :   0 - 0x0
      12'hCEA: dout <= 8'b00000000; // 3306 :   0 - 0x0
      12'hCEB: dout <= 8'b00000000; // 3307 :   0 - 0x0
      12'hCEC: dout <= 8'b00000000; // 3308 :   0 - 0x0
      12'hCED: dout <= 8'b00000000; // 3309 :   0 - 0x0
      12'hCEE: dout <= 8'b00000000; // 3310 :   0 - 0x0
      12'hCEF: dout <= 8'b00000000; // 3311 :   0 - 0x0
      12'hCF0: dout <= 8'b00000000; // 3312 :   0 - 0x0 -- Sprite 0xcf
      12'hCF1: dout <= 8'b00000000; // 3313 :   0 - 0x0
      12'hCF2: dout <= 8'b00000000; // 3314 :   0 - 0x0
      12'hCF3: dout <= 8'b00000000; // 3315 :   0 - 0x0
      12'hCF4: dout <= 8'b00000000; // 3316 :   0 - 0x0
      12'hCF5: dout <= 8'b00000000; // 3317 :   0 - 0x0
      12'hCF6: dout <= 8'b00000000; // 3318 :   0 - 0x0
      12'hCF7: dout <= 8'b00000000; // 3319 :   0 - 0x0
      12'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0 -- plane 1
      12'hCF9: dout <= 8'b00000000; // 3321 :   0 - 0x0
      12'hCFA: dout <= 8'b00000000; // 3322 :   0 - 0x0
      12'hCFB: dout <= 8'b00000000; // 3323 :   0 - 0x0
      12'hCFC: dout <= 8'b00000000; // 3324 :   0 - 0x0
      12'hCFD: dout <= 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout <= 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout <= 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout <= 8'b11111111; // 3328 : 255 - 0xff -- Sprite 0xd0
      12'hD01: dout <= 8'b11111111; // 3329 : 255 - 0xff
      12'hD02: dout <= 8'b11111111; // 3330 : 255 - 0xff
      12'hD03: dout <= 8'b11111111; // 3331 : 255 - 0xff
      12'hD04: dout <= 8'b11111111; // 3332 : 255 - 0xff
      12'hD05: dout <= 8'b11111111; // 3333 : 255 - 0xff
      12'hD06: dout <= 8'b11111111; // 3334 : 255 - 0xff
      12'hD07: dout <= 8'b11111111; // 3335 : 255 - 0xff
      12'hD08: dout <= 8'b11111111; // 3336 : 255 - 0xff -- plane 1
      12'hD09: dout <= 8'b11111111; // 3337 : 255 - 0xff
      12'hD0A: dout <= 8'b11111111; // 3338 : 255 - 0xff
      12'hD0B: dout <= 8'b11111111; // 3339 : 255 - 0xff
      12'hD0C: dout <= 8'b11111111; // 3340 : 255 - 0xff
      12'hD0D: dout <= 8'b11111111; // 3341 : 255 - 0xff
      12'hD0E: dout <= 8'b11111111; // 3342 : 255 - 0xff
      12'hD0F: dout <= 8'b11111111; // 3343 : 255 - 0xff
      12'hD10: dout <= 8'b11111111; // 3344 : 255 - 0xff -- Sprite 0xd1
      12'hD11: dout <= 8'b11111111; // 3345 : 255 - 0xff
      12'hD12: dout <= 8'b11111111; // 3346 : 255 - 0xff
      12'hD13: dout <= 8'b11111111; // 3347 : 255 - 0xff
      12'hD14: dout <= 8'b11111111; // 3348 : 255 - 0xff
      12'hD15: dout <= 8'b11111111; // 3349 : 255 - 0xff
      12'hD16: dout <= 8'b11111111; // 3350 : 255 - 0xff
      12'hD17: dout <= 8'b11111111; // 3351 : 255 - 0xff
      12'hD18: dout <= 8'b11111111; // 3352 : 255 - 0xff -- plane 1
      12'hD19: dout <= 8'b11111111; // 3353 : 255 - 0xff
      12'hD1A: dout <= 8'b11111111; // 3354 : 255 - 0xff
      12'hD1B: dout <= 8'b11111111; // 3355 : 255 - 0xff
      12'hD1C: dout <= 8'b11111111; // 3356 : 255 - 0xff
      12'hD1D: dout <= 8'b11111111; // 3357 : 255 - 0xff
      12'hD1E: dout <= 8'b11111111; // 3358 : 255 - 0xff
      12'hD1F: dout <= 8'b11111111; // 3359 : 255 - 0xff
      12'hD20: dout <= 8'b11111111; // 3360 : 255 - 0xff -- Sprite 0xd2
      12'hD21: dout <= 8'b11111111; // 3361 : 255 - 0xff
      12'hD22: dout <= 8'b11111111; // 3362 : 255 - 0xff
      12'hD23: dout <= 8'b11111111; // 3363 : 255 - 0xff
      12'hD24: dout <= 8'b11111111; // 3364 : 255 - 0xff
      12'hD25: dout <= 8'b11111111; // 3365 : 255 - 0xff
      12'hD26: dout <= 8'b11111111; // 3366 : 255 - 0xff
      12'hD27: dout <= 8'b11111111; // 3367 : 255 - 0xff
      12'hD28: dout <= 8'b11111111; // 3368 : 255 - 0xff -- plane 1
      12'hD29: dout <= 8'b11111111; // 3369 : 255 - 0xff
      12'hD2A: dout <= 8'b11111111; // 3370 : 255 - 0xff
      12'hD2B: dout <= 8'b11111111; // 3371 : 255 - 0xff
      12'hD2C: dout <= 8'b11111111; // 3372 : 255 - 0xff
      12'hD2D: dout <= 8'b11111111; // 3373 : 255 - 0xff
      12'hD2E: dout <= 8'b11111111; // 3374 : 255 - 0xff
      12'hD2F: dout <= 8'b11111111; // 3375 : 255 - 0xff
      12'hD30: dout <= 8'b11111111; // 3376 : 255 - 0xff -- Sprite 0xd3
      12'hD31: dout <= 8'b11111111; // 3377 : 255 - 0xff
      12'hD32: dout <= 8'b11111111; // 3378 : 255 - 0xff
      12'hD33: dout <= 8'b11111111; // 3379 : 255 - 0xff
      12'hD34: dout <= 8'b11111111; // 3380 : 255 - 0xff
      12'hD35: dout <= 8'b11111111; // 3381 : 255 - 0xff
      12'hD36: dout <= 8'b11111111; // 3382 : 255 - 0xff
      12'hD37: dout <= 8'b11111111; // 3383 : 255 - 0xff
      12'hD38: dout <= 8'b11111111; // 3384 : 255 - 0xff -- plane 1
      12'hD39: dout <= 8'b11111111; // 3385 : 255 - 0xff
      12'hD3A: dout <= 8'b11111111; // 3386 : 255 - 0xff
      12'hD3B: dout <= 8'b11111111; // 3387 : 255 - 0xff
      12'hD3C: dout <= 8'b11111111; // 3388 : 255 - 0xff
      12'hD3D: dout <= 8'b11111111; // 3389 : 255 - 0xff
      12'hD3E: dout <= 8'b11111111; // 3390 : 255 - 0xff
      12'hD3F: dout <= 8'b11111111; // 3391 : 255 - 0xff
      12'hD40: dout <= 8'b11111111; // 3392 : 255 - 0xff -- Sprite 0xd4
      12'hD41: dout <= 8'b11111111; // 3393 : 255 - 0xff
      12'hD42: dout <= 8'b11111111; // 3394 : 255 - 0xff
      12'hD43: dout <= 8'b11111111; // 3395 : 255 - 0xff
      12'hD44: dout <= 8'b11111111; // 3396 : 255 - 0xff
      12'hD45: dout <= 8'b11111111; // 3397 : 255 - 0xff
      12'hD46: dout <= 8'b11111111; // 3398 : 255 - 0xff
      12'hD47: dout <= 8'b11111111; // 3399 : 255 - 0xff
      12'hD48: dout <= 8'b11111111; // 3400 : 255 - 0xff -- plane 1
      12'hD49: dout <= 8'b11111111; // 3401 : 255 - 0xff
      12'hD4A: dout <= 8'b11111111; // 3402 : 255 - 0xff
      12'hD4B: dout <= 8'b11111111; // 3403 : 255 - 0xff
      12'hD4C: dout <= 8'b11111111; // 3404 : 255 - 0xff
      12'hD4D: dout <= 8'b11111111; // 3405 : 255 - 0xff
      12'hD4E: dout <= 8'b11111111; // 3406 : 255 - 0xff
      12'hD4F: dout <= 8'b11111111; // 3407 : 255 - 0xff
      12'hD50: dout <= 8'b11111111; // 3408 : 255 - 0xff -- Sprite 0xd5
      12'hD51: dout <= 8'b11111111; // 3409 : 255 - 0xff
      12'hD52: dout <= 8'b11111111; // 3410 : 255 - 0xff
      12'hD53: dout <= 8'b11111111; // 3411 : 255 - 0xff
      12'hD54: dout <= 8'b11111111; // 3412 : 255 - 0xff
      12'hD55: dout <= 8'b11111111; // 3413 : 255 - 0xff
      12'hD56: dout <= 8'b11111111; // 3414 : 255 - 0xff
      12'hD57: dout <= 8'b11111111; // 3415 : 255 - 0xff
      12'hD58: dout <= 8'b11111111; // 3416 : 255 - 0xff -- plane 1
      12'hD59: dout <= 8'b11111111; // 3417 : 255 - 0xff
      12'hD5A: dout <= 8'b11111111; // 3418 : 255 - 0xff
      12'hD5B: dout <= 8'b11111111; // 3419 : 255 - 0xff
      12'hD5C: dout <= 8'b11111111; // 3420 : 255 - 0xff
      12'hD5D: dout <= 8'b11111111; // 3421 : 255 - 0xff
      12'hD5E: dout <= 8'b11111111; // 3422 : 255 - 0xff
      12'hD5F: dout <= 8'b11111111; // 3423 : 255 - 0xff
      12'hD60: dout <= 8'b11111111; // 3424 : 255 - 0xff -- Sprite 0xd6
      12'hD61: dout <= 8'b11111111; // 3425 : 255 - 0xff
      12'hD62: dout <= 8'b11111111; // 3426 : 255 - 0xff
      12'hD63: dout <= 8'b11111111; // 3427 : 255 - 0xff
      12'hD64: dout <= 8'b11111111; // 3428 : 255 - 0xff
      12'hD65: dout <= 8'b11111111; // 3429 : 255 - 0xff
      12'hD66: dout <= 8'b11111111; // 3430 : 255 - 0xff
      12'hD67: dout <= 8'b11111111; // 3431 : 255 - 0xff
      12'hD68: dout <= 8'b11111111; // 3432 : 255 - 0xff -- plane 1
      12'hD69: dout <= 8'b11111111; // 3433 : 255 - 0xff
      12'hD6A: dout <= 8'b11111111; // 3434 : 255 - 0xff
      12'hD6B: dout <= 8'b11111111; // 3435 : 255 - 0xff
      12'hD6C: dout <= 8'b11111111; // 3436 : 255 - 0xff
      12'hD6D: dout <= 8'b11111111; // 3437 : 255 - 0xff
      12'hD6E: dout <= 8'b11111111; // 3438 : 255 - 0xff
      12'hD6F: dout <= 8'b11111111; // 3439 : 255 - 0xff
      12'hD70: dout <= 8'b11111111; // 3440 : 255 - 0xff -- Sprite 0xd7
      12'hD71: dout <= 8'b11111111; // 3441 : 255 - 0xff
      12'hD72: dout <= 8'b11111111; // 3442 : 255 - 0xff
      12'hD73: dout <= 8'b11111111; // 3443 : 255 - 0xff
      12'hD74: dout <= 8'b11111111; // 3444 : 255 - 0xff
      12'hD75: dout <= 8'b11111111; // 3445 : 255 - 0xff
      12'hD76: dout <= 8'b11111111; // 3446 : 255 - 0xff
      12'hD77: dout <= 8'b11111111; // 3447 : 255 - 0xff
      12'hD78: dout <= 8'b11111111; // 3448 : 255 - 0xff -- plane 1
      12'hD79: dout <= 8'b11111111; // 3449 : 255 - 0xff
      12'hD7A: dout <= 8'b11111111; // 3450 : 255 - 0xff
      12'hD7B: dout <= 8'b11111111; // 3451 : 255 - 0xff
      12'hD7C: dout <= 8'b11111111; // 3452 : 255 - 0xff
      12'hD7D: dout <= 8'b11111111; // 3453 : 255 - 0xff
      12'hD7E: dout <= 8'b11111111; // 3454 : 255 - 0xff
      12'hD7F: dout <= 8'b11111111; // 3455 : 255 - 0xff
      12'hD80: dout <= 8'b11111111; // 3456 : 255 - 0xff -- Sprite 0xd8
      12'hD81: dout <= 8'b11111111; // 3457 : 255 - 0xff
      12'hD82: dout <= 8'b11111111; // 3458 : 255 - 0xff
      12'hD83: dout <= 8'b11111111; // 3459 : 255 - 0xff
      12'hD84: dout <= 8'b11111111; // 3460 : 255 - 0xff
      12'hD85: dout <= 8'b11111111; // 3461 : 255 - 0xff
      12'hD86: dout <= 8'b11111111; // 3462 : 255 - 0xff
      12'hD87: dout <= 8'b11111111; // 3463 : 255 - 0xff
      12'hD88: dout <= 8'b11111111; // 3464 : 255 - 0xff -- plane 1
      12'hD89: dout <= 8'b11111111; // 3465 : 255 - 0xff
      12'hD8A: dout <= 8'b11111111; // 3466 : 255 - 0xff
      12'hD8B: dout <= 8'b11111111; // 3467 : 255 - 0xff
      12'hD8C: dout <= 8'b11111111; // 3468 : 255 - 0xff
      12'hD8D: dout <= 8'b11111111; // 3469 : 255 - 0xff
      12'hD8E: dout <= 8'b11111111; // 3470 : 255 - 0xff
      12'hD8F: dout <= 8'b11111111; // 3471 : 255 - 0xff
      12'hD90: dout <= 8'b11111111; // 3472 : 255 - 0xff -- Sprite 0xd9
      12'hD91: dout <= 8'b11111111; // 3473 : 255 - 0xff
      12'hD92: dout <= 8'b11111111; // 3474 : 255 - 0xff
      12'hD93: dout <= 8'b11111111; // 3475 : 255 - 0xff
      12'hD94: dout <= 8'b11111111; // 3476 : 255 - 0xff
      12'hD95: dout <= 8'b11111111; // 3477 : 255 - 0xff
      12'hD96: dout <= 8'b11111111; // 3478 : 255 - 0xff
      12'hD97: dout <= 8'b11111111; // 3479 : 255 - 0xff
      12'hD98: dout <= 8'b11111111; // 3480 : 255 - 0xff -- plane 1
      12'hD99: dout <= 8'b11111111; // 3481 : 255 - 0xff
      12'hD9A: dout <= 8'b11111111; // 3482 : 255 - 0xff
      12'hD9B: dout <= 8'b11111111; // 3483 : 255 - 0xff
      12'hD9C: dout <= 8'b11111111; // 3484 : 255 - 0xff
      12'hD9D: dout <= 8'b11111111; // 3485 : 255 - 0xff
      12'hD9E: dout <= 8'b11111111; // 3486 : 255 - 0xff
      12'hD9F: dout <= 8'b11111111; // 3487 : 255 - 0xff
      12'hDA0: dout <= 8'b11111111; // 3488 : 255 - 0xff -- Sprite 0xda
      12'hDA1: dout <= 8'b11111111; // 3489 : 255 - 0xff
      12'hDA2: dout <= 8'b11111111; // 3490 : 255 - 0xff
      12'hDA3: dout <= 8'b11111111; // 3491 : 255 - 0xff
      12'hDA4: dout <= 8'b11111111; // 3492 : 255 - 0xff
      12'hDA5: dout <= 8'b11111111; // 3493 : 255 - 0xff
      12'hDA6: dout <= 8'b11111111; // 3494 : 255 - 0xff
      12'hDA7: dout <= 8'b11111111; // 3495 : 255 - 0xff
      12'hDA8: dout <= 8'b11111111; // 3496 : 255 - 0xff -- plane 1
      12'hDA9: dout <= 8'b11111111; // 3497 : 255 - 0xff
      12'hDAA: dout <= 8'b11111111; // 3498 : 255 - 0xff
      12'hDAB: dout <= 8'b11111111; // 3499 : 255 - 0xff
      12'hDAC: dout <= 8'b11111111; // 3500 : 255 - 0xff
      12'hDAD: dout <= 8'b11111111; // 3501 : 255 - 0xff
      12'hDAE: dout <= 8'b11111111; // 3502 : 255 - 0xff
      12'hDAF: dout <= 8'b11111111; // 3503 : 255 - 0xff
      12'hDB0: dout <= 8'b11111111; // 3504 : 255 - 0xff -- Sprite 0xdb
      12'hDB1: dout <= 8'b11111111; // 3505 : 255 - 0xff
      12'hDB2: dout <= 8'b11111111; // 3506 : 255 - 0xff
      12'hDB3: dout <= 8'b11111111; // 3507 : 255 - 0xff
      12'hDB4: dout <= 8'b11111111; // 3508 : 255 - 0xff
      12'hDB5: dout <= 8'b11111111; // 3509 : 255 - 0xff
      12'hDB6: dout <= 8'b11111111; // 3510 : 255 - 0xff
      12'hDB7: dout <= 8'b11111111; // 3511 : 255 - 0xff
      12'hDB8: dout <= 8'b11111111; // 3512 : 255 - 0xff -- plane 1
      12'hDB9: dout <= 8'b11111111; // 3513 : 255 - 0xff
      12'hDBA: dout <= 8'b11111111; // 3514 : 255 - 0xff
      12'hDBB: dout <= 8'b11111111; // 3515 : 255 - 0xff
      12'hDBC: dout <= 8'b11111111; // 3516 : 255 - 0xff
      12'hDBD: dout <= 8'b11111111; // 3517 : 255 - 0xff
      12'hDBE: dout <= 8'b11111111; // 3518 : 255 - 0xff
      12'hDBF: dout <= 8'b11111111; // 3519 : 255 - 0xff
      12'hDC0: dout <= 8'b11111111; // 3520 : 255 - 0xff -- Sprite 0xdc
      12'hDC1: dout <= 8'b11111111; // 3521 : 255 - 0xff
      12'hDC2: dout <= 8'b11111111; // 3522 : 255 - 0xff
      12'hDC3: dout <= 8'b11111111; // 3523 : 255 - 0xff
      12'hDC4: dout <= 8'b11111111; // 3524 : 255 - 0xff
      12'hDC5: dout <= 8'b11111111; // 3525 : 255 - 0xff
      12'hDC6: dout <= 8'b11111111; // 3526 : 255 - 0xff
      12'hDC7: dout <= 8'b11111111; // 3527 : 255 - 0xff
      12'hDC8: dout <= 8'b11111111; // 3528 : 255 - 0xff -- plane 1
      12'hDC9: dout <= 8'b11111111; // 3529 : 255 - 0xff
      12'hDCA: dout <= 8'b11111111; // 3530 : 255 - 0xff
      12'hDCB: dout <= 8'b11111111; // 3531 : 255 - 0xff
      12'hDCC: dout <= 8'b11111111; // 3532 : 255 - 0xff
      12'hDCD: dout <= 8'b11111111; // 3533 : 255 - 0xff
      12'hDCE: dout <= 8'b11111111; // 3534 : 255 - 0xff
      12'hDCF: dout <= 8'b11111111; // 3535 : 255 - 0xff
      12'hDD0: dout <= 8'b11111111; // 3536 : 255 - 0xff -- Sprite 0xdd
      12'hDD1: dout <= 8'b11111111; // 3537 : 255 - 0xff
      12'hDD2: dout <= 8'b11111111; // 3538 : 255 - 0xff
      12'hDD3: dout <= 8'b11111111; // 3539 : 255 - 0xff
      12'hDD4: dout <= 8'b11111111; // 3540 : 255 - 0xff
      12'hDD5: dout <= 8'b11111111; // 3541 : 255 - 0xff
      12'hDD6: dout <= 8'b11111111; // 3542 : 255 - 0xff
      12'hDD7: dout <= 8'b11111111; // 3543 : 255 - 0xff
      12'hDD8: dout <= 8'b11111111; // 3544 : 255 - 0xff -- plane 1
      12'hDD9: dout <= 8'b11111111; // 3545 : 255 - 0xff
      12'hDDA: dout <= 8'b11111111; // 3546 : 255 - 0xff
      12'hDDB: dout <= 8'b11111111; // 3547 : 255 - 0xff
      12'hDDC: dout <= 8'b11111111; // 3548 : 255 - 0xff
      12'hDDD: dout <= 8'b11111111; // 3549 : 255 - 0xff
      12'hDDE: dout <= 8'b11111111; // 3550 : 255 - 0xff
      12'hDDF: dout <= 8'b11111111; // 3551 : 255 - 0xff
      12'hDE0: dout <= 8'b11111111; // 3552 : 255 - 0xff -- Sprite 0xde
      12'hDE1: dout <= 8'b11111111; // 3553 : 255 - 0xff
      12'hDE2: dout <= 8'b11111111; // 3554 : 255 - 0xff
      12'hDE3: dout <= 8'b11111111; // 3555 : 255 - 0xff
      12'hDE4: dout <= 8'b11111111; // 3556 : 255 - 0xff
      12'hDE5: dout <= 8'b11111111; // 3557 : 255 - 0xff
      12'hDE6: dout <= 8'b11111111; // 3558 : 255 - 0xff
      12'hDE7: dout <= 8'b11111111; // 3559 : 255 - 0xff
      12'hDE8: dout <= 8'b11111111; // 3560 : 255 - 0xff -- plane 1
      12'hDE9: dout <= 8'b11111111; // 3561 : 255 - 0xff
      12'hDEA: dout <= 8'b11111111; // 3562 : 255 - 0xff
      12'hDEB: dout <= 8'b11111111; // 3563 : 255 - 0xff
      12'hDEC: dout <= 8'b11111111; // 3564 : 255 - 0xff
      12'hDED: dout <= 8'b11111111; // 3565 : 255 - 0xff
      12'hDEE: dout <= 8'b11111111; // 3566 : 255 - 0xff
      12'hDEF: dout <= 8'b11111111; // 3567 : 255 - 0xff
      12'hDF0: dout <= 8'b11111111; // 3568 : 255 - 0xff -- Sprite 0xdf
      12'hDF1: dout <= 8'b11111111; // 3569 : 255 - 0xff
      12'hDF2: dout <= 8'b11111111; // 3570 : 255 - 0xff
      12'hDF3: dout <= 8'b11111111; // 3571 : 255 - 0xff
      12'hDF4: dout <= 8'b11111111; // 3572 : 255 - 0xff
      12'hDF5: dout <= 8'b11111111; // 3573 : 255 - 0xff
      12'hDF6: dout <= 8'b11111111; // 3574 : 255 - 0xff
      12'hDF7: dout <= 8'b11111111; // 3575 : 255 - 0xff
      12'hDF8: dout <= 8'b11111111; // 3576 : 255 - 0xff -- plane 1
      12'hDF9: dout <= 8'b11111111; // 3577 : 255 - 0xff
      12'hDFA: dout <= 8'b11111111; // 3578 : 255 - 0xff
      12'hDFB: dout <= 8'b11111111; // 3579 : 255 - 0xff
      12'hDFC: dout <= 8'b11111111; // 3580 : 255 - 0xff
      12'hDFD: dout <= 8'b11111111; // 3581 : 255 - 0xff
      12'hDFE: dout <= 8'b11111111; // 3582 : 255 - 0xff
      12'hDFF: dout <= 8'b11111111; // 3583 : 255 - 0xff
      12'hE00: dout <= 8'b11111111; // 3584 : 255 - 0xff -- Sprite 0xe0
      12'hE01: dout <= 8'b11111111; // 3585 : 255 - 0xff
      12'hE02: dout <= 8'b11111111; // 3586 : 255 - 0xff
      12'hE03: dout <= 8'b11111111; // 3587 : 255 - 0xff
      12'hE04: dout <= 8'b11111111; // 3588 : 255 - 0xff
      12'hE05: dout <= 8'b11111111; // 3589 : 255 - 0xff
      12'hE06: dout <= 8'b11111111; // 3590 : 255 - 0xff
      12'hE07: dout <= 8'b11111111; // 3591 : 255 - 0xff
      12'hE08: dout <= 8'b11111111; // 3592 : 255 - 0xff -- plane 1
      12'hE09: dout <= 8'b11111111; // 3593 : 255 - 0xff
      12'hE0A: dout <= 8'b11111111; // 3594 : 255 - 0xff
      12'hE0B: dout <= 8'b11111111; // 3595 : 255 - 0xff
      12'hE0C: dout <= 8'b11111111; // 3596 : 255 - 0xff
      12'hE0D: dout <= 8'b11111111; // 3597 : 255 - 0xff
      12'hE0E: dout <= 8'b11111111; // 3598 : 255 - 0xff
      12'hE0F: dout <= 8'b11111111; // 3599 : 255 - 0xff
      12'hE10: dout <= 8'b11111111; // 3600 : 255 - 0xff -- Sprite 0xe1
      12'hE11: dout <= 8'b11111111; // 3601 : 255 - 0xff
      12'hE12: dout <= 8'b11111111; // 3602 : 255 - 0xff
      12'hE13: dout <= 8'b11111111; // 3603 : 255 - 0xff
      12'hE14: dout <= 8'b11111111; // 3604 : 255 - 0xff
      12'hE15: dout <= 8'b11111111; // 3605 : 255 - 0xff
      12'hE16: dout <= 8'b11111111; // 3606 : 255 - 0xff
      12'hE17: dout <= 8'b11111111; // 3607 : 255 - 0xff
      12'hE18: dout <= 8'b11111111; // 3608 : 255 - 0xff -- plane 1
      12'hE19: dout <= 8'b11111111; // 3609 : 255 - 0xff
      12'hE1A: dout <= 8'b11111111; // 3610 : 255 - 0xff
      12'hE1B: dout <= 8'b11111111; // 3611 : 255 - 0xff
      12'hE1C: dout <= 8'b11111111; // 3612 : 255 - 0xff
      12'hE1D: dout <= 8'b11111111; // 3613 : 255 - 0xff
      12'hE1E: dout <= 8'b11111111; // 3614 : 255 - 0xff
      12'hE1F: dout <= 8'b11111111; // 3615 : 255 - 0xff
      12'hE20: dout <= 8'b11111111; // 3616 : 255 - 0xff -- Sprite 0xe2
      12'hE21: dout <= 8'b11111111; // 3617 : 255 - 0xff
      12'hE22: dout <= 8'b11111111; // 3618 : 255 - 0xff
      12'hE23: dout <= 8'b11111111; // 3619 : 255 - 0xff
      12'hE24: dout <= 8'b11111111; // 3620 : 255 - 0xff
      12'hE25: dout <= 8'b11111111; // 3621 : 255 - 0xff
      12'hE26: dout <= 8'b11111111; // 3622 : 255 - 0xff
      12'hE27: dout <= 8'b11111111; // 3623 : 255 - 0xff
      12'hE28: dout <= 8'b11111111; // 3624 : 255 - 0xff -- plane 1
      12'hE29: dout <= 8'b11111111; // 3625 : 255 - 0xff
      12'hE2A: dout <= 8'b11111111; // 3626 : 255 - 0xff
      12'hE2B: dout <= 8'b11111111; // 3627 : 255 - 0xff
      12'hE2C: dout <= 8'b11111111; // 3628 : 255 - 0xff
      12'hE2D: dout <= 8'b11111111; // 3629 : 255 - 0xff
      12'hE2E: dout <= 8'b11111111; // 3630 : 255 - 0xff
      12'hE2F: dout <= 8'b11111111; // 3631 : 255 - 0xff
      12'hE30: dout <= 8'b11111111; // 3632 : 255 - 0xff -- Sprite 0xe3
      12'hE31: dout <= 8'b11111111; // 3633 : 255 - 0xff
      12'hE32: dout <= 8'b11111111; // 3634 : 255 - 0xff
      12'hE33: dout <= 8'b11111111; // 3635 : 255 - 0xff
      12'hE34: dout <= 8'b11111111; // 3636 : 255 - 0xff
      12'hE35: dout <= 8'b11111111; // 3637 : 255 - 0xff
      12'hE36: dout <= 8'b11111111; // 3638 : 255 - 0xff
      12'hE37: dout <= 8'b11111111; // 3639 : 255 - 0xff
      12'hE38: dout <= 8'b11111111; // 3640 : 255 - 0xff -- plane 1
      12'hE39: dout <= 8'b11111111; // 3641 : 255 - 0xff
      12'hE3A: dout <= 8'b11111111; // 3642 : 255 - 0xff
      12'hE3B: dout <= 8'b11111111; // 3643 : 255 - 0xff
      12'hE3C: dout <= 8'b11111111; // 3644 : 255 - 0xff
      12'hE3D: dout <= 8'b11111111; // 3645 : 255 - 0xff
      12'hE3E: dout <= 8'b11111111; // 3646 : 255 - 0xff
      12'hE3F: dout <= 8'b11111111; // 3647 : 255 - 0xff
      12'hE40: dout <= 8'b11111111; // 3648 : 255 - 0xff -- Sprite 0xe4
      12'hE41: dout <= 8'b11111111; // 3649 : 255 - 0xff
      12'hE42: dout <= 8'b11111111; // 3650 : 255 - 0xff
      12'hE43: dout <= 8'b11111111; // 3651 : 255 - 0xff
      12'hE44: dout <= 8'b11111111; // 3652 : 255 - 0xff
      12'hE45: dout <= 8'b11111111; // 3653 : 255 - 0xff
      12'hE46: dout <= 8'b11111111; // 3654 : 255 - 0xff
      12'hE47: dout <= 8'b11111111; // 3655 : 255 - 0xff
      12'hE48: dout <= 8'b11111111; // 3656 : 255 - 0xff -- plane 1
      12'hE49: dout <= 8'b11111111; // 3657 : 255 - 0xff
      12'hE4A: dout <= 8'b11111111; // 3658 : 255 - 0xff
      12'hE4B: dout <= 8'b11111111; // 3659 : 255 - 0xff
      12'hE4C: dout <= 8'b11111111; // 3660 : 255 - 0xff
      12'hE4D: dout <= 8'b11111111; // 3661 : 255 - 0xff
      12'hE4E: dout <= 8'b11111111; // 3662 : 255 - 0xff
      12'hE4F: dout <= 8'b11111111; // 3663 : 255 - 0xff
      12'hE50: dout <= 8'b11111111; // 3664 : 255 - 0xff -- Sprite 0xe5
      12'hE51: dout <= 8'b11111111; // 3665 : 255 - 0xff
      12'hE52: dout <= 8'b11111111; // 3666 : 255 - 0xff
      12'hE53: dout <= 8'b11111111; // 3667 : 255 - 0xff
      12'hE54: dout <= 8'b11111111; // 3668 : 255 - 0xff
      12'hE55: dout <= 8'b11111111; // 3669 : 255 - 0xff
      12'hE56: dout <= 8'b11111111; // 3670 : 255 - 0xff
      12'hE57: dout <= 8'b11111111; // 3671 : 255 - 0xff
      12'hE58: dout <= 8'b11111111; // 3672 : 255 - 0xff -- plane 1
      12'hE59: dout <= 8'b11111111; // 3673 : 255 - 0xff
      12'hE5A: dout <= 8'b11111111; // 3674 : 255 - 0xff
      12'hE5B: dout <= 8'b11111111; // 3675 : 255 - 0xff
      12'hE5C: dout <= 8'b11111111; // 3676 : 255 - 0xff
      12'hE5D: dout <= 8'b11111111; // 3677 : 255 - 0xff
      12'hE5E: dout <= 8'b11111111; // 3678 : 255 - 0xff
      12'hE5F: dout <= 8'b11111111; // 3679 : 255 - 0xff
      12'hE60: dout <= 8'b11111111; // 3680 : 255 - 0xff -- Sprite 0xe6
      12'hE61: dout <= 8'b11111111; // 3681 : 255 - 0xff
      12'hE62: dout <= 8'b11111111; // 3682 : 255 - 0xff
      12'hE63: dout <= 8'b11111111; // 3683 : 255 - 0xff
      12'hE64: dout <= 8'b11111111; // 3684 : 255 - 0xff
      12'hE65: dout <= 8'b11111111; // 3685 : 255 - 0xff
      12'hE66: dout <= 8'b11111111; // 3686 : 255 - 0xff
      12'hE67: dout <= 8'b11111111; // 3687 : 255 - 0xff
      12'hE68: dout <= 8'b11111111; // 3688 : 255 - 0xff -- plane 1
      12'hE69: dout <= 8'b11111111; // 3689 : 255 - 0xff
      12'hE6A: dout <= 8'b11111111; // 3690 : 255 - 0xff
      12'hE6B: dout <= 8'b11111111; // 3691 : 255 - 0xff
      12'hE6C: dout <= 8'b11111111; // 3692 : 255 - 0xff
      12'hE6D: dout <= 8'b11111111; // 3693 : 255 - 0xff
      12'hE6E: dout <= 8'b11111111; // 3694 : 255 - 0xff
      12'hE6F: dout <= 8'b11111111; // 3695 : 255 - 0xff
      12'hE70: dout <= 8'b11111111; // 3696 : 255 - 0xff -- Sprite 0xe7
      12'hE71: dout <= 8'b11111111; // 3697 : 255 - 0xff
      12'hE72: dout <= 8'b11111111; // 3698 : 255 - 0xff
      12'hE73: dout <= 8'b11111111; // 3699 : 255 - 0xff
      12'hE74: dout <= 8'b11111111; // 3700 : 255 - 0xff
      12'hE75: dout <= 8'b11111111; // 3701 : 255 - 0xff
      12'hE76: dout <= 8'b11111111; // 3702 : 255 - 0xff
      12'hE77: dout <= 8'b11111111; // 3703 : 255 - 0xff
      12'hE78: dout <= 8'b11111111; // 3704 : 255 - 0xff -- plane 1
      12'hE79: dout <= 8'b11111111; // 3705 : 255 - 0xff
      12'hE7A: dout <= 8'b11111111; // 3706 : 255 - 0xff
      12'hE7B: dout <= 8'b11111111; // 3707 : 255 - 0xff
      12'hE7C: dout <= 8'b11111111; // 3708 : 255 - 0xff
      12'hE7D: dout <= 8'b11111111; // 3709 : 255 - 0xff
      12'hE7E: dout <= 8'b11111111; // 3710 : 255 - 0xff
      12'hE7F: dout <= 8'b11111111; // 3711 : 255 - 0xff
      12'hE80: dout <= 8'b11111111; // 3712 : 255 - 0xff -- Sprite 0xe8
      12'hE81: dout <= 8'b11111111; // 3713 : 255 - 0xff
      12'hE82: dout <= 8'b11111111; // 3714 : 255 - 0xff
      12'hE83: dout <= 8'b11111111; // 3715 : 255 - 0xff
      12'hE84: dout <= 8'b11111111; // 3716 : 255 - 0xff
      12'hE85: dout <= 8'b11111111; // 3717 : 255 - 0xff
      12'hE86: dout <= 8'b11111111; // 3718 : 255 - 0xff
      12'hE87: dout <= 8'b11111111; // 3719 : 255 - 0xff
      12'hE88: dout <= 8'b11111111; // 3720 : 255 - 0xff -- plane 1
      12'hE89: dout <= 8'b11111111; // 3721 : 255 - 0xff
      12'hE8A: dout <= 8'b11111111; // 3722 : 255 - 0xff
      12'hE8B: dout <= 8'b11111111; // 3723 : 255 - 0xff
      12'hE8C: dout <= 8'b11111111; // 3724 : 255 - 0xff
      12'hE8D: dout <= 8'b11111111; // 3725 : 255 - 0xff
      12'hE8E: dout <= 8'b11111111; // 3726 : 255 - 0xff
      12'hE8F: dout <= 8'b11111111; // 3727 : 255 - 0xff
      12'hE90: dout <= 8'b11111111; // 3728 : 255 - 0xff -- Sprite 0xe9
      12'hE91: dout <= 8'b11111111; // 3729 : 255 - 0xff
      12'hE92: dout <= 8'b11111111; // 3730 : 255 - 0xff
      12'hE93: dout <= 8'b11111111; // 3731 : 255 - 0xff
      12'hE94: dout <= 8'b11111111; // 3732 : 255 - 0xff
      12'hE95: dout <= 8'b11111111; // 3733 : 255 - 0xff
      12'hE96: dout <= 8'b11111111; // 3734 : 255 - 0xff
      12'hE97: dout <= 8'b11111111; // 3735 : 255 - 0xff
      12'hE98: dout <= 8'b11111111; // 3736 : 255 - 0xff -- plane 1
      12'hE99: dout <= 8'b11111111; // 3737 : 255 - 0xff
      12'hE9A: dout <= 8'b11111111; // 3738 : 255 - 0xff
      12'hE9B: dout <= 8'b11111111; // 3739 : 255 - 0xff
      12'hE9C: dout <= 8'b11111111; // 3740 : 255 - 0xff
      12'hE9D: dout <= 8'b11111111; // 3741 : 255 - 0xff
      12'hE9E: dout <= 8'b11111111; // 3742 : 255 - 0xff
      12'hE9F: dout <= 8'b11111111; // 3743 : 255 - 0xff
      12'hEA0: dout <= 8'b11111111; // 3744 : 255 - 0xff -- Sprite 0xea
      12'hEA1: dout <= 8'b11111111; // 3745 : 255 - 0xff
      12'hEA2: dout <= 8'b11111111; // 3746 : 255 - 0xff
      12'hEA3: dout <= 8'b11111111; // 3747 : 255 - 0xff
      12'hEA4: dout <= 8'b11111111; // 3748 : 255 - 0xff
      12'hEA5: dout <= 8'b11111111; // 3749 : 255 - 0xff
      12'hEA6: dout <= 8'b11111111; // 3750 : 255 - 0xff
      12'hEA7: dout <= 8'b11111111; // 3751 : 255 - 0xff
      12'hEA8: dout <= 8'b11111111; // 3752 : 255 - 0xff -- plane 1
      12'hEA9: dout <= 8'b11111111; // 3753 : 255 - 0xff
      12'hEAA: dout <= 8'b11111111; // 3754 : 255 - 0xff
      12'hEAB: dout <= 8'b11111111; // 3755 : 255 - 0xff
      12'hEAC: dout <= 8'b11111111; // 3756 : 255 - 0xff
      12'hEAD: dout <= 8'b11111111; // 3757 : 255 - 0xff
      12'hEAE: dout <= 8'b11111111; // 3758 : 255 - 0xff
      12'hEAF: dout <= 8'b11111111; // 3759 : 255 - 0xff
      12'hEB0: dout <= 8'b11111111; // 3760 : 255 - 0xff -- Sprite 0xeb
      12'hEB1: dout <= 8'b11111111; // 3761 : 255 - 0xff
      12'hEB2: dout <= 8'b11111111; // 3762 : 255 - 0xff
      12'hEB3: dout <= 8'b11111111; // 3763 : 255 - 0xff
      12'hEB4: dout <= 8'b11111111; // 3764 : 255 - 0xff
      12'hEB5: dout <= 8'b11111111; // 3765 : 255 - 0xff
      12'hEB6: dout <= 8'b11111111; // 3766 : 255 - 0xff
      12'hEB7: dout <= 8'b11111111; // 3767 : 255 - 0xff
      12'hEB8: dout <= 8'b11111111; // 3768 : 255 - 0xff -- plane 1
      12'hEB9: dout <= 8'b11111111; // 3769 : 255 - 0xff
      12'hEBA: dout <= 8'b11111111; // 3770 : 255 - 0xff
      12'hEBB: dout <= 8'b11111111; // 3771 : 255 - 0xff
      12'hEBC: dout <= 8'b11111111; // 3772 : 255 - 0xff
      12'hEBD: dout <= 8'b11111111; // 3773 : 255 - 0xff
      12'hEBE: dout <= 8'b11111111; // 3774 : 255 - 0xff
      12'hEBF: dout <= 8'b11111111; // 3775 : 255 - 0xff
      12'hEC0: dout <= 8'b11111111; // 3776 : 255 - 0xff -- Sprite 0xec
      12'hEC1: dout <= 8'b11111111; // 3777 : 255 - 0xff
      12'hEC2: dout <= 8'b11111111; // 3778 : 255 - 0xff
      12'hEC3: dout <= 8'b11111111; // 3779 : 255 - 0xff
      12'hEC4: dout <= 8'b11111111; // 3780 : 255 - 0xff
      12'hEC5: dout <= 8'b11111111; // 3781 : 255 - 0xff
      12'hEC6: dout <= 8'b11111111; // 3782 : 255 - 0xff
      12'hEC7: dout <= 8'b11111111; // 3783 : 255 - 0xff
      12'hEC8: dout <= 8'b11111111; // 3784 : 255 - 0xff -- plane 1
      12'hEC9: dout <= 8'b11111111; // 3785 : 255 - 0xff
      12'hECA: dout <= 8'b11111111; // 3786 : 255 - 0xff
      12'hECB: dout <= 8'b11111111; // 3787 : 255 - 0xff
      12'hECC: dout <= 8'b11111111; // 3788 : 255 - 0xff
      12'hECD: dout <= 8'b11111111; // 3789 : 255 - 0xff
      12'hECE: dout <= 8'b11111111; // 3790 : 255 - 0xff
      12'hECF: dout <= 8'b11111111; // 3791 : 255 - 0xff
      12'hED0: dout <= 8'b11111111; // 3792 : 255 - 0xff -- Sprite 0xed
      12'hED1: dout <= 8'b11111111; // 3793 : 255 - 0xff
      12'hED2: dout <= 8'b11111111; // 3794 : 255 - 0xff
      12'hED3: dout <= 8'b11111111; // 3795 : 255 - 0xff
      12'hED4: dout <= 8'b11111111; // 3796 : 255 - 0xff
      12'hED5: dout <= 8'b11111111; // 3797 : 255 - 0xff
      12'hED6: dout <= 8'b11111111; // 3798 : 255 - 0xff
      12'hED7: dout <= 8'b11111111; // 3799 : 255 - 0xff
      12'hED8: dout <= 8'b11111111; // 3800 : 255 - 0xff -- plane 1
      12'hED9: dout <= 8'b11111111; // 3801 : 255 - 0xff
      12'hEDA: dout <= 8'b11111111; // 3802 : 255 - 0xff
      12'hEDB: dout <= 8'b11111111; // 3803 : 255 - 0xff
      12'hEDC: dout <= 8'b11111111; // 3804 : 255 - 0xff
      12'hEDD: dout <= 8'b11111111; // 3805 : 255 - 0xff
      12'hEDE: dout <= 8'b11111111; // 3806 : 255 - 0xff
      12'hEDF: dout <= 8'b11111111; // 3807 : 255 - 0xff
      12'hEE0: dout <= 8'b11111111; // 3808 : 255 - 0xff -- Sprite 0xee
      12'hEE1: dout <= 8'b11111111; // 3809 : 255 - 0xff
      12'hEE2: dout <= 8'b11111111; // 3810 : 255 - 0xff
      12'hEE3: dout <= 8'b11111111; // 3811 : 255 - 0xff
      12'hEE4: dout <= 8'b11111111; // 3812 : 255 - 0xff
      12'hEE5: dout <= 8'b11111111; // 3813 : 255 - 0xff
      12'hEE6: dout <= 8'b11111111; // 3814 : 255 - 0xff
      12'hEE7: dout <= 8'b11111111; // 3815 : 255 - 0xff
      12'hEE8: dout <= 8'b11111111; // 3816 : 255 - 0xff -- plane 1
      12'hEE9: dout <= 8'b11111111; // 3817 : 255 - 0xff
      12'hEEA: dout <= 8'b11111111; // 3818 : 255 - 0xff
      12'hEEB: dout <= 8'b11111111; // 3819 : 255 - 0xff
      12'hEEC: dout <= 8'b11111111; // 3820 : 255 - 0xff
      12'hEED: dout <= 8'b11111111; // 3821 : 255 - 0xff
      12'hEEE: dout <= 8'b11111111; // 3822 : 255 - 0xff
      12'hEEF: dout <= 8'b11111111; // 3823 : 255 - 0xff
      12'hEF0: dout <= 8'b11111111; // 3824 : 255 - 0xff -- Sprite 0xef
      12'hEF1: dout <= 8'b11111111; // 3825 : 255 - 0xff
      12'hEF2: dout <= 8'b11111111; // 3826 : 255 - 0xff
      12'hEF3: dout <= 8'b11111111; // 3827 : 255 - 0xff
      12'hEF4: dout <= 8'b11111111; // 3828 : 255 - 0xff
      12'hEF5: dout <= 8'b11111111; // 3829 : 255 - 0xff
      12'hEF6: dout <= 8'b11111111; // 3830 : 255 - 0xff
      12'hEF7: dout <= 8'b11111111; // 3831 : 255 - 0xff
      12'hEF8: dout <= 8'b11111111; // 3832 : 255 - 0xff -- plane 1
      12'hEF9: dout <= 8'b11111111; // 3833 : 255 - 0xff
      12'hEFA: dout <= 8'b11111111; // 3834 : 255 - 0xff
      12'hEFB: dout <= 8'b11111111; // 3835 : 255 - 0xff
      12'hEFC: dout <= 8'b11111111; // 3836 : 255 - 0xff
      12'hEFD: dout <= 8'b11111111; // 3837 : 255 - 0xff
      12'hEFE: dout <= 8'b11111111; // 3838 : 255 - 0xff
      12'hEFF: dout <= 8'b11111111; // 3839 : 255 - 0xff
      12'hF00: dout <= 8'b11111111; // 3840 : 255 - 0xff -- Sprite 0xf0
      12'hF01: dout <= 8'b11111111; // 3841 : 255 - 0xff
      12'hF02: dout <= 8'b11111111; // 3842 : 255 - 0xff
      12'hF03: dout <= 8'b11111111; // 3843 : 255 - 0xff
      12'hF04: dout <= 8'b11111111; // 3844 : 255 - 0xff
      12'hF05: dout <= 8'b11111111; // 3845 : 255 - 0xff
      12'hF06: dout <= 8'b11111111; // 3846 : 255 - 0xff
      12'hF07: dout <= 8'b11111111; // 3847 : 255 - 0xff
      12'hF08: dout <= 8'b11111111; // 3848 : 255 - 0xff -- plane 1
      12'hF09: dout <= 8'b11111111; // 3849 : 255 - 0xff
      12'hF0A: dout <= 8'b11111111; // 3850 : 255 - 0xff
      12'hF0B: dout <= 8'b11111111; // 3851 : 255 - 0xff
      12'hF0C: dout <= 8'b11111111; // 3852 : 255 - 0xff
      12'hF0D: dout <= 8'b11111111; // 3853 : 255 - 0xff
      12'hF0E: dout <= 8'b11111111; // 3854 : 255 - 0xff
      12'hF0F: dout <= 8'b11111111; // 3855 : 255 - 0xff
      12'hF10: dout <= 8'b11111111; // 3856 : 255 - 0xff -- Sprite 0xf1
      12'hF11: dout <= 8'b11111111; // 3857 : 255 - 0xff
      12'hF12: dout <= 8'b11111111; // 3858 : 255 - 0xff
      12'hF13: dout <= 8'b11111111; // 3859 : 255 - 0xff
      12'hF14: dout <= 8'b11111111; // 3860 : 255 - 0xff
      12'hF15: dout <= 8'b11111111; // 3861 : 255 - 0xff
      12'hF16: dout <= 8'b11111111; // 3862 : 255 - 0xff
      12'hF17: dout <= 8'b11111111; // 3863 : 255 - 0xff
      12'hF18: dout <= 8'b11111111; // 3864 : 255 - 0xff -- plane 1
      12'hF19: dout <= 8'b11111111; // 3865 : 255 - 0xff
      12'hF1A: dout <= 8'b11111111; // 3866 : 255 - 0xff
      12'hF1B: dout <= 8'b11111111; // 3867 : 255 - 0xff
      12'hF1C: dout <= 8'b11111111; // 3868 : 255 - 0xff
      12'hF1D: dout <= 8'b11111111; // 3869 : 255 - 0xff
      12'hF1E: dout <= 8'b11111111; // 3870 : 255 - 0xff
      12'hF1F: dout <= 8'b11111111; // 3871 : 255 - 0xff
      12'hF20: dout <= 8'b11111111; // 3872 : 255 - 0xff -- Sprite 0xf2
      12'hF21: dout <= 8'b11111111; // 3873 : 255 - 0xff
      12'hF22: dout <= 8'b11111111; // 3874 : 255 - 0xff
      12'hF23: dout <= 8'b11111111; // 3875 : 255 - 0xff
      12'hF24: dout <= 8'b11111111; // 3876 : 255 - 0xff
      12'hF25: dout <= 8'b11111111; // 3877 : 255 - 0xff
      12'hF26: dout <= 8'b11111111; // 3878 : 255 - 0xff
      12'hF27: dout <= 8'b11111111; // 3879 : 255 - 0xff
      12'hF28: dout <= 8'b11111111; // 3880 : 255 - 0xff -- plane 1
      12'hF29: dout <= 8'b11111111; // 3881 : 255 - 0xff
      12'hF2A: dout <= 8'b11111111; // 3882 : 255 - 0xff
      12'hF2B: dout <= 8'b11111111; // 3883 : 255 - 0xff
      12'hF2C: dout <= 8'b11111111; // 3884 : 255 - 0xff
      12'hF2D: dout <= 8'b11111111; // 3885 : 255 - 0xff
      12'hF2E: dout <= 8'b11111111; // 3886 : 255 - 0xff
      12'hF2F: dout <= 8'b11111111; // 3887 : 255 - 0xff
      12'hF30: dout <= 8'b11111111; // 3888 : 255 - 0xff -- Sprite 0xf3
      12'hF31: dout <= 8'b11111111; // 3889 : 255 - 0xff
      12'hF32: dout <= 8'b11111111; // 3890 : 255 - 0xff
      12'hF33: dout <= 8'b11111111; // 3891 : 255 - 0xff
      12'hF34: dout <= 8'b11111111; // 3892 : 255 - 0xff
      12'hF35: dout <= 8'b11111111; // 3893 : 255 - 0xff
      12'hF36: dout <= 8'b11111111; // 3894 : 255 - 0xff
      12'hF37: dout <= 8'b11111111; // 3895 : 255 - 0xff
      12'hF38: dout <= 8'b11111111; // 3896 : 255 - 0xff -- plane 1
      12'hF39: dout <= 8'b11111111; // 3897 : 255 - 0xff
      12'hF3A: dout <= 8'b11111111; // 3898 : 255 - 0xff
      12'hF3B: dout <= 8'b11111111; // 3899 : 255 - 0xff
      12'hF3C: dout <= 8'b11111111; // 3900 : 255 - 0xff
      12'hF3D: dout <= 8'b11111111; // 3901 : 255 - 0xff
      12'hF3E: dout <= 8'b11111111; // 3902 : 255 - 0xff
      12'hF3F: dout <= 8'b11111111; // 3903 : 255 - 0xff
      12'hF40: dout <= 8'b11111111; // 3904 : 255 - 0xff -- Sprite 0xf4
      12'hF41: dout <= 8'b11111111; // 3905 : 255 - 0xff
      12'hF42: dout <= 8'b11111111; // 3906 : 255 - 0xff
      12'hF43: dout <= 8'b11111111; // 3907 : 255 - 0xff
      12'hF44: dout <= 8'b11111111; // 3908 : 255 - 0xff
      12'hF45: dout <= 8'b11111111; // 3909 : 255 - 0xff
      12'hF46: dout <= 8'b11111111; // 3910 : 255 - 0xff
      12'hF47: dout <= 8'b11111111; // 3911 : 255 - 0xff
      12'hF48: dout <= 8'b11111111; // 3912 : 255 - 0xff -- plane 1
      12'hF49: dout <= 8'b11111111; // 3913 : 255 - 0xff
      12'hF4A: dout <= 8'b11111111; // 3914 : 255 - 0xff
      12'hF4B: dout <= 8'b11111111; // 3915 : 255 - 0xff
      12'hF4C: dout <= 8'b11111111; // 3916 : 255 - 0xff
      12'hF4D: dout <= 8'b11111111; // 3917 : 255 - 0xff
      12'hF4E: dout <= 8'b11111111; // 3918 : 255 - 0xff
      12'hF4F: dout <= 8'b11111111; // 3919 : 255 - 0xff
      12'hF50: dout <= 8'b11111111; // 3920 : 255 - 0xff -- Sprite 0xf5
      12'hF51: dout <= 8'b11111111; // 3921 : 255 - 0xff
      12'hF52: dout <= 8'b11111111; // 3922 : 255 - 0xff
      12'hF53: dout <= 8'b11111111; // 3923 : 255 - 0xff
      12'hF54: dout <= 8'b11111111; // 3924 : 255 - 0xff
      12'hF55: dout <= 8'b11111111; // 3925 : 255 - 0xff
      12'hF56: dout <= 8'b11111111; // 3926 : 255 - 0xff
      12'hF57: dout <= 8'b11111111; // 3927 : 255 - 0xff
      12'hF58: dout <= 8'b11111111; // 3928 : 255 - 0xff -- plane 1
      12'hF59: dout <= 8'b11111111; // 3929 : 255 - 0xff
      12'hF5A: dout <= 8'b11111111; // 3930 : 255 - 0xff
      12'hF5B: dout <= 8'b11111111; // 3931 : 255 - 0xff
      12'hF5C: dout <= 8'b11111111; // 3932 : 255 - 0xff
      12'hF5D: dout <= 8'b11111111; // 3933 : 255 - 0xff
      12'hF5E: dout <= 8'b11111111; // 3934 : 255 - 0xff
      12'hF5F: dout <= 8'b11111111; // 3935 : 255 - 0xff
      12'hF60: dout <= 8'b11111111; // 3936 : 255 - 0xff -- Sprite 0xf6
      12'hF61: dout <= 8'b11111111; // 3937 : 255 - 0xff
      12'hF62: dout <= 8'b11111111; // 3938 : 255 - 0xff
      12'hF63: dout <= 8'b11111111; // 3939 : 255 - 0xff
      12'hF64: dout <= 8'b11111111; // 3940 : 255 - 0xff
      12'hF65: dout <= 8'b11111111; // 3941 : 255 - 0xff
      12'hF66: dout <= 8'b11111111; // 3942 : 255 - 0xff
      12'hF67: dout <= 8'b11111111; // 3943 : 255 - 0xff
      12'hF68: dout <= 8'b11111111; // 3944 : 255 - 0xff -- plane 1
      12'hF69: dout <= 8'b11111111; // 3945 : 255 - 0xff
      12'hF6A: dout <= 8'b11111111; // 3946 : 255 - 0xff
      12'hF6B: dout <= 8'b11111111; // 3947 : 255 - 0xff
      12'hF6C: dout <= 8'b11111111; // 3948 : 255 - 0xff
      12'hF6D: dout <= 8'b11111111; // 3949 : 255 - 0xff
      12'hF6E: dout <= 8'b11111111; // 3950 : 255 - 0xff
      12'hF6F: dout <= 8'b11111111; // 3951 : 255 - 0xff
      12'hF70: dout <= 8'b11111111; // 3952 : 255 - 0xff -- Sprite 0xf7
      12'hF71: dout <= 8'b11111111; // 3953 : 255 - 0xff
      12'hF72: dout <= 8'b11111111; // 3954 : 255 - 0xff
      12'hF73: dout <= 8'b11111111; // 3955 : 255 - 0xff
      12'hF74: dout <= 8'b11111111; // 3956 : 255 - 0xff
      12'hF75: dout <= 8'b11111111; // 3957 : 255 - 0xff
      12'hF76: dout <= 8'b11111111; // 3958 : 255 - 0xff
      12'hF77: dout <= 8'b11111111; // 3959 : 255 - 0xff
      12'hF78: dout <= 8'b11111111; // 3960 : 255 - 0xff -- plane 1
      12'hF79: dout <= 8'b11111111; // 3961 : 255 - 0xff
      12'hF7A: dout <= 8'b11111111; // 3962 : 255 - 0xff
      12'hF7B: dout <= 8'b11111111; // 3963 : 255 - 0xff
      12'hF7C: dout <= 8'b11111111; // 3964 : 255 - 0xff
      12'hF7D: dout <= 8'b11111111; // 3965 : 255 - 0xff
      12'hF7E: dout <= 8'b11111111; // 3966 : 255 - 0xff
      12'hF7F: dout <= 8'b11111111; // 3967 : 255 - 0xff
      12'hF80: dout <= 8'b11111111; // 3968 : 255 - 0xff -- Sprite 0xf8
      12'hF81: dout <= 8'b11111111; // 3969 : 255 - 0xff
      12'hF82: dout <= 8'b11111111; // 3970 : 255 - 0xff
      12'hF83: dout <= 8'b11111111; // 3971 : 255 - 0xff
      12'hF84: dout <= 8'b11111111; // 3972 : 255 - 0xff
      12'hF85: dout <= 8'b11111111; // 3973 : 255 - 0xff
      12'hF86: dout <= 8'b11111111; // 3974 : 255 - 0xff
      12'hF87: dout <= 8'b11111111; // 3975 : 255 - 0xff
      12'hF88: dout <= 8'b11111111; // 3976 : 255 - 0xff -- plane 1
      12'hF89: dout <= 8'b11111111; // 3977 : 255 - 0xff
      12'hF8A: dout <= 8'b11111111; // 3978 : 255 - 0xff
      12'hF8B: dout <= 8'b11111111; // 3979 : 255 - 0xff
      12'hF8C: dout <= 8'b11111111; // 3980 : 255 - 0xff
      12'hF8D: dout <= 8'b11111111; // 3981 : 255 - 0xff
      12'hF8E: dout <= 8'b11111111; // 3982 : 255 - 0xff
      12'hF8F: dout <= 8'b11111111; // 3983 : 255 - 0xff
      12'hF90: dout <= 8'b11111111; // 3984 : 255 - 0xff -- Sprite 0xf9
      12'hF91: dout <= 8'b11111111; // 3985 : 255 - 0xff
      12'hF92: dout <= 8'b11111111; // 3986 : 255 - 0xff
      12'hF93: dout <= 8'b11111111; // 3987 : 255 - 0xff
      12'hF94: dout <= 8'b11111111; // 3988 : 255 - 0xff
      12'hF95: dout <= 8'b11111111; // 3989 : 255 - 0xff
      12'hF96: dout <= 8'b11111111; // 3990 : 255 - 0xff
      12'hF97: dout <= 8'b11111111; // 3991 : 255 - 0xff
      12'hF98: dout <= 8'b11111111; // 3992 : 255 - 0xff -- plane 1
      12'hF99: dout <= 8'b11111111; // 3993 : 255 - 0xff
      12'hF9A: dout <= 8'b11111111; // 3994 : 255 - 0xff
      12'hF9B: dout <= 8'b11111111; // 3995 : 255 - 0xff
      12'hF9C: dout <= 8'b11111111; // 3996 : 255 - 0xff
      12'hF9D: dout <= 8'b11111111; // 3997 : 255 - 0xff
      12'hF9E: dout <= 8'b11111111; // 3998 : 255 - 0xff
      12'hF9F: dout <= 8'b11111111; // 3999 : 255 - 0xff
      12'hFA0: dout <= 8'b11111111; // 4000 : 255 - 0xff -- Sprite 0xfa
      12'hFA1: dout <= 8'b11111111; // 4001 : 255 - 0xff
      12'hFA2: dout <= 8'b11111111; // 4002 : 255 - 0xff
      12'hFA3: dout <= 8'b11111111; // 4003 : 255 - 0xff
      12'hFA4: dout <= 8'b11111111; // 4004 : 255 - 0xff
      12'hFA5: dout <= 8'b11111111; // 4005 : 255 - 0xff
      12'hFA6: dout <= 8'b11111111; // 4006 : 255 - 0xff
      12'hFA7: dout <= 8'b11111111; // 4007 : 255 - 0xff
      12'hFA8: dout <= 8'b11111111; // 4008 : 255 - 0xff -- plane 1
      12'hFA9: dout <= 8'b11111111; // 4009 : 255 - 0xff
      12'hFAA: dout <= 8'b11111111; // 4010 : 255 - 0xff
      12'hFAB: dout <= 8'b11111111; // 4011 : 255 - 0xff
      12'hFAC: dout <= 8'b11111111; // 4012 : 255 - 0xff
      12'hFAD: dout <= 8'b11111111; // 4013 : 255 - 0xff
      12'hFAE: dout <= 8'b11111111; // 4014 : 255 - 0xff
      12'hFAF: dout <= 8'b11111111; // 4015 : 255 - 0xff
      12'hFB0: dout <= 8'b11111111; // 4016 : 255 - 0xff -- Sprite 0xfb
      12'hFB1: dout <= 8'b11111111; // 4017 : 255 - 0xff
      12'hFB2: dout <= 8'b11111111; // 4018 : 255 - 0xff
      12'hFB3: dout <= 8'b11111111; // 4019 : 255 - 0xff
      12'hFB4: dout <= 8'b11111111; // 4020 : 255 - 0xff
      12'hFB5: dout <= 8'b11111111; // 4021 : 255 - 0xff
      12'hFB6: dout <= 8'b11111111; // 4022 : 255 - 0xff
      12'hFB7: dout <= 8'b11111111; // 4023 : 255 - 0xff
      12'hFB8: dout <= 8'b11111111; // 4024 : 255 - 0xff -- plane 1
      12'hFB9: dout <= 8'b11111111; // 4025 : 255 - 0xff
      12'hFBA: dout <= 8'b11111111; // 4026 : 255 - 0xff
      12'hFBB: dout <= 8'b11111111; // 4027 : 255 - 0xff
      12'hFBC: dout <= 8'b11111111; // 4028 : 255 - 0xff
      12'hFBD: dout <= 8'b11111111; // 4029 : 255 - 0xff
      12'hFBE: dout <= 8'b11111111; // 4030 : 255 - 0xff
      12'hFBF: dout <= 8'b11111111; // 4031 : 255 - 0xff
      12'hFC0: dout <= 8'b11111111; // 4032 : 255 - 0xff -- Sprite 0xfc
      12'hFC1: dout <= 8'b11111111; // 4033 : 255 - 0xff
      12'hFC2: dout <= 8'b11111111; // 4034 : 255 - 0xff
      12'hFC3: dout <= 8'b11111111; // 4035 : 255 - 0xff
      12'hFC4: dout <= 8'b11111111; // 4036 : 255 - 0xff
      12'hFC5: dout <= 8'b11111111; // 4037 : 255 - 0xff
      12'hFC6: dout <= 8'b11111111; // 4038 : 255 - 0xff
      12'hFC7: dout <= 8'b11111111; // 4039 : 255 - 0xff
      12'hFC8: dout <= 8'b11111111; // 4040 : 255 - 0xff -- plane 1
      12'hFC9: dout <= 8'b11111111; // 4041 : 255 - 0xff
      12'hFCA: dout <= 8'b11111111; // 4042 : 255 - 0xff
      12'hFCB: dout <= 8'b11111111; // 4043 : 255 - 0xff
      12'hFCC: dout <= 8'b11111111; // 4044 : 255 - 0xff
      12'hFCD: dout <= 8'b11111111; // 4045 : 255 - 0xff
      12'hFCE: dout <= 8'b11111111; // 4046 : 255 - 0xff
      12'hFCF: dout <= 8'b11111111; // 4047 : 255 - 0xff
      12'hFD0: dout <= 8'b11111111; // 4048 : 255 - 0xff -- Sprite 0xfd
      12'hFD1: dout <= 8'b11111111; // 4049 : 255 - 0xff
      12'hFD2: dout <= 8'b11111111; // 4050 : 255 - 0xff
      12'hFD3: dout <= 8'b11111111; // 4051 : 255 - 0xff
      12'hFD4: dout <= 8'b11111111; // 4052 : 255 - 0xff
      12'hFD5: dout <= 8'b11111111; // 4053 : 255 - 0xff
      12'hFD6: dout <= 8'b11111111; // 4054 : 255 - 0xff
      12'hFD7: dout <= 8'b11111111; // 4055 : 255 - 0xff
      12'hFD8: dout <= 8'b11111111; // 4056 : 255 - 0xff -- plane 1
      12'hFD9: dout <= 8'b11111111; // 4057 : 255 - 0xff
      12'hFDA: dout <= 8'b11111111; // 4058 : 255 - 0xff
      12'hFDB: dout <= 8'b11111111; // 4059 : 255 - 0xff
      12'hFDC: dout <= 8'b11111111; // 4060 : 255 - 0xff
      12'hFDD: dout <= 8'b11111111; // 4061 : 255 - 0xff
      12'hFDE: dout <= 8'b11111111; // 4062 : 255 - 0xff
      12'hFDF: dout <= 8'b11111111; // 4063 : 255 - 0xff
      12'hFE0: dout <= 8'b11111111; // 4064 : 255 - 0xff -- Sprite 0xfe
      12'hFE1: dout <= 8'b11111111; // 4065 : 255 - 0xff
      12'hFE2: dout <= 8'b11111111; // 4066 : 255 - 0xff
      12'hFE3: dout <= 8'b11111111; // 4067 : 255 - 0xff
      12'hFE4: dout <= 8'b11111111; // 4068 : 255 - 0xff
      12'hFE5: dout <= 8'b11111111; // 4069 : 255 - 0xff
      12'hFE6: dout <= 8'b11111111; // 4070 : 255 - 0xff
      12'hFE7: dout <= 8'b11111111; // 4071 : 255 - 0xff
      12'hFE8: dout <= 8'b11111111; // 4072 : 255 - 0xff -- plane 1
      12'hFE9: dout <= 8'b11111111; // 4073 : 255 - 0xff
      12'hFEA: dout <= 8'b11111111; // 4074 : 255 - 0xff
      12'hFEB: dout <= 8'b11111111; // 4075 : 255 - 0xff
      12'hFEC: dout <= 8'b11111111; // 4076 : 255 - 0xff
      12'hFED: dout <= 8'b11111111; // 4077 : 255 - 0xff
      12'hFEE: dout <= 8'b11111111; // 4078 : 255 - 0xff
      12'hFEF: dout <= 8'b11111111; // 4079 : 255 - 0xff
      12'hFF0: dout <= 8'b11111111; // 4080 : 255 - 0xff -- Sprite 0xff
      12'hFF1: dout <= 8'b11111111; // 4081 : 255 - 0xff
      12'hFF2: dout <= 8'b11111111; // 4082 : 255 - 0xff
      12'hFF3: dout <= 8'b11111111; // 4083 : 255 - 0xff
      12'hFF4: dout <= 8'b11111111; // 4084 : 255 - 0xff
      12'hFF5: dout <= 8'b11111111; // 4085 : 255 - 0xff
      12'hFF6: dout <= 8'b11111111; // 4086 : 255 - 0xff
      12'hFF7: dout <= 8'b11111111; // 4087 : 255 - 0xff
      12'hFF8: dout <= 8'b11111111; // 4088 : 255 - 0xff -- plane 1
      12'hFF9: dout <= 8'b11111111; // 4089 : 255 - 0xff
      12'hFFA: dout <= 8'b11111111; // 4090 : 255 - 0xff
      12'hFFB: dout <= 8'b11111111; // 4091 : 255 - 0xff
      12'hFFC: dout <= 8'b11111111; // 4092 : 255 - 0xff
      12'hFFD: dout <= 8'b11111111; // 4093 : 255 - 0xff
      12'hFFE: dout <= 8'b11111111; // 4094 : 255 - 0xff
      12'hFFF: dout <= 8'b11111111; // 4095 : 255 - 0xff
    endcase
  end

endmodule
