--------------------------------------------------------------------------------
-- Felipe Machado Sanchez
-- Departameto de Tecnologia Electronica
-- Universidad Rey Juan Carlos
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package PKG_ROM_MONSTER_3x4 is

  --signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(4-1 downto 0);
  constant monster_blue : memostruct := (
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1100",
       "1011",
       "1011",
       "1100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0111",
       "0011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0011",
       "0111",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0100",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "1011",
       "1111",
       "1111",
       "1101",
       "0111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "1011",
       "1111",
       "1111",
       "1101",
       "0111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0010",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0010",
       "0010",
       "0010",
       "0010",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0010",
       "0010",
       "0010",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0010",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1100",
       "1011",
       "1011",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0010",
       "0010",
       "0010",
       "0110",
       "1100",
       "1011",
       "1011",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0010",
       "0010",
       "0010",
       "0010",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "1011",
       "1011",
       "1011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0010",
       "0010",
       "0110",
       "1011",
       "1011",
       "1011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "1011",
       "1011",
       "1011",
       "1011",
       "1110",
       "1111",
       "1111",
       "1111",
       "1100",
       "0010",
       "0010",
       "0010",
       "0101",
       "1011",
       "1011",
       "1011",
       "1011",
       "1110",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1111",
       "1111",
       "1111",
       "1101",
       "0100",
       "1011",
       "1011",
       "1011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0010",
       "0010",
       "0010",
       "0100",
       "1011",
       "1011",
       "1011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1101",
       "1111",
       "1111",
       "1100",
       "0010",
       "1100",
       "1011",
       "1011",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0010",
       "0010",
       "0010",
       "0010",
       "1100",
       "1011",
       "1011",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1011",
       "1111",
       "1111",
       "1010",
       "0010",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1010",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0100",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1001",
       "1111",
       "1111",
       "0111",
       "0010",
       "0010",
       "0010",
       "0100",
       "0111",
       "1000",
       "0101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "0111",
       "1000",
       "0101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0111",
       "1111",
       "1111",
       "0110",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0110",
       "1111",
       "1111",
       "0101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0101",
       "1111",
       "1111",
       "0100",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "1111",
       "1111",
       "0011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0011",
       "1111",
       "1111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1111",
       "1111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1111",
       "1111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1110",
       "1110",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1110",
       "1101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1101",
       "1101",
       "0010",
       "0010",
       "0100",
       "1100",
       "1111",
       "1101",
       "0101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0111",
       "1110",
       "1110",
       "1000",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0101",
       "1101",
       "1111",
       "1100",
       "0100",
       "0010",
       "0010",
       "1101",
       "1100",
       "0010",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "0010",
       "0010",
       "0010",
       "0010",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0010",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0010",
       "1100",
       "1101",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0011",
       "0100",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0100",
       "0011",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111"
        );

  constant  monster_green : memostruct := (
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1100",
       "1011",
       "1011",
       "1100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0111",
       "0011",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "0110",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0100",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "1011",
       "1111",
       "1111",
       "1101",
       "0111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "1011",
       "1111",
       "1111",
       "1101",
       "0111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0001",
       "0001",
       "0001",
       "0001",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0001",
       "0001",
       "0001",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0001",
       "0001",
       "0001",
       "0011",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1001",
       "0111",
       "0111",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0001",
       "0001",
       "0001",
       "0110",
       "1001",
       "0111",
       "0111",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0001",
       "0001",
       "0001",
       "0001",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0111",
       "0111",
       "0111",
       "0111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1101",
       "0001",
       "0001",
       "0001",
       "0101",
       "0111",
       "0111",
       "0111",
       "0111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0111",
       "0111",
       "0111",
       "0111",
       "1101",
       "1111",
       "1111",
       "1111",
       "1100",
       "0001",
       "0001",
       "0001",
       "0011",
       "0111",
       "0111",
       "0111",
       "0111",
       "1101",
       "1111",
       "1111",
       "1111",
       "1100",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1111",
       "1111",
       "1111",
       "1101",
       "0011",
       "0111",
       "0111",
       "0111",
       "0111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1010",
       "0001",
       "0001",
       "0001",
       "0011",
       "0111",
       "0111",
       "0111",
       "0111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1011",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1101",
       "1111",
       "1111",
       "1011",
       "0010",
       "1001",
       "0111",
       "0111",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0001",
       "0001",
       "0001",
       "0010",
       "1001",
       "0111",
       "0111",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1011",
       "1111",
       "1111",
       "1010",
       "0001",
       "1000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0001",
       "0001",
       "0001",
       "0001",
       "1000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1010",
       "1111",
       "1111",
       "1001",
       "0001",
       "0001",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0011",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0011",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1000",
       "1111",
       "1111",
       "0111",
       "0001",
       "0001",
       "0001",
       "0011",
       "0111",
       "0111",
       "0101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "0111",
       "0111",
       "0101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0111",
       "1111",
       "1111",
       "0110",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0110",
       "1111",
       "1111",
       "0101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0101",
       "1111",
       "1111",
       "0100",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0100",
       "1111",
       "1111",
       "0011",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "1111",
       "1111",
       "0010",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0010",
       "1111",
       "1111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1111",
       "1111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1110",
       "1110",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1110",
       "1101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1101",
       "1101",
       "0001",
       "0001",
       "0011",
       "1011",
       "1111",
       "1101",
       "0101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0111",
       "1110",
       "1110",
       "0111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0101",
       "1101",
       "1111",
       "1100",
       "0100",
       "0001",
       "0001",
       "1100",
       "1100",
       "0001",
       "0100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "0001",
       "0001",
       "0001",
       "0001",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0001",
       "0001",
       "0001",
       "0001",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0001",
       "1100",
       "1101",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0011",
       "0011",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0011",
       "0011",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111"
        );


  constant monster_red : memostruct := (
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1100",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0000",
       "0000",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "0100",
       "0000",
       "0000",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0000",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1011",
       "0000",
       "0000",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0000",
       "0000",
       "0000",
       "0000",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1001",
       "0000",
       "0000",
       "0000",
       "0000",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0000",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1011",
       "0000",
       "0000",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "0110",
       "0000",
       "0000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "0110",
       "0000",
       "0000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111"
        );



end PKG_ROM_MONSTER_3x4;

