//-   Sprites Pattern table COLOR PLANE 0
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: smario_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_SMARIO_SPR_PLN0
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table COLOR PLANE 0
      11'h0: dout  = 8'b00000011; //    0 :   3 - 0x3 -- Sprite 0x0
      11'h1: dout  = 8'b00001111; //    1 :  15 - 0xf
      11'h2: dout  = 8'b00011111; //    2 :  31 - 0x1f
      11'h3: dout  = 8'b00011111; //    3 :  31 - 0x1f
      11'h4: dout  = 8'b00011100; //    4 :  28 - 0x1c
      11'h5: dout  = 8'b00100100; //    5 :  36 - 0x24
      11'h6: dout  = 8'b00100110; //    6 :  38 - 0x26
      11'h7: dout  = 8'b01100110; //    7 : 102 - 0x66
      11'h8: dout  = 8'b11100000; //    8 : 224 - 0xe0 -- Sprite 0x1
      11'h9: dout  = 8'b11000000; //    9 : 192 - 0xc0
      11'hA: dout  = 8'b10000000; //   10 : 128 - 0x80
      11'hB: dout  = 8'b11111100; //   11 : 252 - 0xfc
      11'hC: dout  = 8'b10000000; //   12 : 128 - 0x80
      11'hD: dout  = 8'b11000000; //   13 : 192 - 0xc0
      11'hE: dout  = 8'b00000000; //   14 :   0 - 0x0
      11'hF: dout  = 8'b00100000; //   15 :  32 - 0x20
      11'h10: dout  = 8'b01100000; //   16 :  96 - 0x60 -- Sprite 0x2
      11'h11: dout  = 8'b01110000; //   17 : 112 - 0x70
      11'h12: dout  = 8'b00011000; //   18 :  24 - 0x18
      11'h13: dout  = 8'b00000111; //   19 :   7 - 0x7
      11'h14: dout  = 8'b00001111; //   20 :  15 - 0xf
      11'h15: dout  = 8'b00011111; //   21 :  31 - 0x1f
      11'h16: dout  = 8'b00111111; //   22 :  63 - 0x3f
      11'h17: dout  = 8'b01111111; //   23 : 127 - 0x7f
      11'h18: dout  = 8'b11111100; //   24 : 252 - 0xfc -- Sprite 0x3
      11'h19: dout  = 8'b01111100; //   25 : 124 - 0x7c
      11'h1A: dout  = 8'b00000000; //   26 :   0 - 0x0
      11'h1B: dout  = 8'b00000000; //   27 :   0 - 0x0
      11'h1C: dout  = 8'b11100000; //   28 : 224 - 0xe0
      11'h1D: dout  = 8'b11110000; //   29 : 240 - 0xf0
      11'h1E: dout  = 8'b11111000; //   30 : 248 - 0xf8
      11'h1F: dout  = 8'b11111000; //   31 : 248 - 0xf8
      11'h20: dout  = 8'b01111111; //   32 : 127 - 0x7f -- Sprite 0x4
      11'h21: dout  = 8'b01111111; //   33 : 127 - 0x7f
      11'h22: dout  = 8'b11111111; //   34 : 255 - 0xff
      11'h23: dout  = 8'b11111111; //   35 : 255 - 0xff
      11'h24: dout  = 8'b00000111; //   36 :   7 - 0x7
      11'h25: dout  = 8'b00000111; //   37 :   7 - 0x7
      11'h26: dout  = 8'b00001111; //   38 :  15 - 0xf
      11'h27: dout  = 8'b00001111; //   39 :  15 - 0xf
      11'h28: dout  = 8'b11111101; //   40 : 253 - 0xfd -- Sprite 0x5
      11'h29: dout  = 8'b11111110; //   41 : 254 - 0xfe
      11'h2A: dout  = 8'b10110100; //   42 : 180 - 0xb4
      11'h2B: dout  = 8'b11111000; //   43 : 248 - 0xf8
      11'h2C: dout  = 8'b11111000; //   44 : 248 - 0xf8
      11'h2D: dout  = 8'b11111001; //   45 : 249 - 0xf9
      11'h2E: dout  = 8'b11111011; //   46 : 251 - 0xfb
      11'h2F: dout  = 8'b11111111; //   47 : 255 - 0xff
      11'h30: dout  = 8'b00011111; //   48 :  31 - 0x1f -- Sprite 0x6
      11'h31: dout  = 8'b00111111; //   49 :  63 - 0x3f
      11'h32: dout  = 8'b11111111; //   50 : 255 - 0xff
      11'h33: dout  = 8'b11111111; //   51 : 255 - 0xff
      11'h34: dout  = 8'b11111100; //   52 : 252 - 0xfc
      11'h35: dout  = 8'b01110000; //   53 : 112 - 0x70
      11'h36: dout  = 8'b01110000; //   54 : 112 - 0x70
      11'h37: dout  = 8'b00111000; //   55 :  56 - 0x38
      11'h38: dout  = 8'b11111111; //   56 : 255 - 0xff -- Sprite 0x7
      11'h39: dout  = 8'b11111111; //   57 : 255 - 0xff
      11'h3A: dout  = 8'b11111111; //   58 : 255 - 0xff
      11'h3B: dout  = 8'b00011111; //   59 :  31 - 0x1f
      11'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      11'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      11'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      11'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      11'h40: dout  = 8'b00000000; //   64 :   0 - 0x0 -- Sprite 0x8
      11'h41: dout  = 8'b00000000; //   65 :   0 - 0x0
      11'h42: dout  = 8'b00000001; //   66 :   1 - 0x1
      11'h43: dout  = 8'b00000111; //   67 :   7 - 0x7
      11'h44: dout  = 8'b00001111; //   68 :  15 - 0xf
      11'h45: dout  = 8'b00001111; //   69 :  15 - 0xf
      11'h46: dout  = 8'b00001110; //   70 :  14 - 0xe
      11'h47: dout  = 8'b00010010; //   71 :  18 - 0x12
      11'h48: dout  = 8'b00000000; //   72 :   0 - 0x0 -- Sprite 0x9
      11'h49: dout  = 8'b00000000; //   73 :   0 - 0x0
      11'h4A: dout  = 8'b11110000; //   74 : 240 - 0xf0
      11'h4B: dout  = 8'b11100000; //   75 : 224 - 0xe0
      11'h4C: dout  = 8'b11000000; //   76 : 192 - 0xc0
      11'h4D: dout  = 8'b11111110; //   77 : 254 - 0xfe
      11'h4E: dout  = 8'b01000000; //   78 :  64 - 0x40
      11'h4F: dout  = 8'b01100000; //   79 :  96 - 0x60
      11'h50: dout  = 8'b00010011; //   80 :  19 - 0x13 -- Sprite 0xa
      11'h51: dout  = 8'b00110011; //   81 :  51 - 0x33
      11'h52: dout  = 8'b00110000; //   82 :  48 - 0x30
      11'h53: dout  = 8'b00011000; //   83 :  24 - 0x18
      11'h54: dout  = 8'b00000100; //   84 :   4 - 0x4
      11'h55: dout  = 8'b00001111; //   85 :  15 - 0xf
      11'h56: dout  = 8'b00011111; //   86 :  31 - 0x1f
      11'h57: dout  = 8'b00011111; //   87 :  31 - 0x1f
      11'h58: dout  = 8'b00000000; //   88 :   0 - 0x0 -- Sprite 0xb
      11'h59: dout  = 8'b00010000; //   89 :  16 - 0x10
      11'h5A: dout  = 8'b01111110; //   90 : 126 - 0x7e
      11'h5B: dout  = 8'b00111110; //   91 :  62 - 0x3e
      11'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      11'h5D: dout  = 8'b00000000; //   93 :   0 - 0x0
      11'h5E: dout  = 8'b11000000; //   94 : 192 - 0xc0
      11'h5F: dout  = 8'b11100000; //   95 : 224 - 0xe0
      11'h60: dout  = 8'b00111111; //   96 :  63 - 0x3f -- Sprite 0xc
      11'h61: dout  = 8'b00111111; //   97 :  63 - 0x3f
      11'h62: dout  = 8'b00111111; //   98 :  63 - 0x3f
      11'h63: dout  = 8'b00011111; //   99 :  31 - 0x1f
      11'h64: dout  = 8'b00011111; //  100 :  31 - 0x1f
      11'h65: dout  = 8'b00011111; //  101 :  31 - 0x1f
      11'h66: dout  = 8'b00011111; //  102 :  31 - 0x1f
      11'h67: dout  = 8'b00011111; //  103 :  31 - 0x1f
      11'h68: dout  = 8'b11110000; //  104 : 240 - 0xf0 -- Sprite 0xd
      11'h69: dout  = 8'b11110000; //  105 : 240 - 0xf0
      11'h6A: dout  = 8'b11110000; //  106 : 240 - 0xf0
      11'h6B: dout  = 8'b11111000; //  107 : 248 - 0xf8
      11'h6C: dout  = 8'b11111000; //  108 : 248 - 0xf8
      11'h6D: dout  = 8'b11111000; //  109 : 248 - 0xf8
      11'h6E: dout  = 8'b11111000; //  110 : 248 - 0xf8
      11'h6F: dout  = 8'b11111000; //  111 : 248 - 0xf8
      11'h70: dout  = 8'b11111111; //  112 : 255 - 0xff -- Sprite 0xe
      11'h71: dout  = 8'b11111111; //  113 : 255 - 0xff
      11'h72: dout  = 8'b11111111; //  114 : 255 - 0xff
      11'h73: dout  = 8'b11111110; //  115 : 254 - 0xfe
      11'h74: dout  = 8'b11110000; //  116 : 240 - 0xf0
      11'h75: dout  = 8'b11000000; //  117 : 192 - 0xc0
      11'h76: dout  = 8'b10000000; //  118 : 128 - 0x80
      11'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      11'h78: dout  = 8'b11111100; //  120 : 252 - 0xfc -- Sprite 0xf
      11'h79: dout  = 8'b11111100; //  121 : 252 - 0xfc
      11'h7A: dout  = 8'b11111000; //  122 : 248 - 0xf8
      11'h7B: dout  = 8'b01111000; //  123 : 120 - 0x78
      11'h7C: dout  = 8'b01111000; //  124 : 120 - 0x78
      11'h7D: dout  = 8'b01111000; //  125 : 120 - 0x78
      11'h7E: dout  = 8'b01111110; //  126 : 126 - 0x7e
      11'h7F: dout  = 8'b01111110; //  127 : 126 - 0x7e
      11'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      11'h81: dout  = 8'b00000011; //  129 :   3 - 0x3
      11'h82: dout  = 8'b00001111; //  130 :  15 - 0xf
      11'h83: dout  = 8'b00011111; //  131 :  31 - 0x1f
      11'h84: dout  = 8'b00011111; //  132 :  31 - 0x1f
      11'h85: dout  = 8'b00011100; //  133 :  28 - 0x1c
      11'h86: dout  = 8'b00100100; //  134 :  36 - 0x24
      11'h87: dout  = 8'b00100110; //  135 :  38 - 0x26
      11'h88: dout  = 8'b00000000; //  136 :   0 - 0x0 -- Sprite 0x11
      11'h89: dout  = 8'b11100000; //  137 : 224 - 0xe0
      11'h8A: dout  = 8'b11000000; //  138 : 192 - 0xc0
      11'h8B: dout  = 8'b10000000; //  139 : 128 - 0x80
      11'h8C: dout  = 8'b11111100; //  140 : 252 - 0xfc
      11'h8D: dout  = 8'b10000000; //  141 : 128 - 0x80
      11'h8E: dout  = 8'b11000000; //  142 : 192 - 0xc0
      11'h8F: dout  = 8'b00000000; //  143 :   0 - 0x0
      11'h90: dout  = 8'b01100110; //  144 : 102 - 0x66 -- Sprite 0x12
      11'h91: dout  = 8'b01100000; //  145 :  96 - 0x60
      11'h92: dout  = 8'b00110000; //  146 :  48 - 0x30
      11'h93: dout  = 8'b00011000; //  147 :  24 - 0x18
      11'h94: dout  = 8'b00001111; //  148 :  15 - 0xf
      11'h95: dout  = 8'b00011111; //  149 :  31 - 0x1f
      11'h96: dout  = 8'b00111111; //  150 :  63 - 0x3f
      11'h97: dout  = 8'b00111111; //  151 :  63 - 0x3f
      11'h98: dout  = 8'b00100000; //  152 :  32 - 0x20 -- Sprite 0x13
      11'h99: dout  = 8'b11111100; //  153 : 252 - 0xfc
      11'h9A: dout  = 8'b01111100; //  154 : 124 - 0x7c
      11'h9B: dout  = 8'b00000000; //  155 :   0 - 0x0
      11'h9C: dout  = 8'b00000000; //  156 :   0 - 0x0
      11'h9D: dout  = 8'b11100000; //  157 : 224 - 0xe0
      11'h9E: dout  = 8'b11100000; //  158 : 224 - 0xe0
      11'h9F: dout  = 8'b11110000; //  159 : 240 - 0xf0
      11'hA0: dout  = 8'b00111111; //  160 :  63 - 0x3f -- Sprite 0x14
      11'hA1: dout  = 8'b00111111; //  161 :  63 - 0x3f
      11'hA2: dout  = 8'b00111111; //  162 :  63 - 0x3f
      11'hA3: dout  = 8'b00111111; //  163 :  63 - 0x3f
      11'hA4: dout  = 8'b00111111; //  164 :  63 - 0x3f
      11'hA5: dout  = 8'b00111111; //  165 :  63 - 0x3f
      11'hA6: dout  = 8'b00111111; //  166 :  63 - 0x3f
      11'hA7: dout  = 8'b00011111; //  167 :  31 - 0x1f
      11'hA8: dout  = 8'b11110000; //  168 : 240 - 0xf0 -- Sprite 0x15
      11'hA9: dout  = 8'b10010000; //  169 : 144 - 0x90
      11'hAA: dout  = 8'b00000000; //  170 :   0 - 0x0
      11'hAB: dout  = 8'b00001000; //  171 :   8 - 0x8
      11'hAC: dout  = 8'b00001100; //  172 :  12 - 0xc
      11'hAD: dout  = 8'b00011100; //  173 :  28 - 0x1c
      11'hAE: dout  = 8'b11111100; //  174 : 252 - 0xfc
      11'hAF: dout  = 8'b11111000; //  175 : 248 - 0xf8
      11'hB0: dout  = 8'b00001111; //  176 :  15 - 0xf -- Sprite 0x16
      11'hB1: dout  = 8'b00001111; //  177 :  15 - 0xf
      11'hB2: dout  = 8'b00000111; //  178 :   7 - 0x7
      11'hB3: dout  = 8'b00000111; //  179 :   7 - 0x7
      11'hB4: dout  = 8'b00000111; //  180 :   7 - 0x7
      11'hB5: dout  = 8'b00001111; //  181 :  15 - 0xf
      11'hB6: dout  = 8'b00001111; //  182 :  15 - 0xf
      11'hB7: dout  = 8'b00000011; //  183 :   3 - 0x3
      11'hB8: dout  = 8'b11111000; //  184 : 248 - 0xf8 -- Sprite 0x17
      11'hB9: dout  = 8'b11110000; //  185 : 240 - 0xf0
      11'hBA: dout  = 8'b11100000; //  186 : 224 - 0xe0
      11'hBB: dout  = 8'b11110000; //  187 : 240 - 0xf0
      11'hBC: dout  = 8'b10110000; //  188 : 176 - 0xb0
      11'hBD: dout  = 8'b10000000; //  189 : 128 - 0x80
      11'hBE: dout  = 8'b11100000; //  190 : 224 - 0xe0
      11'hBF: dout  = 8'b11100000; //  191 : 224 - 0xe0
      11'hC0: dout  = 8'b00000011; //  192 :   3 - 0x3 -- Sprite 0x18
      11'hC1: dout  = 8'b00111111; //  193 :  63 - 0x3f
      11'hC2: dout  = 8'b01111111; //  194 : 127 - 0x7f
      11'hC3: dout  = 8'b00011001; //  195 :  25 - 0x19
      11'hC4: dout  = 8'b00001001; //  196 :   9 - 0x9
      11'hC5: dout  = 8'b00001001; //  197 :   9 - 0x9
      11'hC6: dout  = 8'b00101000; //  198 :  40 - 0x28
      11'hC7: dout  = 8'b01011100; //  199 :  92 - 0x5c
      11'hC8: dout  = 8'b11111000; //  200 : 248 - 0xf8 -- Sprite 0x19
      11'hC9: dout  = 8'b11100000; //  201 : 224 - 0xe0
      11'hCA: dout  = 8'b11100000; //  202 : 224 - 0xe0
      11'hCB: dout  = 8'b11111100; //  203 : 252 - 0xfc
      11'hCC: dout  = 8'b00100110; //  204 :  38 - 0x26
      11'hCD: dout  = 8'b00110000; //  205 :  48 - 0x30
      11'hCE: dout  = 8'b10000000; //  206 : 128 - 0x80
      11'hCF: dout  = 8'b00010000; //  207 :  16 - 0x10
      11'hD0: dout  = 8'b00111110; //  208 :  62 - 0x3e -- Sprite 0x1a
      11'hD1: dout  = 8'b00011110; //  209 :  30 - 0x1e
      11'hD2: dout  = 8'b00111111; //  210 :  63 - 0x3f
      11'hD3: dout  = 8'b00111000; //  211 :  56 - 0x38
      11'hD4: dout  = 8'b00110000; //  212 :  48 - 0x30
      11'hD5: dout  = 8'b00110000; //  213 :  48 - 0x30
      11'hD6: dout  = 8'b00000000; //  214 :   0 - 0x0
      11'hD7: dout  = 8'b00111010; //  215 :  58 - 0x3a
      11'hD8: dout  = 8'b01111000; //  216 : 120 - 0x78 -- Sprite 0x1b
      11'hD9: dout  = 8'b00011110; //  217 :  30 - 0x1e
      11'hDA: dout  = 8'b10000000; //  218 : 128 - 0x80
      11'hDB: dout  = 8'b11111110; //  219 : 254 - 0xfe
      11'hDC: dout  = 8'b01111110; //  220 : 126 - 0x7e
      11'hDD: dout  = 8'b01111110; //  221 : 126 - 0x7e
      11'hDE: dout  = 8'b01111111; //  222 : 127 - 0x7f
      11'hDF: dout  = 8'b01111111; //  223 : 127 - 0x7f
      11'hE0: dout  = 8'b00111100; //  224 :  60 - 0x3c -- Sprite 0x1c
      11'hE1: dout  = 8'b00111111; //  225 :  63 - 0x3f
      11'hE2: dout  = 8'b00011111; //  226 :  31 - 0x1f
      11'hE3: dout  = 8'b00001111; //  227 :  15 - 0xf
      11'hE4: dout  = 8'b00000111; //  228 :   7 - 0x7
      11'hE5: dout  = 8'b00111111; //  229 :  63 - 0x3f
      11'hE6: dout  = 8'b00100001; //  230 :  33 - 0x21
      11'hE7: dout  = 8'b00100000; //  231 :  32 - 0x20
      11'hE8: dout  = 8'b11111111; //  232 : 255 - 0xff -- Sprite 0x1d
      11'hE9: dout  = 8'b11111111; //  233 : 255 - 0xff
      11'hEA: dout  = 8'b11111111; //  234 : 255 - 0xff
      11'hEB: dout  = 8'b11111110; //  235 : 254 - 0xfe
      11'hEC: dout  = 8'b11111110; //  236 : 254 - 0xfe
      11'hED: dout  = 8'b11111110; //  237 : 254 - 0xfe
      11'hEE: dout  = 8'b11111100; //  238 : 252 - 0xfc
      11'hEF: dout  = 8'b01110000; //  239 : 112 - 0x70
      11'hF0: dout  = 8'b00001111; //  240 :  15 - 0xf -- Sprite 0x1e
      11'hF1: dout  = 8'b10011111; //  241 : 159 - 0x9f
      11'hF2: dout  = 8'b11001111; //  242 : 207 - 0xcf
      11'hF3: dout  = 8'b11111111; //  243 : 255 - 0xff
      11'hF4: dout  = 8'b01111111; //  244 : 127 - 0x7f
      11'hF5: dout  = 8'b00111111; //  245 :  63 - 0x3f
      11'hF6: dout  = 8'b00011110; //  246 :  30 - 0x1e
      11'hF7: dout  = 8'b00001110; //  247 :  14 - 0xe
      11'hF8: dout  = 8'b00100000; //  248 :  32 - 0x20 -- Sprite 0x1f
      11'hF9: dout  = 8'b11000000; //  249 : 192 - 0xc0
      11'hFA: dout  = 8'b10000000; //  250 : 128 - 0x80
      11'hFB: dout  = 8'b10000000; //  251 : 128 - 0x80
      11'hFC: dout  = 8'b00000000; //  252 :   0 - 0x0
      11'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      11'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      11'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      11'h101: dout  = 8'b00000000; //  257 :   0 - 0x0
      11'h102: dout  = 8'b00000011; //  258 :   3 - 0x3
      11'h103: dout  = 8'b00001111; //  259 :  15 - 0xf
      11'h104: dout  = 8'b00011111; //  260 :  31 - 0x1f
      11'h105: dout  = 8'b00011111; //  261 :  31 - 0x1f
      11'h106: dout  = 8'b00011100; //  262 :  28 - 0x1c
      11'h107: dout  = 8'b00100100; //  263 :  36 - 0x24
      11'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- Sprite 0x21
      11'h109: dout  = 8'b00000100; //  265 :   4 - 0x4
      11'h10A: dout  = 8'b11100110; //  266 : 230 - 0xe6
      11'h10B: dout  = 8'b11100000; //  267 : 224 - 0xe0
      11'h10C: dout  = 8'b11111111; //  268 : 255 - 0xff
      11'h10D: dout  = 8'b11111111; //  269 : 255 - 0xff
      11'h10E: dout  = 8'b10001111; //  270 : 143 - 0x8f
      11'h10F: dout  = 8'b10000011; //  271 : 131 - 0x83
      11'h110: dout  = 8'b00100110; //  272 :  38 - 0x26 -- Sprite 0x22
      11'h111: dout  = 8'b00100110; //  273 :  38 - 0x26
      11'h112: dout  = 8'b01100000; //  274 :  96 - 0x60
      11'h113: dout  = 8'b01111000; //  275 : 120 - 0x78
      11'h114: dout  = 8'b00011000; //  276 :  24 - 0x18
      11'h115: dout  = 8'b00001111; //  277 :  15 - 0xf
      11'h116: dout  = 8'b01111111; //  278 : 127 - 0x7f
      11'h117: dout  = 8'b11111111; //  279 : 255 - 0xff
      11'h118: dout  = 8'b00000001; //  280 :   1 - 0x1 -- Sprite 0x23
      11'h119: dout  = 8'b00100001; //  281 :  33 - 0x21
      11'h11A: dout  = 8'b11111110; //  282 : 254 - 0xfe
      11'h11B: dout  = 8'b01111010; //  283 : 122 - 0x7a
      11'h11C: dout  = 8'b00000110; //  284 :   6 - 0x6
      11'h11D: dout  = 8'b11111110; //  285 : 254 - 0xfe
      11'h11E: dout  = 8'b11111100; //  286 : 252 - 0xfc
      11'h11F: dout  = 8'b11111100; //  287 : 252 - 0xfc
      11'h120: dout  = 8'b11111111; //  288 : 255 - 0xff -- Sprite 0x24
      11'h121: dout  = 8'b11001111; //  289 : 207 - 0xcf
      11'h122: dout  = 8'b10000111; //  290 : 135 - 0x87
      11'h123: dout  = 8'b00000111; //  291 :   7 - 0x7
      11'h124: dout  = 8'b00000111; //  292 :   7 - 0x7
      11'h125: dout  = 8'b00001111; //  293 :  15 - 0xf
      11'h126: dout  = 8'b00011111; //  294 :  31 - 0x1f
      11'h127: dout  = 8'b00011111; //  295 :  31 - 0x1f
      11'h128: dout  = 8'b11111000; //  296 : 248 - 0xf8 -- Sprite 0x25
      11'h129: dout  = 8'b11111000; //  297 : 248 - 0xf8
      11'h12A: dout  = 8'b11110000; //  298 : 240 - 0xf0
      11'h12B: dout  = 8'b10111000; //  299 : 184 - 0xb8
      11'h12C: dout  = 8'b11111000; //  300 : 248 - 0xf8
      11'h12D: dout  = 8'b11111001; //  301 : 249 - 0xf9
      11'h12E: dout  = 8'b11111011; //  302 : 251 - 0xfb
      11'h12F: dout  = 8'b11111111; //  303 : 255 - 0xff
      11'h130: dout  = 8'b00011111; //  304 :  31 - 0x1f -- Sprite 0x26
      11'h131: dout  = 8'b11111111; //  305 : 255 - 0xff
      11'h132: dout  = 8'b11111111; //  306 : 255 - 0xff
      11'h133: dout  = 8'b11111111; //  307 : 255 - 0xff
      11'h134: dout  = 8'b11111111; //  308 : 255 - 0xff
      11'h135: dout  = 8'b11111110; //  309 : 254 - 0xfe
      11'h136: dout  = 8'b11000000; //  310 : 192 - 0xc0
      11'h137: dout  = 8'b10000000; //  311 : 128 - 0x80
      11'h138: dout  = 8'b11111111; //  312 : 255 - 0xff -- Sprite 0x27
      11'h139: dout  = 8'b11111111; //  313 : 255 - 0xff
      11'h13A: dout  = 8'b11111111; //  314 : 255 - 0xff
      11'h13B: dout  = 8'b00111111; //  315 :  63 - 0x3f
      11'h13C: dout  = 8'b00000000; //  316 :   0 - 0x0
      11'h13D: dout  = 8'b00000000; //  317 :   0 - 0x0
      11'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      11'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      11'h140: dout  = 8'b00010011; //  320 :  19 - 0x13 -- Sprite 0x28
      11'h141: dout  = 8'b00110011; //  321 :  51 - 0x33
      11'h142: dout  = 8'b00110000; //  322 :  48 - 0x30
      11'h143: dout  = 8'b00011000; //  323 :  24 - 0x18
      11'h144: dout  = 8'b00000100; //  324 :   4 - 0x4
      11'h145: dout  = 8'b00001111; //  325 :  15 - 0xf
      11'h146: dout  = 8'b00011111; //  326 :  31 - 0x1f
      11'h147: dout  = 8'b00011111; //  327 :  31 - 0x1f
      11'h148: dout  = 8'b00000000; //  328 :   0 - 0x0 -- Sprite 0x29
      11'h149: dout  = 8'b00010000; //  329 :  16 - 0x10
      11'h14A: dout  = 8'b01111110; //  330 : 126 - 0x7e
      11'h14B: dout  = 8'b00110000; //  331 :  48 - 0x30
      11'h14C: dout  = 8'b11100000; //  332 : 224 - 0xe0
      11'h14D: dout  = 8'b11110000; //  333 : 240 - 0xf0
      11'h14E: dout  = 8'b11110000; //  334 : 240 - 0xf0
      11'h14F: dout  = 8'b11100000; //  335 : 224 - 0xe0
      11'h150: dout  = 8'b00011111; //  336 :  31 - 0x1f -- Sprite 0x2a
      11'h151: dout  = 8'b00011111; //  337 :  31 - 0x1f
      11'h152: dout  = 8'b00001111; //  338 :  15 - 0xf
      11'h153: dout  = 8'b00001111; //  339 :  15 - 0xf
      11'h154: dout  = 8'b00001111; //  340 :  15 - 0xf
      11'h155: dout  = 8'b00011111; //  341 :  31 - 0x1f
      11'h156: dout  = 8'b00011111; //  342 :  31 - 0x1f
      11'h157: dout  = 8'b00011111; //  343 :  31 - 0x1f
      11'h158: dout  = 8'b11110000; //  344 : 240 - 0xf0 -- Sprite 0x2b
      11'h159: dout  = 8'b11110000; //  345 : 240 - 0xf0
      11'h15A: dout  = 8'b11111000; //  346 : 248 - 0xf8
      11'h15B: dout  = 8'b11111000; //  347 : 248 - 0xf8
      11'h15C: dout  = 8'b10111000; //  348 : 184 - 0xb8
      11'h15D: dout  = 8'b11111000; //  349 : 248 - 0xf8
      11'h15E: dout  = 8'b11111000; //  350 : 248 - 0xf8
      11'h15F: dout  = 8'b11111000; //  351 : 248 - 0xf8
      11'h160: dout  = 8'b00111111; //  352 :  63 - 0x3f -- Sprite 0x2c
      11'h161: dout  = 8'b11111111; //  353 : 255 - 0xff
      11'h162: dout  = 8'b11111111; //  354 : 255 - 0xff
      11'h163: dout  = 8'b11111111; //  355 : 255 - 0xff
      11'h164: dout  = 8'b11110110; //  356 : 246 - 0xf6
      11'h165: dout  = 8'b11000110; //  357 : 198 - 0xc6
      11'h166: dout  = 8'b10000100; //  358 : 132 - 0x84
      11'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      11'h168: dout  = 8'b11110000; //  360 : 240 - 0xf0 -- Sprite 0x2d
      11'h169: dout  = 8'b11100000; //  361 : 224 - 0xe0
      11'h16A: dout  = 8'b10000000; //  362 : 128 - 0x80
      11'h16B: dout  = 8'b00000000; //  363 :   0 - 0x0
      11'h16C: dout  = 8'b00000000; //  364 :   0 - 0x0
      11'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      11'h16E: dout  = 8'b00000000; //  366 :   0 - 0x0
      11'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      11'h170: dout  = 8'b00011111; //  368 :  31 - 0x1f -- Sprite 0x2e
      11'h171: dout  = 8'b00011111; //  369 :  31 - 0x1f
      11'h172: dout  = 8'b00111111; //  370 :  63 - 0x3f
      11'h173: dout  = 8'b00111111; //  371 :  63 - 0x3f
      11'h174: dout  = 8'b00011111; //  372 :  31 - 0x1f
      11'h175: dout  = 8'b00001111; //  373 :  15 - 0xf
      11'h176: dout  = 8'b00001111; //  374 :  15 - 0xf
      11'h177: dout  = 8'b00011111; //  375 :  31 - 0x1f
      11'h178: dout  = 8'b11110000; //  376 : 240 - 0xf0 -- Sprite 0x2f
      11'h179: dout  = 8'b11110000; //  377 : 240 - 0xf0
      11'h17A: dout  = 8'b11111000; //  378 : 248 - 0xf8
      11'h17B: dout  = 8'b11111000; //  379 : 248 - 0xf8
      11'h17C: dout  = 8'b10111000; //  380 : 184 - 0xb8
      11'h17D: dout  = 8'b11111000; //  381 : 248 - 0xf8
      11'h17E: dout  = 8'b11111000; //  382 : 248 - 0xf8
      11'h17F: dout  = 8'b11110000; //  383 : 240 - 0xf0
      11'h180: dout  = 8'b11100000; //  384 : 224 - 0xe0 -- Sprite 0x30
      11'h181: dout  = 8'b11110000; //  385 : 240 - 0xf0
      11'h182: dout  = 8'b11110000; //  386 : 240 - 0xf0
      11'h183: dout  = 8'b11110000; //  387 : 240 - 0xf0
      11'h184: dout  = 8'b11110000; //  388 : 240 - 0xf0
      11'h185: dout  = 8'b11110000; //  389 : 240 - 0xf0
      11'h186: dout  = 8'b11111000; //  390 : 248 - 0xf8
      11'h187: dout  = 8'b11110000; //  391 : 240 - 0xf0
      11'h188: dout  = 8'b00011111; //  392 :  31 - 0x1f -- Sprite 0x31
      11'h189: dout  = 8'b00011111; //  393 :  31 - 0x1f
      11'h18A: dout  = 8'b00011111; //  394 :  31 - 0x1f
      11'h18B: dout  = 8'b00111111; //  395 :  63 - 0x3f
      11'h18C: dout  = 8'b00111110; //  396 :  62 - 0x3e
      11'h18D: dout  = 8'b00111100; //  397 :  60 - 0x3c
      11'h18E: dout  = 8'b00111000; //  398 :  56 - 0x38
      11'h18F: dout  = 8'b00011000; //  399 :  24 - 0x18
      11'h190: dout  = 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      11'h191: dout  = 8'b00000011; //  401 :   3 - 0x3
      11'h192: dout  = 8'b00000111; //  402 :   7 - 0x7
      11'h193: dout  = 8'b00000111; //  403 :   7 - 0x7
      11'h194: dout  = 8'b00001010; //  404 :  10 - 0xa
      11'h195: dout  = 8'b00001011; //  405 :  11 - 0xb
      11'h196: dout  = 8'b00001100; //  406 :  12 - 0xc
      11'h197: dout  = 8'b00000000; //  407 :   0 - 0x0
      11'h198: dout  = 8'b00000000; //  408 :   0 - 0x0 -- Sprite 0x33
      11'h199: dout  = 8'b11100000; //  409 : 224 - 0xe0
      11'h19A: dout  = 8'b11111100; //  410 : 252 - 0xfc
      11'h19B: dout  = 8'b00100000; //  411 :  32 - 0x20
      11'h19C: dout  = 8'b00100000; //  412 :  32 - 0x20
      11'h19D: dout  = 8'b00010000; //  413 :  16 - 0x10
      11'h19E: dout  = 8'b00111100; //  414 :  60 - 0x3c
      11'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      11'h1A0: dout  = 8'b00000111; //  416 :   7 - 0x7 -- Sprite 0x34
      11'h1A1: dout  = 8'b00000111; //  417 :   7 - 0x7
      11'h1A2: dout  = 8'b00000111; //  418 :   7 - 0x7
      11'h1A3: dout  = 8'b00011111; //  419 :  31 - 0x1f
      11'h1A4: dout  = 8'b00011111; //  420 :  31 - 0x1f
      11'h1A5: dout  = 8'b00111110; //  421 :  62 - 0x3e
      11'h1A6: dout  = 8'b00100001; //  422 :  33 - 0x21
      11'h1A7: dout  = 8'b00000001; //  423 :   1 - 0x1
      11'h1A8: dout  = 8'b11100000; //  424 : 224 - 0xe0 -- Sprite 0x35
      11'h1A9: dout  = 8'b11100000; //  425 : 224 - 0xe0
      11'h1AA: dout  = 8'b11100000; //  426 : 224 - 0xe0
      11'h1AB: dout  = 8'b11110000; //  427 : 240 - 0xf0
      11'h1AC: dout  = 8'b11110000; //  428 : 240 - 0xf0
      11'h1AD: dout  = 8'b11100000; //  429 : 224 - 0xe0
      11'h1AE: dout  = 8'b11000000; //  430 : 192 - 0xc0
      11'h1AF: dout  = 8'b11100000; //  431 : 224 - 0xe0
      11'h1B0: dout  = 8'b00000111; //  432 :   7 - 0x7 -- Sprite 0x36
      11'h1B1: dout  = 8'b00001111; //  433 :  15 - 0xf
      11'h1B2: dout  = 8'b00001110; //  434 :  14 - 0xe
      11'h1B3: dout  = 8'b00010100; //  435 :  20 - 0x14
      11'h1B4: dout  = 8'b00010110; //  436 :  22 - 0x16
      11'h1B5: dout  = 8'b00011000; //  437 :  24 - 0x18
      11'h1B6: dout  = 8'b00000000; //  438 :   0 - 0x0
      11'h1B7: dout  = 8'b00111111; //  439 :  63 - 0x3f
      11'h1B8: dout  = 8'b11000000; //  440 : 192 - 0xc0 -- Sprite 0x37
      11'h1B9: dout  = 8'b11111000; //  441 : 248 - 0xf8
      11'h1BA: dout  = 8'b01000000; //  442 :  64 - 0x40
      11'h1BB: dout  = 8'b01000000; //  443 :  64 - 0x40
      11'h1BC: dout  = 8'b00100000; //  444 :  32 - 0x20
      11'h1BD: dout  = 8'b01111000; //  445 : 120 - 0x78
      11'h1BE: dout  = 8'b00000000; //  446 :   0 - 0x0
      11'h1BF: dout  = 8'b11000000; //  447 : 192 - 0xc0
      11'h1C0: dout  = 8'b00111111; //  448 :  63 - 0x3f -- Sprite 0x38
      11'h1C1: dout  = 8'b00001110; //  449 :  14 - 0xe
      11'h1C2: dout  = 8'b00001111; //  450 :  15 - 0xf
      11'h1C3: dout  = 8'b00011111; //  451 :  31 - 0x1f
      11'h1C4: dout  = 8'b00111111; //  452 :  63 - 0x3f
      11'h1C5: dout  = 8'b01111100; //  453 : 124 - 0x7c
      11'h1C6: dout  = 8'b01110000; //  454 : 112 - 0x70
      11'h1C7: dout  = 8'b00111000; //  455 :  56 - 0x38
      11'h1C8: dout  = 8'b11110000; //  456 : 240 - 0xf0 -- Sprite 0x39
      11'h1C9: dout  = 8'b11111000; //  457 : 248 - 0xf8
      11'h1CA: dout  = 8'b11100100; //  458 : 228 - 0xe4
      11'h1CB: dout  = 8'b11111100; //  459 : 252 - 0xfc
      11'h1CC: dout  = 8'b11111100; //  460 : 252 - 0xfc
      11'h1CD: dout  = 8'b01111100; //  461 : 124 - 0x7c
      11'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout  = 8'b00000111; //  464 :   7 - 0x7 -- Sprite 0x3a
      11'h1D1: dout  = 8'b00001111; //  465 :  15 - 0xf
      11'h1D2: dout  = 8'b00001110; //  466 :  14 - 0xe
      11'h1D3: dout  = 8'b00010100; //  467 :  20 - 0x14
      11'h1D4: dout  = 8'b00010110; //  468 :  22 - 0x16
      11'h1D5: dout  = 8'b00011000; //  469 :  24 - 0x18
      11'h1D6: dout  = 8'b00000000; //  470 :   0 - 0x0
      11'h1D7: dout  = 8'b00001111; //  471 :  15 - 0xf
      11'h1D8: dout  = 8'b00011111; //  472 :  31 - 0x1f -- Sprite 0x3b
      11'h1D9: dout  = 8'b00011111; //  473 :  31 - 0x1f
      11'h1DA: dout  = 8'b00011111; //  474 :  31 - 0x1f
      11'h1DB: dout  = 8'b00011100; //  475 :  28 - 0x1c
      11'h1DC: dout  = 8'b00001100; //  476 :  12 - 0xc
      11'h1DD: dout  = 8'b00000111; //  477 :   7 - 0x7
      11'h1DE: dout  = 8'b00000111; //  478 :   7 - 0x7
      11'h1DF: dout  = 8'b00000111; //  479 :   7 - 0x7
      11'h1E0: dout  = 8'b11100000; //  480 : 224 - 0xe0 -- Sprite 0x3c
      11'h1E1: dout  = 8'b01100000; //  481 :  96 - 0x60
      11'h1E2: dout  = 8'b11110000; //  482 : 240 - 0xf0
      11'h1E3: dout  = 8'b01110000; //  483 : 112 - 0x70
      11'h1E4: dout  = 8'b11100000; //  484 : 224 - 0xe0
      11'h1E5: dout  = 8'b11100000; //  485 : 224 - 0xe0
      11'h1E6: dout  = 8'b11110000; //  486 : 240 - 0xf0
      11'h1E7: dout  = 8'b10000000; //  487 : 128 - 0x80
      11'h1E8: dout  = 8'b00000111; //  488 :   7 - 0x7 -- Sprite 0x3d
      11'h1E9: dout  = 8'b00011111; //  489 :  31 - 0x1f
      11'h1EA: dout  = 8'b00111111; //  490 :  63 - 0x3f
      11'h1EB: dout  = 8'b00010010; //  491 :  18 - 0x12
      11'h1EC: dout  = 8'b00010011; //  492 :  19 - 0x13
      11'h1ED: dout  = 8'b00001000; //  493 :   8 - 0x8
      11'h1EE: dout  = 8'b00011111; //  494 :  31 - 0x1f
      11'h1EF: dout  = 8'b00110001; //  495 :  49 - 0x31
      11'h1F0: dout  = 8'b11000000; //  496 : 192 - 0xc0 -- Sprite 0x3e
      11'h1F1: dout  = 8'b11110000; //  497 : 240 - 0xf0
      11'h1F2: dout  = 8'b01000000; //  498 :  64 - 0x40
      11'h1F3: dout  = 8'b00000000; //  499 :   0 - 0x0
      11'h1F4: dout  = 8'b00110000; //  500 :  48 - 0x30
      11'h1F5: dout  = 8'b00011000; //  501 :  24 - 0x18
      11'h1F6: dout  = 8'b11000000; //  502 : 192 - 0xc0
      11'h1F7: dout  = 8'b11111000; //  503 : 248 - 0xf8
      11'h1F8: dout  = 8'b00110001; //  504 :  49 - 0x31 -- Sprite 0x3f
      11'h1F9: dout  = 8'b00111001; //  505 :  57 - 0x39
      11'h1FA: dout  = 8'b00011111; //  506 :  31 - 0x1f
      11'h1FB: dout  = 8'b00011111; //  507 :  31 - 0x1f
      11'h1FC: dout  = 8'b00001111; //  508 :  15 - 0xf
      11'h1FD: dout  = 8'b01011111; //  509 :  95 - 0x5f
      11'h1FE: dout  = 8'b01111110; //  510 : 126 - 0x7e
      11'h1FF: dout  = 8'b00111100; //  511 :  60 - 0x3c
      11'h200: dout  = 8'b11111000; //  512 : 248 - 0xf8 -- Sprite 0x40
      11'h201: dout  = 8'b11111000; //  513 : 248 - 0xf8
      11'h202: dout  = 8'b11110000; //  514 : 240 - 0xf0
      11'h203: dout  = 8'b11100000; //  515 : 224 - 0xe0
      11'h204: dout  = 8'b11100000; //  516 : 224 - 0xe0
      11'h205: dout  = 8'b11000000; //  517 : 192 - 0xc0
      11'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      11'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      11'h208: dout  = 8'b00000000; //  520 :   0 - 0x0 -- Sprite 0x41
      11'h209: dout  = 8'b11100000; //  521 : 224 - 0xe0
      11'h20A: dout  = 8'b11111100; //  522 : 252 - 0xfc
      11'h20B: dout  = 8'b00100111; //  523 :  39 - 0x27
      11'h20C: dout  = 8'b00100111; //  524 :  39 - 0x27
      11'h20D: dout  = 8'b00010001; //  525 :  17 - 0x11
      11'h20E: dout  = 8'b00111110; //  526 :  62 - 0x3e
      11'h20F: dout  = 8'b00000100; //  527 :   4 - 0x4
      11'h210: dout  = 8'b00111111; //  528 :  63 - 0x3f -- Sprite 0x42
      11'h211: dout  = 8'b01111111; //  529 : 127 - 0x7f
      11'h212: dout  = 8'b00111111; //  530 :  63 - 0x3f
      11'h213: dout  = 8'b00001111; //  531 :  15 - 0xf
      11'h214: dout  = 8'b00011111; //  532 :  31 - 0x1f
      11'h215: dout  = 8'b00111111; //  533 :  63 - 0x3f
      11'h216: dout  = 8'b01111111; //  534 : 127 - 0x7f
      11'h217: dout  = 8'b01001111; //  535 :  79 - 0x4f
      11'h218: dout  = 8'b11111000; //  536 : 248 - 0xf8 -- Sprite 0x43
      11'h219: dout  = 8'b11111001; //  537 : 249 - 0xf9
      11'h21A: dout  = 8'b11111001; //  538 : 249 - 0xf9
      11'h21B: dout  = 8'b10110111; //  539 : 183 - 0xb7
      11'h21C: dout  = 8'b11111111; //  540 : 255 - 0xff
      11'h21D: dout  = 8'b11111111; //  541 : 255 - 0xff
      11'h21E: dout  = 8'b11100000; //  542 : 224 - 0xe0
      11'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      11'h220: dout  = 8'b00000111; //  544 :   7 - 0x7 -- Sprite 0x44
      11'h221: dout  = 8'b00000111; //  545 :   7 - 0x7
      11'h222: dout  = 8'b00001111; //  546 :  15 - 0xf
      11'h223: dout  = 8'b00111111; //  547 :  63 - 0x3f
      11'h224: dout  = 8'b00111111; //  548 :  63 - 0x3f
      11'h225: dout  = 8'b00111111; //  549 :  63 - 0x3f
      11'h226: dout  = 8'b00100110; //  550 :  38 - 0x26
      11'h227: dout  = 8'b00000100; //  551 :   4 - 0x4
      11'h228: dout  = 8'b11110000; //  552 : 240 - 0xf0 -- Sprite 0x45
      11'h229: dout  = 8'b11110000; //  553 : 240 - 0xf0
      11'h22A: dout  = 8'b11110000; //  554 : 240 - 0xf0
      11'h22B: dout  = 8'b11100000; //  555 : 224 - 0xe0
      11'h22C: dout  = 8'b11000000; //  556 : 192 - 0xc0
      11'h22D: dout  = 8'b00000000; //  557 :   0 - 0x0
      11'h22E: dout  = 8'b00000000; //  558 :   0 - 0x0
      11'h22F: dout  = 8'b00000000; //  559 :   0 - 0x0
      11'h230: dout  = 8'b00000111; //  560 :   7 - 0x7 -- Sprite 0x46
      11'h231: dout  = 8'b00000111; //  561 :   7 - 0x7
      11'h232: dout  = 8'b00001111; //  562 :  15 - 0xf
      11'h233: dout  = 8'b00011111; //  563 :  31 - 0x1f
      11'h234: dout  = 8'b00111111; //  564 :  63 - 0x3f
      11'h235: dout  = 8'b00001111; //  565 :  15 - 0xf
      11'h236: dout  = 8'b00011100; //  566 :  28 - 0x1c
      11'h237: dout  = 8'b00011000; //  567 :  24 - 0x18
      11'h238: dout  = 8'b11100000; //  568 : 224 - 0xe0 -- Sprite 0x47
      11'h239: dout  = 8'b11100000; //  569 : 224 - 0xe0
      11'h23A: dout  = 8'b11100000; //  570 : 224 - 0xe0
      11'h23B: dout  = 8'b11100000; //  571 : 224 - 0xe0
      11'h23C: dout  = 8'b11000000; //  572 : 192 - 0xc0
      11'h23D: dout  = 8'b10000000; //  573 : 128 - 0x80
      11'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      11'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout  = 8'b00000111; //  576 :   7 - 0x7 -- Sprite 0x48
      11'h241: dout  = 8'b00001111; //  577 :  15 - 0xf
      11'h242: dout  = 8'b00011111; //  578 :  31 - 0x1f
      11'h243: dout  = 8'b00001111; //  579 :  15 - 0xf
      11'h244: dout  = 8'b00111111; //  580 :  63 - 0x3f
      11'h245: dout  = 8'b00001111; //  581 :  15 - 0xf
      11'h246: dout  = 8'b00011100; //  582 :  28 - 0x1c
      11'h247: dout  = 8'b00011000; //  583 :  24 - 0x18
      11'h248: dout  = 8'b11100000; //  584 : 224 - 0xe0 -- Sprite 0x49
      11'h249: dout  = 8'b11100000; //  585 : 224 - 0xe0
      11'h24A: dout  = 8'b11100000; //  586 : 224 - 0xe0
      11'h24B: dout  = 8'b01000000; //  587 :  64 - 0x40
      11'h24C: dout  = 8'b11000000; //  588 : 192 - 0xc0
      11'h24D: dout  = 8'b10000000; //  589 : 128 - 0x80
      11'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      11'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      11'h250: dout  = 8'b01111111; //  592 : 127 - 0x7f -- Sprite 0x4a
      11'h251: dout  = 8'b11111111; //  593 : 255 - 0xff
      11'h252: dout  = 8'b11111111; //  594 : 255 - 0xff
      11'h253: dout  = 8'b11111011; //  595 : 251 - 0xfb
      11'h254: dout  = 8'b00001111; //  596 :  15 - 0xf
      11'h255: dout  = 8'b00001111; //  597 :  15 - 0xf
      11'h256: dout  = 8'b00001111; //  598 :  15 - 0xf
      11'h257: dout  = 8'b00011111; //  599 :  31 - 0x1f
      11'h258: dout  = 8'b00111111; //  600 :  63 - 0x3f -- Sprite 0x4b
      11'h259: dout  = 8'b01111110; //  601 : 126 - 0x7e
      11'h25A: dout  = 8'b01111100; //  602 : 124 - 0x7c
      11'h25B: dout  = 8'b01111100; //  603 : 124 - 0x7c
      11'h25C: dout  = 8'b00111100; //  604 :  60 - 0x3c
      11'h25D: dout  = 8'b00111100; //  605 :  60 - 0x3c
      11'h25E: dout  = 8'b11111100; //  606 : 252 - 0xfc
      11'h25F: dout  = 8'b11111100; //  607 : 252 - 0xfc
      11'h260: dout  = 8'b01100000; //  608 :  96 - 0x60 -- Sprite 0x4c
      11'h261: dout  = 8'b01110000; //  609 : 112 - 0x70
      11'h262: dout  = 8'b00011000; //  610 :  24 - 0x18
      11'h263: dout  = 8'b00001000; //  611 :   8 - 0x8
      11'h264: dout  = 8'b00001111; //  612 :  15 - 0xf
      11'h265: dout  = 8'b00011111; //  613 :  31 - 0x1f
      11'h266: dout  = 8'b00111111; //  614 :  63 - 0x3f
      11'h267: dout  = 8'b01111111; //  615 : 127 - 0x7f
      11'h268: dout  = 8'b11111100; //  616 : 252 - 0xfc -- Sprite 0x4d
      11'h269: dout  = 8'b01111100; //  617 : 124 - 0x7c
      11'h26A: dout  = 8'b00000000; //  618 :   0 - 0x0
      11'h26B: dout  = 8'b00100000; //  619 :  32 - 0x20
      11'h26C: dout  = 8'b11110000; //  620 : 240 - 0xf0
      11'h26D: dout  = 8'b11111000; //  621 : 248 - 0xf8
      11'h26E: dout  = 8'b11111100; //  622 : 252 - 0xfc
      11'h26F: dout  = 8'b11111110; //  623 : 254 - 0xfe
      11'h270: dout  = 8'b00001011; //  624 :  11 - 0xb -- Sprite 0x4e
      11'h271: dout  = 8'b00001111; //  625 :  15 - 0xf
      11'h272: dout  = 8'b00011111; //  626 :  31 - 0x1f
      11'h273: dout  = 8'b00011110; //  627 :  30 - 0x1e
      11'h274: dout  = 8'b00111100; //  628 :  60 - 0x3c
      11'h275: dout  = 8'b00111100; //  629 :  60 - 0x3c
      11'h276: dout  = 8'b00111100; //  630 :  60 - 0x3c
      11'h277: dout  = 8'b01111100; //  631 : 124 - 0x7c
      11'h278: dout  = 8'b00011111; //  632 :  31 - 0x1f -- Sprite 0x4f
      11'h279: dout  = 8'b00111111; //  633 :  63 - 0x3f
      11'h27A: dout  = 8'b00001101; //  634 :  13 - 0xd
      11'h27B: dout  = 8'b00000111; //  635 :   7 - 0x7
      11'h27C: dout  = 8'b00001111; //  636 :  15 - 0xf
      11'h27D: dout  = 8'b00001110; //  637 :  14 - 0xe
      11'h27E: dout  = 8'b00011100; //  638 :  28 - 0x1c
      11'h27F: dout  = 8'b00111100; //  639 :  60 - 0x3c
      11'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x50
      11'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      11'h282: dout  = 8'b00000000; //  642 :   0 - 0x0
      11'h283: dout  = 8'b00000000; //  643 :   0 - 0x0
      11'h284: dout  = 8'b00000000; //  644 :   0 - 0x0
      11'h285: dout  = 8'b00000000; //  645 :   0 - 0x0
      11'h286: dout  = 8'b00000000; //  646 :   0 - 0x0
      11'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      11'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- Sprite 0x51
      11'h289: dout  = 8'b00000111; //  649 :   7 - 0x7
      11'h28A: dout  = 8'b00011111; //  650 :  31 - 0x1f
      11'h28B: dout  = 8'b11111111; //  651 : 255 - 0xff
      11'h28C: dout  = 8'b00000111; //  652 :   7 - 0x7
      11'h28D: dout  = 8'b00011111; //  653 :  31 - 0x1f
      11'h28E: dout  = 8'b00001111; //  654 :  15 - 0xf
      11'h28F: dout  = 8'b00000110; //  655 :   6 - 0x6
      11'h290: dout  = 8'b00111111; //  656 :  63 - 0x3f -- Sprite 0x52
      11'h291: dout  = 8'b11111111; //  657 : 255 - 0xff
      11'h292: dout  = 8'b11111111; //  658 : 255 - 0xff
      11'h293: dout  = 8'b11111111; //  659 : 255 - 0xff
      11'h294: dout  = 8'b11111111; //  660 : 255 - 0xff
      11'h295: dout  = 8'b11111111; //  661 : 255 - 0xff
      11'h296: dout  = 8'b11111011; //  662 : 251 - 0xfb
      11'h297: dout  = 8'b01110110; //  663 : 118 - 0x76
      11'h298: dout  = 8'b00100000; //  664 :  32 - 0x20 -- Sprite 0x53
      11'h299: dout  = 8'b11111000; //  665 : 248 - 0xf8
      11'h29A: dout  = 8'b11111111; //  666 : 255 - 0xff
      11'h29B: dout  = 8'b11000011; //  667 : 195 - 0xc3
      11'h29C: dout  = 8'b11111101; //  668 : 253 - 0xfd
      11'h29D: dout  = 8'b11111110; //  669 : 254 - 0xfe
      11'h29E: dout  = 8'b11110000; //  670 : 240 - 0xf0
      11'h29F: dout  = 8'b01000000; //  671 :  64 - 0x40
      11'h2A0: dout  = 8'b01000000; //  672 :  64 - 0x40 -- Sprite 0x54
      11'h2A1: dout  = 8'b11100000; //  673 : 224 - 0xe0
      11'h2A2: dout  = 8'b01000000; //  674 :  64 - 0x40
      11'h2A3: dout  = 8'b01000000; //  675 :  64 - 0x40
      11'h2A4: dout  = 8'b01000001; //  676 :  65 - 0x41
      11'h2A5: dout  = 8'b01000001; //  677 :  65 - 0x41
      11'h2A6: dout  = 8'b01001111; //  678 :  79 - 0x4f
      11'h2A7: dout  = 8'b01000111; //  679 :  71 - 0x47
      11'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      11'h2A9: dout  = 8'b00000000; //  681 :   0 - 0x0
      11'h2AA: dout  = 8'b00000000; //  682 :   0 - 0x0
      11'h2AB: dout  = 8'b00000000; //  683 :   0 - 0x0
      11'h2AC: dout  = 8'b00000000; //  684 :   0 - 0x0
      11'h2AD: dout  = 8'b00000000; //  685 :   0 - 0x0
      11'h2AE: dout  = 8'b11100000; //  686 : 224 - 0xe0
      11'h2AF: dout  = 8'b11000000; //  687 : 192 - 0xc0
      11'h2B0: dout  = 8'b01000011; //  688 :  67 - 0x43 -- Sprite 0x56
      11'h2B1: dout  = 8'b01000110; //  689 :  70 - 0x46
      11'h2B2: dout  = 8'b01000100; //  690 :  68 - 0x44
      11'h2B3: dout  = 8'b01000000; //  691 :  64 - 0x40
      11'h2B4: dout  = 8'b01000000; //  692 :  64 - 0x40
      11'h2B5: dout  = 8'b01000000; //  693 :  64 - 0x40
      11'h2B6: dout  = 8'b01000000; //  694 :  64 - 0x40
      11'h2B7: dout  = 8'b01000000; //  695 :  64 - 0x40
      11'h2B8: dout  = 8'b10000000; //  696 : 128 - 0x80 -- Sprite 0x57
      11'h2B9: dout  = 8'b11000000; //  697 : 192 - 0xc0
      11'h2BA: dout  = 8'b01000000; //  698 :  64 - 0x40
      11'h2BB: dout  = 8'b00000000; //  699 :   0 - 0x0
      11'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      11'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      11'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      11'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      11'h2C0: dout  = 8'b00110001; //  704 :  49 - 0x31 -- Sprite 0x58
      11'h2C1: dout  = 8'b00110000; //  705 :  48 - 0x30
      11'h2C2: dout  = 8'b00111000; //  706 :  56 - 0x38
      11'h2C3: dout  = 8'b01111100; //  707 : 124 - 0x7c
      11'h2C4: dout  = 8'b01111111; //  708 : 127 - 0x7f
      11'h2C5: dout  = 8'b11111111; //  709 : 255 - 0xff
      11'h2C6: dout  = 8'b11111111; //  710 : 255 - 0xff
      11'h2C7: dout  = 8'b11111011; //  711 : 251 - 0xfb
      11'h2C8: dout  = 8'b00010000; //  712 :  16 - 0x10 -- Sprite 0x59
      11'h2C9: dout  = 8'b01111110; //  713 : 126 - 0x7e
      11'h2CA: dout  = 8'b00111110; //  714 :  62 - 0x3e
      11'h2CB: dout  = 8'b00000000; //  715 :   0 - 0x0
      11'h2CC: dout  = 8'b00011110; //  716 :  30 - 0x1e
      11'h2CD: dout  = 8'b11111110; //  717 : 254 - 0xfe
      11'h2CE: dout  = 8'b11111111; //  718 : 255 - 0xff
      11'h2CF: dout  = 8'b11111111; //  719 : 255 - 0xff
      11'h2D0: dout  = 8'b11111111; //  720 : 255 - 0xff -- Sprite 0x5a
      11'h2D1: dout  = 8'b11111111; //  721 : 255 - 0xff
      11'h2D2: dout  = 8'b11100011; //  722 : 227 - 0xe3
      11'h2D3: dout  = 8'b11000011; //  723 : 195 - 0xc3
      11'h2D4: dout  = 8'b10000111; //  724 : 135 - 0x87
      11'h2D5: dout  = 8'b01001000; //  725 :  72 - 0x48
      11'h2D6: dout  = 8'b00111100; //  726 :  60 - 0x3c
      11'h2D7: dout  = 8'b11111100; //  727 : 252 - 0xfc
      11'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- Sprite 0x5b
      11'h2D9: dout  = 8'b11111111; //  729 : 255 - 0xff
      11'h2DA: dout  = 8'b11000011; //  730 : 195 - 0xc3
      11'h2DB: dout  = 8'b10000011; //  731 : 131 - 0x83
      11'h2DC: dout  = 8'b10000011; //  732 : 131 - 0x83
      11'h2DD: dout  = 8'b11111111; //  733 : 255 - 0xff
      11'h2DE: dout  = 8'b11111111; //  734 : 255 - 0xff
      11'h2DF: dout  = 8'b11111111; //  735 : 255 - 0xff
      11'h2E0: dout  = 8'b00011111; //  736 :  31 - 0x1f -- Sprite 0x5c
      11'h2E1: dout  = 8'b00011111; //  737 :  31 - 0x1f
      11'h2E2: dout  = 8'b00001111; //  738 :  15 - 0xf
      11'h2E3: dout  = 8'b00000111; //  739 :   7 - 0x7
      11'h2E4: dout  = 8'b00000001; //  740 :   1 - 0x1
      11'h2E5: dout  = 8'b00000000; //  741 :   0 - 0x0
      11'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      11'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      11'h2E8: dout  = 8'b11110000; //  744 : 240 - 0xf0 -- Sprite 0x5d
      11'h2E9: dout  = 8'b11111011; //  745 : 251 - 0xfb
      11'h2EA: dout  = 8'b11111111; //  746 : 255 - 0xff
      11'h2EB: dout  = 8'b11111111; //  747 : 255 - 0xff
      11'h2EC: dout  = 8'b11111110; //  748 : 254 - 0xfe
      11'h2ED: dout  = 8'b00111110; //  749 :  62 - 0x3e
      11'h2EE: dout  = 8'b00001100; //  750 :  12 - 0xc
      11'h2EF: dout  = 8'b00000100; //  751 :   4 - 0x4
      11'h2F0: dout  = 8'b00011111; //  752 :  31 - 0x1f -- Sprite 0x5e
      11'h2F1: dout  = 8'b00011111; //  753 :  31 - 0x1f
      11'h2F2: dout  = 8'b00001111; //  754 :  15 - 0xf
      11'h2F3: dout  = 8'b00001111; //  755 :  15 - 0xf
      11'h2F4: dout  = 8'b00000111; //  756 :   7 - 0x7
      11'h2F5: dout  = 8'b00000000; //  757 :   0 - 0x0
      11'h2F6: dout  = 8'b00000000; //  758 :   0 - 0x0
      11'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      11'h2F8: dout  = 8'b11111011; //  760 : 251 - 0xfb -- Sprite 0x5f
      11'h2F9: dout  = 8'b11111111; //  761 : 255 - 0xff
      11'h2FA: dout  = 8'b11111111; //  762 : 255 - 0xff
      11'h2FB: dout  = 8'b11111111; //  763 : 255 - 0xff
      11'h2FC: dout  = 8'b11111111; //  764 : 255 - 0xff
      11'h2FD: dout  = 8'b00000000; //  765 :   0 - 0x0
      11'h2FE: dout  = 8'b00000000; //  766 :   0 - 0x0
      11'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      11'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      11'h301: dout  = 8'b00011000; //  769 :  24 - 0x18
      11'h302: dout  = 8'b00111100; //  770 :  60 - 0x3c
      11'h303: dout  = 8'b01111110; //  771 : 126 - 0x7e
      11'h304: dout  = 8'b01101110; //  772 : 110 - 0x6e
      11'h305: dout  = 8'b11011111; //  773 : 223 - 0xdf
      11'h306: dout  = 8'b11011111; //  774 : 223 - 0xdf
      11'h307: dout  = 8'b11011111; //  775 : 223 - 0xdf
      11'h308: dout  = 8'b00000000; //  776 :   0 - 0x0 -- Sprite 0x61
      11'h309: dout  = 8'b00011000; //  777 :  24 - 0x18
      11'h30A: dout  = 8'b00011000; //  778 :  24 - 0x18
      11'h30B: dout  = 8'b00111100; //  779 :  60 - 0x3c
      11'h30C: dout  = 8'b00111100; //  780 :  60 - 0x3c
      11'h30D: dout  = 8'b00111100; //  781 :  60 - 0x3c
      11'h30E: dout  = 8'b00111100; //  782 :  60 - 0x3c
      11'h30F: dout  = 8'b00011100; //  783 :  28 - 0x1c
      11'h310: dout  = 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x62
      11'h311: dout  = 8'b00001000; //  785 :   8 - 0x8
      11'h312: dout  = 8'b00001000; //  786 :   8 - 0x8
      11'h313: dout  = 8'b00001000; //  787 :   8 - 0x8
      11'h314: dout  = 8'b00001000; //  788 :   8 - 0x8
      11'h315: dout  = 8'b00001000; //  789 :   8 - 0x8
      11'h316: dout  = 8'b00001000; //  790 :   8 - 0x8
      11'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      11'h318: dout  = 8'b00000000; //  792 :   0 - 0x0 -- Sprite 0x63
      11'h319: dout  = 8'b00001000; //  793 :   8 - 0x8
      11'h31A: dout  = 8'b00001000; //  794 :   8 - 0x8
      11'h31B: dout  = 8'b00000100; //  795 :   4 - 0x4
      11'h31C: dout  = 8'b00000100; //  796 :   4 - 0x4
      11'h31D: dout  = 8'b00000100; //  797 :   4 - 0x4
      11'h31E: dout  = 8'b00000100; //  798 :   4 - 0x4
      11'h31F: dout  = 8'b00000100; //  799 :   4 - 0x4
      11'h320: dout  = 8'b00111100; //  800 :  60 - 0x3c -- Sprite 0x64
      11'h321: dout  = 8'b01111110; //  801 : 126 - 0x7e
      11'h322: dout  = 8'b01110111; //  802 : 119 - 0x77
      11'h323: dout  = 8'b11111011; //  803 : 251 - 0xfb
      11'h324: dout  = 8'b10011111; //  804 : 159 - 0x9f
      11'h325: dout  = 8'b01011111; //  805 :  95 - 0x5f
      11'h326: dout  = 8'b10001110; //  806 : 142 - 0x8e
      11'h327: dout  = 8'b00100000; //  807 :  32 - 0x20
      11'h328: dout  = 8'b01011100; //  808 :  92 - 0x5c -- Sprite 0x65
      11'h329: dout  = 8'b00101110; //  809 :  46 - 0x2e
      11'h32A: dout  = 8'b10001111; //  810 : 143 - 0x8f
      11'h32B: dout  = 8'b00111111; //  811 :  63 - 0x3f
      11'h32C: dout  = 8'b01111011; //  812 : 123 - 0x7b
      11'h32D: dout  = 8'b01110111; //  813 : 119 - 0x77
      11'h32E: dout  = 8'b01111110; //  814 : 126 - 0x7e
      11'h32F: dout  = 8'b00111100; //  815 :  60 - 0x3c
      11'h330: dout  = 8'b00010011; //  816 :  19 - 0x13 -- Sprite 0x66
      11'h331: dout  = 8'b01001111; //  817 :  79 - 0x4f
      11'h332: dout  = 8'b00111111; //  818 :  63 - 0x3f
      11'h333: dout  = 8'b10111111; //  819 : 191 - 0xbf
      11'h334: dout  = 8'b00111111; //  820 :  63 - 0x3f
      11'h335: dout  = 8'b01111010; //  821 : 122 - 0x7a
      11'h336: dout  = 8'b11111000; //  822 : 248 - 0xf8
      11'h337: dout  = 8'b11111000; //  823 : 248 - 0xf8
      11'h338: dout  = 8'b00000000; //  824 :   0 - 0x0 -- Sprite 0x67
      11'h339: dout  = 8'b00001000; //  825 :   8 - 0x8
      11'h33A: dout  = 8'b00000101; //  826 :   5 - 0x5
      11'h33B: dout  = 8'b00001111; //  827 :  15 - 0xf
      11'h33C: dout  = 8'b00101111; //  828 :  47 - 0x2f
      11'h33D: dout  = 8'b00011101; //  829 :  29 - 0x1d
      11'h33E: dout  = 8'b00011100; //  830 :  28 - 0x1c
      11'h33F: dout  = 8'b00111100; //  831 :  60 - 0x3c
      11'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      11'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      11'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      11'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      11'h344: dout  = 8'b00000010; //  836 :   2 - 0x2
      11'h345: dout  = 8'b00001011; //  837 :  11 - 0xb
      11'h346: dout  = 8'b00000111; //  838 :   7 - 0x7
      11'h347: dout  = 8'b00001111; //  839 :  15 - 0xf
      11'h348: dout  = 8'b00000000; //  840 :   0 - 0x0 -- Sprite 0x69
      11'h349: dout  = 8'b00000000; //  841 :   0 - 0x0
      11'h34A: dout  = 8'b00000000; //  842 :   0 - 0x0
      11'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      11'h34C: dout  = 8'b00000000; //  844 :   0 - 0x0
      11'h34D: dout  = 8'b00001000; //  845 :   8 - 0x8
      11'h34E: dout  = 8'b00000100; //  846 :   4 - 0x4
      11'h34F: dout  = 8'b00000100; //  847 :   4 - 0x4
      11'h350: dout  = 8'b00000010; //  848 :   2 - 0x2 -- Sprite 0x6a
      11'h351: dout  = 8'b00000010; //  849 :   2 - 0x2
      11'h352: dout  = 8'b00000010; //  850 :   2 - 0x2
      11'h353: dout  = 8'b00000101; //  851 :   5 - 0x5
      11'h354: dout  = 8'b01110001; //  852 : 113 - 0x71
      11'h355: dout  = 8'b01111111; //  853 : 127 - 0x7f
      11'h356: dout  = 8'b01111111; //  854 : 127 - 0x7f
      11'h357: dout  = 8'b01111111; //  855 : 127 - 0x7f
      11'h358: dout  = 8'b00000000; //  856 :   0 - 0x0 -- Sprite 0x6b
      11'h359: dout  = 8'b00000000; //  857 :   0 - 0x0
      11'h35A: dout  = 8'b00000000; //  858 :   0 - 0x0
      11'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      11'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      11'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      11'h35E: dout  = 8'b00000000; //  862 :   0 - 0x0
      11'h35F: dout  = 8'b00000100; //  863 :   4 - 0x4
      11'h360: dout  = 8'b00000010; //  864 :   2 - 0x2 -- Sprite 0x6c
      11'h361: dout  = 8'b00000010; //  865 :   2 - 0x2
      11'h362: dout  = 8'b00000000; //  866 :   0 - 0x0
      11'h363: dout  = 8'b00000001; //  867 :   1 - 0x1
      11'h364: dout  = 8'b00010011; //  868 :  19 - 0x13
      11'h365: dout  = 8'b00111111; //  869 :  63 - 0x3f
      11'h366: dout  = 8'b01111111; //  870 : 127 - 0x7f
      11'h367: dout  = 8'b01111111; //  871 : 127 - 0x7f
      11'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      11'h369: dout  = 8'b01000000; //  873 :  64 - 0x40
      11'h36A: dout  = 8'b01100000; //  874 :  96 - 0x60
      11'h36B: dout  = 8'b01110000; //  875 : 112 - 0x70
      11'h36C: dout  = 8'b01110011; //  876 : 115 - 0x73
      11'h36D: dout  = 8'b00100111; //  877 :  39 - 0x27
      11'h36E: dout  = 8'b00001111; //  878 :  15 - 0xf
      11'h36F: dout  = 8'b00011111; //  879 :  31 - 0x1f
      11'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      11'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout  = 8'b00000000; //  882 :   0 - 0x0
      11'h373: dout  = 8'b00000000; //  883 :   0 - 0x0
      11'h374: dout  = 8'b00000011; //  884 :   3 - 0x3
      11'h375: dout  = 8'b00000111; //  885 :   7 - 0x7
      11'h376: dout  = 8'b00001111; //  886 :  15 - 0xf
      11'h377: dout  = 8'b00011111; //  887 :  31 - 0x1f
      11'h378: dout  = 8'b01111111; //  888 : 127 - 0x7f -- Sprite 0x6f
      11'h379: dout  = 8'b01111111; //  889 : 127 - 0x7f
      11'h37A: dout  = 8'b00111111; //  890 :  63 - 0x3f
      11'h37B: dout  = 8'b00111111; //  891 :  63 - 0x3f
      11'h37C: dout  = 8'b00011111; //  892 :  31 - 0x1f
      11'h37D: dout  = 8'b00011111; //  893 :  31 - 0x1f
      11'h37E: dout  = 8'b00001111; //  894 :  15 - 0xf
      11'h37F: dout  = 8'b00000111; //  895 :   7 - 0x7
      11'h380: dout  = 8'b00000011; //  896 :   3 - 0x3 -- Sprite 0x70
      11'h381: dout  = 8'b00000111; //  897 :   7 - 0x7
      11'h382: dout  = 8'b00001111; //  898 :  15 - 0xf
      11'h383: dout  = 8'b00011111; //  899 :  31 - 0x1f
      11'h384: dout  = 8'b00111111; //  900 :  63 - 0x3f
      11'h385: dout  = 8'b01110111; //  901 : 119 - 0x77
      11'h386: dout  = 8'b01110111; //  902 : 119 - 0x77
      11'h387: dout  = 8'b11110101; //  903 : 245 - 0xf5
      11'h388: dout  = 8'b11000000; //  904 : 192 - 0xc0 -- Sprite 0x71
      11'h389: dout  = 8'b11100000; //  905 : 224 - 0xe0
      11'h38A: dout  = 8'b11110000; //  906 : 240 - 0xf0
      11'h38B: dout  = 8'b11111000; //  907 : 248 - 0xf8
      11'h38C: dout  = 8'b11111100; //  908 : 252 - 0xfc
      11'h38D: dout  = 8'b11101110; //  909 : 238 - 0xee
      11'h38E: dout  = 8'b11101110; //  910 : 238 - 0xee
      11'h38F: dout  = 8'b10101111; //  911 : 175 - 0xaf
      11'h390: dout  = 8'b11110001; //  912 : 241 - 0xf1 -- Sprite 0x72
      11'h391: dout  = 8'b11111111; //  913 : 255 - 0xff
      11'h392: dout  = 8'b01111000; //  914 : 120 - 0x78
      11'h393: dout  = 8'b00000000; //  915 :   0 - 0x0
      11'h394: dout  = 8'b00000000; //  916 :   0 - 0x0
      11'h395: dout  = 8'b00011000; //  917 :  24 - 0x18
      11'h396: dout  = 8'b00011100; //  918 :  28 - 0x1c
      11'h397: dout  = 8'b00001110; //  919 :  14 - 0xe
      11'h398: dout  = 8'b10001111; //  920 : 143 - 0x8f -- Sprite 0x73
      11'h399: dout  = 8'b11111111; //  921 : 255 - 0xff
      11'h39A: dout  = 8'b00011110; //  922 :  30 - 0x1e
      11'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      11'h39C: dout  = 8'b00001100; //  924 :  12 - 0xc
      11'h39D: dout  = 8'b00111110; //  925 :  62 - 0x3e
      11'h39E: dout  = 8'b01111110; //  926 : 126 - 0x7e
      11'h39F: dout  = 8'b01111100; //  927 : 124 - 0x7c
      11'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x74
      11'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      11'h3A2: dout  = 8'b00000000; //  930 :   0 - 0x0
      11'h3A3: dout  = 8'b00000000; //  931 :   0 - 0x0
      11'h3A4: dout  = 8'b00000000; //  932 :   0 - 0x0
      11'h3A5: dout  = 8'b00000000; //  933 :   0 - 0x0
      11'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      11'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      11'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0 -- Sprite 0x75
      11'h3A9: dout  = 8'b00000010; //  937 :   2 - 0x2
      11'h3AA: dout  = 8'b01000001; //  938 :  65 - 0x41
      11'h3AB: dout  = 8'b01000001; //  939 :  65 - 0x41
      11'h3AC: dout  = 8'b01100001; //  940 :  97 - 0x61
      11'h3AD: dout  = 8'b00110011; //  941 :  51 - 0x33
      11'h3AE: dout  = 8'b00000110; //  942 :   6 - 0x6
      11'h3AF: dout  = 8'b00111100; //  943 :  60 - 0x3c
      11'h3B0: dout  = 8'b00000011; //  944 :   3 - 0x3 -- Sprite 0x76
      11'h3B1: dout  = 8'b00000111; //  945 :   7 - 0x7
      11'h3B2: dout  = 8'b00001111; //  946 :  15 - 0xf
      11'h3B3: dout  = 8'b00011111; //  947 :  31 - 0x1f
      11'h3B4: dout  = 8'b00111111; //  948 :  63 - 0x3f
      11'h3B5: dout  = 8'b01111111; //  949 : 127 - 0x7f
      11'h3B6: dout  = 8'b01111111; //  950 : 127 - 0x7f
      11'h3B7: dout  = 8'b11111111; //  951 : 255 - 0xff
      11'h3B8: dout  = 8'b11000000; //  952 : 192 - 0xc0 -- Sprite 0x77
      11'h3B9: dout  = 8'b11100000; //  953 : 224 - 0xe0
      11'h3BA: dout  = 8'b11110000; //  954 : 240 - 0xf0
      11'h3BB: dout  = 8'b11111000; //  955 : 248 - 0xf8
      11'h3BC: dout  = 8'b11111100; //  956 : 252 - 0xfc
      11'h3BD: dout  = 8'b11111110; //  957 : 254 - 0xfe
      11'h3BE: dout  = 8'b11111110; //  958 : 254 - 0xfe
      11'h3BF: dout  = 8'b11111111; //  959 : 255 - 0xff
      11'h3C0: dout  = 8'b11111111; //  960 : 255 - 0xff -- Sprite 0x78
      11'h3C1: dout  = 8'b11111111; //  961 : 255 - 0xff
      11'h3C2: dout  = 8'b11111111; //  962 : 255 - 0xff
      11'h3C3: dout  = 8'b01111000; //  963 : 120 - 0x78
      11'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      11'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      11'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      11'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      11'h3C8: dout  = 8'b11111111; //  968 : 255 - 0xff -- Sprite 0x79
      11'h3C9: dout  = 8'b11111111; //  969 : 255 - 0xff
      11'h3CA: dout  = 8'b11111111; //  970 : 255 - 0xff
      11'h3CB: dout  = 8'b00011110; //  971 :  30 - 0x1e
      11'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      11'h3CD: dout  = 8'b00100000; //  973 :  32 - 0x20
      11'h3CE: dout  = 8'b00100000; //  974 :  32 - 0x20
      11'h3CF: dout  = 8'b01000000; //  975 :  64 - 0x40
      11'h3D0: dout  = 8'b00010110; //  976 :  22 - 0x16 -- Sprite 0x7a
      11'h3D1: dout  = 8'b00011111; //  977 :  31 - 0x1f
      11'h3D2: dout  = 8'b00111111; //  978 :  63 - 0x3f
      11'h3D3: dout  = 8'b01111111; //  979 : 127 - 0x7f
      11'h3D4: dout  = 8'b00111101; //  980 :  61 - 0x3d
      11'h3D5: dout  = 8'b00011101; //  981 :  29 - 0x1d
      11'h3D6: dout  = 8'b00111111; //  982 :  63 - 0x3f
      11'h3D7: dout  = 8'b00011111; //  983 :  31 - 0x1f
      11'h3D8: dout  = 8'b10000000; //  984 : 128 - 0x80 -- Sprite 0x7b
      11'h3D9: dout  = 8'b10000000; //  985 : 128 - 0x80
      11'h3DA: dout  = 8'b11000000; //  986 : 192 - 0xc0
      11'h3DB: dout  = 8'b11100000; //  987 : 224 - 0xe0
      11'h3DC: dout  = 8'b11110000; //  988 : 240 - 0xf0
      11'h3DD: dout  = 8'b11110000; //  989 : 240 - 0xf0
      11'h3DE: dout  = 8'b11110000; //  990 : 240 - 0xf0
      11'h3DF: dout  = 8'b11111000; //  991 : 248 - 0xf8
      11'h3E0: dout  = 8'b00111100; //  992 :  60 - 0x3c -- Sprite 0x7c
      11'h3E1: dout  = 8'b11111010; //  993 : 250 - 0xfa
      11'h3E2: dout  = 8'b10110001; //  994 : 177 - 0xb1
      11'h3E3: dout  = 8'b01110010; //  995 : 114 - 0x72
      11'h3E4: dout  = 8'b11110010; //  996 : 242 - 0xf2
      11'h3E5: dout  = 8'b11011011; //  997 : 219 - 0xdb
      11'h3E6: dout  = 8'b11011111; //  998 : 223 - 0xdf
      11'h3E7: dout  = 8'b01011111; //  999 :  95 - 0x5f
      11'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- Sprite 0x7d
      11'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      11'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      11'h3EB: dout  = 8'b00000001; // 1003 :   1 - 0x1
      11'h3EC: dout  = 8'b00000001; // 1004 :   1 - 0x1
      11'h3ED: dout  = 8'b00000001; // 1005 :   1 - 0x1
      11'h3EE: dout  = 8'b00000110; // 1006 :   6 - 0x6
      11'h3EF: dout  = 8'b00011110; // 1007 :  30 - 0x1e
      11'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x7e
      11'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      11'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      11'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      11'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      11'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      11'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      11'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      11'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0 -- Sprite 0x7f
      11'h3F9: dout  = 8'b01111100; // 1017 : 124 - 0x7c
      11'h3FA: dout  = 8'b11010110; // 1018 : 214 - 0xd6
      11'h3FB: dout  = 8'b10010010; // 1019 : 146 - 0x92
      11'h3FC: dout  = 8'b10111010; // 1020 : 186 - 0xba
      11'h3FD: dout  = 8'b11101110; // 1021 : 238 - 0xee
      11'h3FE: dout  = 8'b11111110; // 1022 : 254 - 0xfe
      11'h3FF: dout  = 8'b00111000; // 1023 :  56 - 0x38
      11'h400: dout  = 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x80
      11'h401: dout  = 8'b00010101; // 1025 :  21 - 0x15
      11'h402: dout  = 8'b00111111; // 1026 :  63 - 0x3f
      11'h403: dout  = 8'b01100010; // 1027 :  98 - 0x62
      11'h404: dout  = 8'b01011111; // 1028 :  95 - 0x5f
      11'h405: dout  = 8'b11111111; // 1029 : 255 - 0xff
      11'h406: dout  = 8'b10011111; // 1030 : 159 - 0x9f
      11'h407: dout  = 8'b01111101; // 1031 : 125 - 0x7d
      11'h408: dout  = 8'b00000000; // 1032 :   0 - 0x0 -- Sprite 0x81
      11'h409: dout  = 8'b00000000; // 1033 :   0 - 0x0
      11'h40A: dout  = 8'b00000000; // 1034 :   0 - 0x0
      11'h40B: dout  = 8'b00000000; // 1035 :   0 - 0x0
      11'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      11'h40D: dout  = 8'b00000000; // 1037 :   0 - 0x0
      11'h40E: dout  = 8'b00000000; // 1038 :   0 - 0x0
      11'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      11'h410: dout  = 8'b00101111; // 1040 :  47 - 0x2f -- Sprite 0x82
      11'h411: dout  = 8'b00011110; // 1041 :  30 - 0x1e
      11'h412: dout  = 8'b00101111; // 1042 :  47 - 0x2f
      11'h413: dout  = 8'b00101111; // 1043 :  47 - 0x2f
      11'h414: dout  = 8'b00101111; // 1044 :  47 - 0x2f
      11'h415: dout  = 8'b00010101; // 1045 :  21 - 0x15
      11'h416: dout  = 8'b00001101; // 1046 :  13 - 0xd
      11'h417: dout  = 8'b00001110; // 1047 :  14 - 0xe
      11'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0 -- Sprite 0x83
      11'h419: dout  = 8'b00000000; // 1049 :   0 - 0x0
      11'h41A: dout  = 8'b00000000; // 1050 :   0 - 0x0
      11'h41B: dout  = 8'b00000000; // 1051 :   0 - 0x0
      11'h41C: dout  = 8'b00000000; // 1052 :   0 - 0x0
      11'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      11'h41E: dout  = 8'b00000000; // 1054 :   0 - 0x0
      11'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      11'h420: dout  = 8'b00011100; // 1056 :  28 - 0x1c -- Sprite 0x84
      11'h421: dout  = 8'b00111110; // 1057 :  62 - 0x3e
      11'h422: dout  = 8'b01111111; // 1058 : 127 - 0x7f
      11'h423: dout  = 8'b11111111; // 1059 : 255 - 0xff
      11'h424: dout  = 8'b11111111; // 1060 : 255 - 0xff
      11'h425: dout  = 8'b11111110; // 1061 : 254 - 0xfe
      11'h426: dout  = 8'b01111100; // 1062 : 124 - 0x7c
      11'h427: dout  = 8'b00111000; // 1063 :  56 - 0x38
      11'h428: dout  = 8'b00000000; // 1064 :   0 - 0x0 -- Sprite 0x85
      11'h429: dout  = 8'b11111111; // 1065 : 255 - 0xff
      11'h42A: dout  = 8'b11111111; // 1066 : 255 - 0xff
      11'h42B: dout  = 8'b11111111; // 1067 : 255 - 0xff
      11'h42C: dout  = 8'b11111111; // 1068 : 255 - 0xff
      11'h42D: dout  = 8'b11111111; // 1069 : 255 - 0xff
      11'h42E: dout  = 8'b11111111; // 1070 : 255 - 0xff
      11'h42F: dout  = 8'b11111111; // 1071 : 255 - 0xff
      11'h430: dout  = 8'b11111111; // 1072 : 255 - 0xff -- Sprite 0x86
      11'h431: dout  = 8'b11111111; // 1073 : 255 - 0xff
      11'h432: dout  = 8'b11111111; // 1074 : 255 - 0xff
      11'h433: dout  = 8'b11111111; // 1075 : 255 - 0xff
      11'h434: dout  = 8'b11111111; // 1076 : 255 - 0xff
      11'h435: dout  = 8'b11111111; // 1077 : 255 - 0xff
      11'h436: dout  = 8'b11111111; // 1078 : 255 - 0xff
      11'h437: dout  = 8'b11111111; // 1079 : 255 - 0xff
      11'h438: dout  = 8'b01111111; // 1080 : 127 - 0x7f -- Sprite 0x87
      11'h439: dout  = 8'b11111111; // 1081 : 255 - 0xff
      11'h43A: dout  = 8'b11111111; // 1082 : 255 - 0xff
      11'h43B: dout  = 8'b11111111; // 1083 : 255 - 0xff
      11'h43C: dout  = 8'b11111111; // 1084 : 255 - 0xff
      11'h43D: dout  = 8'b11111111; // 1085 : 255 - 0xff
      11'h43E: dout  = 8'b11111111; // 1086 : 255 - 0xff
      11'h43F: dout  = 8'b11111111; // 1087 : 255 - 0xff
      11'h440: dout  = 8'b01101000; // 1088 : 104 - 0x68 -- Sprite 0x88
      11'h441: dout  = 8'b01001110; // 1089 :  78 - 0x4e
      11'h442: dout  = 8'b11100000; // 1090 : 224 - 0xe0
      11'h443: dout  = 8'b11100000; // 1091 : 224 - 0xe0
      11'h444: dout  = 8'b11100000; // 1092 : 224 - 0xe0
      11'h445: dout  = 8'b11110000; // 1093 : 240 - 0xf0
      11'h446: dout  = 8'b11111000; // 1094 : 248 - 0xf8
      11'h447: dout  = 8'b11111100; // 1095 : 252 - 0xfc
      11'h448: dout  = 8'b00111111; // 1096 :  63 - 0x3f -- Sprite 0x89
      11'h449: dout  = 8'b01011100; // 1097 :  92 - 0x5c
      11'h44A: dout  = 8'b00111001; // 1098 :  57 - 0x39
      11'h44B: dout  = 8'b00111011; // 1099 :  59 - 0x3b
      11'h44C: dout  = 8'b10111011; // 1100 : 187 - 0xbb
      11'h44D: dout  = 8'b11111001; // 1101 : 249 - 0xf9
      11'h44E: dout  = 8'b11111100; // 1102 : 252 - 0xfc
      11'h44F: dout  = 8'b11111110; // 1103 : 254 - 0xfe
      11'h450: dout  = 8'b11000000; // 1104 : 192 - 0xc0 -- Sprite 0x8a
      11'h451: dout  = 8'b11110000; // 1105 : 240 - 0xf0
      11'h452: dout  = 8'b11110000; // 1106 : 240 - 0xf0
      11'h453: dout  = 8'b11110000; // 1107 : 240 - 0xf0
      11'h454: dout  = 8'b11110000; // 1108 : 240 - 0xf0
      11'h455: dout  = 8'b11100000; // 1109 : 224 - 0xe0
      11'h456: dout  = 8'b11000000; // 1110 : 192 - 0xc0
      11'h457: dout  = 8'b00000000; // 1111 :   0 - 0x0
      11'h458: dout  = 8'b11111110; // 1112 : 254 - 0xfe -- Sprite 0x8b
      11'h459: dout  = 8'b11111100; // 1113 : 252 - 0xfc
      11'h45A: dout  = 8'b01100001; // 1114 :  97 - 0x61
      11'h45B: dout  = 8'b00001111; // 1115 :  15 - 0xf
      11'h45C: dout  = 8'b11111111; // 1116 : 255 - 0xff
      11'h45D: dout  = 8'b11111110; // 1117 : 254 - 0xfe
      11'h45E: dout  = 8'b11110000; // 1118 : 240 - 0xf0
      11'h45F: dout  = 8'b11100000; // 1119 : 224 - 0xe0
      11'h460: dout  = 8'b01101110; // 1120 : 110 - 0x6e -- Sprite 0x8c
      11'h461: dout  = 8'b01000000; // 1121 :  64 - 0x40
      11'h462: dout  = 8'b11100000; // 1122 : 224 - 0xe0
      11'h463: dout  = 8'b11100000; // 1123 : 224 - 0xe0
      11'h464: dout  = 8'b11100000; // 1124 : 224 - 0xe0
      11'h465: dout  = 8'b11100000; // 1125 : 224 - 0xe0
      11'h466: dout  = 8'b11100000; // 1126 : 224 - 0xe0
      11'h467: dout  = 8'b11000000; // 1127 : 192 - 0xc0
      11'h468: dout  = 8'b00000001; // 1128 :   1 - 0x1 -- Sprite 0x8d
      11'h469: dout  = 8'b00000001; // 1129 :   1 - 0x1
      11'h46A: dout  = 8'b00000011; // 1130 :   3 - 0x3
      11'h46B: dout  = 8'b00000011; // 1131 :   3 - 0x3
      11'h46C: dout  = 8'b00000111; // 1132 :   7 - 0x7
      11'h46D: dout  = 8'b01111111; // 1133 : 127 - 0x7f
      11'h46E: dout  = 8'b01111111; // 1134 : 127 - 0x7f
      11'h46F: dout  = 8'b00111111; // 1135 :  63 - 0x3f
      11'h470: dout  = 8'b00000110; // 1136 :   6 - 0x6 -- Sprite 0x8e
      11'h471: dout  = 8'b00000111; // 1137 :   7 - 0x7
      11'h472: dout  = 8'b00111111; // 1138 :  63 - 0x3f
      11'h473: dout  = 8'b00111100; // 1139 :  60 - 0x3c
      11'h474: dout  = 8'b00011001; // 1140 :  25 - 0x19
      11'h475: dout  = 8'b01111011; // 1141 : 123 - 0x7b
      11'h476: dout  = 8'b01111111; // 1142 : 127 - 0x7f
      11'h477: dout  = 8'b00111111; // 1143 :  63 - 0x3f
      11'h478: dout  = 8'b00111111; // 1144 :  63 - 0x3f -- Sprite 0x8f
      11'h479: dout  = 8'b01111111; // 1145 : 127 - 0x7f
      11'h47A: dout  = 8'b01111111; // 1146 : 127 - 0x7f
      11'h47B: dout  = 8'b00011111; // 1147 :  31 - 0x1f
      11'h47C: dout  = 8'b00111111; // 1148 :  63 - 0x3f
      11'h47D: dout  = 8'b00111111; // 1149 :  63 - 0x3f
      11'h47E: dout  = 8'b00000111; // 1150 :   7 - 0x7
      11'h47F: dout  = 8'b00000110; // 1151 :   6 - 0x6
      11'h480: dout  = 8'b00000011; // 1152 :   3 - 0x3 -- Sprite 0x90
      11'h481: dout  = 8'b00000111; // 1153 :   7 - 0x7
      11'h482: dout  = 8'b00001111; // 1154 :  15 - 0xf
      11'h483: dout  = 8'b00001111; // 1155 :  15 - 0xf
      11'h484: dout  = 8'b00001111; // 1156 :  15 - 0xf
      11'h485: dout  = 8'b00001111; // 1157 :  15 - 0xf
      11'h486: dout  = 8'b00000111; // 1158 :   7 - 0x7
      11'h487: dout  = 8'b00000011; // 1159 :   3 - 0x3
      11'h488: dout  = 8'b11111000; // 1160 : 248 - 0xf8 -- Sprite 0x91
      11'h489: dout  = 8'b11111000; // 1161 : 248 - 0xf8
      11'h48A: dout  = 8'b11111000; // 1162 : 248 - 0xf8
      11'h48B: dout  = 8'b10100000; // 1163 : 160 - 0xa0
      11'h48C: dout  = 8'b11100001; // 1164 : 225 - 0xe1
      11'h48D: dout  = 8'b11111111; // 1165 : 255 - 0xff
      11'h48E: dout  = 8'b11111111; // 1166 : 255 - 0xff
      11'h48F: dout  = 8'b11111111; // 1167 : 255 - 0xff
      11'h490: dout  = 8'b00001111; // 1168 :  15 - 0xf -- Sprite 0x92
      11'h491: dout  = 8'b00001111; // 1169 :  15 - 0xf
      11'h492: dout  = 8'b00001111; // 1170 :  15 - 0xf
      11'h493: dout  = 8'b00011111; // 1171 :  31 - 0x1f
      11'h494: dout  = 8'b00011111; // 1172 :  31 - 0x1f
      11'h495: dout  = 8'b00011111; // 1173 :  31 - 0x1f
      11'h496: dout  = 8'b00001111; // 1174 :  15 - 0xf
      11'h497: dout  = 8'b00000111; // 1175 :   7 - 0x7
      11'h498: dout  = 8'b11100000; // 1176 : 224 - 0xe0 -- Sprite 0x93
      11'h499: dout  = 8'b11111000; // 1177 : 248 - 0xf8
      11'h49A: dout  = 8'b11111000; // 1178 : 248 - 0xf8
      11'h49B: dout  = 8'b11111000; // 1179 : 248 - 0xf8
      11'h49C: dout  = 8'b11111111; // 1180 : 255 - 0xff
      11'h49D: dout  = 8'b11111110; // 1181 : 254 - 0xfe
      11'h49E: dout  = 8'b11110000; // 1182 : 240 - 0xf0
      11'h49F: dout  = 8'b11000000; // 1183 : 192 - 0xc0
      11'h4A0: dout  = 8'b00000001; // 1184 :   1 - 0x1 -- Sprite 0x94
      11'h4A1: dout  = 8'b00001111; // 1185 :  15 - 0xf
      11'h4A2: dout  = 8'b00001111; // 1186 :  15 - 0xf
      11'h4A3: dout  = 8'b00011111; // 1187 :  31 - 0x1f
      11'h4A4: dout  = 8'b00111001; // 1188 :  57 - 0x39
      11'h4A5: dout  = 8'b00110011; // 1189 :  51 - 0x33
      11'h4A6: dout  = 8'b00110111; // 1190 :  55 - 0x37
      11'h4A7: dout  = 8'b01111111; // 1191 : 127 - 0x7f
      11'h4A8: dout  = 8'b01111111; // 1192 : 127 - 0x7f -- Sprite 0x95
      11'h4A9: dout  = 8'b00111111; // 1193 :  63 - 0x3f
      11'h4AA: dout  = 8'b00111111; // 1194 :  63 - 0x3f
      11'h4AB: dout  = 8'b00111111; // 1195 :  63 - 0x3f
      11'h4AC: dout  = 8'b00011111; // 1196 :  31 - 0x1f
      11'h4AD: dout  = 8'b00001111; // 1197 :  15 - 0xf
      11'h4AE: dout  = 8'b00001111; // 1198 :  15 - 0xf
      11'h4AF: dout  = 8'b00000001; // 1199 :   1 - 0x1
      11'h4B0: dout  = 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x96
      11'h4B1: dout  = 8'b00000000; // 1201 :   0 - 0x0
      11'h4B2: dout  = 8'b00000011; // 1202 :   3 - 0x3
      11'h4B3: dout  = 8'b00000011; // 1203 :   3 - 0x3
      11'h4B4: dout  = 8'b01000111; // 1204 :  71 - 0x47
      11'h4B5: dout  = 8'b01100111; // 1205 : 103 - 0x67
      11'h4B6: dout  = 8'b01110111; // 1206 : 119 - 0x77
      11'h4B7: dout  = 8'b01110111; // 1207 : 119 - 0x77
      11'h4B8: dout  = 8'b00000000; // 1208 :   0 - 0x0 -- Sprite 0x97
      11'h4B9: dout  = 8'b00000000; // 1209 :   0 - 0x0
      11'h4BA: dout  = 8'b00000000; // 1210 :   0 - 0x0
      11'h4BB: dout  = 8'b00000000; // 1211 :   0 - 0x0
      11'h4BC: dout  = 8'b10001000; // 1212 : 136 - 0x88
      11'h4BD: dout  = 8'b10011000; // 1213 : 152 - 0x98
      11'h4BE: dout  = 8'b11111000; // 1214 : 248 - 0xf8
      11'h4BF: dout  = 8'b11110000; // 1215 : 240 - 0xf0
      11'h4C0: dout  = 8'b01111110; // 1216 : 126 - 0x7e -- Sprite 0x98
      11'h4C1: dout  = 8'b01111111; // 1217 : 127 - 0x7f
      11'h4C2: dout  = 8'b11111111; // 1218 : 255 - 0xff
      11'h4C3: dout  = 8'b00011111; // 1219 :  31 - 0x1f
      11'h4C4: dout  = 8'b00000111; // 1220 :   7 - 0x7
      11'h4C5: dout  = 8'b00110000; // 1221 :  48 - 0x30
      11'h4C6: dout  = 8'b00011100; // 1222 :  28 - 0x1c
      11'h4C7: dout  = 8'b00001100; // 1223 :  12 - 0xc
      11'h4C8: dout  = 8'b01111110; // 1224 : 126 - 0x7e -- Sprite 0x99
      11'h4C9: dout  = 8'b00111000; // 1225 :  56 - 0x38
      11'h4CA: dout  = 8'b11110110; // 1226 : 246 - 0xf6
      11'h4CB: dout  = 8'b11101101; // 1227 : 237 - 0xed
      11'h4CC: dout  = 8'b11011111; // 1228 : 223 - 0xdf
      11'h4CD: dout  = 8'b00111000; // 1229 :  56 - 0x38
      11'h4CE: dout  = 8'b01110000; // 1230 : 112 - 0x70
      11'h4CF: dout  = 8'b01100000; // 1231 :  96 - 0x60
      11'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      11'h4D1: dout  = 8'b00000000; // 1233 :   0 - 0x0
      11'h4D2: dout  = 8'b00000000; // 1234 :   0 - 0x0
      11'h4D3: dout  = 8'b00000011; // 1235 :   3 - 0x3
      11'h4D4: dout  = 8'b00000011; // 1236 :   3 - 0x3
      11'h4D5: dout  = 8'b01000111; // 1237 :  71 - 0x47
      11'h4D6: dout  = 8'b01100111; // 1238 : 103 - 0x67
      11'h4D7: dout  = 8'b01110111; // 1239 : 119 - 0x77
      11'h4D8: dout  = 8'b00000000; // 1240 :   0 - 0x0 -- Sprite 0x9b
      11'h4D9: dout  = 8'b00000000; // 1241 :   0 - 0x0
      11'h4DA: dout  = 8'b00000000; // 1242 :   0 - 0x0
      11'h4DB: dout  = 8'b00000000; // 1243 :   0 - 0x0
      11'h4DC: dout  = 8'b00000000; // 1244 :   0 - 0x0
      11'h4DD: dout  = 8'b10001000; // 1245 : 136 - 0x88
      11'h4DE: dout  = 8'b10011000; // 1246 : 152 - 0x98
      11'h4DF: dout  = 8'b11111000; // 1247 : 248 - 0xf8
      11'h4E0: dout  = 8'b01110111; // 1248 : 119 - 0x77 -- Sprite 0x9c
      11'h4E1: dout  = 8'b01111110; // 1249 : 126 - 0x7e
      11'h4E2: dout  = 8'b01111111; // 1250 : 127 - 0x7f
      11'h4E3: dout  = 8'b11111111; // 1251 : 255 - 0xff
      11'h4E4: dout  = 8'b00011111; // 1252 :  31 - 0x1f
      11'h4E5: dout  = 8'b00000111; // 1253 :   7 - 0x7
      11'h4E6: dout  = 8'b01110000; // 1254 : 112 - 0x70
      11'h4E7: dout  = 8'b11110000; // 1255 : 240 - 0xf0
      11'h4E8: dout  = 8'b11110000; // 1256 : 240 - 0xf0 -- Sprite 0x9d
      11'h4E9: dout  = 8'b01111110; // 1257 : 126 - 0x7e
      11'h4EA: dout  = 8'b00111000; // 1258 :  56 - 0x38
      11'h4EB: dout  = 8'b11110110; // 1259 : 246 - 0xf6
      11'h4EC: dout  = 8'b11101101; // 1260 : 237 - 0xed
      11'h4ED: dout  = 8'b11011111; // 1261 : 223 - 0xdf
      11'h4EE: dout  = 8'b00111000; // 1262 :  56 - 0x38
      11'h4EF: dout  = 8'b00111100; // 1263 :  60 - 0x3c
      11'h4F0: dout  = 8'b00000011; // 1264 :   3 - 0x3 -- Sprite 0x9e
      11'h4F1: dout  = 8'b00000111; // 1265 :   7 - 0x7
      11'h4F2: dout  = 8'b00001010; // 1266 :  10 - 0xa
      11'h4F3: dout  = 8'b00011010; // 1267 :  26 - 0x1a
      11'h4F4: dout  = 8'b00011100; // 1268 :  28 - 0x1c
      11'h4F5: dout  = 8'b00011110; // 1269 :  30 - 0x1e
      11'h4F6: dout  = 8'b00001011; // 1270 :  11 - 0xb
      11'h4F7: dout  = 8'b00001000; // 1271 :   8 - 0x8
      11'h4F8: dout  = 8'b00011100; // 1272 :  28 - 0x1c -- Sprite 0x9f
      11'h4F9: dout  = 8'b00111111; // 1273 :  63 - 0x3f
      11'h4FA: dout  = 8'b00111111; // 1274 :  63 - 0x3f
      11'h4FB: dout  = 8'b00111101; // 1275 :  61 - 0x3d
      11'h4FC: dout  = 8'b00111111; // 1276 :  63 - 0x3f
      11'h4FD: dout  = 8'b00011111; // 1277 :  31 - 0x1f
      11'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      11'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0xa0
      11'h501: dout  = 8'b00000000; // 1281 :   0 - 0x0
      11'h502: dout  = 8'b00000100; // 1282 :   4 - 0x4
      11'h503: dout  = 8'b01001100; // 1283 :  76 - 0x4c
      11'h504: dout  = 8'b01001110; // 1284 :  78 - 0x4e
      11'h505: dout  = 8'b01001110; // 1285 :  78 - 0x4e
      11'h506: dout  = 8'b01000110; // 1286 :  70 - 0x46
      11'h507: dout  = 8'b01101111; // 1287 : 111 - 0x6f
      11'h508: dout  = 8'b00000000; // 1288 :   0 - 0x0 -- Sprite 0xa1
      11'h509: dout  = 8'b00011111; // 1289 :  31 - 0x1f
      11'h50A: dout  = 8'b00111111; // 1290 :  63 - 0x3f
      11'h50B: dout  = 8'b00111111; // 1291 :  63 - 0x3f
      11'h50C: dout  = 8'b01001111; // 1292 :  79 - 0x4f
      11'h50D: dout  = 8'b01011111; // 1293 :  95 - 0x5f
      11'h50E: dout  = 8'b01111111; // 1294 : 127 - 0x7f
      11'h50F: dout  = 8'b01111111; // 1295 : 127 - 0x7f
      11'h510: dout  = 8'b01111111; // 1296 : 127 - 0x7f -- Sprite 0xa2
      11'h511: dout  = 8'b01100111; // 1297 : 103 - 0x67
      11'h512: dout  = 8'b10100011; // 1298 : 163 - 0xa3
      11'h513: dout  = 8'b10110000; // 1299 : 176 - 0xb0
      11'h514: dout  = 8'b11011000; // 1300 : 216 - 0xd8
      11'h515: dout  = 8'b11011110; // 1301 : 222 - 0xde
      11'h516: dout  = 8'b11011100; // 1302 : 220 - 0xdc
      11'h517: dout  = 8'b11001000; // 1303 : 200 - 0xc8
      11'h518: dout  = 8'b01111111; // 1304 : 127 - 0x7f -- Sprite 0xa3
      11'h519: dout  = 8'b01111111; // 1305 : 127 - 0x7f
      11'h51A: dout  = 8'b01111111; // 1306 : 127 - 0x7f
      11'h51B: dout  = 8'b00011111; // 1307 :  31 - 0x1f
      11'h51C: dout  = 8'b01000111; // 1308 :  71 - 0x47
      11'h51D: dout  = 8'b01110000; // 1309 : 112 - 0x70
      11'h51E: dout  = 8'b01110000; // 1310 : 112 - 0x70
      11'h51F: dout  = 8'b00111001; // 1311 :  57 - 0x39
      11'h520: dout  = 8'b11101000; // 1312 : 232 - 0xe8 -- Sprite 0xa4
      11'h521: dout  = 8'b11101000; // 1313 : 232 - 0xe8
      11'h522: dout  = 8'b11100000; // 1314 : 224 - 0xe0
      11'h523: dout  = 8'b11000000; // 1315 : 192 - 0xc0
      11'h524: dout  = 8'b00010000; // 1316 :  16 - 0x10
      11'h525: dout  = 8'b01110000; // 1317 : 112 - 0x70
      11'h526: dout  = 8'b11100000; // 1318 : 224 - 0xe0
      11'h527: dout  = 8'b11000000; // 1319 : 192 - 0xc0
      11'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- Sprite 0xa5
      11'h529: dout  = 8'b00000000; // 1321 :   0 - 0x0
      11'h52A: dout  = 8'b00000000; // 1322 :   0 - 0x0
      11'h52B: dout  = 8'b00100000; // 1323 :  32 - 0x20
      11'h52C: dout  = 8'b01100110; // 1324 : 102 - 0x66
      11'h52D: dout  = 8'b01100110; // 1325 : 102 - 0x66
      11'h52E: dout  = 8'b01100110; // 1326 : 102 - 0x66
      11'h52F: dout  = 8'b01100010; // 1327 :  98 - 0x62
      11'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0xa6
      11'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      11'h532: dout  = 8'b00011111; // 1330 :  31 - 0x1f
      11'h533: dout  = 8'b00111111; // 1331 :  63 - 0x3f
      11'h534: dout  = 8'b01111111; // 1332 : 127 - 0x7f
      11'h535: dout  = 8'b01001111; // 1333 :  79 - 0x4f
      11'h536: dout  = 8'b01011111; // 1334 :  95 - 0x5f
      11'h537: dout  = 8'b01111111; // 1335 : 127 - 0x7f
      11'h538: dout  = 8'b01110111; // 1336 : 119 - 0x77 -- Sprite 0xa7
      11'h539: dout  = 8'b01111111; // 1337 : 127 - 0x7f
      11'h53A: dout  = 8'b00111111; // 1338 :  63 - 0x3f
      11'h53B: dout  = 8'b10110111; // 1339 : 183 - 0xb7
      11'h53C: dout  = 8'b10110011; // 1340 : 179 - 0xb3
      11'h53D: dout  = 8'b11011011; // 1341 : 219 - 0xdb
      11'h53E: dout  = 8'b11011010; // 1342 : 218 - 0xda
      11'h53F: dout  = 8'b11011000; // 1343 : 216 - 0xd8
      11'h540: dout  = 8'b01111111; // 1344 : 127 - 0x7f -- Sprite 0xa8
      11'h541: dout  = 8'b01111111; // 1345 : 127 - 0x7f
      11'h542: dout  = 8'b01111111; // 1346 : 127 - 0x7f
      11'h543: dout  = 8'b01111111; // 1347 : 127 - 0x7f
      11'h544: dout  = 8'b00011111; // 1348 :  31 - 0x1f
      11'h545: dout  = 8'b00000111; // 1349 :   7 - 0x7
      11'h546: dout  = 8'b01110000; // 1350 : 112 - 0x70
      11'h547: dout  = 8'b11110000; // 1351 : 240 - 0xf0
      11'h548: dout  = 8'b11001100; // 1352 : 204 - 0xcc -- Sprite 0xa9
      11'h549: dout  = 8'b11101000; // 1353 : 232 - 0xe8
      11'h54A: dout  = 8'b11101000; // 1354 : 232 - 0xe8
      11'h54B: dout  = 8'b11100000; // 1355 : 224 - 0xe0
      11'h54C: dout  = 8'b11000000; // 1356 : 192 - 0xc0
      11'h54D: dout  = 8'b00011000; // 1357 :  24 - 0x18
      11'h54E: dout  = 8'b01111100; // 1358 : 124 - 0x7c
      11'h54F: dout  = 8'b00111110; // 1359 :  62 - 0x3e
      11'h550: dout  = 8'b00000011; // 1360 :   3 - 0x3 -- Sprite 0xaa
      11'h551: dout  = 8'b00001111; // 1361 :  15 - 0xf
      11'h552: dout  = 8'b00011111; // 1362 :  31 - 0x1f
      11'h553: dout  = 8'b00111111; // 1363 :  63 - 0x3f
      11'h554: dout  = 8'b00111011; // 1364 :  59 - 0x3b
      11'h555: dout  = 8'b00111111; // 1365 :  63 - 0x3f
      11'h556: dout  = 8'b01111111; // 1366 : 127 - 0x7f
      11'h557: dout  = 8'b01111111; // 1367 : 127 - 0x7f
      11'h558: dout  = 8'b10000000; // 1368 : 128 - 0x80 -- Sprite 0xab
      11'h559: dout  = 8'b11110000; // 1369 : 240 - 0xf0
      11'h55A: dout  = 8'b11111000; // 1370 : 248 - 0xf8
      11'h55B: dout  = 8'b11111100; // 1371 : 252 - 0xfc
      11'h55C: dout  = 8'b11111110; // 1372 : 254 - 0xfe
      11'h55D: dout  = 8'b11111110; // 1373 : 254 - 0xfe
      11'h55E: dout  = 8'b11111111; // 1374 : 255 - 0xff
      11'h55F: dout  = 8'b11111110; // 1375 : 254 - 0xfe
      11'h560: dout  = 8'b01111111; // 1376 : 127 - 0x7f -- Sprite 0xac
      11'h561: dout  = 8'b01111111; // 1377 : 127 - 0x7f
      11'h562: dout  = 8'b01111111; // 1378 : 127 - 0x7f
      11'h563: dout  = 8'b01111111; // 1379 : 127 - 0x7f
      11'h564: dout  = 8'b11111111; // 1380 : 255 - 0xff
      11'h565: dout  = 8'b00001111; // 1381 :  15 - 0xf
      11'h566: dout  = 8'b00000011; // 1382 :   3 - 0x3
      11'h567: dout  = 8'b00000000; // 1383 :   0 - 0x0
      11'h568: dout  = 8'b11111110; // 1384 : 254 - 0xfe -- Sprite 0xad
      11'h569: dout  = 8'b11111011; // 1385 : 251 - 0xfb
      11'h56A: dout  = 8'b11111111; // 1386 : 255 - 0xff
      11'h56B: dout  = 8'b11111111; // 1387 : 255 - 0xff
      11'h56C: dout  = 8'b11110110; // 1388 : 246 - 0xf6
      11'h56D: dout  = 8'b11100000; // 1389 : 224 - 0xe0
      11'h56E: dout  = 8'b11000000; // 1390 : 192 - 0xc0
      11'h56F: dout  = 8'b00000000; // 1391 :   0 - 0x0
      11'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      11'h571: dout  = 8'b00000011; // 1393 :   3 - 0x3
      11'h572: dout  = 8'b00001111; // 1394 :  15 - 0xf
      11'h573: dout  = 8'b00011111; // 1395 :  31 - 0x1f
      11'h574: dout  = 8'b00111111; // 1396 :  63 - 0x3f
      11'h575: dout  = 8'b00111011; // 1397 :  59 - 0x3b
      11'h576: dout  = 8'b00111111; // 1398 :  63 - 0x3f
      11'h577: dout  = 8'b01111111; // 1399 : 127 - 0x7f
      11'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Sprite 0xaf
      11'h579: dout  = 8'b11000000; // 1401 : 192 - 0xc0
      11'h57A: dout  = 8'b11110000; // 1402 : 240 - 0xf0
      11'h57B: dout  = 8'b11111000; // 1403 : 248 - 0xf8
      11'h57C: dout  = 8'b11111100; // 1404 : 252 - 0xfc
      11'h57D: dout  = 8'b11111110; // 1405 : 254 - 0xfe
      11'h57E: dout  = 8'b11111110; // 1406 : 254 - 0xfe
      11'h57F: dout  = 8'b11111111; // 1407 : 255 - 0xff
      11'h580: dout  = 8'b01111111; // 1408 : 127 - 0x7f -- Sprite 0xb0
      11'h581: dout  = 8'b01111111; // 1409 : 127 - 0x7f
      11'h582: dout  = 8'b01111111; // 1410 : 127 - 0x7f
      11'h583: dout  = 8'b01111111; // 1411 : 127 - 0x7f
      11'h584: dout  = 8'b01111111; // 1412 : 127 - 0x7f
      11'h585: dout  = 8'b11111111; // 1413 : 255 - 0xff
      11'h586: dout  = 8'b00001111; // 1414 :  15 - 0xf
      11'h587: dout  = 8'b00000011; // 1415 :   3 - 0x3
      11'h588: dout  = 8'b11111110; // 1416 : 254 - 0xfe -- Sprite 0xb1
      11'h589: dout  = 8'b11111110; // 1417 : 254 - 0xfe
      11'h58A: dout  = 8'b11111011; // 1418 : 251 - 0xfb
      11'h58B: dout  = 8'b11111111; // 1419 : 255 - 0xff
      11'h58C: dout  = 8'b11111111; // 1420 : 255 - 0xff
      11'h58D: dout  = 8'b11110110; // 1421 : 246 - 0xf6
      11'h58E: dout  = 8'b11100000; // 1422 : 224 - 0xe0
      11'h58F: dout  = 8'b11000000; // 1423 : 192 - 0xc0
      11'h590: dout  = 8'b00000000; // 1424 :   0 - 0x0 -- Sprite 0xb2
      11'h591: dout  = 8'b00000001; // 1425 :   1 - 0x1
      11'h592: dout  = 8'b00000001; // 1426 :   1 - 0x1
      11'h593: dout  = 8'b00000001; // 1427 :   1 - 0x1
      11'h594: dout  = 8'b00000001; // 1428 :   1 - 0x1
      11'h595: dout  = 8'b00000000; // 1429 :   0 - 0x0
      11'h596: dout  = 8'b00000000; // 1430 :   0 - 0x0
      11'h597: dout  = 8'b00001000; // 1431 :   8 - 0x8
      11'h598: dout  = 8'b01111000; // 1432 : 120 - 0x78 -- Sprite 0xb3
      11'h599: dout  = 8'b11110000; // 1433 : 240 - 0xf0
      11'h59A: dout  = 8'b11111000; // 1434 : 248 - 0xf8
      11'h59B: dout  = 8'b11100100; // 1435 : 228 - 0xe4
      11'h59C: dout  = 8'b11000000; // 1436 : 192 - 0xc0
      11'h59D: dout  = 8'b11001010; // 1437 : 202 - 0xca
      11'h59E: dout  = 8'b11001010; // 1438 : 202 - 0xca
      11'h59F: dout  = 8'b11000000; // 1439 : 192 - 0xc0
      11'h5A0: dout  = 8'b00001111; // 1440 :  15 - 0xf -- Sprite 0xb4
      11'h5A1: dout  = 8'b00011111; // 1441 :  31 - 0x1f
      11'h5A2: dout  = 8'b10011111; // 1442 : 159 - 0x9f
      11'h5A3: dout  = 8'b11111111; // 1443 : 255 - 0xff
      11'h5A4: dout  = 8'b11111111; // 1444 : 255 - 0xff
      11'h5A5: dout  = 8'b01111111; // 1445 : 127 - 0x7f
      11'h5A6: dout  = 8'b01110100; // 1446 : 116 - 0x74
      11'h5A7: dout  = 8'b00100000; // 1447 :  32 - 0x20
      11'h5A8: dout  = 8'b11100100; // 1448 : 228 - 0xe4 -- Sprite 0xb5
      11'h5A9: dout  = 8'b11111111; // 1449 : 255 - 0xff
      11'h5AA: dout  = 8'b11111110; // 1450 : 254 - 0xfe
      11'h5AB: dout  = 8'b11111100; // 1451 : 252 - 0xfc
      11'h5AC: dout  = 8'b10011100; // 1452 : 156 - 0x9c
      11'h5AD: dout  = 8'b00011110; // 1453 :  30 - 0x1e
      11'h5AE: dout  = 8'b00000000; // 1454 :   0 - 0x0
      11'h5AF: dout  = 8'b00000000; // 1455 :   0 - 0x0
      11'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0xb6
      11'h5B1: dout  = 8'b00000001; // 1457 :   1 - 0x1
      11'h5B2: dout  = 8'b00000011; // 1458 :   3 - 0x3
      11'h5B3: dout  = 8'b00000011; // 1459 :   3 - 0x3
      11'h5B4: dout  = 8'b00000111; // 1460 :   7 - 0x7
      11'h5B5: dout  = 8'b00000011; // 1461 :   3 - 0x3
      11'h5B6: dout  = 8'b00000001; // 1462 :   1 - 0x1
      11'h5B7: dout  = 8'b00000000; // 1463 :   0 - 0x0
      11'h5B8: dout  = 8'b00000000; // 1464 :   0 - 0x0 -- Sprite 0xb7
      11'h5B9: dout  = 8'b01011111; // 1465 :  95 - 0x5f
      11'h5BA: dout  = 8'b01111111; // 1466 : 127 - 0x7f
      11'h5BB: dout  = 8'b01111111; // 1467 : 127 - 0x7f
      11'h5BC: dout  = 8'b00111111; // 1468 :  63 - 0x3f
      11'h5BD: dout  = 8'b00111111; // 1469 :  63 - 0x3f
      11'h5BE: dout  = 8'b00010100; // 1470 :  20 - 0x14
      11'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      11'h5C0: dout  = 8'b11000000; // 1472 : 192 - 0xc0 -- Sprite 0xb8
      11'h5C1: dout  = 8'b11100000; // 1473 : 224 - 0xe0
      11'h5C2: dout  = 8'b11110000; // 1474 : 240 - 0xf0
      11'h5C3: dout  = 8'b00110000; // 1475 :  48 - 0x30
      11'h5C4: dout  = 8'b00111000; // 1476 :  56 - 0x38
      11'h5C5: dout  = 8'b00111100; // 1477 :  60 - 0x3c
      11'h5C6: dout  = 8'b00111100; // 1478 :  60 - 0x3c
      11'h5C7: dout  = 8'b11111100; // 1479 : 252 - 0xfc
      11'h5C8: dout  = 8'b00000111; // 1480 :   7 - 0x7 -- Sprite 0xb9
      11'h5C9: dout  = 8'b00001111; // 1481 :  15 - 0xf
      11'h5CA: dout  = 8'b00011111; // 1482 :  31 - 0x1f
      11'h5CB: dout  = 8'b00100010; // 1483 :  34 - 0x22
      11'h5CC: dout  = 8'b00100000; // 1484 :  32 - 0x20
      11'h5CD: dout  = 8'b00100101; // 1485 :  37 - 0x25
      11'h5CE: dout  = 8'b00100101; // 1486 :  37 - 0x25
      11'h5CF: dout  = 8'b00011111; // 1487 :  31 - 0x1f
      11'h5D0: dout  = 8'b11111110; // 1488 : 254 - 0xfe -- Sprite 0xba
      11'h5D1: dout  = 8'b11111110; // 1489 : 254 - 0xfe
      11'h5D2: dout  = 8'b01111110; // 1490 : 126 - 0x7e
      11'h5D3: dout  = 8'b00111010; // 1491 :  58 - 0x3a
      11'h5D4: dout  = 8'b00000010; // 1492 :   2 - 0x2
      11'h5D5: dout  = 8'b00000001; // 1493 :   1 - 0x1
      11'h5D6: dout  = 8'b01000001; // 1494 :  65 - 0x41
      11'h5D7: dout  = 8'b01000001; // 1495 :  65 - 0x41
      11'h5D8: dout  = 8'b00011111; // 1496 :  31 - 0x1f -- Sprite 0xbb
      11'h5D9: dout  = 8'b00111111; // 1497 :  63 - 0x3f
      11'h5DA: dout  = 8'b01111110; // 1498 : 126 - 0x7e
      11'h5DB: dout  = 8'b01011100; // 1499 :  92 - 0x5c
      11'h5DC: dout  = 8'b01000000; // 1500 :  64 - 0x40
      11'h5DD: dout  = 8'b10000000; // 1501 : 128 - 0x80
      11'h5DE: dout  = 8'b10000010; // 1502 : 130 - 0x82
      11'h5DF: dout  = 8'b10000010; // 1503 : 130 - 0x82
      11'h5E0: dout  = 8'b10000010; // 1504 : 130 - 0x82 -- Sprite 0xbc
      11'h5E1: dout  = 8'b10000000; // 1505 : 128 - 0x80
      11'h5E2: dout  = 8'b10100000; // 1506 : 160 - 0xa0
      11'h5E3: dout  = 8'b01000100; // 1507 :  68 - 0x44
      11'h5E4: dout  = 8'b01000011; // 1508 :  67 - 0x43
      11'h5E5: dout  = 8'b01000000; // 1509 :  64 - 0x40
      11'h5E6: dout  = 8'b00100001; // 1510 :  33 - 0x21
      11'h5E7: dout  = 8'b00011110; // 1511 :  30 - 0x1e
      11'h5E8: dout  = 8'b00011100; // 1512 :  28 - 0x1c -- Sprite 0xbd
      11'h5E9: dout  = 8'b00111111; // 1513 :  63 - 0x3f
      11'h5EA: dout  = 8'b00111110; // 1514 :  62 - 0x3e
      11'h5EB: dout  = 8'b00111100; // 1515 :  60 - 0x3c
      11'h5EC: dout  = 8'b01000000; // 1516 :  64 - 0x40
      11'h5ED: dout  = 8'b10000000; // 1517 : 128 - 0x80
      11'h5EE: dout  = 8'b10000010; // 1518 : 130 - 0x82
      11'h5EF: dout  = 8'b10000010; // 1519 : 130 - 0x82
      11'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      11'h5F1: dout  = 8'b00000000; // 1521 :   0 - 0x0
      11'h5F2: dout  = 8'b10000000; // 1522 : 128 - 0x80
      11'h5F3: dout  = 8'b10000000; // 1523 : 128 - 0x80
      11'h5F4: dout  = 8'b10010010; // 1524 : 146 - 0x92
      11'h5F5: dout  = 8'b10011101; // 1525 : 157 - 0x9d
      11'h5F6: dout  = 8'b11000111; // 1526 : 199 - 0xc7
      11'h5F7: dout  = 8'b11101111; // 1527 : 239 - 0xef
      11'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      11'h5F9: dout  = 8'b00100011; // 1529 :  35 - 0x23
      11'h5FA: dout  = 8'b00110011; // 1530 :  51 - 0x33
      11'h5FB: dout  = 8'b00111111; // 1531 :  63 - 0x3f
      11'h5FC: dout  = 8'b00111111; // 1532 :  63 - 0x3f
      11'h5FD: dout  = 8'b01111111; // 1533 : 127 - 0x7f
      11'h5FE: dout  = 8'b01111111; // 1534 : 127 - 0x7f
      11'h5FF: dout  = 8'b01111111; // 1535 : 127 - 0x7f
      11'h600: dout  = 8'b11111110; // 1536 : 254 - 0xfe -- Sprite 0xc0
      11'h601: dout  = 8'b11111000; // 1537 : 248 - 0xf8
      11'h602: dout  = 8'b10100000; // 1538 : 160 - 0xa0
      11'h603: dout  = 8'b00000000; // 1539 :   0 - 0x0
      11'h604: dout  = 8'b00000000; // 1540 :   0 - 0x0
      11'h605: dout  = 8'b00000000; // 1541 :   0 - 0x0
      11'h606: dout  = 8'b10000000; // 1542 : 128 - 0x80
      11'h607: dout  = 8'b10000000; // 1543 : 128 - 0x80
      11'h608: dout  = 8'b01111110; // 1544 : 126 - 0x7e -- Sprite 0xc1
      11'h609: dout  = 8'b01111111; // 1545 : 127 - 0x7f
      11'h60A: dout  = 8'b01111101; // 1546 : 125 - 0x7d
      11'h60B: dout  = 8'b00111111; // 1547 :  63 - 0x3f
      11'h60C: dout  = 8'b00011110; // 1548 :  30 - 0x1e
      11'h60D: dout  = 8'b10001111; // 1549 : 143 - 0x8f
      11'h60E: dout  = 8'b10001111; // 1550 : 143 - 0x8f
      11'h60F: dout  = 8'b00011001; // 1551 :  25 - 0x19
      11'h610: dout  = 8'b11100000; // 1552 : 224 - 0xe0 -- Sprite 0xc2
      11'h611: dout  = 8'b00001110; // 1553 :  14 - 0xe
      11'h612: dout  = 8'b01110011; // 1554 : 115 - 0x73
      11'h613: dout  = 8'b11110011; // 1555 : 243 - 0xf3
      11'h614: dout  = 8'b11111001; // 1556 : 249 - 0xf9
      11'h615: dout  = 8'b11111001; // 1557 : 249 - 0xf9
      11'h616: dout  = 8'b11111000; // 1558 : 248 - 0xf8
      11'h617: dout  = 8'b01110000; // 1559 : 112 - 0x70
      11'h618: dout  = 8'b00001110; // 1560 :  14 - 0xe -- Sprite 0xc3
      11'h619: dout  = 8'b01100110; // 1561 : 102 - 0x66
      11'h61A: dout  = 8'b11100010; // 1562 : 226 - 0xe2
      11'h61B: dout  = 8'b11110110; // 1563 : 246 - 0xf6
      11'h61C: dout  = 8'b11111111; // 1564 : 255 - 0xff
      11'h61D: dout  = 8'b11111111; // 1565 : 255 - 0xff
      11'h61E: dout  = 8'b00011111; // 1566 :  31 - 0x1f
      11'h61F: dout  = 8'b10011000; // 1567 : 152 - 0x98
      11'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      11'h621: dout  = 8'b00000000; // 1569 :   0 - 0x0
      11'h622: dout  = 8'b00000000; // 1570 :   0 - 0x0
      11'h623: dout  = 8'b00000100; // 1571 :   4 - 0x4
      11'h624: dout  = 8'b00001111; // 1572 :  15 - 0xf
      11'h625: dout  = 8'b00001111; // 1573 :  15 - 0xf
      11'h626: dout  = 8'b00011111; // 1574 :  31 - 0x1f
      11'h627: dout  = 8'b00000111; // 1575 :   7 - 0x7
      11'h628: dout  = 8'b11110011; // 1576 : 243 - 0xf3 -- Sprite 0xc5
      11'h629: dout  = 8'b11100111; // 1577 : 231 - 0xe7
      11'h62A: dout  = 8'b11101110; // 1578 : 238 - 0xee
      11'h62B: dout  = 8'b11101100; // 1579 : 236 - 0xec
      11'h62C: dout  = 8'b11001101; // 1580 : 205 - 0xcd
      11'h62D: dout  = 8'b11001111; // 1581 : 207 - 0xcf
      11'h62E: dout  = 8'b11001111; // 1582 : 207 - 0xcf
      11'h62F: dout  = 8'b11011111; // 1583 : 223 - 0xdf
      11'h630: dout  = 8'b00100111; // 1584 :  39 - 0x27 -- Sprite 0xc6
      11'h631: dout  = 8'b00111111; // 1585 :  63 - 0x3f
      11'h632: dout  = 8'b00111111; // 1586 :  63 - 0x3f
      11'h633: dout  = 8'b01111000; // 1587 : 120 - 0x78
      11'h634: dout  = 8'b00111100; // 1588 :  60 - 0x3c
      11'h635: dout  = 8'b00011111; // 1589 :  31 - 0x1f
      11'h636: dout  = 8'b00011111; // 1590 :  31 - 0x1f
      11'h637: dout  = 8'b01110011; // 1591 : 115 - 0x73
      11'h638: dout  = 8'b10011111; // 1592 : 159 - 0x9f -- Sprite 0xc7
      11'h639: dout  = 8'b00111110; // 1593 :  62 - 0x3e
      11'h63A: dout  = 8'b01111100; // 1594 : 124 - 0x7c
      11'h63B: dout  = 8'b11111100; // 1595 : 252 - 0xfc
      11'h63C: dout  = 8'b11111000; // 1596 : 248 - 0xf8
      11'h63D: dout  = 8'b11111000; // 1597 : 248 - 0xf8
      11'h63E: dout  = 8'b11000000; // 1598 : 192 - 0xc0
      11'h63F: dout  = 8'b01000000; // 1599 :  64 - 0x40
      11'h640: dout  = 8'b01111111; // 1600 : 127 - 0x7f -- Sprite 0xc8
      11'h641: dout  = 8'b01111110; // 1601 : 126 - 0x7e
      11'h642: dout  = 8'b01111000; // 1602 : 120 - 0x78
      11'h643: dout  = 8'b00000001; // 1603 :   1 - 0x1
      11'h644: dout  = 8'b00000111; // 1604 :   7 - 0x7
      11'h645: dout  = 8'b00011111; // 1605 :  31 - 0x1f
      11'h646: dout  = 8'b00111100; // 1606 :  60 - 0x3c
      11'h647: dout  = 8'b01111100; // 1607 : 124 - 0x7c
      11'h648: dout  = 8'b11111100; // 1608 : 252 - 0xfc -- Sprite 0xc9
      11'h649: dout  = 8'b11111000; // 1609 : 248 - 0xf8
      11'h64A: dout  = 8'b10100000; // 1610 : 160 - 0xa0
      11'h64B: dout  = 8'b11111110; // 1611 : 254 - 0xfe
      11'h64C: dout  = 8'b11111100; // 1612 : 252 - 0xfc
      11'h64D: dout  = 8'b11110000; // 1613 : 240 - 0xf0
      11'h64E: dout  = 8'b10000000; // 1614 : 128 - 0x80
      11'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      11'h650: dout  = 8'b01111110; // 1616 : 126 - 0x7e -- Sprite 0xca
      11'h651: dout  = 8'b01111111; // 1617 : 127 - 0x7f
      11'h652: dout  = 8'b01111111; // 1618 : 127 - 0x7f
      11'h653: dout  = 8'b00111111; // 1619 :  63 - 0x3f
      11'h654: dout  = 8'b00011111; // 1620 :  31 - 0x1f
      11'h655: dout  = 8'b10001111; // 1621 : 143 - 0x8f
      11'h656: dout  = 8'b10001111; // 1622 : 143 - 0x8f
      11'h657: dout  = 8'b00011000; // 1623 :  24 - 0x18
      11'h658: dout  = 8'b10011111; // 1624 : 159 - 0x9f -- Sprite 0xcb
      11'h659: dout  = 8'b00111110; // 1625 :  62 - 0x3e
      11'h65A: dout  = 8'b01111100; // 1626 : 124 - 0x7c
      11'h65B: dout  = 8'b11111000; // 1627 : 248 - 0xf8
      11'h65C: dout  = 8'b11111000; // 1628 : 248 - 0xf8
      11'h65D: dout  = 8'b00111100; // 1629 :  60 - 0x3c
      11'h65E: dout  = 8'b00011000; // 1630 :  24 - 0x18
      11'h65F: dout  = 8'b11111000; // 1631 : 248 - 0xf8
      11'h660: dout  = 8'b01111111; // 1632 : 127 - 0x7f -- Sprite 0xcc
      11'h661: dout  = 8'b01111111; // 1633 : 127 - 0x7f
      11'h662: dout  = 8'b01111000; // 1634 : 120 - 0x78
      11'h663: dout  = 8'b00000001; // 1635 :   1 - 0x1
      11'h664: dout  = 8'b00000111; // 1636 :   7 - 0x7
      11'h665: dout  = 8'b00010011; // 1637 :  19 - 0x13
      11'h666: dout  = 8'b11110001; // 1638 : 241 - 0xf1
      11'h667: dout  = 8'b00000011; // 1639 :   3 - 0x3
      11'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0 -- Sprite 0xcd
      11'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      11'h66A: dout  = 8'b00011100; // 1642 :  28 - 0x1c
      11'h66B: dout  = 8'b00011101; // 1643 :  29 - 0x1d
      11'h66C: dout  = 8'b00011011; // 1644 :  27 - 0x1b
      11'h66D: dout  = 8'b11000011; // 1645 : 195 - 0xc3
      11'h66E: dout  = 8'b11100011; // 1646 : 227 - 0xe3
      11'h66F: dout  = 8'b11100001; // 1647 : 225 - 0xe1
      11'h670: dout  = 8'b11100000; // 1648 : 224 - 0xe0 -- Sprite 0xce
      11'h671: dout  = 8'b11001101; // 1649 : 205 - 0xcd
      11'h672: dout  = 8'b00011101; // 1650 :  29 - 0x1d
      11'h673: dout  = 8'b01001111; // 1651 :  79 - 0x4f
      11'h674: dout  = 8'b11101110; // 1652 : 238 - 0xee
      11'h675: dout  = 8'b11111111; // 1653 : 255 - 0xff
      11'h676: dout  = 8'b00111111; // 1654 :  63 - 0x3f
      11'h677: dout  = 8'b00111111; // 1655 :  63 - 0x3f
      11'h678: dout  = 8'b00111111; // 1656 :  63 - 0x3f -- Sprite 0xcf
      11'h679: dout  = 8'b00111111; // 1657 :  63 - 0x3f
      11'h67A: dout  = 8'b00000000; // 1658 :   0 - 0x0
      11'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      11'h67C: dout  = 8'b01110000; // 1660 : 112 - 0x70
      11'h67D: dout  = 8'b10111000; // 1661 : 184 - 0xb8
      11'h67E: dout  = 8'b11111100; // 1662 : 252 - 0xfc
      11'h67F: dout  = 8'b11111100; // 1663 : 252 - 0xfc
      11'h680: dout  = 8'b00000111; // 1664 :   7 - 0x7 -- Sprite 0xd0
      11'h681: dout  = 8'b00001111; // 1665 :  15 - 0xf
      11'h682: dout  = 8'b00011111; // 1666 :  31 - 0x1f
      11'h683: dout  = 8'b00111111; // 1667 :  63 - 0x3f
      11'h684: dout  = 8'b00111110; // 1668 :  62 - 0x3e
      11'h685: dout  = 8'b01111100; // 1669 : 124 - 0x7c
      11'h686: dout  = 8'b01111000; // 1670 : 120 - 0x78
      11'h687: dout  = 8'b01111000; // 1671 : 120 - 0x78
      11'h688: dout  = 8'b00111111; // 1672 :  63 - 0x3f -- Sprite 0xd1
      11'h689: dout  = 8'b01011100; // 1673 :  92 - 0x5c
      11'h68A: dout  = 8'b00111001; // 1674 :  57 - 0x39
      11'h68B: dout  = 8'b00111011; // 1675 :  59 - 0x3b
      11'h68C: dout  = 8'b10111111; // 1676 : 191 - 0xbf
      11'h68D: dout  = 8'b11111111; // 1677 : 255 - 0xff
      11'h68E: dout  = 8'b11111110; // 1678 : 254 - 0xfe
      11'h68F: dout  = 8'b11111110; // 1679 : 254 - 0xfe
      11'h690: dout  = 8'b11000000; // 1680 : 192 - 0xc0 -- Sprite 0xd2
      11'h691: dout  = 8'b11000000; // 1681 : 192 - 0xc0
      11'h692: dout  = 8'b10000000; // 1682 : 128 - 0x80
      11'h693: dout  = 8'b10000000; // 1683 : 128 - 0x80
      11'h694: dout  = 8'b10000000; // 1684 : 128 - 0x80
      11'h695: dout  = 8'b10000000; // 1685 : 128 - 0x80
      11'h696: dout  = 8'b00000000; // 1686 :   0 - 0x0
      11'h697: dout  = 8'b00000000; // 1687 :   0 - 0x0
      11'h698: dout  = 8'b11111110; // 1688 : 254 - 0xfe -- Sprite 0xd3
      11'h699: dout  = 8'b11111100; // 1689 : 252 - 0xfc
      11'h69A: dout  = 8'b01100001; // 1690 :  97 - 0x61
      11'h69B: dout  = 8'b00001111; // 1691 :  15 - 0xf
      11'h69C: dout  = 8'b01111111; // 1692 : 127 - 0x7f
      11'h69D: dout  = 8'b00111111; // 1693 :  63 - 0x3f
      11'h69E: dout  = 8'b00011111; // 1694 :  31 - 0x1f
      11'h69F: dout  = 8'b00011110; // 1695 :  30 - 0x1e
      11'h6A0: dout  = 8'b11110000; // 1696 : 240 - 0xf0 -- Sprite 0xd4
      11'h6A1: dout  = 8'b01111000; // 1697 : 120 - 0x78
      11'h6A2: dout  = 8'b11100100; // 1698 : 228 - 0xe4
      11'h6A3: dout  = 8'b11001000; // 1699 : 200 - 0xc8
      11'h6A4: dout  = 8'b11001100; // 1700 : 204 - 0xcc
      11'h6A5: dout  = 8'b10111110; // 1701 : 190 - 0xbe
      11'h6A6: dout  = 8'b10111110; // 1702 : 190 - 0xbe
      11'h6A7: dout  = 8'b00111110; // 1703 :  62 - 0x3e
      11'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0 -- Sprite 0xd5
      11'h6A9: dout  = 8'b00000001; // 1705 :   1 - 0x1
      11'h6AA: dout  = 8'b00000000; // 1706 :   0 - 0x0
      11'h6AB: dout  = 8'b00000111; // 1707 :   7 - 0x7
      11'h6AC: dout  = 8'b00000111; // 1708 :   7 - 0x7
      11'h6AD: dout  = 8'b00000111; // 1709 :   7 - 0x7
      11'h6AE: dout  = 8'b00000111; // 1710 :   7 - 0x7
      11'h6AF: dout  = 8'b00011111; // 1711 :  31 - 0x1f
      11'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      11'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      11'h6B2: dout  = 8'b00001111; // 1714 :  15 - 0xf
      11'h6B3: dout  = 8'b00111111; // 1715 :  63 - 0x3f
      11'h6B4: dout  = 8'b00111111; // 1716 :  63 - 0x3f
      11'h6B5: dout  = 8'b00001111; // 1717 :  15 - 0xf
      11'h6B6: dout  = 8'b00000000; // 1718 :   0 - 0x0
      11'h6B7: dout  = 8'b00000000; // 1719 :   0 - 0x0
      11'h6B8: dout  = 8'b01111000; // 1720 : 120 - 0x78 -- Sprite 0xd7
      11'h6B9: dout  = 8'b01111100; // 1721 : 124 - 0x7c
      11'h6BA: dout  = 8'b01111110; // 1722 : 126 - 0x7e
      11'h6BB: dout  = 8'b01111111; // 1723 : 127 - 0x7f
      11'h6BC: dout  = 8'b00111111; // 1724 :  63 - 0x3f
      11'h6BD: dout  = 8'b00111111; // 1725 :  63 - 0x3f
      11'h6BE: dout  = 8'b00011011; // 1726 :  27 - 0x1b
      11'h6BF: dout  = 8'b00001001; // 1727 :   9 - 0x9
      11'h6C0: dout  = 8'b00001100; // 1728 :  12 - 0xc -- Sprite 0xd8
      11'h6C1: dout  = 8'b00000000; // 1729 :   0 - 0x0
      11'h6C2: dout  = 8'b00000000; // 1730 :   0 - 0x0
      11'h6C3: dout  = 8'b00000000; // 1731 :   0 - 0x0
      11'h6C4: dout  = 8'b00000111; // 1732 :   7 - 0x7
      11'h6C5: dout  = 8'b01111111; // 1733 : 127 - 0x7f
      11'h6C6: dout  = 8'b01111100; // 1734 : 124 - 0x7c
      11'h6C7: dout  = 8'b00000000; // 1735 :   0 - 0x0
      11'h6C8: dout  = 8'b00000001; // 1736 :   1 - 0x1 -- Sprite 0xd9
      11'h6C9: dout  = 8'b11100001; // 1737 : 225 - 0xe1
      11'h6CA: dout  = 8'b01110001; // 1738 : 113 - 0x71
      11'h6CB: dout  = 8'b01111001; // 1739 : 121 - 0x79
      11'h6CC: dout  = 8'b00111101; // 1740 :  61 - 0x3d
      11'h6CD: dout  = 8'b00111101; // 1741 :  61 - 0x3d
      11'h6CE: dout  = 8'b00011111; // 1742 :  31 - 0x1f
      11'h6CF: dout  = 8'b00000011; // 1743 :   3 - 0x3
      11'h6D0: dout  = 8'b00111111; // 1744 :  63 - 0x3f -- Sprite 0xda
      11'h6D1: dout  = 8'b00111111; // 1745 :  63 - 0x3f
      11'h6D2: dout  = 8'b00011111; // 1746 :  31 - 0x1f
      11'h6D3: dout  = 8'b00011011; // 1747 :  27 - 0x1b
      11'h6D4: dout  = 8'b00110110; // 1748 :  54 - 0x36
      11'h6D5: dout  = 8'b00110000; // 1749 :  48 - 0x30
      11'h6D6: dout  = 8'b01111111; // 1750 : 127 - 0x7f
      11'h6D7: dout  = 8'b00111111; // 1751 :  63 - 0x3f
      11'h6D8: dout  = 8'b11111000; // 1752 : 248 - 0xf8 -- Sprite 0xdb
      11'h6D9: dout  = 8'b11111000; // 1753 : 248 - 0xf8
      11'h6DA: dout  = 8'b11111000; // 1754 : 248 - 0xf8
      11'h6DB: dout  = 8'b10111000; // 1755 : 184 - 0xb8
      11'h6DC: dout  = 8'b00011000; // 1756 :  24 - 0x18
      11'h6DD: dout  = 8'b11011000; // 1757 : 216 - 0xd8
      11'h6DE: dout  = 8'b11011000; // 1758 : 216 - 0xd8
      11'h6DF: dout  = 8'b10111000; // 1759 : 184 - 0xb8
      11'h6E0: dout  = 8'b00000001; // 1760 :   1 - 0x1 -- Sprite 0xdc
      11'h6E1: dout  = 8'b00000010; // 1761 :   2 - 0x2
      11'h6E2: dout  = 8'b00000100; // 1762 :   4 - 0x4
      11'h6E3: dout  = 8'b00000100; // 1763 :   4 - 0x4
      11'h6E4: dout  = 8'b00001000; // 1764 :   8 - 0x8
      11'h6E5: dout  = 8'b00001000; // 1765 :   8 - 0x8
      11'h6E6: dout  = 8'b00010000; // 1766 :  16 - 0x10
      11'h6E7: dout  = 8'b00010000; // 1767 :  16 - 0x10
      11'h6E8: dout  = 8'b00000000; // 1768 :   0 - 0x0 -- Sprite 0xdd
      11'h6E9: dout  = 8'b00001111; // 1769 :  15 - 0xf
      11'h6EA: dout  = 8'b00010011; // 1770 :  19 - 0x13
      11'h6EB: dout  = 8'b00001101; // 1771 :  13 - 0xd
      11'h6EC: dout  = 8'b00001101; // 1772 :  13 - 0xd
      11'h6ED: dout  = 8'b00010011; // 1773 :  19 - 0x13
      11'h6EE: dout  = 8'b00001100; // 1774 :  12 - 0xc
      11'h6EF: dout  = 8'b00100000; // 1775 :  32 - 0x20
      11'h6F0: dout  = 8'b00000000; // 1776 :   0 - 0x0 -- Sprite 0xde
      11'h6F1: dout  = 8'b00100100; // 1777 :  36 - 0x24
      11'h6F2: dout  = 8'b00000000; // 1778 :   0 - 0x0
      11'h6F3: dout  = 8'b00100100; // 1779 :  36 - 0x24
      11'h6F4: dout  = 8'b00000000; // 1780 :   0 - 0x0
      11'h6F5: dout  = 8'b00000100; // 1781 :   4 - 0x4
      11'h6F6: dout  = 8'b00000000; // 1782 :   0 - 0x0
      11'h6F7: dout  = 8'b00000000; // 1783 :   0 - 0x0
      11'h6F8: dout  = 8'b00001111; // 1784 :  15 - 0xf -- Sprite 0xdf
      11'h6F9: dout  = 8'b01000001; // 1785 :  65 - 0x41
      11'h6FA: dout  = 8'b00000000; // 1786 :   0 - 0x0
      11'h6FB: dout  = 8'b10001000; // 1787 : 136 - 0x88
      11'h6FC: dout  = 8'b00000000; // 1788 :   0 - 0x0
      11'h6FD: dout  = 8'b01000100; // 1789 :  68 - 0x44
      11'h6FE: dout  = 8'b00000000; // 1790 :   0 - 0x0
      11'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      11'h700: dout  = 8'b00111000; // 1792 :  56 - 0x38 -- Sprite 0xe0
      11'h701: dout  = 8'b01111100; // 1793 : 124 - 0x7c
      11'h702: dout  = 8'b11111110; // 1794 : 254 - 0xfe
      11'h703: dout  = 8'b11111110; // 1795 : 254 - 0xfe
      11'h704: dout  = 8'b00111011; // 1796 :  59 - 0x3b
      11'h705: dout  = 8'b00000011; // 1797 :   3 - 0x3
      11'h706: dout  = 8'b00000011; // 1798 :   3 - 0x3
      11'h707: dout  = 8'b00000011; // 1799 :   3 - 0x3
      11'h708: dout  = 8'b00000011; // 1800 :   3 - 0x3 -- Sprite 0xe1
      11'h709: dout  = 8'b00110011; // 1801 :  51 - 0x33
      11'h70A: dout  = 8'b01111011; // 1802 : 123 - 0x7b
      11'h70B: dout  = 8'b01111111; // 1803 : 127 - 0x7f
      11'h70C: dout  = 8'b11111111; // 1804 : 255 - 0xff
      11'h70D: dout  = 8'b11111011; // 1805 : 251 - 0xfb
      11'h70E: dout  = 8'b00000011; // 1806 :   3 - 0x3
      11'h70F: dout  = 8'b00000011; // 1807 :   3 - 0x3
      11'h710: dout  = 8'b11011100; // 1808 : 220 - 0xdc -- Sprite 0xe2
      11'h711: dout  = 8'b11000000; // 1809 : 192 - 0xc0
      11'h712: dout  = 8'b11100000; // 1810 : 224 - 0xe0
      11'h713: dout  = 8'b11100000; // 1811 : 224 - 0xe0
      11'h714: dout  = 8'b11100000; // 1812 : 224 - 0xe0
      11'h715: dout  = 8'b11100000; // 1813 : 224 - 0xe0
      11'h716: dout  = 8'b11100000; // 1814 : 224 - 0xe0
      11'h717: dout  = 8'b11000000; // 1815 : 192 - 0xc0
      11'h718: dout  = 8'b00111111; // 1816 :  63 - 0x3f -- Sprite 0xe3
      11'h719: dout  = 8'b01011111; // 1817 :  95 - 0x5f
      11'h71A: dout  = 8'b00111111; // 1818 :  63 - 0x3f
      11'h71B: dout  = 8'b00111111; // 1819 :  63 - 0x3f
      11'h71C: dout  = 8'b10111011; // 1820 : 187 - 0xbb
      11'h71D: dout  = 8'b11111000; // 1821 : 248 - 0xf8
      11'h71E: dout  = 8'b11111110; // 1822 : 254 - 0xfe
      11'h71F: dout  = 8'b11111110; // 1823 : 254 - 0xfe
      11'h720: dout  = 8'b00011111; // 1824 :  31 - 0x1f -- Sprite 0xe4
      11'h721: dout  = 8'b00001111; // 1825 :  15 - 0xf
      11'h722: dout  = 8'b00001111; // 1826 :  15 - 0xf
      11'h723: dout  = 8'b00011111; // 1827 :  31 - 0x1f
      11'h724: dout  = 8'b00011111; // 1828 :  31 - 0x1f
      11'h725: dout  = 8'b00011110; // 1829 :  30 - 0x1e
      11'h726: dout  = 8'b00111000; // 1830 :  56 - 0x38
      11'h727: dout  = 8'b00110000; // 1831 :  48 - 0x30
      11'h728: dout  = 8'b00000000; // 1832 :   0 - 0x0 -- Sprite 0xe5
      11'h729: dout  = 8'b00100000; // 1833 :  32 - 0x20
      11'h72A: dout  = 8'b01100000; // 1834 :  96 - 0x60
      11'h72B: dout  = 8'b01100000; // 1835 :  96 - 0x60
      11'h72C: dout  = 8'b01110000; // 1836 : 112 - 0x70
      11'h72D: dout  = 8'b11110000; // 1837 : 240 - 0xf0
      11'h72E: dout  = 8'b11111000; // 1838 : 248 - 0xf8
      11'h72F: dout  = 8'b11111000; // 1839 : 248 - 0xf8
      11'h730: dout  = 8'b11111000; // 1840 : 248 - 0xf8 -- Sprite 0xe6
      11'h731: dout  = 8'b11111100; // 1841 : 252 - 0xfc
      11'h732: dout  = 8'b11111100; // 1842 : 252 - 0xfc
      11'h733: dout  = 8'b01111110; // 1843 : 126 - 0x7e
      11'h734: dout  = 8'b01111110; // 1844 : 126 - 0x7e
      11'h735: dout  = 8'b00111110; // 1845 :  62 - 0x3e
      11'h736: dout  = 8'b00011111; // 1846 :  31 - 0x1f
      11'h737: dout  = 8'b00000111; // 1847 :   7 - 0x7
      11'h738: dout  = 8'b00000000; // 1848 :   0 - 0x0 -- Sprite 0xe7
      11'h739: dout  = 8'b11000000; // 1849 : 192 - 0xc0
      11'h73A: dout  = 8'b01110000; // 1850 : 112 - 0x70
      11'h73B: dout  = 8'b10111000; // 1851 : 184 - 0xb8
      11'h73C: dout  = 8'b11110100; // 1852 : 244 - 0xf4
      11'h73D: dout  = 8'b11110010; // 1853 : 242 - 0xf2
      11'h73E: dout  = 8'b11110101; // 1854 : 245 - 0xf5
      11'h73F: dout  = 8'b01111011; // 1855 : 123 - 0x7b
      11'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0xe8
      11'h741: dout  = 8'b11011111; // 1857 : 223 - 0xdf
      11'h742: dout  = 8'b00010000; // 1858 :  16 - 0x10
      11'h743: dout  = 8'b11111111; // 1859 : 255 - 0xff
      11'h744: dout  = 8'b11011111; // 1860 : 223 - 0xdf
      11'h745: dout  = 8'b11111111; // 1861 : 255 - 0xff
      11'h746: dout  = 8'b11111111; // 1862 : 255 - 0xff
      11'h747: dout  = 8'b11111001; // 1863 : 249 - 0xf9
      11'h748: dout  = 8'b00011111; // 1864 :  31 - 0x1f -- Sprite 0xe9
      11'h749: dout  = 8'b00011111; // 1865 :  31 - 0x1f
      11'h74A: dout  = 8'b00111110; // 1866 :  62 - 0x3e
      11'h74B: dout  = 8'b11111100; // 1867 : 252 - 0xfc
      11'h74C: dout  = 8'b11111000; // 1868 : 248 - 0xf8
      11'h74D: dout  = 8'b11110000; // 1869 : 240 - 0xf0
      11'h74E: dout  = 8'b11000000; // 1870 : 192 - 0xc0
      11'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      11'h750: dout  = 8'b11111000; // 1872 : 248 - 0xf8 -- Sprite 0xea
      11'h751: dout  = 8'b11111100; // 1873 : 252 - 0xfc
      11'h752: dout  = 8'b11111110; // 1874 : 254 - 0xfe
      11'h753: dout  = 8'b11111111; // 1875 : 255 - 0xff
      11'h754: dout  = 8'b11111111; // 1876 : 255 - 0xff
      11'h755: dout  = 8'b11011111; // 1877 : 223 - 0xdf
      11'h756: dout  = 8'b11011111; // 1878 : 223 - 0xdf
      11'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      11'h758: dout  = 8'b11000001; // 1880 : 193 - 0xc1 -- Sprite 0xeb
      11'h759: dout  = 8'b11110001; // 1881 : 241 - 0xf1
      11'h75A: dout  = 8'b01111001; // 1882 : 121 - 0x79
      11'h75B: dout  = 8'b01111101; // 1883 : 125 - 0x7d
      11'h75C: dout  = 8'b00111101; // 1884 :  61 - 0x3d
      11'h75D: dout  = 8'b00111111; // 1885 :  63 - 0x3f
      11'h75E: dout  = 8'b00011111; // 1886 :  31 - 0x1f
      11'h75F: dout  = 8'b00000011; // 1887 :   3 - 0x3
      11'h760: dout  = 8'b00000010; // 1888 :   2 - 0x2 -- Sprite 0xec
      11'h761: dout  = 8'b00000110; // 1889 :   6 - 0x6
      11'h762: dout  = 8'b00001110; // 1890 :  14 - 0xe
      11'h763: dout  = 8'b00001110; // 1891 :  14 - 0xe
      11'h764: dout  = 8'b00011110; // 1892 :  30 - 0x1e
      11'h765: dout  = 8'b00011110; // 1893 :  30 - 0x1e
      11'h766: dout  = 8'b00111110; // 1894 :  62 - 0x3e
      11'h767: dout  = 8'b00111110; // 1895 :  62 - 0x3e
      11'h768: dout  = 8'b00111110; // 1896 :  62 - 0x3e -- Sprite 0xed
      11'h769: dout  = 8'b00111110; // 1897 :  62 - 0x3e
      11'h76A: dout  = 8'b00111110; // 1898 :  62 - 0x3e
      11'h76B: dout  = 8'b00111110; // 1899 :  62 - 0x3e
      11'h76C: dout  = 8'b00011110; // 1900 :  30 - 0x1e
      11'h76D: dout  = 8'b00011110; // 1901 :  30 - 0x1e
      11'h76E: dout  = 8'b00001110; // 1902 :  14 - 0xe
      11'h76F: dout  = 8'b00000010; // 1903 :   2 - 0x2
      11'h770: dout  = 8'b11000001; // 1904 : 193 - 0xc1 -- Sprite 0xee
      11'h771: dout  = 8'b11110001; // 1905 : 241 - 0xf1
      11'h772: dout  = 8'b01111001; // 1906 : 121 - 0x79
      11'h773: dout  = 8'b01111101; // 1907 : 125 - 0x7d
      11'h774: dout  = 8'b00111101; // 1908 :  61 - 0x3d
      11'h775: dout  = 8'b00111111; // 1909 :  63 - 0x3f
      11'h776: dout  = 8'b00011111; // 1910 :  31 - 0x1f
      11'h777: dout  = 8'b00000011; // 1911 :   3 - 0x3
      11'h778: dout  = 8'b01111100; // 1912 : 124 - 0x7c -- Sprite 0xef
      11'h779: dout  = 8'b00000000; // 1913 :   0 - 0x0
      11'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      11'h77B: dout  = 8'b11111111; // 1915 : 255 - 0xff
      11'h77C: dout  = 8'b11000011; // 1916 : 195 - 0xc3
      11'h77D: dout  = 8'b01111111; // 1917 : 127 - 0x7f
      11'h77E: dout  = 8'b00011111; // 1918 :  31 - 0x1f
      11'h77F: dout  = 8'b00000011; // 1919 :   3 - 0x3
      11'h780: dout  = 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0xf0
      11'h781: dout  = 8'b11111111; // 1921 : 255 - 0xff
      11'h782: dout  = 8'b01111100; // 1922 : 124 - 0x7c
      11'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      11'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      11'h785: dout  = 8'b01111100; // 1925 : 124 - 0x7c
      11'h786: dout  = 8'b11111111; // 1926 : 255 - 0xff
      11'h787: dout  = 8'b11111111; // 1927 : 255 - 0xff
      11'h788: dout  = 8'b11111111; // 1928 : 255 - 0xff -- Sprite 0xf1
      11'h789: dout  = 8'b11111111; // 1929 : 255 - 0xff
      11'h78A: dout  = 8'b00000000; // 1930 :   0 - 0x0
      11'h78B: dout  = 8'b00000100; // 1931 :   4 - 0x4
      11'h78C: dout  = 8'b00001100; // 1932 :  12 - 0xc
      11'h78D: dout  = 8'b00011000; // 1933 :  24 - 0x18
      11'h78E: dout  = 8'b00110000; // 1934 :  48 - 0x30
      11'h78F: dout  = 8'b00000000; // 1935 :   0 - 0x0
      11'h790: dout  = 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0xf2
      11'h791: dout  = 8'b11111111; // 1937 : 255 - 0xff
      11'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      11'h793: dout  = 8'b00000100; // 1939 :   4 - 0x4
      11'h794: dout  = 8'b00000100; // 1940 :   4 - 0x4
      11'h795: dout  = 8'b00000100; // 1941 :   4 - 0x4
      11'h796: dout  = 8'b00001000; // 1942 :   8 - 0x8
      11'h797: dout  = 8'b00001000; // 1943 :   8 - 0x8
      11'h798: dout  = 8'b00001000; // 1944 :   8 - 0x8 -- Sprite 0xf3
      11'h799: dout  = 8'b00010000; // 1945 :  16 - 0x10
      11'h79A: dout  = 8'b00010000; // 1946 :  16 - 0x10
      11'h79B: dout  = 8'b00000000; // 1947 :   0 - 0x0
      11'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      11'h79D: dout  = 8'b00010000; // 1949 :  16 - 0x10
      11'h79E: dout  = 8'b00010000; // 1950 :  16 - 0x10
      11'h79F: dout  = 8'b00001000; // 1951 :   8 - 0x8
      11'h7A0: dout  = 8'b01111111; // 1952 : 127 - 0x7f -- Sprite 0xf4
      11'h7A1: dout  = 8'b00111111; // 1953 :  63 - 0x3f
      11'h7A2: dout  = 8'b00111111; // 1954 :  63 - 0x3f
      11'h7A3: dout  = 8'b00111110; // 1955 :  62 - 0x3e
      11'h7A4: dout  = 8'b00011111; // 1956 :  31 - 0x1f
      11'h7A5: dout  = 8'b00001111; // 1957 :  15 - 0xf
      11'h7A6: dout  = 8'b00000011; // 1958 :   3 - 0x3
      11'h7A7: dout  = 8'b00000000; // 1959 :   0 - 0x0
      11'h7A8: dout  = 8'b00000011; // 1960 :   3 - 0x3 -- Sprite 0xf5
      11'h7A9: dout  = 8'b00001111; // 1961 :  15 - 0xf
      11'h7AA: dout  = 8'b11111111; // 1962 : 255 - 0xff
      11'h7AB: dout  = 8'b01111111; // 1963 : 127 - 0x7f
      11'h7AC: dout  = 8'b01111111; // 1964 : 127 - 0x7f
      11'h7AD: dout  = 8'b01111111; // 1965 : 127 - 0x7f
      11'h7AE: dout  = 8'b01111111; // 1966 : 127 - 0x7f
      11'h7AF: dout  = 8'b01111111; // 1967 : 127 - 0x7f
      11'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      11'h7B1: dout  = 8'b00000000; // 1969 :   0 - 0x0
      11'h7B2: dout  = 8'b00000000; // 1970 :   0 - 0x0
      11'h7B3: dout  = 8'b00000000; // 1971 :   0 - 0x0
      11'h7B4: dout  = 8'b00000000; // 1972 :   0 - 0x0
      11'h7B5: dout  = 8'b00000000; // 1973 :   0 - 0x0
      11'h7B6: dout  = 8'b00000000; // 1974 :   0 - 0x0
      11'h7B7: dout  = 8'b00000000; // 1975 :   0 - 0x0
      11'h7B8: dout  = 8'b00000000; // 1976 :   0 - 0x0 -- Sprite 0xf7
      11'h7B9: dout  = 8'b00000000; // 1977 :   0 - 0x0
      11'h7BA: dout  = 8'b00000000; // 1978 :   0 - 0x0
      11'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      11'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      11'h7BD: dout  = 8'b00000000; // 1981 :   0 - 0x0
      11'h7BE: dout  = 8'b00000000; // 1982 :   0 - 0x0
      11'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      11'h7C0: dout  = 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0xf8
      11'h7C1: dout  = 8'b00000000; // 1985 :   0 - 0x0
      11'h7C2: dout  = 8'b00000000; // 1986 :   0 - 0x0
      11'h7C3: dout  = 8'b00000000; // 1987 :   0 - 0x0
      11'h7C4: dout  = 8'b00000000; // 1988 :   0 - 0x0
      11'h7C5: dout  = 8'b00000000; // 1989 :   0 - 0x0
      11'h7C6: dout  = 8'b00000000; // 1990 :   0 - 0x0
      11'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0 -- Sprite 0xf9
      11'h7C9: dout  = 8'b00000000; // 1993 :   0 - 0x0
      11'h7CA: dout  = 8'b00000000; // 1994 :   0 - 0x0
      11'h7CB: dout  = 8'b00000000; // 1995 :   0 - 0x0
      11'h7CC: dout  = 8'b00000000; // 1996 :   0 - 0x0
      11'h7CD: dout  = 8'b00000000; // 1997 :   0 - 0x0
      11'h7CE: dout  = 8'b00000000; // 1998 :   0 - 0x0
      11'h7CF: dout  = 8'b00000000; // 1999 :   0 - 0x0
      11'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0xfa
      11'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      11'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      11'h7D3: dout  = 8'b00000000; // 2003 :   0 - 0x0
      11'h7D4: dout  = 8'b00000000; // 2004 :   0 - 0x0
      11'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout  = 8'b00000000; // 2006 :   0 - 0x0
      11'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0 -- Sprite 0xfb
      11'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      11'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      11'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      11'h7DC: dout  = 8'b00000000; // 2012 :   0 - 0x0
      11'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      11'h7DE: dout  = 8'b00000000; // 2014 :   0 - 0x0
      11'h7DF: dout  = 8'b00000000; // 2015 :   0 - 0x0
      11'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      11'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      11'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      11'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      11'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      11'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      11'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      11'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      11'h7E8: dout  = 8'b00000000; // 2024 :   0 - 0x0 -- Sprite 0xfd
      11'h7E9: dout  = 8'b00000000; // 2025 :   0 - 0x0
      11'h7EA: dout  = 8'b00000000; // 2026 :   0 - 0x0
      11'h7EB: dout  = 8'b00000000; // 2027 :   0 - 0x0
      11'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      11'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      11'h7EE: dout  = 8'b00000000; // 2030 :   0 - 0x0
      11'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0xfe
      11'h7F1: dout  = 8'b00000000; // 2033 :   0 - 0x0
      11'h7F2: dout  = 8'b00000000; // 2034 :   0 - 0x0
      11'h7F3: dout  = 8'b00000000; // 2035 :   0 - 0x0
      11'h7F4: dout  = 8'b00000000; // 2036 :   0 - 0x0
      11'h7F5: dout  = 8'b00000000; // 2037 :   0 - 0x0
      11'h7F6: dout  = 8'b00000000; // 2038 :   0 - 0x0
      11'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      11'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      11'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      11'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      11'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      11'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      11'h7FD: dout  = 8'b01111100; // 2045 : 124 - 0x7c
      11'h7FE: dout  = 8'b00111000; // 2046 :  56 - 0x38
      11'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
    endcase
  end

endmodule
