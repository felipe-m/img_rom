--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: sprilo_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_SPRILO is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(13-1 downto 0);  --8192 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_SPRILO;

architecture BEHAVIORAL of ROM_PTABLE_SPRILO is
  signal addr_int  : natural range 0 to 2**13-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Pattern Table 0---------
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Sprite 0x1
    "00000000", --   17 - 0x11  :    0 - 0x0
    "00000000", --   18 - 0x12  :    0 - 0x0
    "00000000", --   19 - 0x13  :    0 - 0x0
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00000000", --   21 - 0x15  :    0 - 0x0
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Sprite 0x2
    "00000000", --   33 - 0x21  :    0 - 0x0
    "00000000", --   34 - 0x22  :    0 - 0x0
    "00000000", --   35 - 0x23  :    0 - 0x0
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Sprite 0x3
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00000000", --   51 - 0x33  :    0 - 0x0
    "00000000", --   52 - 0x34  :    0 - 0x0
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000000", --   54 - 0x36  :    0 - 0x0
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Sprite 0x4
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Sprite 0x5
    "00000000", --   81 - 0x51  :    0 - 0x0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00000000", --   88 - 0x58  :    0 - 0x0
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Sprite 0x6
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Sprite 0x7
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x8
    "01111110", --  129 - 0x81  :  126 - 0x7e
    "01111110", --  130 - 0x82  :  126 - 0x7e
    "00111100", --  131 - 0x83  :   60 - 0x3c
    "00111100", --  132 - 0x84  :   60 - 0x3c
    "01111110", --  133 - 0x85  :  126 - 0x7e
    "01011010", --  134 - 0x86  :   90 - 0x5a
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0
    "01000010", --  137 - 0x89  :   66 - 0x42
    "01000010", --  138 - 0x8a  :   66 - 0x42
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "01000010", --  141 - 0x8d  :   66 - 0x42
    "01100110", --  142 - 0x8e  :  102 - 0x66
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Sprite 0x9
    "01100110", --  145 - 0x91  :  102 - 0x66
    "01111100", --  146 - 0x92  :  124 - 0x7c
    "01111110", --  147 - 0x93  :  126 - 0x7e
    "01111110", --  148 - 0x94  :  126 - 0x7e
    "01111100", --  149 - 0x95  :  124 - 0x7c
    "01100110", --  150 - 0x96  :  102 - 0x66
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0
    "01100110", --  153 - 0x99  :  102 - 0x66
    "00000010", --  154 - 0x9a  :    2 - 0x2
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "00000010", --  157 - 0x9d  :    2 - 0x2
    "01100110", --  158 - 0x9e  :  102 - 0x66
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00010000", --  160 - 0xa0  :   16 - 0x10 -- Sprite 0xa
    "00011000", --  161 - 0xa1  :   24 - 0x18
    "00111000", --  162 - 0xa2  :   56 - 0x38
    "11111110", --  163 - 0xa3  :  254 - 0xfe
    "01111101", --  164 - 0xa4  :  125 - 0x7d
    "00011100", --  165 - 0xa5  :   28 - 0x1c
    "00010000", --  166 - 0xa6  :   16 - 0x10
    "00001000", --  167 - 0xa7  :    8 - 0x8
    "00010000", --  168 - 0xa8  :   16 - 0x10
    "00001000", --  169 - 0xa9  :    8 - 0x8
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "10000010", --  171 - 0xab  :  130 - 0x82
    "01000011", --  172 - 0xac  :   67 - 0x43
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00011000", --  174 - 0xae  :   24 - 0x18
    "00001000", --  175 - 0xaf  :    8 - 0x8
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0xb
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0xc
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "00000000", --  194 - 0xc2  :    0 - 0x0
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00000000", --  196 - 0xc4  :    0 - 0x0
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Sprite 0xd
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00000000", --  211 - 0xd3  :    0 - 0x0
    "00000000", --  212 - 0xd4  :    0 - 0x0
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Sprite 0xe
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00000000", --  228 - 0xe4  :    0 - 0x0
    "00000000", --  229 - 0xe5  :    0 - 0x0
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Sprite 0xf
    "00000000", --  241 - 0xf1  :    0 - 0x0
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "00000000", --  243 - 0xf3  :    0 - 0x0
    "00000000", --  244 - 0xf4  :    0 - 0x0
    "00000000", --  245 - 0xf5  :    0 - 0x0
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x10
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00000000", --  272 - 0x110  :    0 - 0x0 -- Sprite 0x11
    "00000000", --  273 - 0x111  :    0 - 0x0
    "00000000", --  274 - 0x112  :    0 - 0x0
    "00000000", --  275 - 0x113  :    0 - 0x0
    "00000000", --  276 - 0x114  :    0 - 0x0
    "00000000", --  277 - 0x115  :    0 - 0x0
    "00000000", --  278 - 0x116  :    0 - 0x0
    "00000000", --  279 - 0x117  :    0 - 0x0
    "00000000", --  280 - 0x118  :    0 - 0x0
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00000000", --  283 - 0x11b  :    0 - 0x0
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Sprite 0x12
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000000", --  298 - 0x12a  :    0 - 0x0
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x13
    "00000000", --  305 - 0x131  :    0 - 0x0
    "00000000", --  306 - 0x132  :    0 - 0x0
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "00000000", --  309 - 0x135  :    0 - 0x0
    "00000000", --  310 - 0x136  :    0 - 0x0
    "00000000", --  311 - 0x137  :    0 - 0x0
    "00000000", --  312 - 0x138  :    0 - 0x0
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Sprite 0x14
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "00000000", --  324 - 0x144  :    0 - 0x0
    "00000000", --  325 - 0x145  :    0 - 0x0
    "00000000", --  326 - 0x146  :    0 - 0x0
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00000000", --  328 - 0x148  :    0 - 0x0
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000000", --  330 - 0x14a  :    0 - 0x0
    "00000000", --  331 - 0x14b  :    0 - 0x0
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00000000", --  336 - 0x150  :    0 - 0x0 -- Sprite 0x15
    "00000000", --  337 - 0x151  :    0 - 0x0
    "00000000", --  338 - 0x152  :    0 - 0x0
    "00000000", --  339 - 0x153  :    0 - 0x0
    "00000000", --  340 - 0x154  :    0 - 0x0
    "00000000", --  341 - 0x155  :    0 - 0x0
    "00000000", --  342 - 0x156  :    0 - 0x0
    "00000000", --  343 - 0x157  :    0 - 0x0
    "00000000", --  344 - 0x158  :    0 - 0x0
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x16
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Sprite 0x17
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000000", --  376 - 0x178  :    0 - 0x0
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00000000", --  379 - 0x17b  :    0 - 0x0
    "00000000", --  380 - 0x17c  :    0 - 0x0
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000000", --  384 - 0x180  :    0 - 0x0 -- Sprite 0x18
    "00000000", --  385 - 0x181  :    0 - 0x0
    "00000000", --  386 - 0x182  :    0 - 0x0
    "00000000", --  387 - 0x183  :    0 - 0x0
    "00000000", --  388 - 0x184  :    0 - 0x0
    "00000000", --  389 - 0x185  :    0 - 0x0
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Sprite 0x19
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000000", --  403 - 0x193  :    0 - 0x0
    "00000000", --  404 - 0x194  :    0 - 0x0
    "00000000", --  405 - 0x195  :    0 - 0x0
    "00000000", --  406 - 0x196  :    0 - 0x0
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00000000", --  408 - 0x198  :    0 - 0x0
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "00000000", --  411 - 0x19b  :    0 - 0x0
    "00000000", --  412 - 0x19c  :    0 - 0x0
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- Sprite 0x1a
    "00000000", --  417 - 0x1a1  :    0 - 0x0
    "00000000", --  418 - 0x1a2  :    0 - 0x0
    "00000000", --  419 - 0x1a3  :    0 - 0x0
    "00000000", --  420 - 0x1a4  :    0 - 0x0
    "00000000", --  421 - 0x1a5  :    0 - 0x0
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "00000000", --  424 - 0x1a8  :    0 - 0x0
    "00000000", --  425 - 0x1a9  :    0 - 0x0
    "00000000", --  426 - 0x1aa  :    0 - 0x0
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x1b
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00000000", --  434 - 0x1b2  :    0 - 0x0
    "00000000", --  435 - 0x1b3  :    0 - 0x0
    "00000000", --  436 - 0x1b4  :    0 - 0x0
    "00000000", --  437 - 0x1b5  :    0 - 0x0
    "00000000", --  438 - 0x1b6  :    0 - 0x0
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "00000000", --  440 - 0x1b8  :    0 - 0x0
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Sprite 0x1c
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "00000000", --  453 - 0x1c5  :    0 - 0x0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x1d
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "00000000", --  467 - 0x1d3  :    0 - 0x0
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "00000000", --  469 - 0x1d5  :    0 - 0x0
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x1e
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "00000000", --  485 - 0x1e5  :    0 - 0x0
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Sprite 0x1f
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00000000", --  500 - 0x1f4  :    0 - 0x0
    "00000000", --  501 - 0x1f5  :    0 - 0x0
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "00000000", --  504 - 0x1f8  :    0 - 0x0
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Sprite 0x20
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Sprite 0x21
    "00000000", --  529 - 0x211  :    0 - 0x0
    "00000000", --  530 - 0x212  :    0 - 0x0
    "00000000", --  531 - 0x213  :    0 - 0x0
    "00000000", --  532 - 0x214  :    0 - 0x0
    "00000000", --  533 - 0x215  :    0 - 0x0
    "00000000", --  534 - 0x216  :    0 - 0x0
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00000000", --  536 - 0x218  :    0 - 0x0
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Sprite 0x22
    "00000000", --  545 - 0x221  :    0 - 0x0
    "00000000", --  546 - 0x222  :    0 - 0x0
    "00000000", --  547 - 0x223  :    0 - 0x0
    "00000000", --  548 - 0x224  :    0 - 0x0
    "00000000", --  549 - 0x225  :    0 - 0x0
    "00000000", --  550 - 0x226  :    0 - 0x0
    "00000000", --  551 - 0x227  :    0 - 0x0
    "00000000", --  552 - 0x228  :    0 - 0x0
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000000", --  560 - 0x230  :    0 - 0x0 -- Sprite 0x23
    "00000000", --  561 - 0x231  :    0 - 0x0
    "00000000", --  562 - 0x232  :    0 - 0x0
    "00000000", --  563 - 0x233  :    0 - 0x0
    "00000000", --  564 - 0x234  :    0 - 0x0
    "00000000", --  565 - 0x235  :    0 - 0x0
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00000000", --  568 - 0x238  :    0 - 0x0
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Sprite 0x24
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00000000", --  584 - 0x248  :    0 - 0x0
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000000", --  592 - 0x250  :    0 - 0x0 -- Sprite 0x25
    "00000000", --  593 - 0x251  :    0 - 0x0
    "00000000", --  594 - 0x252  :    0 - 0x0
    "00000000", --  595 - 0x253  :    0 - 0x0
    "00000000", --  596 - 0x254  :    0 - 0x0
    "00000000", --  597 - 0x255  :    0 - 0x0
    "00000000", --  598 - 0x256  :    0 - 0x0
    "00000000", --  599 - 0x257  :    0 - 0x0
    "00000000", --  600 - 0x258  :    0 - 0x0
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Sprite 0x26
    "00000000", --  609 - 0x261  :    0 - 0x0
    "00000000", --  610 - 0x262  :    0 - 0x0
    "00000000", --  611 - 0x263  :    0 - 0x0
    "00000000", --  612 - 0x264  :    0 - 0x0
    "00000000", --  613 - 0x265  :    0 - 0x0
    "00000000", --  614 - 0x266  :    0 - 0x0
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Sprite 0x27
    "00000000", --  625 - 0x271  :    0 - 0x0
    "00000000", --  626 - 0x272  :    0 - 0x0
    "00000000", --  627 - 0x273  :    0 - 0x0
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000000", --  629 - 0x275  :    0 - 0x0
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0
    "00000000", --  633 - 0x279  :    0 - 0x0
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "00000000", --  635 - 0x27b  :    0 - 0x0
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x28
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Sprite 0x29
    "00000000", --  657 - 0x291  :    0 - 0x0
    "00000000", --  658 - 0x292  :    0 - 0x0
    "00000000", --  659 - 0x293  :    0 - 0x0
    "00000000", --  660 - 0x294  :    0 - 0x0
    "00000000", --  661 - 0x295  :    0 - 0x0
    "00000000", --  662 - 0x296  :    0 - 0x0
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Sprite 0x2a
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "00000000", --  674 - 0x2a2  :    0 - 0x0
    "00000000", --  675 - 0x2a3  :    0 - 0x0
    "00000000", --  676 - 0x2a4  :    0 - 0x0
    "00000000", --  677 - 0x2a5  :    0 - 0x0
    "00000000", --  678 - 0x2a6  :    0 - 0x0
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "00000000", --  680 - 0x2a8  :    0 - 0x0
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "00000000", --  686 - 0x2ae  :    0 - 0x0
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "00000000", --  688 - 0x2b0  :    0 - 0x0 -- Sprite 0x2b
    "00000000", --  689 - 0x2b1  :    0 - 0x0
    "00000000", --  690 - 0x2b2  :    0 - 0x0
    "00000000", --  691 - 0x2b3  :    0 - 0x0
    "00000000", --  692 - 0x2b4  :    0 - 0x0
    "00000000", --  693 - 0x2b5  :    0 - 0x0
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "00000000", --  696 - 0x2b8  :    0 - 0x0
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "00000000", --  707 - 0x2c3  :    0 - 0x0
    "00000000", --  708 - 0x2c4  :    0 - 0x0
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x2d
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x2f
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00000000", --  754 - 0x2f2  :    0 - 0x0
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "00000000", --  756 - 0x2f4  :    0 - 0x0
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "00000000", --  764 - 0x2fc  :    0 - 0x0
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x30
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00000000", --  770 - 0x302  :    0 - 0x0
    "00000000", --  771 - 0x303  :    0 - 0x0
    "00000000", --  772 - 0x304  :    0 - 0x0
    "00000000", --  773 - 0x305  :    0 - 0x0
    "00000000", --  774 - 0x306  :    0 - 0x0
    "00000000", --  775 - 0x307  :    0 - 0x0
    "00000000", --  776 - 0x308  :    0 - 0x0
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000000", --  779 - 0x30b  :    0 - 0x0
    "00000000", --  780 - 0x30c  :    0 - 0x0
    "00000000", --  781 - 0x30d  :    0 - 0x0
    "00000000", --  782 - 0x30e  :    0 - 0x0
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Sprite 0x31
    "00000000", --  785 - 0x311  :    0 - 0x0
    "00000000", --  786 - 0x312  :    0 - 0x0
    "00000000", --  787 - 0x313  :    0 - 0x0
    "00000000", --  788 - 0x314  :    0 - 0x0
    "00000000", --  789 - 0x315  :    0 - 0x0
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Sprite 0x32
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "00000000", --  804 - 0x324  :    0 - 0x0
    "00000000", --  805 - 0x325  :    0 - 0x0
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "00000000", --  813 - 0x32d  :    0 - 0x0
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Sprite 0x33
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000000", --  818 - 0x332  :    0 - 0x0
    "00000000", --  819 - 0x333  :    0 - 0x0
    "00000000", --  820 - 0x334  :    0 - 0x0
    "00000000", --  821 - 0x335  :    0 - 0x0
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000000", --  824 - 0x338  :    0 - 0x0
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x34
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Sprite 0x35
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Sprite 0x36
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "00000000", --  868 - 0x364  :    0 - 0x0
    "00000000", --  869 - 0x365  :    0 - 0x0
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x37
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00000000", --  888 - 0x378  :    0 - 0x0
    "00000000", --  889 - 0x379  :    0 - 0x0
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Sprite 0x38
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Sprite 0x39
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Sprite 0x3b
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Sprite 0x3d
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x3e
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Sprite 0x3f
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Sprite 0x40
    "00000000", -- 1025 - 0x401  :    0 - 0x0
    "00000000", -- 1026 - 0x402  :    0 - 0x0
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00000000", -- 1029 - 0x405  :    0 - 0x0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00000000", -- 1032 - 0x408  :    0 - 0x0
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Sprite 0x41
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "00000000", -- 1045 - 0x415  :    0 - 0x0
    "00000000", -- 1046 - 0x416  :    0 - 0x0
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- Sprite 0x42
    "00000000", -- 1057 - 0x421  :    0 - 0x0
    "00000000", -- 1058 - 0x422  :    0 - 0x0
    "00000000", -- 1059 - 0x423  :    0 - 0x0
    "00000000", -- 1060 - 0x424  :    0 - 0x0
    "00000000", -- 1061 - 0x425  :    0 - 0x0
    "00000000", -- 1062 - 0x426  :    0 - 0x0
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Sprite 0x43
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Sprite 0x44
    "00000000", -- 1089 - 0x441  :    0 - 0x0
    "00000000", -- 1090 - 0x442  :    0 - 0x0
    "00000000", -- 1091 - 0x443  :    0 - 0x0
    "00000000", -- 1092 - 0x444  :    0 - 0x0
    "00000000", -- 1093 - 0x445  :    0 - 0x0
    "00000000", -- 1094 - 0x446  :    0 - 0x0
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00000000", -- 1096 - 0x448  :    0 - 0x0
    "00000000", -- 1097 - 0x449  :    0 - 0x0
    "00000000", -- 1098 - 0x44a  :    0 - 0x0
    "00000000", -- 1099 - 0x44b  :    0 - 0x0
    "00000000", -- 1100 - 0x44c  :    0 - 0x0
    "00000000", -- 1101 - 0x44d  :    0 - 0x0
    "00000000", -- 1102 - 0x44e  :    0 - 0x0
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Sprite 0x45
    "00000000", -- 1105 - 0x451  :    0 - 0x0
    "00000000", -- 1106 - 0x452  :    0 - 0x0
    "00000000", -- 1107 - 0x453  :    0 - 0x0
    "00000000", -- 1108 - 0x454  :    0 - 0x0
    "00000000", -- 1109 - 0x455  :    0 - 0x0
    "00000000", -- 1110 - 0x456  :    0 - 0x0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00000000", -- 1112 - 0x458  :    0 - 0x0
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "00000000", -- 1114 - 0x45a  :    0 - 0x0
    "00000000", -- 1115 - 0x45b  :    0 - 0x0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00000000", -- 1117 - 0x45d  :    0 - 0x0
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Sprite 0x46
    "00000000", -- 1121 - 0x461  :    0 - 0x0
    "00000000", -- 1122 - 0x462  :    0 - 0x0
    "00000000", -- 1123 - 0x463  :    0 - 0x0
    "00000000", -- 1124 - 0x464  :    0 - 0x0
    "00000000", -- 1125 - 0x465  :    0 - 0x0
    "00000000", -- 1126 - 0x466  :    0 - 0x0
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000000", -- 1128 - 0x468  :    0 - 0x0
    "00000000", -- 1129 - 0x469  :    0 - 0x0
    "00000000", -- 1130 - 0x46a  :    0 - 0x0
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0 -- Sprite 0x47
    "00000000", -- 1137 - 0x471  :    0 - 0x0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "00000000", -- 1140 - 0x474  :    0 - 0x0
    "00000000", -- 1141 - 0x475  :    0 - 0x0
    "00000000", -- 1142 - 0x476  :    0 - 0x0
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000000", -- 1144 - 0x478  :    0 - 0x0
    "00000000", -- 1145 - 0x479  :    0 - 0x0
    "00000000", -- 1146 - 0x47a  :    0 - 0x0
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x48
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00000000", -- 1156 - 0x484  :    0 - 0x0
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "00000000", -- 1158 - 0x486  :    0 - 0x0
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0 -- Sprite 0x49
    "00000000", -- 1169 - 0x491  :    0 - 0x0
    "00000000", -- 1170 - 0x492  :    0 - 0x0
    "00000000", -- 1171 - 0x493  :    0 - 0x0
    "00000000", -- 1172 - 0x494  :    0 - 0x0
    "00000000", -- 1173 - 0x495  :    0 - 0x0
    "00000000", -- 1174 - 0x496  :    0 - 0x0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "00000000", -- 1176 - 0x498  :    0 - 0x0
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- Sprite 0x4a
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000000", -- 1186 - 0x4a2  :    0 - 0x0
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00000000", -- 1188 - 0x4a4  :    0 - 0x0
    "00000000", -- 1189 - 0x4a5  :    0 - 0x0
    "00000000", -- 1190 - 0x4a6  :    0 - 0x0
    "00000000", -- 1191 - 0x4a7  :    0 - 0x0
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00000000", -- 1194 - 0x4aa  :    0 - 0x0
    "00000000", -- 1195 - 0x4ab  :    0 - 0x0
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0 -- Sprite 0x4b
    "00000000", -- 1201 - 0x4b1  :    0 - 0x0
    "00000000", -- 1202 - 0x4b2  :    0 - 0x0
    "00000000", -- 1203 - 0x4b3  :    0 - 0x0
    "00000000", -- 1204 - 0x4b4  :    0 - 0x0
    "00000000", -- 1205 - 0x4b5  :    0 - 0x0
    "00000000", -- 1206 - 0x4b6  :    0 - 0x0
    "00000000", -- 1207 - 0x4b7  :    0 - 0x0
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- Sprite 0x4c
    "00000000", -- 1217 - 0x4c1  :    0 - 0x0
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000000", -- 1219 - 0x4c3  :    0 - 0x0
    "00000000", -- 1220 - 0x4c4  :    0 - 0x0
    "00000000", -- 1221 - 0x4c5  :    0 - 0x0
    "00000000", -- 1222 - 0x4c6  :    0 - 0x0
    "00000000", -- 1223 - 0x4c7  :    0 - 0x0
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "00000000", -- 1228 - 0x4cc  :    0 - 0x0
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Sprite 0x4d
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00000000", -- 1235 - 0x4d3  :    0 - 0x0
    "00000000", -- 1236 - 0x4d4  :    0 - 0x0
    "00000000", -- 1237 - 0x4d5  :    0 - 0x0
    "00000000", -- 1238 - 0x4d6  :    0 - 0x0
    "00000000", -- 1239 - 0x4d7  :    0 - 0x0
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0 -- Sprite 0x4e
    "00000000", -- 1249 - 0x4e1  :    0 - 0x0
    "00000000", -- 1250 - 0x4e2  :    0 - 0x0
    "00000000", -- 1251 - 0x4e3  :    0 - 0x0
    "00000000", -- 1252 - 0x4e4  :    0 - 0x0
    "00000000", -- 1253 - 0x4e5  :    0 - 0x0
    "00000000", -- 1254 - 0x4e6  :    0 - 0x0
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0
    "00000000", -- 1257 - 0x4e9  :    0 - 0x0
    "00000000", -- 1258 - 0x4ea  :    0 - 0x0
    "00000000", -- 1259 - 0x4eb  :    0 - 0x0
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00000000", -- 1261 - 0x4ed  :    0 - 0x0
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0 -- Sprite 0x4f
    "00000000", -- 1265 - 0x4f1  :    0 - 0x0
    "00000000", -- 1266 - 0x4f2  :    0 - 0x0
    "00000000", -- 1267 - 0x4f3  :    0 - 0x0
    "00000000", -- 1268 - 0x4f4  :    0 - 0x0
    "00000000", -- 1269 - 0x4f5  :    0 - 0x0
    "00000000", -- 1270 - 0x4f6  :    0 - 0x0
    "00000000", -- 1271 - 0x4f7  :    0 - 0x0
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- Sprite 0x50
    "00000000", -- 1281 - 0x501  :    0 - 0x0
    "00000000", -- 1282 - 0x502  :    0 - 0x0
    "00000000", -- 1283 - 0x503  :    0 - 0x0
    "00000000", -- 1284 - 0x504  :    0 - 0x0
    "00000000", -- 1285 - 0x505  :    0 - 0x0
    "00000000", -- 1286 - 0x506  :    0 - 0x0
    "00000000", -- 1287 - 0x507  :    0 - 0x0
    "00000000", -- 1288 - 0x508  :    0 - 0x0
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00000000", -- 1290 - 0x50a  :    0 - 0x0
    "00000000", -- 1291 - 0x50b  :    0 - 0x0
    "00000000", -- 1292 - 0x50c  :    0 - 0x0
    "00000000", -- 1293 - 0x50d  :    0 - 0x0
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00000000", -- 1296 - 0x510  :    0 - 0x0 -- Sprite 0x51
    "00000000", -- 1297 - 0x511  :    0 - 0x0
    "00000000", -- 1298 - 0x512  :    0 - 0x0
    "00000000", -- 1299 - 0x513  :    0 - 0x0
    "00000000", -- 1300 - 0x514  :    0 - 0x0
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "00000000", -- 1302 - 0x516  :    0 - 0x0
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "00000000", -- 1304 - 0x518  :    0 - 0x0
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "00000000", -- 1306 - 0x51a  :    0 - 0x0
    "00000000", -- 1307 - 0x51b  :    0 - 0x0
    "00000000", -- 1308 - 0x51c  :    0 - 0x0
    "00000000", -- 1309 - 0x51d  :    0 - 0x0
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Sprite 0x52
    "00000000", -- 1313 - 0x521  :    0 - 0x0
    "00000000", -- 1314 - 0x522  :    0 - 0x0
    "00000000", -- 1315 - 0x523  :    0 - 0x0
    "00000000", -- 1316 - 0x524  :    0 - 0x0
    "00000000", -- 1317 - 0x525  :    0 - 0x0
    "00000000", -- 1318 - 0x526  :    0 - 0x0
    "00000000", -- 1319 - 0x527  :    0 - 0x0
    "00000000", -- 1320 - 0x528  :    0 - 0x0
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "00000000", -- 1324 - 0x52c  :    0 - 0x0
    "00000000", -- 1325 - 0x52d  :    0 - 0x0
    "00000000", -- 1326 - 0x52e  :    0 - 0x0
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Sprite 0x53
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "00000000", -- 1331 - 0x533  :    0 - 0x0
    "00000000", -- 1332 - 0x534  :    0 - 0x0
    "00000000", -- 1333 - 0x535  :    0 - 0x0
    "00000000", -- 1334 - 0x536  :    0 - 0x0
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "00000000", -- 1336 - 0x538  :    0 - 0x0
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "00000000", -- 1338 - 0x53a  :    0 - 0x0
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Sprite 0x54
    "00000000", -- 1345 - 0x541  :    0 - 0x0
    "00000000", -- 1346 - 0x542  :    0 - 0x0
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00000000", -- 1349 - 0x545  :    0 - 0x0
    "00000000", -- 1350 - 0x546  :    0 - 0x0
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "00000000", -- 1352 - 0x548  :    0 - 0x0
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "00000000", -- 1354 - 0x54a  :    0 - 0x0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "00000000", -- 1357 - 0x54d  :    0 - 0x0
    "00000000", -- 1358 - 0x54e  :    0 - 0x0
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0x55
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Sprite 0x56
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "00000000", -- 1380 - 0x564  :    0 - 0x0
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "00000000", -- 1386 - 0x56a  :    0 - 0x0
    "00000000", -- 1387 - 0x56b  :    0 - 0x0
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0x57
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000000", -- 1396 - 0x574  :    0 - 0x0
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Sprite 0x58
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "00000000", -- 1410 - 0x582  :    0 - 0x0
    "00000000", -- 1411 - 0x583  :    0 - 0x0
    "00000000", -- 1412 - 0x584  :    0 - 0x0
    "00000000", -- 1413 - 0x585  :    0 - 0x0
    "00000000", -- 1414 - 0x586  :    0 - 0x0
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00000000", -- 1416 - 0x588  :    0 - 0x0
    "00000000", -- 1417 - 0x589  :    0 - 0x0
    "00000000", -- 1418 - 0x58a  :    0 - 0x0
    "00000000", -- 1419 - 0x58b  :    0 - 0x0
    "00000000", -- 1420 - 0x58c  :    0 - 0x0
    "00000000", -- 1421 - 0x58d  :    0 - 0x0
    "00000000", -- 1422 - 0x58e  :    0 - 0x0
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "00000000", -- 1424 - 0x590  :    0 - 0x0 -- Sprite 0x59
    "00000000", -- 1425 - 0x591  :    0 - 0x0
    "00000000", -- 1426 - 0x592  :    0 - 0x0
    "00000000", -- 1427 - 0x593  :    0 - 0x0
    "00000000", -- 1428 - 0x594  :    0 - 0x0
    "00000000", -- 1429 - 0x595  :    0 - 0x0
    "00000000", -- 1430 - 0x596  :    0 - 0x0
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00000000", -- 1432 - 0x598  :    0 - 0x0
    "00000000", -- 1433 - 0x599  :    0 - 0x0
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00000000", -- 1435 - 0x59b  :    0 - 0x0
    "00000000", -- 1436 - 0x59c  :    0 - 0x0
    "00000000", -- 1437 - 0x59d  :    0 - 0x0
    "00000000", -- 1438 - 0x59e  :    0 - 0x0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0 -- Sprite 0x5a
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "00000000", -- 1442 - 0x5a2  :    0 - 0x0
    "00000000", -- 1443 - 0x5a3  :    0 - 0x0
    "00000000", -- 1444 - 0x5a4  :    0 - 0x0
    "00000000", -- 1445 - 0x5a5  :    0 - 0x0
    "00000000", -- 1446 - 0x5a6  :    0 - 0x0
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "00000000", -- 1450 - 0x5aa  :    0 - 0x0
    "00000000", -- 1451 - 0x5ab  :    0 - 0x0
    "00000000", -- 1452 - 0x5ac  :    0 - 0x0
    "00000000", -- 1453 - 0x5ad  :    0 - 0x0
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0x5b
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00000000", -- 1461 - 0x5b5  :    0 - 0x0
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "00000000", -- 1466 - 0x5ba  :    0 - 0x0
    "00000000", -- 1467 - 0x5bb  :    0 - 0x0
    "00000000", -- 1468 - 0x5bc  :    0 - 0x0
    "00000000", -- 1469 - 0x5bd  :    0 - 0x0
    "00000000", -- 1470 - 0x5be  :    0 - 0x0
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Sprite 0x5c
    "00000000", -- 1473 - 0x5c1  :    0 - 0x0
    "00000000", -- 1474 - 0x5c2  :    0 - 0x0
    "00000000", -- 1475 - 0x5c3  :    0 - 0x0
    "00000000", -- 1476 - 0x5c4  :    0 - 0x0
    "00000000", -- 1477 - 0x5c5  :    0 - 0x0
    "00000000", -- 1478 - 0x5c6  :    0 - 0x0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "00000000", -- 1482 - 0x5ca  :    0 - 0x0
    "00000000", -- 1483 - 0x5cb  :    0 - 0x0
    "00000000", -- 1484 - 0x5cc  :    0 - 0x0
    "00000000", -- 1485 - 0x5cd  :    0 - 0x0
    "00000000", -- 1486 - 0x5ce  :    0 - 0x0
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Sprite 0x5d
    "00000000", -- 1489 - 0x5d1  :    0 - 0x0
    "00000000", -- 1490 - 0x5d2  :    0 - 0x0
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "00000000", -- 1492 - 0x5d4  :    0 - 0x0
    "00000000", -- 1493 - 0x5d5  :    0 - 0x0
    "00000000", -- 1494 - 0x5d6  :    0 - 0x0
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Sprite 0x5e
    "00000000", -- 1505 - 0x5e1  :    0 - 0x0
    "00000000", -- 1506 - 0x5e2  :    0 - 0x0
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "00000000", -- 1508 - 0x5e4  :    0 - 0x0
    "00000000", -- 1509 - 0x5e5  :    0 - 0x0
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00000000", -- 1514 - 0x5ea  :    0 - 0x0
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "00000000", -- 1516 - 0x5ec  :    0 - 0x0
    "00000000", -- 1517 - 0x5ed  :    0 - 0x0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Sprite 0x5f
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0x60
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000000", -- 1542 - 0x606  :    0 - 0x0
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00000000", -- 1544 - 0x608  :    0 - 0x0
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0x61
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0x62
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000000", -- 1578 - 0x62a  :    0 - 0x0
    "00000000", -- 1579 - 0x62b  :    0 - 0x0
    "00000000", -- 1580 - 0x62c  :    0 - 0x0
    "00000000", -- 1581 - 0x62d  :    0 - 0x0
    "00000000", -- 1582 - 0x62e  :    0 - 0x0
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "00000000", -- 1584 - 0x630  :    0 - 0x0 -- Sprite 0x63
    "00000000", -- 1585 - 0x631  :    0 - 0x0
    "00000000", -- 1586 - 0x632  :    0 - 0x0
    "00000000", -- 1587 - 0x633  :    0 - 0x0
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "00000000", -- 1589 - 0x635  :    0 - 0x0
    "00000000", -- 1590 - 0x636  :    0 - 0x0
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00000000", -- 1592 - 0x638  :    0 - 0x0
    "00000000", -- 1593 - 0x639  :    0 - 0x0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "00000000", -- 1596 - 0x63c  :    0 - 0x0
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0x64
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00000000", -- 1608 - 0x648  :    0 - 0x0
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0x65
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "00000000", -- 1622 - 0x656  :    0 - 0x0
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Sprite 0x66
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Sprite 0x67
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0x68
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00000000", -- 1680 - 0x690  :    0 - 0x0 -- Sprite 0x69
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00000000", -- 1685 - 0x695  :    0 - 0x0
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00000000", -- 1688 - 0x698  :    0 - 0x0
    "00000000", -- 1689 - 0x699  :    0 - 0x0
    "00000000", -- 1690 - 0x69a  :    0 - 0x0
    "00000000", -- 1691 - 0x69b  :    0 - 0x0
    "00000000", -- 1692 - 0x69c  :    0 - 0x0
    "00000000", -- 1693 - 0x69d  :    0 - 0x0
    "00000000", -- 1694 - 0x69e  :    0 - 0x0
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0x6a
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0
    "00000000", -- 1705 - 0x6a9  :    0 - 0x0
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0x6b
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "00000000", -- 1715 - 0x6b3  :    0 - 0x0
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "00000000", -- 1720 - 0x6b8  :    0 - 0x0
    "00000000", -- 1721 - 0x6b9  :    0 - 0x0
    "00000000", -- 1722 - 0x6ba  :    0 - 0x0
    "00000000", -- 1723 - 0x6bb  :    0 - 0x0
    "00000000", -- 1724 - 0x6bc  :    0 - 0x0
    "00000000", -- 1725 - 0x6bd  :    0 - 0x0
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Sprite 0x6c
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000000", -- 1734 - 0x6c6  :    0 - 0x0
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "00000000", -- 1738 - 0x6ca  :    0 - 0x0
    "00000000", -- 1739 - 0x6cb  :    0 - 0x0
    "00000000", -- 1740 - 0x6cc  :    0 - 0x0
    "00000000", -- 1741 - 0x6cd  :    0 - 0x0
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Sprite 0x6d
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0
    "00000000", -- 1753 - 0x6d9  :    0 - 0x0
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "00000000", -- 1755 - 0x6db  :    0 - 0x0
    "00000000", -- 1756 - 0x6dc  :    0 - 0x0
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Sprite 0x6e
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00000000", -- 1773 - 0x6ed  :    0 - 0x0
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0 -- Sprite 0x6f
    "00000000", -- 1777 - 0x6f1  :    0 - 0x0
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00000000", -- 1779 - 0x6f3  :    0 - 0x0
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "00000000", -- 1781 - 0x6f5  :    0 - 0x0
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "00000000", -- 1784 - 0x6f8  :    0 - 0x0
    "00000000", -- 1785 - 0x6f9  :    0 - 0x0
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "00000000", -- 1787 - 0x6fb  :    0 - 0x0
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "00000000", -- 1789 - 0x6fd  :    0 - 0x0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Sprite 0x70
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0 -- Sprite 0x71
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000000", -- 1816 - 0x718  :    0 - 0x0
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Sprite 0x72
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000000", -- 1828 - 0x724  :    0 - 0x0
    "00000000", -- 1829 - 0x725  :    0 - 0x0
    "00000000", -- 1830 - 0x726  :    0 - 0x0
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "00000000", -- 1840 - 0x730  :    0 - 0x0 -- Sprite 0x73
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "00000000", -- 1845 - 0x735  :    0 - 0x0
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0x74
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Sprite 0x75
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0x76
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Sprite 0x77
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0x78
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Sprite 0x79
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Sprite 0x7a
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0x7b
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0x7c
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Sprite 0x7d
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0x7e
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Sprite 0x7f
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000", -- 2047 - 0x7ff  :    0 - 0x0
    "00000000", -- 2048 - 0x800  :    0 - 0x0 -- Sprite 0x80
    "00000000", -- 2049 - 0x801  :    0 - 0x0
    "00000000", -- 2050 - 0x802  :    0 - 0x0
    "00000000", -- 2051 - 0x803  :    0 - 0x0
    "00000000", -- 2052 - 0x804  :    0 - 0x0
    "00000000", -- 2053 - 0x805  :    0 - 0x0
    "00000000", -- 2054 - 0x806  :    0 - 0x0
    "00000000", -- 2055 - 0x807  :    0 - 0x0
    "00000000", -- 2056 - 0x808  :    0 - 0x0
    "00000000", -- 2057 - 0x809  :    0 - 0x0
    "00000000", -- 2058 - 0x80a  :    0 - 0x0
    "00000000", -- 2059 - 0x80b  :    0 - 0x0
    "00000000", -- 2060 - 0x80c  :    0 - 0x0
    "00000000", -- 2061 - 0x80d  :    0 - 0x0
    "00000000", -- 2062 - 0x80e  :    0 - 0x0
    "00000000", -- 2063 - 0x80f  :    0 - 0x0
    "00000000", -- 2064 - 0x810  :    0 - 0x0 -- Sprite 0x81
    "00000000", -- 2065 - 0x811  :    0 - 0x0
    "00000000", -- 2066 - 0x812  :    0 - 0x0
    "00000000", -- 2067 - 0x813  :    0 - 0x0
    "00000000", -- 2068 - 0x814  :    0 - 0x0
    "00000000", -- 2069 - 0x815  :    0 - 0x0
    "00000000", -- 2070 - 0x816  :    0 - 0x0
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "00000000", -- 2072 - 0x818  :    0 - 0x0
    "00000000", -- 2073 - 0x819  :    0 - 0x0
    "00000000", -- 2074 - 0x81a  :    0 - 0x0
    "00000000", -- 2075 - 0x81b  :    0 - 0x0
    "00000000", -- 2076 - 0x81c  :    0 - 0x0
    "00000000", -- 2077 - 0x81d  :    0 - 0x0
    "00000000", -- 2078 - 0x81e  :    0 - 0x0
    "00000000", -- 2079 - 0x81f  :    0 - 0x0
    "00000000", -- 2080 - 0x820  :    0 - 0x0 -- Sprite 0x82
    "00000000", -- 2081 - 0x821  :    0 - 0x0
    "00000000", -- 2082 - 0x822  :    0 - 0x0
    "00000000", -- 2083 - 0x823  :    0 - 0x0
    "00000000", -- 2084 - 0x824  :    0 - 0x0
    "00000000", -- 2085 - 0x825  :    0 - 0x0
    "00000000", -- 2086 - 0x826  :    0 - 0x0
    "00000000", -- 2087 - 0x827  :    0 - 0x0
    "00000000", -- 2088 - 0x828  :    0 - 0x0
    "00000000", -- 2089 - 0x829  :    0 - 0x0
    "00000000", -- 2090 - 0x82a  :    0 - 0x0
    "00000000", -- 2091 - 0x82b  :    0 - 0x0
    "00000000", -- 2092 - 0x82c  :    0 - 0x0
    "00000000", -- 2093 - 0x82d  :    0 - 0x0
    "00000000", -- 2094 - 0x82e  :    0 - 0x0
    "00000000", -- 2095 - 0x82f  :    0 - 0x0
    "00000000", -- 2096 - 0x830  :    0 - 0x0 -- Sprite 0x83
    "00000000", -- 2097 - 0x831  :    0 - 0x0
    "00000000", -- 2098 - 0x832  :    0 - 0x0
    "00000000", -- 2099 - 0x833  :    0 - 0x0
    "00000000", -- 2100 - 0x834  :    0 - 0x0
    "00000000", -- 2101 - 0x835  :    0 - 0x0
    "00000000", -- 2102 - 0x836  :    0 - 0x0
    "00000000", -- 2103 - 0x837  :    0 - 0x0
    "00000000", -- 2104 - 0x838  :    0 - 0x0
    "00000000", -- 2105 - 0x839  :    0 - 0x0
    "00000000", -- 2106 - 0x83a  :    0 - 0x0
    "00000000", -- 2107 - 0x83b  :    0 - 0x0
    "00000000", -- 2108 - 0x83c  :    0 - 0x0
    "00000000", -- 2109 - 0x83d  :    0 - 0x0
    "00000000", -- 2110 - 0x83e  :    0 - 0x0
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "00000000", -- 2112 - 0x840  :    0 - 0x0 -- Sprite 0x84
    "00000000", -- 2113 - 0x841  :    0 - 0x0
    "00000000", -- 2114 - 0x842  :    0 - 0x0
    "00000000", -- 2115 - 0x843  :    0 - 0x0
    "00000000", -- 2116 - 0x844  :    0 - 0x0
    "00000000", -- 2117 - 0x845  :    0 - 0x0
    "00000000", -- 2118 - 0x846  :    0 - 0x0
    "00000000", -- 2119 - 0x847  :    0 - 0x0
    "00000000", -- 2120 - 0x848  :    0 - 0x0
    "00000000", -- 2121 - 0x849  :    0 - 0x0
    "00000000", -- 2122 - 0x84a  :    0 - 0x0
    "00000000", -- 2123 - 0x84b  :    0 - 0x0
    "00000000", -- 2124 - 0x84c  :    0 - 0x0
    "00000000", -- 2125 - 0x84d  :    0 - 0x0
    "00000000", -- 2126 - 0x84e  :    0 - 0x0
    "00000000", -- 2127 - 0x84f  :    0 - 0x0
    "00000000", -- 2128 - 0x850  :    0 - 0x0 -- Sprite 0x85
    "00000000", -- 2129 - 0x851  :    0 - 0x0
    "00000000", -- 2130 - 0x852  :    0 - 0x0
    "00000000", -- 2131 - 0x853  :    0 - 0x0
    "00000000", -- 2132 - 0x854  :    0 - 0x0
    "00000000", -- 2133 - 0x855  :    0 - 0x0
    "00000000", -- 2134 - 0x856  :    0 - 0x0
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "00000000", -- 2136 - 0x858  :    0 - 0x0
    "00000000", -- 2137 - 0x859  :    0 - 0x0
    "00000000", -- 2138 - 0x85a  :    0 - 0x0
    "00000000", -- 2139 - 0x85b  :    0 - 0x0
    "00000000", -- 2140 - 0x85c  :    0 - 0x0
    "00000000", -- 2141 - 0x85d  :    0 - 0x0
    "00000000", -- 2142 - 0x85e  :    0 - 0x0
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "00000000", -- 2144 - 0x860  :    0 - 0x0 -- Sprite 0x86
    "00000000", -- 2145 - 0x861  :    0 - 0x0
    "00000000", -- 2146 - 0x862  :    0 - 0x0
    "00000000", -- 2147 - 0x863  :    0 - 0x0
    "00000000", -- 2148 - 0x864  :    0 - 0x0
    "00000000", -- 2149 - 0x865  :    0 - 0x0
    "00000000", -- 2150 - 0x866  :    0 - 0x0
    "00000000", -- 2151 - 0x867  :    0 - 0x0
    "00000000", -- 2152 - 0x868  :    0 - 0x0
    "00000000", -- 2153 - 0x869  :    0 - 0x0
    "00000000", -- 2154 - 0x86a  :    0 - 0x0
    "00000000", -- 2155 - 0x86b  :    0 - 0x0
    "00000000", -- 2156 - 0x86c  :    0 - 0x0
    "00000000", -- 2157 - 0x86d  :    0 - 0x0
    "00000000", -- 2158 - 0x86e  :    0 - 0x0
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "00000000", -- 2160 - 0x870  :    0 - 0x0 -- Sprite 0x87
    "00000000", -- 2161 - 0x871  :    0 - 0x0
    "00000000", -- 2162 - 0x872  :    0 - 0x0
    "00000000", -- 2163 - 0x873  :    0 - 0x0
    "00000000", -- 2164 - 0x874  :    0 - 0x0
    "00000000", -- 2165 - 0x875  :    0 - 0x0
    "00000000", -- 2166 - 0x876  :    0 - 0x0
    "00000000", -- 2167 - 0x877  :    0 - 0x0
    "00000000", -- 2168 - 0x878  :    0 - 0x0
    "00000000", -- 2169 - 0x879  :    0 - 0x0
    "00000000", -- 2170 - 0x87a  :    0 - 0x0
    "00000000", -- 2171 - 0x87b  :    0 - 0x0
    "00000000", -- 2172 - 0x87c  :    0 - 0x0
    "00000000", -- 2173 - 0x87d  :    0 - 0x0
    "00000000", -- 2174 - 0x87e  :    0 - 0x0
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "00000000", -- 2176 - 0x880  :    0 - 0x0 -- Sprite 0x88
    "00000000", -- 2177 - 0x881  :    0 - 0x0
    "00000000", -- 2178 - 0x882  :    0 - 0x0
    "00000000", -- 2179 - 0x883  :    0 - 0x0
    "00000000", -- 2180 - 0x884  :    0 - 0x0
    "00000000", -- 2181 - 0x885  :    0 - 0x0
    "00000000", -- 2182 - 0x886  :    0 - 0x0
    "00000000", -- 2183 - 0x887  :    0 - 0x0
    "00000000", -- 2184 - 0x888  :    0 - 0x0
    "00000000", -- 2185 - 0x889  :    0 - 0x0
    "00000000", -- 2186 - 0x88a  :    0 - 0x0
    "00000000", -- 2187 - 0x88b  :    0 - 0x0
    "00000000", -- 2188 - 0x88c  :    0 - 0x0
    "00000000", -- 2189 - 0x88d  :    0 - 0x0
    "00000000", -- 2190 - 0x88e  :    0 - 0x0
    "00000000", -- 2191 - 0x88f  :    0 - 0x0
    "00000000", -- 2192 - 0x890  :    0 - 0x0 -- Sprite 0x89
    "00000000", -- 2193 - 0x891  :    0 - 0x0
    "00000000", -- 2194 - 0x892  :    0 - 0x0
    "00000000", -- 2195 - 0x893  :    0 - 0x0
    "00000000", -- 2196 - 0x894  :    0 - 0x0
    "00000000", -- 2197 - 0x895  :    0 - 0x0
    "00000000", -- 2198 - 0x896  :    0 - 0x0
    "00000000", -- 2199 - 0x897  :    0 - 0x0
    "00000000", -- 2200 - 0x898  :    0 - 0x0
    "00000000", -- 2201 - 0x899  :    0 - 0x0
    "00000000", -- 2202 - 0x89a  :    0 - 0x0
    "00000000", -- 2203 - 0x89b  :    0 - 0x0
    "00000000", -- 2204 - 0x89c  :    0 - 0x0
    "00000000", -- 2205 - 0x89d  :    0 - 0x0
    "00000000", -- 2206 - 0x89e  :    0 - 0x0
    "00000000", -- 2207 - 0x89f  :    0 - 0x0
    "00000000", -- 2208 - 0x8a0  :    0 - 0x0 -- Sprite 0x8a
    "00000000", -- 2209 - 0x8a1  :    0 - 0x0
    "00000000", -- 2210 - 0x8a2  :    0 - 0x0
    "00000000", -- 2211 - 0x8a3  :    0 - 0x0
    "00000000", -- 2212 - 0x8a4  :    0 - 0x0
    "00000000", -- 2213 - 0x8a5  :    0 - 0x0
    "00000000", -- 2214 - 0x8a6  :    0 - 0x0
    "00000000", -- 2215 - 0x8a7  :    0 - 0x0
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0
    "00000000", -- 2217 - 0x8a9  :    0 - 0x0
    "00000000", -- 2218 - 0x8aa  :    0 - 0x0
    "00000000", -- 2219 - 0x8ab  :    0 - 0x0
    "00000000", -- 2220 - 0x8ac  :    0 - 0x0
    "00000000", -- 2221 - 0x8ad  :    0 - 0x0
    "00000000", -- 2222 - 0x8ae  :    0 - 0x0
    "00000000", -- 2223 - 0x8af  :    0 - 0x0
    "00000000", -- 2224 - 0x8b0  :    0 - 0x0 -- Sprite 0x8b
    "00000000", -- 2225 - 0x8b1  :    0 - 0x0
    "00000000", -- 2226 - 0x8b2  :    0 - 0x0
    "00000000", -- 2227 - 0x8b3  :    0 - 0x0
    "00000000", -- 2228 - 0x8b4  :    0 - 0x0
    "00000000", -- 2229 - 0x8b5  :    0 - 0x0
    "00000000", -- 2230 - 0x8b6  :    0 - 0x0
    "00000000", -- 2231 - 0x8b7  :    0 - 0x0
    "00000000", -- 2232 - 0x8b8  :    0 - 0x0
    "00000000", -- 2233 - 0x8b9  :    0 - 0x0
    "00000000", -- 2234 - 0x8ba  :    0 - 0x0
    "00000000", -- 2235 - 0x8bb  :    0 - 0x0
    "00000000", -- 2236 - 0x8bc  :    0 - 0x0
    "00000000", -- 2237 - 0x8bd  :    0 - 0x0
    "00000000", -- 2238 - 0x8be  :    0 - 0x0
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "00000000", -- 2240 - 0x8c0  :    0 - 0x0 -- Sprite 0x8c
    "00000000", -- 2241 - 0x8c1  :    0 - 0x0
    "00000000", -- 2242 - 0x8c2  :    0 - 0x0
    "00000000", -- 2243 - 0x8c3  :    0 - 0x0
    "00000000", -- 2244 - 0x8c4  :    0 - 0x0
    "00000000", -- 2245 - 0x8c5  :    0 - 0x0
    "00000000", -- 2246 - 0x8c6  :    0 - 0x0
    "00000000", -- 2247 - 0x8c7  :    0 - 0x0
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0
    "00000000", -- 2249 - 0x8c9  :    0 - 0x0
    "00000000", -- 2250 - 0x8ca  :    0 - 0x0
    "00000000", -- 2251 - 0x8cb  :    0 - 0x0
    "00000000", -- 2252 - 0x8cc  :    0 - 0x0
    "00000000", -- 2253 - 0x8cd  :    0 - 0x0
    "00000000", -- 2254 - 0x8ce  :    0 - 0x0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "00000000", -- 2256 - 0x8d0  :    0 - 0x0 -- Sprite 0x8d
    "00000000", -- 2257 - 0x8d1  :    0 - 0x0
    "00000000", -- 2258 - 0x8d2  :    0 - 0x0
    "00000000", -- 2259 - 0x8d3  :    0 - 0x0
    "00000000", -- 2260 - 0x8d4  :    0 - 0x0
    "00000000", -- 2261 - 0x8d5  :    0 - 0x0
    "00000000", -- 2262 - 0x8d6  :    0 - 0x0
    "00000000", -- 2263 - 0x8d7  :    0 - 0x0
    "00000000", -- 2264 - 0x8d8  :    0 - 0x0
    "00000000", -- 2265 - 0x8d9  :    0 - 0x0
    "00000000", -- 2266 - 0x8da  :    0 - 0x0
    "00000000", -- 2267 - 0x8db  :    0 - 0x0
    "00000000", -- 2268 - 0x8dc  :    0 - 0x0
    "00000000", -- 2269 - 0x8dd  :    0 - 0x0
    "00000000", -- 2270 - 0x8de  :    0 - 0x0
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "00000000", -- 2272 - 0x8e0  :    0 - 0x0 -- Sprite 0x8e
    "00000000", -- 2273 - 0x8e1  :    0 - 0x0
    "00000000", -- 2274 - 0x8e2  :    0 - 0x0
    "00000000", -- 2275 - 0x8e3  :    0 - 0x0
    "00000000", -- 2276 - 0x8e4  :    0 - 0x0
    "00000000", -- 2277 - 0x8e5  :    0 - 0x0
    "00000000", -- 2278 - 0x8e6  :    0 - 0x0
    "00000000", -- 2279 - 0x8e7  :    0 - 0x0
    "00000000", -- 2280 - 0x8e8  :    0 - 0x0
    "00000000", -- 2281 - 0x8e9  :    0 - 0x0
    "00000000", -- 2282 - 0x8ea  :    0 - 0x0
    "00000000", -- 2283 - 0x8eb  :    0 - 0x0
    "00000000", -- 2284 - 0x8ec  :    0 - 0x0
    "00000000", -- 2285 - 0x8ed  :    0 - 0x0
    "00000000", -- 2286 - 0x8ee  :    0 - 0x0
    "00000000", -- 2287 - 0x8ef  :    0 - 0x0
    "00000000", -- 2288 - 0x8f0  :    0 - 0x0 -- Sprite 0x8f
    "00000000", -- 2289 - 0x8f1  :    0 - 0x0
    "00000000", -- 2290 - 0x8f2  :    0 - 0x0
    "00000000", -- 2291 - 0x8f3  :    0 - 0x0
    "00000000", -- 2292 - 0x8f4  :    0 - 0x0
    "00000000", -- 2293 - 0x8f5  :    0 - 0x0
    "00000000", -- 2294 - 0x8f6  :    0 - 0x0
    "00000000", -- 2295 - 0x8f7  :    0 - 0x0
    "00000000", -- 2296 - 0x8f8  :    0 - 0x0
    "00000000", -- 2297 - 0x8f9  :    0 - 0x0
    "00000000", -- 2298 - 0x8fa  :    0 - 0x0
    "00000000", -- 2299 - 0x8fb  :    0 - 0x0
    "00000000", -- 2300 - 0x8fc  :    0 - 0x0
    "00000000", -- 2301 - 0x8fd  :    0 - 0x0
    "00000000", -- 2302 - 0x8fe  :    0 - 0x0
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "00000000", -- 2304 - 0x900  :    0 - 0x0 -- Sprite 0x90
    "00000000", -- 2305 - 0x901  :    0 - 0x0
    "00000000", -- 2306 - 0x902  :    0 - 0x0
    "00000000", -- 2307 - 0x903  :    0 - 0x0
    "00000000", -- 2308 - 0x904  :    0 - 0x0
    "00000000", -- 2309 - 0x905  :    0 - 0x0
    "00000000", -- 2310 - 0x906  :    0 - 0x0
    "00000000", -- 2311 - 0x907  :    0 - 0x0
    "00000000", -- 2312 - 0x908  :    0 - 0x0
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "00000000", -- 2315 - 0x90b  :    0 - 0x0
    "00000000", -- 2316 - 0x90c  :    0 - 0x0
    "00000000", -- 2317 - 0x90d  :    0 - 0x0
    "00000000", -- 2318 - 0x90e  :    0 - 0x0
    "00000000", -- 2319 - 0x90f  :    0 - 0x0
    "00000000", -- 2320 - 0x910  :    0 - 0x0 -- Sprite 0x91
    "00000000", -- 2321 - 0x911  :    0 - 0x0
    "00000000", -- 2322 - 0x912  :    0 - 0x0
    "00000000", -- 2323 - 0x913  :    0 - 0x0
    "00000000", -- 2324 - 0x914  :    0 - 0x0
    "00000000", -- 2325 - 0x915  :    0 - 0x0
    "00000000", -- 2326 - 0x916  :    0 - 0x0
    "00000000", -- 2327 - 0x917  :    0 - 0x0
    "00000000", -- 2328 - 0x918  :    0 - 0x0
    "00000000", -- 2329 - 0x919  :    0 - 0x0
    "00000000", -- 2330 - 0x91a  :    0 - 0x0
    "00000000", -- 2331 - 0x91b  :    0 - 0x0
    "00000000", -- 2332 - 0x91c  :    0 - 0x0
    "00000000", -- 2333 - 0x91d  :    0 - 0x0
    "00000000", -- 2334 - 0x91e  :    0 - 0x0
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "00000000", -- 2336 - 0x920  :    0 - 0x0 -- Sprite 0x92
    "00000000", -- 2337 - 0x921  :    0 - 0x0
    "00000000", -- 2338 - 0x922  :    0 - 0x0
    "00000000", -- 2339 - 0x923  :    0 - 0x0
    "00000000", -- 2340 - 0x924  :    0 - 0x0
    "00000000", -- 2341 - 0x925  :    0 - 0x0
    "00000000", -- 2342 - 0x926  :    0 - 0x0
    "00000000", -- 2343 - 0x927  :    0 - 0x0
    "00000000", -- 2344 - 0x928  :    0 - 0x0
    "00000000", -- 2345 - 0x929  :    0 - 0x0
    "00000000", -- 2346 - 0x92a  :    0 - 0x0
    "00000000", -- 2347 - 0x92b  :    0 - 0x0
    "00000000", -- 2348 - 0x92c  :    0 - 0x0
    "00000000", -- 2349 - 0x92d  :    0 - 0x0
    "00000000", -- 2350 - 0x92e  :    0 - 0x0
    "00000000", -- 2351 - 0x92f  :    0 - 0x0
    "00000000", -- 2352 - 0x930  :    0 - 0x0 -- Sprite 0x93
    "00000000", -- 2353 - 0x931  :    0 - 0x0
    "00000000", -- 2354 - 0x932  :    0 - 0x0
    "00000000", -- 2355 - 0x933  :    0 - 0x0
    "00000000", -- 2356 - 0x934  :    0 - 0x0
    "00000000", -- 2357 - 0x935  :    0 - 0x0
    "00000000", -- 2358 - 0x936  :    0 - 0x0
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "00000000", -- 2360 - 0x938  :    0 - 0x0
    "00000000", -- 2361 - 0x939  :    0 - 0x0
    "00000000", -- 2362 - 0x93a  :    0 - 0x0
    "00000000", -- 2363 - 0x93b  :    0 - 0x0
    "00000000", -- 2364 - 0x93c  :    0 - 0x0
    "00000000", -- 2365 - 0x93d  :    0 - 0x0
    "00000000", -- 2366 - 0x93e  :    0 - 0x0
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Sprite 0x94
    "00000000", -- 2369 - 0x941  :    0 - 0x0
    "00000000", -- 2370 - 0x942  :    0 - 0x0
    "00000000", -- 2371 - 0x943  :    0 - 0x0
    "00000000", -- 2372 - 0x944  :    0 - 0x0
    "00000000", -- 2373 - 0x945  :    0 - 0x0
    "00000000", -- 2374 - 0x946  :    0 - 0x0
    "00000000", -- 2375 - 0x947  :    0 - 0x0
    "00000000", -- 2376 - 0x948  :    0 - 0x0
    "00000000", -- 2377 - 0x949  :    0 - 0x0
    "00000000", -- 2378 - 0x94a  :    0 - 0x0
    "00000000", -- 2379 - 0x94b  :    0 - 0x0
    "00000000", -- 2380 - 0x94c  :    0 - 0x0
    "00000000", -- 2381 - 0x94d  :    0 - 0x0
    "00000000", -- 2382 - 0x94e  :    0 - 0x0
    "00000000", -- 2383 - 0x94f  :    0 - 0x0
    "00000000", -- 2384 - 0x950  :    0 - 0x0 -- Sprite 0x95
    "00000000", -- 2385 - 0x951  :    0 - 0x0
    "00000000", -- 2386 - 0x952  :    0 - 0x0
    "00000000", -- 2387 - 0x953  :    0 - 0x0
    "00000000", -- 2388 - 0x954  :    0 - 0x0
    "00000000", -- 2389 - 0x955  :    0 - 0x0
    "00000000", -- 2390 - 0x956  :    0 - 0x0
    "00000000", -- 2391 - 0x957  :    0 - 0x0
    "00000000", -- 2392 - 0x958  :    0 - 0x0
    "00000000", -- 2393 - 0x959  :    0 - 0x0
    "00000000", -- 2394 - 0x95a  :    0 - 0x0
    "00000000", -- 2395 - 0x95b  :    0 - 0x0
    "00000000", -- 2396 - 0x95c  :    0 - 0x0
    "00000000", -- 2397 - 0x95d  :    0 - 0x0
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "00000000", -- 2400 - 0x960  :    0 - 0x0 -- Sprite 0x96
    "00000000", -- 2401 - 0x961  :    0 - 0x0
    "00000000", -- 2402 - 0x962  :    0 - 0x0
    "00000000", -- 2403 - 0x963  :    0 - 0x0
    "00000000", -- 2404 - 0x964  :    0 - 0x0
    "00000000", -- 2405 - 0x965  :    0 - 0x0
    "00000000", -- 2406 - 0x966  :    0 - 0x0
    "00000000", -- 2407 - 0x967  :    0 - 0x0
    "00000000", -- 2408 - 0x968  :    0 - 0x0
    "00000000", -- 2409 - 0x969  :    0 - 0x0
    "00000000", -- 2410 - 0x96a  :    0 - 0x0
    "00000000", -- 2411 - 0x96b  :    0 - 0x0
    "00000000", -- 2412 - 0x96c  :    0 - 0x0
    "00000000", -- 2413 - 0x96d  :    0 - 0x0
    "00000000", -- 2414 - 0x96e  :    0 - 0x0
    "00000000", -- 2415 - 0x96f  :    0 - 0x0
    "00000000", -- 2416 - 0x970  :    0 - 0x0 -- Sprite 0x97
    "00000000", -- 2417 - 0x971  :    0 - 0x0
    "00000000", -- 2418 - 0x972  :    0 - 0x0
    "00000000", -- 2419 - 0x973  :    0 - 0x0
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "00000000", -- 2424 - 0x978  :    0 - 0x0
    "00000000", -- 2425 - 0x979  :    0 - 0x0
    "00000000", -- 2426 - 0x97a  :    0 - 0x0
    "00000000", -- 2427 - 0x97b  :    0 - 0x0
    "00000000", -- 2428 - 0x97c  :    0 - 0x0
    "00000000", -- 2429 - 0x97d  :    0 - 0x0
    "00000000", -- 2430 - 0x97e  :    0 - 0x0
    "00000000", -- 2431 - 0x97f  :    0 - 0x0
    "00000000", -- 2432 - 0x980  :    0 - 0x0 -- Sprite 0x98
    "00000000", -- 2433 - 0x981  :    0 - 0x0
    "00000000", -- 2434 - 0x982  :    0 - 0x0
    "00000000", -- 2435 - 0x983  :    0 - 0x0
    "00000000", -- 2436 - 0x984  :    0 - 0x0
    "00000000", -- 2437 - 0x985  :    0 - 0x0
    "00000000", -- 2438 - 0x986  :    0 - 0x0
    "00000000", -- 2439 - 0x987  :    0 - 0x0
    "00000000", -- 2440 - 0x988  :    0 - 0x0
    "00000000", -- 2441 - 0x989  :    0 - 0x0
    "00000000", -- 2442 - 0x98a  :    0 - 0x0
    "00000000", -- 2443 - 0x98b  :    0 - 0x0
    "00000000", -- 2444 - 0x98c  :    0 - 0x0
    "00000000", -- 2445 - 0x98d  :    0 - 0x0
    "00000000", -- 2446 - 0x98e  :    0 - 0x0
    "00000000", -- 2447 - 0x98f  :    0 - 0x0
    "00000000", -- 2448 - 0x990  :    0 - 0x0 -- Sprite 0x99
    "00000000", -- 2449 - 0x991  :    0 - 0x0
    "00000000", -- 2450 - 0x992  :    0 - 0x0
    "00000000", -- 2451 - 0x993  :    0 - 0x0
    "00000000", -- 2452 - 0x994  :    0 - 0x0
    "00000000", -- 2453 - 0x995  :    0 - 0x0
    "00000000", -- 2454 - 0x996  :    0 - 0x0
    "00000000", -- 2455 - 0x997  :    0 - 0x0
    "00000000", -- 2456 - 0x998  :    0 - 0x0
    "00000000", -- 2457 - 0x999  :    0 - 0x0
    "00000000", -- 2458 - 0x99a  :    0 - 0x0
    "00000000", -- 2459 - 0x99b  :    0 - 0x0
    "00000000", -- 2460 - 0x99c  :    0 - 0x0
    "00000000", -- 2461 - 0x99d  :    0 - 0x0
    "00000000", -- 2462 - 0x99e  :    0 - 0x0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "00000000", -- 2464 - 0x9a0  :    0 - 0x0 -- Sprite 0x9a
    "00000000", -- 2465 - 0x9a1  :    0 - 0x0
    "00000000", -- 2466 - 0x9a2  :    0 - 0x0
    "00000000", -- 2467 - 0x9a3  :    0 - 0x0
    "00000000", -- 2468 - 0x9a4  :    0 - 0x0
    "00000000", -- 2469 - 0x9a5  :    0 - 0x0
    "00000000", -- 2470 - 0x9a6  :    0 - 0x0
    "00000000", -- 2471 - 0x9a7  :    0 - 0x0
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "00000000", -- 2474 - 0x9aa  :    0 - 0x0
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00000000", -- 2476 - 0x9ac  :    0 - 0x0
    "00000000", -- 2477 - 0x9ad  :    0 - 0x0
    "00000000", -- 2478 - 0x9ae  :    0 - 0x0
    "00000000", -- 2479 - 0x9af  :    0 - 0x0
    "00000000", -- 2480 - 0x9b0  :    0 - 0x0 -- Sprite 0x9b
    "00000000", -- 2481 - 0x9b1  :    0 - 0x0
    "00000000", -- 2482 - 0x9b2  :    0 - 0x0
    "00000000", -- 2483 - 0x9b3  :    0 - 0x0
    "00000000", -- 2484 - 0x9b4  :    0 - 0x0
    "00000000", -- 2485 - 0x9b5  :    0 - 0x0
    "00000000", -- 2486 - 0x9b6  :    0 - 0x0
    "00000000", -- 2487 - 0x9b7  :    0 - 0x0
    "00000000", -- 2488 - 0x9b8  :    0 - 0x0
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "00000000", -- 2490 - 0x9ba  :    0 - 0x0
    "00000000", -- 2491 - 0x9bb  :    0 - 0x0
    "00000000", -- 2492 - 0x9bc  :    0 - 0x0
    "00000000", -- 2493 - 0x9bd  :    0 - 0x0
    "00000000", -- 2494 - 0x9be  :    0 - 0x0
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0 -- Sprite 0x9c
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000000", -- 2498 - 0x9c2  :    0 - 0x0
    "00000000", -- 2499 - 0x9c3  :    0 - 0x0
    "00000000", -- 2500 - 0x9c4  :    0 - 0x0
    "00000000", -- 2501 - 0x9c5  :    0 - 0x0
    "00000000", -- 2502 - 0x9c6  :    0 - 0x0
    "00000000", -- 2503 - 0x9c7  :    0 - 0x0
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0 -- Sprite 0x9d
    "00000000", -- 2513 - 0x9d1  :    0 - 0x0
    "00000000", -- 2514 - 0x9d2  :    0 - 0x0
    "00000000", -- 2515 - 0x9d3  :    0 - 0x0
    "00000000", -- 2516 - 0x9d4  :    0 - 0x0
    "00000000", -- 2517 - 0x9d5  :    0 - 0x0
    "00000000", -- 2518 - 0x9d6  :    0 - 0x0
    "00000000", -- 2519 - 0x9d7  :    0 - 0x0
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0
    "00000000", -- 2521 - 0x9d9  :    0 - 0x0
    "00000000", -- 2522 - 0x9da  :    0 - 0x0
    "00000000", -- 2523 - 0x9db  :    0 - 0x0
    "00000000", -- 2524 - 0x9dc  :    0 - 0x0
    "00000000", -- 2525 - 0x9dd  :    0 - 0x0
    "00000000", -- 2526 - 0x9de  :    0 - 0x0
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0 -- Sprite 0x9e
    "00000000", -- 2529 - 0x9e1  :    0 - 0x0
    "00000000", -- 2530 - 0x9e2  :    0 - 0x0
    "00000000", -- 2531 - 0x9e3  :    0 - 0x0
    "00000000", -- 2532 - 0x9e4  :    0 - 0x0
    "00000000", -- 2533 - 0x9e5  :    0 - 0x0
    "00000000", -- 2534 - 0x9e6  :    0 - 0x0
    "00000000", -- 2535 - 0x9e7  :    0 - 0x0
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0
    "00000000", -- 2537 - 0x9e9  :    0 - 0x0
    "00000000", -- 2538 - 0x9ea  :    0 - 0x0
    "00000000", -- 2539 - 0x9eb  :    0 - 0x0
    "00000000", -- 2540 - 0x9ec  :    0 - 0x0
    "00000000", -- 2541 - 0x9ed  :    0 - 0x0
    "00000000", -- 2542 - 0x9ee  :    0 - 0x0
    "00000000", -- 2543 - 0x9ef  :    0 - 0x0
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0 -- Sprite 0x9f
    "00000000", -- 2545 - 0x9f1  :    0 - 0x0
    "00000000", -- 2546 - 0x9f2  :    0 - 0x0
    "00000000", -- 2547 - 0x9f3  :    0 - 0x0
    "00000000", -- 2548 - 0x9f4  :    0 - 0x0
    "00000000", -- 2549 - 0x9f5  :    0 - 0x0
    "00000000", -- 2550 - 0x9f6  :    0 - 0x0
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00000000", -- 2560 - 0xa00  :    0 - 0x0 -- Sprite 0xa0
    "00000000", -- 2561 - 0xa01  :    0 - 0x0
    "00000000", -- 2562 - 0xa02  :    0 - 0x0
    "00000000", -- 2563 - 0xa03  :    0 - 0x0
    "00000000", -- 2564 - 0xa04  :    0 - 0x0
    "00000000", -- 2565 - 0xa05  :    0 - 0x0
    "00000000", -- 2566 - 0xa06  :    0 - 0x0
    "00000000", -- 2567 - 0xa07  :    0 - 0x0
    "00000000", -- 2568 - 0xa08  :    0 - 0x0
    "00000000", -- 2569 - 0xa09  :    0 - 0x0
    "00000000", -- 2570 - 0xa0a  :    0 - 0x0
    "00000000", -- 2571 - 0xa0b  :    0 - 0x0
    "00000000", -- 2572 - 0xa0c  :    0 - 0x0
    "00000000", -- 2573 - 0xa0d  :    0 - 0x0
    "00000000", -- 2574 - 0xa0e  :    0 - 0x0
    "00000000", -- 2575 - 0xa0f  :    0 - 0x0
    "00000000", -- 2576 - 0xa10  :    0 - 0x0 -- Sprite 0xa1
    "00000000", -- 2577 - 0xa11  :    0 - 0x0
    "00000000", -- 2578 - 0xa12  :    0 - 0x0
    "00000000", -- 2579 - 0xa13  :    0 - 0x0
    "00000000", -- 2580 - 0xa14  :    0 - 0x0
    "00000000", -- 2581 - 0xa15  :    0 - 0x0
    "00000000", -- 2582 - 0xa16  :    0 - 0x0
    "00000000", -- 2583 - 0xa17  :    0 - 0x0
    "00000000", -- 2584 - 0xa18  :    0 - 0x0
    "00000000", -- 2585 - 0xa19  :    0 - 0x0
    "00000000", -- 2586 - 0xa1a  :    0 - 0x0
    "00000000", -- 2587 - 0xa1b  :    0 - 0x0
    "00000000", -- 2588 - 0xa1c  :    0 - 0x0
    "00000000", -- 2589 - 0xa1d  :    0 - 0x0
    "00000000", -- 2590 - 0xa1e  :    0 - 0x0
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "00000000", -- 2592 - 0xa20  :    0 - 0x0 -- Sprite 0xa2
    "00000000", -- 2593 - 0xa21  :    0 - 0x0
    "00000000", -- 2594 - 0xa22  :    0 - 0x0
    "00000000", -- 2595 - 0xa23  :    0 - 0x0
    "00000000", -- 2596 - 0xa24  :    0 - 0x0
    "00000000", -- 2597 - 0xa25  :    0 - 0x0
    "00000000", -- 2598 - 0xa26  :    0 - 0x0
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00000000", -- 2600 - 0xa28  :    0 - 0x0
    "00000000", -- 2601 - 0xa29  :    0 - 0x0
    "00000000", -- 2602 - 0xa2a  :    0 - 0x0
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "00000000", -- 2608 - 0xa30  :    0 - 0x0 -- Sprite 0xa3
    "00000000", -- 2609 - 0xa31  :    0 - 0x0
    "00000000", -- 2610 - 0xa32  :    0 - 0x0
    "00000000", -- 2611 - 0xa33  :    0 - 0x0
    "00000000", -- 2612 - 0xa34  :    0 - 0x0
    "00000000", -- 2613 - 0xa35  :    0 - 0x0
    "00000000", -- 2614 - 0xa36  :    0 - 0x0
    "00000000", -- 2615 - 0xa37  :    0 - 0x0
    "00000000", -- 2616 - 0xa38  :    0 - 0x0
    "00000000", -- 2617 - 0xa39  :    0 - 0x0
    "00000000", -- 2618 - 0xa3a  :    0 - 0x0
    "00000000", -- 2619 - 0xa3b  :    0 - 0x0
    "00000000", -- 2620 - 0xa3c  :    0 - 0x0
    "00000000", -- 2621 - 0xa3d  :    0 - 0x0
    "00000000", -- 2622 - 0xa3e  :    0 - 0x0
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "00000000", -- 2624 - 0xa40  :    0 - 0x0 -- Sprite 0xa4
    "00000000", -- 2625 - 0xa41  :    0 - 0x0
    "00000000", -- 2626 - 0xa42  :    0 - 0x0
    "00000000", -- 2627 - 0xa43  :    0 - 0x0
    "00000000", -- 2628 - 0xa44  :    0 - 0x0
    "00000000", -- 2629 - 0xa45  :    0 - 0x0
    "00000000", -- 2630 - 0xa46  :    0 - 0x0
    "00000000", -- 2631 - 0xa47  :    0 - 0x0
    "00000000", -- 2632 - 0xa48  :    0 - 0x0
    "00000000", -- 2633 - 0xa49  :    0 - 0x0
    "00000000", -- 2634 - 0xa4a  :    0 - 0x0
    "00000000", -- 2635 - 0xa4b  :    0 - 0x0
    "00000000", -- 2636 - 0xa4c  :    0 - 0x0
    "00000000", -- 2637 - 0xa4d  :    0 - 0x0
    "00000000", -- 2638 - 0xa4e  :    0 - 0x0
    "00000000", -- 2639 - 0xa4f  :    0 - 0x0
    "00000000", -- 2640 - 0xa50  :    0 - 0x0 -- Sprite 0xa5
    "00000000", -- 2641 - 0xa51  :    0 - 0x0
    "00000000", -- 2642 - 0xa52  :    0 - 0x0
    "00000000", -- 2643 - 0xa53  :    0 - 0x0
    "00000000", -- 2644 - 0xa54  :    0 - 0x0
    "00000000", -- 2645 - 0xa55  :    0 - 0x0
    "00000000", -- 2646 - 0xa56  :    0 - 0x0
    "00000000", -- 2647 - 0xa57  :    0 - 0x0
    "00000000", -- 2648 - 0xa58  :    0 - 0x0
    "00000000", -- 2649 - 0xa59  :    0 - 0x0
    "00000000", -- 2650 - 0xa5a  :    0 - 0x0
    "00000000", -- 2651 - 0xa5b  :    0 - 0x0
    "00000000", -- 2652 - 0xa5c  :    0 - 0x0
    "00000000", -- 2653 - 0xa5d  :    0 - 0x0
    "00000000", -- 2654 - 0xa5e  :    0 - 0x0
    "00000000", -- 2655 - 0xa5f  :    0 - 0x0
    "00000000", -- 2656 - 0xa60  :    0 - 0x0 -- Sprite 0xa6
    "00000000", -- 2657 - 0xa61  :    0 - 0x0
    "00000000", -- 2658 - 0xa62  :    0 - 0x0
    "00000000", -- 2659 - 0xa63  :    0 - 0x0
    "00000000", -- 2660 - 0xa64  :    0 - 0x0
    "00000000", -- 2661 - 0xa65  :    0 - 0x0
    "00000000", -- 2662 - 0xa66  :    0 - 0x0
    "00000000", -- 2663 - 0xa67  :    0 - 0x0
    "00000000", -- 2664 - 0xa68  :    0 - 0x0
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "00000000", -- 2666 - 0xa6a  :    0 - 0x0
    "00000000", -- 2667 - 0xa6b  :    0 - 0x0
    "00000000", -- 2668 - 0xa6c  :    0 - 0x0
    "00000000", -- 2669 - 0xa6d  :    0 - 0x0
    "00000000", -- 2670 - 0xa6e  :    0 - 0x0
    "00000000", -- 2671 - 0xa6f  :    0 - 0x0
    "00000000", -- 2672 - 0xa70  :    0 - 0x0 -- Sprite 0xa7
    "00000000", -- 2673 - 0xa71  :    0 - 0x0
    "00000000", -- 2674 - 0xa72  :    0 - 0x0
    "00000000", -- 2675 - 0xa73  :    0 - 0x0
    "00000000", -- 2676 - 0xa74  :    0 - 0x0
    "00000000", -- 2677 - 0xa75  :    0 - 0x0
    "00000000", -- 2678 - 0xa76  :    0 - 0x0
    "00000000", -- 2679 - 0xa77  :    0 - 0x0
    "00000000", -- 2680 - 0xa78  :    0 - 0x0
    "00000000", -- 2681 - 0xa79  :    0 - 0x0
    "00000000", -- 2682 - 0xa7a  :    0 - 0x0
    "00000000", -- 2683 - 0xa7b  :    0 - 0x0
    "00000000", -- 2684 - 0xa7c  :    0 - 0x0
    "00000000", -- 2685 - 0xa7d  :    0 - 0x0
    "00000000", -- 2686 - 0xa7e  :    0 - 0x0
    "00000000", -- 2687 - 0xa7f  :    0 - 0x0
    "00000000", -- 2688 - 0xa80  :    0 - 0x0 -- Sprite 0xa8
    "00000000", -- 2689 - 0xa81  :    0 - 0x0
    "00000000", -- 2690 - 0xa82  :    0 - 0x0
    "00000000", -- 2691 - 0xa83  :    0 - 0x0
    "00000000", -- 2692 - 0xa84  :    0 - 0x0
    "00000000", -- 2693 - 0xa85  :    0 - 0x0
    "00000000", -- 2694 - 0xa86  :    0 - 0x0
    "00000000", -- 2695 - 0xa87  :    0 - 0x0
    "00000000", -- 2696 - 0xa88  :    0 - 0x0
    "00000000", -- 2697 - 0xa89  :    0 - 0x0
    "00000000", -- 2698 - 0xa8a  :    0 - 0x0
    "00000000", -- 2699 - 0xa8b  :    0 - 0x0
    "00000000", -- 2700 - 0xa8c  :    0 - 0x0
    "00000000", -- 2701 - 0xa8d  :    0 - 0x0
    "00000000", -- 2702 - 0xa8e  :    0 - 0x0
    "00000000", -- 2703 - 0xa8f  :    0 - 0x0
    "00000000", -- 2704 - 0xa90  :    0 - 0x0 -- Sprite 0xa9
    "00000000", -- 2705 - 0xa91  :    0 - 0x0
    "00000000", -- 2706 - 0xa92  :    0 - 0x0
    "00000000", -- 2707 - 0xa93  :    0 - 0x0
    "00000000", -- 2708 - 0xa94  :    0 - 0x0
    "00000000", -- 2709 - 0xa95  :    0 - 0x0
    "00000000", -- 2710 - 0xa96  :    0 - 0x0
    "00000000", -- 2711 - 0xa97  :    0 - 0x0
    "00000000", -- 2712 - 0xa98  :    0 - 0x0
    "00000000", -- 2713 - 0xa99  :    0 - 0x0
    "00000000", -- 2714 - 0xa9a  :    0 - 0x0
    "00000000", -- 2715 - 0xa9b  :    0 - 0x0
    "00000000", -- 2716 - 0xa9c  :    0 - 0x0
    "00000000", -- 2717 - 0xa9d  :    0 - 0x0
    "00000000", -- 2718 - 0xa9e  :    0 - 0x0
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "00000000", -- 2720 - 0xaa0  :    0 - 0x0 -- Sprite 0xaa
    "00000000", -- 2721 - 0xaa1  :    0 - 0x0
    "00000000", -- 2722 - 0xaa2  :    0 - 0x0
    "00000000", -- 2723 - 0xaa3  :    0 - 0x0
    "00000000", -- 2724 - 0xaa4  :    0 - 0x0
    "00000000", -- 2725 - 0xaa5  :    0 - 0x0
    "00000000", -- 2726 - 0xaa6  :    0 - 0x0
    "00000000", -- 2727 - 0xaa7  :    0 - 0x0
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "00000000", -- 2730 - 0xaaa  :    0 - 0x0
    "00000000", -- 2731 - 0xaab  :    0 - 0x0
    "00000000", -- 2732 - 0xaac  :    0 - 0x0
    "00000000", -- 2733 - 0xaad  :    0 - 0x0
    "00000000", -- 2734 - 0xaae  :    0 - 0x0
    "00000000", -- 2735 - 0xaaf  :    0 - 0x0
    "00000000", -- 2736 - 0xab0  :    0 - 0x0 -- Sprite 0xab
    "00000000", -- 2737 - 0xab1  :    0 - 0x0
    "00000000", -- 2738 - 0xab2  :    0 - 0x0
    "00000000", -- 2739 - 0xab3  :    0 - 0x0
    "00000000", -- 2740 - 0xab4  :    0 - 0x0
    "00000000", -- 2741 - 0xab5  :    0 - 0x0
    "00000000", -- 2742 - 0xab6  :    0 - 0x0
    "00000000", -- 2743 - 0xab7  :    0 - 0x0
    "00000000", -- 2744 - 0xab8  :    0 - 0x0
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "00000000", -- 2747 - 0xabb  :    0 - 0x0
    "00000000", -- 2748 - 0xabc  :    0 - 0x0
    "00000000", -- 2749 - 0xabd  :    0 - 0x0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "00000000", -- 2752 - 0xac0  :    0 - 0x0 -- Sprite 0xac
    "00000000", -- 2753 - 0xac1  :    0 - 0x0
    "00000000", -- 2754 - 0xac2  :    0 - 0x0
    "00000000", -- 2755 - 0xac3  :    0 - 0x0
    "00000000", -- 2756 - 0xac4  :    0 - 0x0
    "00000000", -- 2757 - 0xac5  :    0 - 0x0
    "00000000", -- 2758 - 0xac6  :    0 - 0x0
    "00000000", -- 2759 - 0xac7  :    0 - 0x0
    "00000000", -- 2760 - 0xac8  :    0 - 0x0
    "00000000", -- 2761 - 0xac9  :    0 - 0x0
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000000", -- 2763 - 0xacb  :    0 - 0x0
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "00000000", -- 2768 - 0xad0  :    0 - 0x0 -- Sprite 0xad
    "00000000", -- 2769 - 0xad1  :    0 - 0x0
    "00000000", -- 2770 - 0xad2  :    0 - 0x0
    "00000000", -- 2771 - 0xad3  :    0 - 0x0
    "00000000", -- 2772 - 0xad4  :    0 - 0x0
    "00000000", -- 2773 - 0xad5  :    0 - 0x0
    "00000000", -- 2774 - 0xad6  :    0 - 0x0
    "00000000", -- 2775 - 0xad7  :    0 - 0x0
    "00000000", -- 2776 - 0xad8  :    0 - 0x0
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "00000000", -- 2778 - 0xada  :    0 - 0x0
    "00000000", -- 2779 - 0xadb  :    0 - 0x0
    "00000000", -- 2780 - 0xadc  :    0 - 0x0
    "00000000", -- 2781 - 0xadd  :    0 - 0x0
    "00000000", -- 2782 - 0xade  :    0 - 0x0
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "00000000", -- 2784 - 0xae0  :    0 - 0x0 -- Sprite 0xae
    "00000000", -- 2785 - 0xae1  :    0 - 0x0
    "00000000", -- 2786 - 0xae2  :    0 - 0x0
    "00000000", -- 2787 - 0xae3  :    0 - 0x0
    "00000000", -- 2788 - 0xae4  :    0 - 0x0
    "00000000", -- 2789 - 0xae5  :    0 - 0x0
    "00000000", -- 2790 - 0xae6  :    0 - 0x0
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "00000000", -- 2792 - 0xae8  :    0 - 0x0
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000000", -- 2794 - 0xaea  :    0 - 0x0
    "00000000", -- 2795 - 0xaeb  :    0 - 0x0
    "00000000", -- 2796 - 0xaec  :    0 - 0x0
    "00000000", -- 2797 - 0xaed  :    0 - 0x0
    "00000000", -- 2798 - 0xaee  :    0 - 0x0
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "00000000", -- 2800 - 0xaf0  :    0 - 0x0 -- Sprite 0xaf
    "00000000", -- 2801 - 0xaf1  :    0 - 0x0
    "00000000", -- 2802 - 0xaf2  :    0 - 0x0
    "00000000", -- 2803 - 0xaf3  :    0 - 0x0
    "00000000", -- 2804 - 0xaf4  :    0 - 0x0
    "00000000", -- 2805 - 0xaf5  :    0 - 0x0
    "00000000", -- 2806 - 0xaf6  :    0 - 0x0
    "00000000", -- 2807 - 0xaf7  :    0 - 0x0
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0
    "00000000", -- 2809 - 0xaf9  :    0 - 0x0
    "00000000", -- 2810 - 0xafa  :    0 - 0x0
    "00000000", -- 2811 - 0xafb  :    0 - 0x0
    "00000000", -- 2812 - 0xafc  :    0 - 0x0
    "00000000", -- 2813 - 0xafd  :    0 - 0x0
    "00000000", -- 2814 - 0xafe  :    0 - 0x0
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "00000000", -- 2816 - 0xb00  :    0 - 0x0 -- Sprite 0xb0
    "00000000", -- 2817 - 0xb01  :    0 - 0x0
    "00000000", -- 2818 - 0xb02  :    0 - 0x0
    "00000000", -- 2819 - 0xb03  :    0 - 0x0
    "00000000", -- 2820 - 0xb04  :    0 - 0x0
    "00000000", -- 2821 - 0xb05  :    0 - 0x0
    "00000000", -- 2822 - 0xb06  :    0 - 0x0
    "00000000", -- 2823 - 0xb07  :    0 - 0x0
    "00000000", -- 2824 - 0xb08  :    0 - 0x0
    "00000000", -- 2825 - 0xb09  :    0 - 0x0
    "00000000", -- 2826 - 0xb0a  :    0 - 0x0
    "00000000", -- 2827 - 0xb0b  :    0 - 0x0
    "00000000", -- 2828 - 0xb0c  :    0 - 0x0
    "00000000", -- 2829 - 0xb0d  :    0 - 0x0
    "00000000", -- 2830 - 0xb0e  :    0 - 0x0
    "00000000", -- 2831 - 0xb0f  :    0 - 0x0
    "00000000", -- 2832 - 0xb10  :    0 - 0x0 -- Sprite 0xb1
    "00000000", -- 2833 - 0xb11  :    0 - 0x0
    "00000000", -- 2834 - 0xb12  :    0 - 0x0
    "00000000", -- 2835 - 0xb13  :    0 - 0x0
    "00000000", -- 2836 - 0xb14  :    0 - 0x0
    "00000000", -- 2837 - 0xb15  :    0 - 0x0
    "00000000", -- 2838 - 0xb16  :    0 - 0x0
    "00000000", -- 2839 - 0xb17  :    0 - 0x0
    "00000000", -- 2840 - 0xb18  :    0 - 0x0
    "00000000", -- 2841 - 0xb19  :    0 - 0x0
    "00000000", -- 2842 - 0xb1a  :    0 - 0x0
    "00000000", -- 2843 - 0xb1b  :    0 - 0x0
    "00000000", -- 2844 - 0xb1c  :    0 - 0x0
    "00000000", -- 2845 - 0xb1d  :    0 - 0x0
    "00000000", -- 2846 - 0xb1e  :    0 - 0x0
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "00000000", -- 2848 - 0xb20  :    0 - 0x0 -- Sprite 0xb2
    "00000000", -- 2849 - 0xb21  :    0 - 0x0
    "00000000", -- 2850 - 0xb22  :    0 - 0x0
    "00000000", -- 2851 - 0xb23  :    0 - 0x0
    "00000000", -- 2852 - 0xb24  :    0 - 0x0
    "00000000", -- 2853 - 0xb25  :    0 - 0x0
    "00000000", -- 2854 - 0xb26  :    0 - 0x0
    "00000000", -- 2855 - 0xb27  :    0 - 0x0
    "00000000", -- 2856 - 0xb28  :    0 - 0x0
    "00000000", -- 2857 - 0xb29  :    0 - 0x0
    "00000000", -- 2858 - 0xb2a  :    0 - 0x0
    "00000000", -- 2859 - 0xb2b  :    0 - 0x0
    "00000000", -- 2860 - 0xb2c  :    0 - 0x0
    "00000000", -- 2861 - 0xb2d  :    0 - 0x0
    "00000000", -- 2862 - 0xb2e  :    0 - 0x0
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "00000000", -- 2864 - 0xb30  :    0 - 0x0 -- Sprite 0xb3
    "00000000", -- 2865 - 0xb31  :    0 - 0x0
    "00000000", -- 2866 - 0xb32  :    0 - 0x0
    "00000000", -- 2867 - 0xb33  :    0 - 0x0
    "00000000", -- 2868 - 0xb34  :    0 - 0x0
    "00000000", -- 2869 - 0xb35  :    0 - 0x0
    "00000000", -- 2870 - 0xb36  :    0 - 0x0
    "00000000", -- 2871 - 0xb37  :    0 - 0x0
    "00000000", -- 2872 - 0xb38  :    0 - 0x0
    "00000000", -- 2873 - 0xb39  :    0 - 0x0
    "00000000", -- 2874 - 0xb3a  :    0 - 0x0
    "00000000", -- 2875 - 0xb3b  :    0 - 0x0
    "00000000", -- 2876 - 0xb3c  :    0 - 0x0
    "00000000", -- 2877 - 0xb3d  :    0 - 0x0
    "00000000", -- 2878 - 0xb3e  :    0 - 0x0
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "00000000", -- 2880 - 0xb40  :    0 - 0x0 -- Sprite 0xb4
    "00000000", -- 2881 - 0xb41  :    0 - 0x0
    "00000000", -- 2882 - 0xb42  :    0 - 0x0
    "00000000", -- 2883 - 0xb43  :    0 - 0x0
    "00000000", -- 2884 - 0xb44  :    0 - 0x0
    "00000000", -- 2885 - 0xb45  :    0 - 0x0
    "00000000", -- 2886 - 0xb46  :    0 - 0x0
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "00000000", -- 2888 - 0xb48  :    0 - 0x0
    "00000000", -- 2889 - 0xb49  :    0 - 0x0
    "00000000", -- 2890 - 0xb4a  :    0 - 0x0
    "00000000", -- 2891 - 0xb4b  :    0 - 0x0
    "00000000", -- 2892 - 0xb4c  :    0 - 0x0
    "00000000", -- 2893 - 0xb4d  :    0 - 0x0
    "00000000", -- 2894 - 0xb4e  :    0 - 0x0
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "00000000", -- 2896 - 0xb50  :    0 - 0x0 -- Sprite 0xb5
    "00000000", -- 2897 - 0xb51  :    0 - 0x0
    "00000000", -- 2898 - 0xb52  :    0 - 0x0
    "00000000", -- 2899 - 0xb53  :    0 - 0x0
    "00000000", -- 2900 - 0xb54  :    0 - 0x0
    "00000000", -- 2901 - 0xb55  :    0 - 0x0
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "00000000", -- 2904 - 0xb58  :    0 - 0x0
    "00000000", -- 2905 - 0xb59  :    0 - 0x0
    "00000000", -- 2906 - 0xb5a  :    0 - 0x0
    "00000000", -- 2907 - 0xb5b  :    0 - 0x0
    "00000000", -- 2908 - 0xb5c  :    0 - 0x0
    "00000000", -- 2909 - 0xb5d  :    0 - 0x0
    "00000000", -- 2910 - 0xb5e  :    0 - 0x0
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "00000000", -- 2912 - 0xb60  :    0 - 0x0 -- Sprite 0xb6
    "00000000", -- 2913 - 0xb61  :    0 - 0x0
    "00000000", -- 2914 - 0xb62  :    0 - 0x0
    "00000000", -- 2915 - 0xb63  :    0 - 0x0
    "00000000", -- 2916 - 0xb64  :    0 - 0x0
    "00000000", -- 2917 - 0xb65  :    0 - 0x0
    "00000000", -- 2918 - 0xb66  :    0 - 0x0
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "00000000", -- 2920 - 0xb68  :    0 - 0x0
    "00000000", -- 2921 - 0xb69  :    0 - 0x0
    "00000000", -- 2922 - 0xb6a  :    0 - 0x0
    "00000000", -- 2923 - 0xb6b  :    0 - 0x0
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00000000", -- 2928 - 0xb70  :    0 - 0x0 -- Sprite 0xb7
    "00000000", -- 2929 - 0xb71  :    0 - 0x0
    "00000000", -- 2930 - 0xb72  :    0 - 0x0
    "00000000", -- 2931 - 0xb73  :    0 - 0x0
    "00000000", -- 2932 - 0xb74  :    0 - 0x0
    "00000000", -- 2933 - 0xb75  :    0 - 0x0
    "00000000", -- 2934 - 0xb76  :    0 - 0x0
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "00000000", -- 2936 - 0xb78  :    0 - 0x0
    "00000000", -- 2937 - 0xb79  :    0 - 0x0
    "00000000", -- 2938 - 0xb7a  :    0 - 0x0
    "00000000", -- 2939 - 0xb7b  :    0 - 0x0
    "00000000", -- 2940 - 0xb7c  :    0 - 0x0
    "00000000", -- 2941 - 0xb7d  :    0 - 0x0
    "00000000", -- 2942 - 0xb7e  :    0 - 0x0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "00000000", -- 2944 - 0xb80  :    0 - 0x0 -- Sprite 0xb8
    "00000000", -- 2945 - 0xb81  :    0 - 0x0
    "00000000", -- 2946 - 0xb82  :    0 - 0x0
    "00000000", -- 2947 - 0xb83  :    0 - 0x0
    "00000000", -- 2948 - 0xb84  :    0 - 0x0
    "00000000", -- 2949 - 0xb85  :    0 - 0x0
    "00000000", -- 2950 - 0xb86  :    0 - 0x0
    "00000000", -- 2951 - 0xb87  :    0 - 0x0
    "00000000", -- 2952 - 0xb88  :    0 - 0x0
    "00000000", -- 2953 - 0xb89  :    0 - 0x0
    "00000000", -- 2954 - 0xb8a  :    0 - 0x0
    "00000000", -- 2955 - 0xb8b  :    0 - 0x0
    "00000000", -- 2956 - 0xb8c  :    0 - 0x0
    "00000000", -- 2957 - 0xb8d  :    0 - 0x0
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00000000", -- 2960 - 0xb90  :    0 - 0x0 -- Sprite 0xb9
    "00000000", -- 2961 - 0xb91  :    0 - 0x0
    "00000000", -- 2962 - 0xb92  :    0 - 0x0
    "00000000", -- 2963 - 0xb93  :    0 - 0x0
    "00000000", -- 2964 - 0xb94  :    0 - 0x0
    "00000000", -- 2965 - 0xb95  :    0 - 0x0
    "00000000", -- 2966 - 0xb96  :    0 - 0x0
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "00000000", -- 2968 - 0xb98  :    0 - 0x0
    "00000000", -- 2969 - 0xb99  :    0 - 0x0
    "00000000", -- 2970 - 0xb9a  :    0 - 0x0
    "00000000", -- 2971 - 0xb9b  :    0 - 0x0
    "00000000", -- 2972 - 0xb9c  :    0 - 0x0
    "00000000", -- 2973 - 0xb9d  :    0 - 0x0
    "00000000", -- 2974 - 0xb9e  :    0 - 0x0
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "00000000", -- 2976 - 0xba0  :    0 - 0x0 -- Sprite 0xba
    "00000000", -- 2977 - 0xba1  :    0 - 0x0
    "00000000", -- 2978 - 0xba2  :    0 - 0x0
    "00000000", -- 2979 - 0xba3  :    0 - 0x0
    "00000000", -- 2980 - 0xba4  :    0 - 0x0
    "00000000", -- 2981 - 0xba5  :    0 - 0x0
    "00000000", -- 2982 - 0xba6  :    0 - 0x0
    "00000000", -- 2983 - 0xba7  :    0 - 0x0
    "00000000", -- 2984 - 0xba8  :    0 - 0x0
    "00000000", -- 2985 - 0xba9  :    0 - 0x0
    "00000000", -- 2986 - 0xbaa  :    0 - 0x0
    "00000000", -- 2987 - 0xbab  :    0 - 0x0
    "00000000", -- 2988 - 0xbac  :    0 - 0x0
    "00000000", -- 2989 - 0xbad  :    0 - 0x0
    "00000000", -- 2990 - 0xbae  :    0 - 0x0
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "00000000", -- 2992 - 0xbb0  :    0 - 0x0 -- Sprite 0xbb
    "00000000", -- 2993 - 0xbb1  :    0 - 0x0
    "00000000", -- 2994 - 0xbb2  :    0 - 0x0
    "00000000", -- 2995 - 0xbb3  :    0 - 0x0
    "00000000", -- 2996 - 0xbb4  :    0 - 0x0
    "00000000", -- 2997 - 0xbb5  :    0 - 0x0
    "00000000", -- 2998 - 0xbb6  :    0 - 0x0
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "00000000", -- 3000 - 0xbb8  :    0 - 0x0
    "00000000", -- 3001 - 0xbb9  :    0 - 0x0
    "00000000", -- 3002 - 0xbba  :    0 - 0x0
    "00000000", -- 3003 - 0xbbb  :    0 - 0x0
    "00000000", -- 3004 - 0xbbc  :    0 - 0x0
    "00000000", -- 3005 - 0xbbd  :    0 - 0x0
    "00000000", -- 3006 - 0xbbe  :    0 - 0x0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Sprite 0xbc
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000000", -- 3011 - 0xbc3  :    0 - 0x0
    "00000000", -- 3012 - 0xbc4  :    0 - 0x0
    "00000000", -- 3013 - 0xbc5  :    0 - 0x0
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000000", -- 3022 - 0xbce  :    0 - 0x0
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0 -- Sprite 0xbd
    "00000000", -- 3025 - 0xbd1  :    0 - 0x0
    "00000000", -- 3026 - 0xbd2  :    0 - 0x0
    "00000000", -- 3027 - 0xbd3  :    0 - 0x0
    "00000000", -- 3028 - 0xbd4  :    0 - 0x0
    "00000000", -- 3029 - 0xbd5  :    0 - 0x0
    "00000000", -- 3030 - 0xbd6  :    0 - 0x0
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0
    "00000000", -- 3033 - 0xbd9  :    0 - 0x0
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00000000", -- 3035 - 0xbdb  :    0 - 0x0
    "00000000", -- 3036 - 0xbdc  :    0 - 0x0
    "00000000", -- 3037 - 0xbdd  :    0 - 0x0
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0 -- Sprite 0xbe
    "00000000", -- 3041 - 0xbe1  :    0 - 0x0
    "00000000", -- 3042 - 0xbe2  :    0 - 0x0
    "00000000", -- 3043 - 0xbe3  :    0 - 0x0
    "00000000", -- 3044 - 0xbe4  :    0 - 0x0
    "00000000", -- 3045 - 0xbe5  :    0 - 0x0
    "00000000", -- 3046 - 0xbe6  :    0 - 0x0
    "00000000", -- 3047 - 0xbe7  :    0 - 0x0
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0
    "00000000", -- 3049 - 0xbe9  :    0 - 0x0
    "00000000", -- 3050 - 0xbea  :    0 - 0x0
    "00000000", -- 3051 - 0xbeb  :    0 - 0x0
    "00000000", -- 3052 - 0xbec  :    0 - 0x0
    "00000000", -- 3053 - 0xbed  :    0 - 0x0
    "00000000", -- 3054 - 0xbee  :    0 - 0x0
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0 -- Sprite 0xbf
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00000000", -- 3058 - 0xbf2  :    0 - 0x0
    "00000000", -- 3059 - 0xbf3  :    0 - 0x0
    "00000000", -- 3060 - 0xbf4  :    0 - 0x0
    "00000000", -- 3061 - 0xbf5  :    0 - 0x0
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0
    "00000000", -- 3065 - 0xbf9  :    0 - 0x0
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00000000", -- 3068 - 0xbfc  :    0 - 0x0
    "00000000", -- 3069 - 0xbfd  :    0 - 0x0
    "00000000", -- 3070 - 0xbfe  :    0 - 0x0
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00000000", -- 3072 - 0xc00  :    0 - 0x0 -- Sprite 0xc0
    "00000000", -- 3073 - 0xc01  :    0 - 0x0
    "00000000", -- 3074 - 0xc02  :    0 - 0x0
    "00000000", -- 3075 - 0xc03  :    0 - 0x0
    "00000000", -- 3076 - 0xc04  :    0 - 0x0
    "00000000", -- 3077 - 0xc05  :    0 - 0x0
    "00000000", -- 3078 - 0xc06  :    0 - 0x0
    "00000000", -- 3079 - 0xc07  :    0 - 0x0
    "00000000", -- 3080 - 0xc08  :    0 - 0x0
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "00000000", -- 3083 - 0xc0b  :    0 - 0x0
    "00000000", -- 3084 - 0xc0c  :    0 - 0x0
    "00000000", -- 3085 - 0xc0d  :    0 - 0x0
    "00000000", -- 3086 - 0xc0e  :    0 - 0x0
    "00000000", -- 3087 - 0xc0f  :    0 - 0x0
    "00000000", -- 3088 - 0xc10  :    0 - 0x0 -- Sprite 0xc1
    "00000000", -- 3089 - 0xc11  :    0 - 0x0
    "00000000", -- 3090 - 0xc12  :    0 - 0x0
    "00000000", -- 3091 - 0xc13  :    0 - 0x0
    "00000000", -- 3092 - 0xc14  :    0 - 0x0
    "00000000", -- 3093 - 0xc15  :    0 - 0x0
    "00000000", -- 3094 - 0xc16  :    0 - 0x0
    "00000000", -- 3095 - 0xc17  :    0 - 0x0
    "00000000", -- 3096 - 0xc18  :    0 - 0x0
    "00000000", -- 3097 - 0xc19  :    0 - 0x0
    "00000000", -- 3098 - 0xc1a  :    0 - 0x0
    "00000000", -- 3099 - 0xc1b  :    0 - 0x0
    "00000000", -- 3100 - 0xc1c  :    0 - 0x0
    "00000000", -- 3101 - 0xc1d  :    0 - 0x0
    "00000000", -- 3102 - 0xc1e  :    0 - 0x0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00000000", -- 3104 - 0xc20  :    0 - 0x0 -- Sprite 0xc2
    "00000000", -- 3105 - 0xc21  :    0 - 0x0
    "00000000", -- 3106 - 0xc22  :    0 - 0x0
    "00000000", -- 3107 - 0xc23  :    0 - 0x0
    "00000000", -- 3108 - 0xc24  :    0 - 0x0
    "00000000", -- 3109 - 0xc25  :    0 - 0x0
    "00000000", -- 3110 - 0xc26  :    0 - 0x0
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "00000000", -- 3115 - 0xc2b  :    0 - 0x0
    "00000000", -- 3116 - 0xc2c  :    0 - 0x0
    "00000000", -- 3117 - 0xc2d  :    0 - 0x0
    "00000000", -- 3118 - 0xc2e  :    0 - 0x0
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "00000000", -- 3120 - 0xc30  :    0 - 0x0 -- Sprite 0xc3
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "00000000", -- 3122 - 0xc32  :    0 - 0x0
    "00000000", -- 3123 - 0xc33  :    0 - 0x0
    "00000000", -- 3124 - 0xc34  :    0 - 0x0
    "00000000", -- 3125 - 0xc35  :    0 - 0x0
    "00000000", -- 3126 - 0xc36  :    0 - 0x0
    "00000000", -- 3127 - 0xc37  :    0 - 0x0
    "00000000", -- 3128 - 0xc38  :    0 - 0x0
    "00000000", -- 3129 - 0xc39  :    0 - 0x0
    "00000000", -- 3130 - 0xc3a  :    0 - 0x0
    "00000000", -- 3131 - 0xc3b  :    0 - 0x0
    "00000000", -- 3132 - 0xc3c  :    0 - 0x0
    "00000000", -- 3133 - 0xc3d  :    0 - 0x0
    "00000000", -- 3134 - 0xc3e  :    0 - 0x0
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 3137 - 0xc41  :    0 - 0x0
    "00000000", -- 3138 - 0xc42  :    0 - 0x0
    "00000000", -- 3139 - 0xc43  :    0 - 0x0
    "00000000", -- 3140 - 0xc44  :    0 - 0x0
    "00000000", -- 3141 - 0xc45  :    0 - 0x0
    "00000000", -- 3142 - 0xc46  :    0 - 0x0
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00000000", -- 3144 - 0xc48  :    0 - 0x0
    "00000000", -- 3145 - 0xc49  :    0 - 0x0
    "00000000", -- 3146 - 0xc4a  :    0 - 0x0
    "00000000", -- 3147 - 0xc4b  :    0 - 0x0
    "00000000", -- 3148 - 0xc4c  :    0 - 0x0
    "00000000", -- 3149 - 0xc4d  :    0 - 0x0
    "00000000", -- 3150 - 0xc4e  :    0 - 0x0
    "00000000", -- 3151 - 0xc4f  :    0 - 0x0
    "00000000", -- 3152 - 0xc50  :    0 - 0x0 -- Sprite 0xc5
    "00000000", -- 3153 - 0xc51  :    0 - 0x0
    "00000000", -- 3154 - 0xc52  :    0 - 0x0
    "00000000", -- 3155 - 0xc53  :    0 - 0x0
    "00000000", -- 3156 - 0xc54  :    0 - 0x0
    "00000000", -- 3157 - 0xc55  :    0 - 0x0
    "00000000", -- 3158 - 0xc56  :    0 - 0x0
    "00000000", -- 3159 - 0xc57  :    0 - 0x0
    "00000000", -- 3160 - 0xc58  :    0 - 0x0
    "00000000", -- 3161 - 0xc59  :    0 - 0x0
    "00000000", -- 3162 - 0xc5a  :    0 - 0x0
    "00000000", -- 3163 - 0xc5b  :    0 - 0x0
    "00000000", -- 3164 - 0xc5c  :    0 - 0x0
    "00000000", -- 3165 - 0xc5d  :    0 - 0x0
    "00000000", -- 3166 - 0xc5e  :    0 - 0x0
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "00000000", -- 3168 - 0xc60  :    0 - 0x0 -- Sprite 0xc6
    "00000000", -- 3169 - 0xc61  :    0 - 0x0
    "00000000", -- 3170 - 0xc62  :    0 - 0x0
    "00000000", -- 3171 - 0xc63  :    0 - 0x0
    "00000000", -- 3172 - 0xc64  :    0 - 0x0
    "00000000", -- 3173 - 0xc65  :    0 - 0x0
    "00000000", -- 3174 - 0xc66  :    0 - 0x0
    "00000000", -- 3175 - 0xc67  :    0 - 0x0
    "00000000", -- 3176 - 0xc68  :    0 - 0x0
    "00000000", -- 3177 - 0xc69  :    0 - 0x0
    "00000000", -- 3178 - 0xc6a  :    0 - 0x0
    "00000000", -- 3179 - 0xc6b  :    0 - 0x0
    "00000000", -- 3180 - 0xc6c  :    0 - 0x0
    "00000000", -- 3181 - 0xc6d  :    0 - 0x0
    "00000000", -- 3182 - 0xc6e  :    0 - 0x0
    "00000000", -- 3183 - 0xc6f  :    0 - 0x0
    "00000000", -- 3184 - 0xc70  :    0 - 0x0 -- Sprite 0xc7
    "00000000", -- 3185 - 0xc71  :    0 - 0x0
    "00000000", -- 3186 - 0xc72  :    0 - 0x0
    "00000000", -- 3187 - 0xc73  :    0 - 0x0
    "00000000", -- 3188 - 0xc74  :    0 - 0x0
    "00000000", -- 3189 - 0xc75  :    0 - 0x0
    "00000000", -- 3190 - 0xc76  :    0 - 0x0
    "00000000", -- 3191 - 0xc77  :    0 - 0x0
    "00000000", -- 3192 - 0xc78  :    0 - 0x0
    "00000000", -- 3193 - 0xc79  :    0 - 0x0
    "00000000", -- 3194 - 0xc7a  :    0 - 0x0
    "00000000", -- 3195 - 0xc7b  :    0 - 0x0
    "00000000", -- 3196 - 0xc7c  :    0 - 0x0
    "00000000", -- 3197 - 0xc7d  :    0 - 0x0
    "00000000", -- 3198 - 0xc7e  :    0 - 0x0
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Sprite 0xc8
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000000", -- 3204 - 0xc84  :    0 - 0x0
    "00000000", -- 3205 - 0xc85  :    0 - 0x0
    "00000000", -- 3206 - 0xc86  :    0 - 0x0
    "00000000", -- 3207 - 0xc87  :    0 - 0x0
    "00000000", -- 3208 - 0xc88  :    0 - 0x0
    "00000000", -- 3209 - 0xc89  :    0 - 0x0
    "00000000", -- 3210 - 0xc8a  :    0 - 0x0
    "00000000", -- 3211 - 0xc8b  :    0 - 0x0
    "00000000", -- 3212 - 0xc8c  :    0 - 0x0
    "00000000", -- 3213 - 0xc8d  :    0 - 0x0
    "00000000", -- 3214 - 0xc8e  :    0 - 0x0
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00000000", -- 3216 - 0xc90  :    0 - 0x0 -- Sprite 0xc9
    "00000000", -- 3217 - 0xc91  :    0 - 0x0
    "00000000", -- 3218 - 0xc92  :    0 - 0x0
    "00000000", -- 3219 - 0xc93  :    0 - 0x0
    "00000000", -- 3220 - 0xc94  :    0 - 0x0
    "00000000", -- 3221 - 0xc95  :    0 - 0x0
    "00000000", -- 3222 - 0xc96  :    0 - 0x0
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "00000000", -- 3224 - 0xc98  :    0 - 0x0
    "00000000", -- 3225 - 0xc99  :    0 - 0x0
    "00000000", -- 3226 - 0xc9a  :    0 - 0x0
    "00000000", -- 3227 - 0xc9b  :    0 - 0x0
    "00000000", -- 3228 - 0xc9c  :    0 - 0x0
    "00000000", -- 3229 - 0xc9d  :    0 - 0x0
    "00000000", -- 3230 - 0xc9e  :    0 - 0x0
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00000000", -- 3232 - 0xca0  :    0 - 0x0 -- Sprite 0xca
    "00000000", -- 3233 - 0xca1  :    0 - 0x0
    "00000000", -- 3234 - 0xca2  :    0 - 0x0
    "00000000", -- 3235 - 0xca3  :    0 - 0x0
    "00000000", -- 3236 - 0xca4  :    0 - 0x0
    "00000000", -- 3237 - 0xca5  :    0 - 0x0
    "00000000", -- 3238 - 0xca6  :    0 - 0x0
    "00000000", -- 3239 - 0xca7  :    0 - 0x0
    "00000000", -- 3240 - 0xca8  :    0 - 0x0
    "00000000", -- 3241 - 0xca9  :    0 - 0x0
    "00000000", -- 3242 - 0xcaa  :    0 - 0x0
    "00000000", -- 3243 - 0xcab  :    0 - 0x0
    "00000000", -- 3244 - 0xcac  :    0 - 0x0
    "00000000", -- 3245 - 0xcad  :    0 - 0x0
    "00000000", -- 3246 - 0xcae  :    0 - 0x0
    "00000000", -- 3247 - 0xcaf  :    0 - 0x0
    "00000000", -- 3248 - 0xcb0  :    0 - 0x0 -- Sprite 0xcb
    "00000000", -- 3249 - 0xcb1  :    0 - 0x0
    "00000000", -- 3250 - 0xcb2  :    0 - 0x0
    "00000000", -- 3251 - 0xcb3  :    0 - 0x0
    "00000000", -- 3252 - 0xcb4  :    0 - 0x0
    "00000000", -- 3253 - 0xcb5  :    0 - 0x0
    "00000000", -- 3254 - 0xcb6  :    0 - 0x0
    "00000000", -- 3255 - 0xcb7  :    0 - 0x0
    "00000000", -- 3256 - 0xcb8  :    0 - 0x0
    "00000000", -- 3257 - 0xcb9  :    0 - 0x0
    "00000000", -- 3258 - 0xcba  :    0 - 0x0
    "00000000", -- 3259 - 0xcbb  :    0 - 0x0
    "00000000", -- 3260 - 0xcbc  :    0 - 0x0
    "00000000", -- 3261 - 0xcbd  :    0 - 0x0
    "00000000", -- 3262 - 0xcbe  :    0 - 0x0
    "00000000", -- 3263 - 0xcbf  :    0 - 0x0
    "00000000", -- 3264 - 0xcc0  :    0 - 0x0 -- Sprite 0xcc
    "00000000", -- 3265 - 0xcc1  :    0 - 0x0
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "00000000", -- 3267 - 0xcc3  :    0 - 0x0
    "00000000", -- 3268 - 0xcc4  :    0 - 0x0
    "00000000", -- 3269 - 0xcc5  :    0 - 0x0
    "00000000", -- 3270 - 0xcc6  :    0 - 0x0
    "00000000", -- 3271 - 0xcc7  :    0 - 0x0
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000000", -- 3274 - 0xcca  :    0 - 0x0
    "00000000", -- 3275 - 0xccb  :    0 - 0x0
    "00000000", -- 3276 - 0xccc  :    0 - 0x0
    "00000000", -- 3277 - 0xccd  :    0 - 0x0
    "00000000", -- 3278 - 0xcce  :    0 - 0x0
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00000000", -- 3282 - 0xcd2  :    0 - 0x0
    "00000000", -- 3283 - 0xcd3  :    0 - 0x0
    "00000000", -- 3284 - 0xcd4  :    0 - 0x0
    "00000000", -- 3285 - 0xcd5  :    0 - 0x0
    "00000000", -- 3286 - 0xcd6  :    0 - 0x0
    "00000000", -- 3287 - 0xcd7  :    0 - 0x0
    "00000000", -- 3288 - 0xcd8  :    0 - 0x0
    "00000000", -- 3289 - 0xcd9  :    0 - 0x0
    "00000000", -- 3290 - 0xcda  :    0 - 0x0
    "00000000", -- 3291 - 0xcdb  :    0 - 0x0
    "00000000", -- 3292 - 0xcdc  :    0 - 0x0
    "00000000", -- 3293 - 0xcdd  :    0 - 0x0
    "00000000", -- 3294 - 0xcde  :    0 - 0x0
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "00000000", -- 3299 - 0xce3  :    0 - 0x0
    "00000000", -- 3300 - 0xce4  :    0 - 0x0
    "00000000", -- 3301 - 0xce5  :    0 - 0x0
    "00000000", -- 3302 - 0xce6  :    0 - 0x0
    "00000000", -- 3303 - 0xce7  :    0 - 0x0
    "00000000", -- 3304 - 0xce8  :    0 - 0x0
    "00000000", -- 3305 - 0xce9  :    0 - 0x0
    "00000000", -- 3306 - 0xcea  :    0 - 0x0
    "00000000", -- 3307 - 0xceb  :    0 - 0x0
    "00000000", -- 3308 - 0xcec  :    0 - 0x0
    "00000000", -- 3309 - 0xced  :    0 - 0x0
    "00000000", -- 3310 - 0xcee  :    0 - 0x0
    "00000000", -- 3311 - 0xcef  :    0 - 0x0
    "00000000", -- 3312 - 0xcf0  :    0 - 0x0 -- Sprite 0xcf
    "00000000", -- 3313 - 0xcf1  :    0 - 0x0
    "00000000", -- 3314 - 0xcf2  :    0 - 0x0
    "00000000", -- 3315 - 0xcf3  :    0 - 0x0
    "00000000", -- 3316 - 0xcf4  :    0 - 0x0
    "00000000", -- 3317 - 0xcf5  :    0 - 0x0
    "00000000", -- 3318 - 0xcf6  :    0 - 0x0
    "00000000", -- 3319 - 0xcf7  :    0 - 0x0
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0
    "00000000", -- 3321 - 0xcf9  :    0 - 0x0
    "00000000", -- 3322 - 0xcfa  :    0 - 0x0
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00000000", -- 3328 - 0xd00  :    0 - 0x0 -- Sprite 0xd0
    "00000000", -- 3329 - 0xd01  :    0 - 0x0
    "00000000", -- 3330 - 0xd02  :    0 - 0x0
    "00000000", -- 3331 - 0xd03  :    0 - 0x0
    "00000000", -- 3332 - 0xd04  :    0 - 0x0
    "00000000", -- 3333 - 0xd05  :    0 - 0x0
    "00000000", -- 3334 - 0xd06  :    0 - 0x0
    "00000000", -- 3335 - 0xd07  :    0 - 0x0
    "00000000", -- 3336 - 0xd08  :    0 - 0x0
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "00000000", -- 3338 - 0xd0a  :    0 - 0x0
    "00000000", -- 3339 - 0xd0b  :    0 - 0x0
    "00000000", -- 3340 - 0xd0c  :    0 - 0x0
    "00000000", -- 3341 - 0xd0d  :    0 - 0x0
    "00000000", -- 3342 - 0xd0e  :    0 - 0x0
    "00000000", -- 3343 - 0xd0f  :    0 - 0x0
    "00000000", -- 3344 - 0xd10  :    0 - 0x0 -- Sprite 0xd1
    "00000000", -- 3345 - 0xd11  :    0 - 0x0
    "00000000", -- 3346 - 0xd12  :    0 - 0x0
    "00000000", -- 3347 - 0xd13  :    0 - 0x0
    "00000000", -- 3348 - 0xd14  :    0 - 0x0
    "00000000", -- 3349 - 0xd15  :    0 - 0x0
    "00000000", -- 3350 - 0xd16  :    0 - 0x0
    "00000000", -- 3351 - 0xd17  :    0 - 0x0
    "00000000", -- 3352 - 0xd18  :    0 - 0x0
    "00000000", -- 3353 - 0xd19  :    0 - 0x0
    "00000000", -- 3354 - 0xd1a  :    0 - 0x0
    "00000000", -- 3355 - 0xd1b  :    0 - 0x0
    "00000000", -- 3356 - 0xd1c  :    0 - 0x0
    "00000000", -- 3357 - 0xd1d  :    0 - 0x0
    "00000000", -- 3358 - 0xd1e  :    0 - 0x0
    "00000000", -- 3359 - 0xd1f  :    0 - 0x0
    "00000000", -- 3360 - 0xd20  :    0 - 0x0 -- Sprite 0xd2
    "00000000", -- 3361 - 0xd21  :    0 - 0x0
    "00000000", -- 3362 - 0xd22  :    0 - 0x0
    "00000000", -- 3363 - 0xd23  :    0 - 0x0
    "00000000", -- 3364 - 0xd24  :    0 - 0x0
    "00000000", -- 3365 - 0xd25  :    0 - 0x0
    "00000000", -- 3366 - 0xd26  :    0 - 0x0
    "00000000", -- 3367 - 0xd27  :    0 - 0x0
    "00000000", -- 3368 - 0xd28  :    0 - 0x0
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "00000000", -- 3370 - 0xd2a  :    0 - 0x0
    "00000000", -- 3371 - 0xd2b  :    0 - 0x0
    "00000000", -- 3372 - 0xd2c  :    0 - 0x0
    "00000000", -- 3373 - 0xd2d  :    0 - 0x0
    "00000000", -- 3374 - 0xd2e  :    0 - 0x0
    "00000000", -- 3375 - 0xd2f  :    0 - 0x0
    "00000000", -- 3376 - 0xd30  :    0 - 0x0 -- Sprite 0xd3
    "00000000", -- 3377 - 0xd31  :    0 - 0x0
    "00000000", -- 3378 - 0xd32  :    0 - 0x0
    "00000000", -- 3379 - 0xd33  :    0 - 0x0
    "00000000", -- 3380 - 0xd34  :    0 - 0x0
    "00000000", -- 3381 - 0xd35  :    0 - 0x0
    "00000000", -- 3382 - 0xd36  :    0 - 0x0
    "00000000", -- 3383 - 0xd37  :    0 - 0x0
    "00000000", -- 3384 - 0xd38  :    0 - 0x0
    "00000000", -- 3385 - 0xd39  :    0 - 0x0
    "00000000", -- 3386 - 0xd3a  :    0 - 0x0
    "00000000", -- 3387 - 0xd3b  :    0 - 0x0
    "00000000", -- 3388 - 0xd3c  :    0 - 0x0
    "00000000", -- 3389 - 0xd3d  :    0 - 0x0
    "00000000", -- 3390 - 0xd3e  :    0 - 0x0
    "00000000", -- 3391 - 0xd3f  :    0 - 0x0
    "00000000", -- 3392 - 0xd40  :    0 - 0x0 -- Sprite 0xd4
    "00000000", -- 3393 - 0xd41  :    0 - 0x0
    "00000000", -- 3394 - 0xd42  :    0 - 0x0
    "00000000", -- 3395 - 0xd43  :    0 - 0x0
    "00000000", -- 3396 - 0xd44  :    0 - 0x0
    "00000000", -- 3397 - 0xd45  :    0 - 0x0
    "00000000", -- 3398 - 0xd46  :    0 - 0x0
    "00000000", -- 3399 - 0xd47  :    0 - 0x0
    "00000000", -- 3400 - 0xd48  :    0 - 0x0
    "00000000", -- 3401 - 0xd49  :    0 - 0x0
    "00000000", -- 3402 - 0xd4a  :    0 - 0x0
    "00000000", -- 3403 - 0xd4b  :    0 - 0x0
    "00000000", -- 3404 - 0xd4c  :    0 - 0x0
    "00000000", -- 3405 - 0xd4d  :    0 - 0x0
    "00000000", -- 3406 - 0xd4e  :    0 - 0x0
    "00000000", -- 3407 - 0xd4f  :    0 - 0x0
    "00000000", -- 3408 - 0xd50  :    0 - 0x0 -- Sprite 0xd5
    "00000000", -- 3409 - 0xd51  :    0 - 0x0
    "00000000", -- 3410 - 0xd52  :    0 - 0x0
    "00000000", -- 3411 - 0xd53  :    0 - 0x0
    "00000000", -- 3412 - 0xd54  :    0 - 0x0
    "00000000", -- 3413 - 0xd55  :    0 - 0x0
    "00000000", -- 3414 - 0xd56  :    0 - 0x0
    "00000000", -- 3415 - 0xd57  :    0 - 0x0
    "00000000", -- 3416 - 0xd58  :    0 - 0x0
    "00000000", -- 3417 - 0xd59  :    0 - 0x0
    "00000000", -- 3418 - 0xd5a  :    0 - 0x0
    "00000000", -- 3419 - 0xd5b  :    0 - 0x0
    "00000000", -- 3420 - 0xd5c  :    0 - 0x0
    "00000000", -- 3421 - 0xd5d  :    0 - 0x0
    "00000000", -- 3422 - 0xd5e  :    0 - 0x0
    "00000000", -- 3423 - 0xd5f  :    0 - 0x0
    "00000000", -- 3424 - 0xd60  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 3425 - 0xd61  :    0 - 0x0
    "00000000", -- 3426 - 0xd62  :    0 - 0x0
    "00000000", -- 3427 - 0xd63  :    0 - 0x0
    "00000000", -- 3428 - 0xd64  :    0 - 0x0
    "00000000", -- 3429 - 0xd65  :    0 - 0x0
    "00000000", -- 3430 - 0xd66  :    0 - 0x0
    "00000000", -- 3431 - 0xd67  :    0 - 0x0
    "00000000", -- 3432 - 0xd68  :    0 - 0x0
    "00000000", -- 3433 - 0xd69  :    0 - 0x0
    "00000000", -- 3434 - 0xd6a  :    0 - 0x0
    "00000000", -- 3435 - 0xd6b  :    0 - 0x0
    "00000000", -- 3436 - 0xd6c  :    0 - 0x0
    "00000000", -- 3437 - 0xd6d  :    0 - 0x0
    "00000000", -- 3438 - 0xd6e  :    0 - 0x0
    "00000000", -- 3439 - 0xd6f  :    0 - 0x0
    "00000000", -- 3440 - 0xd70  :    0 - 0x0 -- Sprite 0xd7
    "00000000", -- 3441 - 0xd71  :    0 - 0x0
    "00000000", -- 3442 - 0xd72  :    0 - 0x0
    "00000000", -- 3443 - 0xd73  :    0 - 0x0
    "00000000", -- 3444 - 0xd74  :    0 - 0x0
    "00000000", -- 3445 - 0xd75  :    0 - 0x0
    "00000000", -- 3446 - 0xd76  :    0 - 0x0
    "00000000", -- 3447 - 0xd77  :    0 - 0x0
    "00000000", -- 3448 - 0xd78  :    0 - 0x0
    "00000000", -- 3449 - 0xd79  :    0 - 0x0
    "00000000", -- 3450 - 0xd7a  :    0 - 0x0
    "00000000", -- 3451 - 0xd7b  :    0 - 0x0
    "00000000", -- 3452 - 0xd7c  :    0 - 0x0
    "00000000", -- 3453 - 0xd7d  :    0 - 0x0
    "00000000", -- 3454 - 0xd7e  :    0 - 0x0
    "00000000", -- 3455 - 0xd7f  :    0 - 0x0
    "00000000", -- 3456 - 0xd80  :    0 - 0x0 -- Sprite 0xd8
    "00000000", -- 3457 - 0xd81  :    0 - 0x0
    "00000000", -- 3458 - 0xd82  :    0 - 0x0
    "00000000", -- 3459 - 0xd83  :    0 - 0x0
    "00000000", -- 3460 - 0xd84  :    0 - 0x0
    "00000000", -- 3461 - 0xd85  :    0 - 0x0
    "00000000", -- 3462 - 0xd86  :    0 - 0x0
    "00000000", -- 3463 - 0xd87  :    0 - 0x0
    "00000000", -- 3464 - 0xd88  :    0 - 0x0
    "00000000", -- 3465 - 0xd89  :    0 - 0x0
    "00000000", -- 3466 - 0xd8a  :    0 - 0x0
    "00000000", -- 3467 - 0xd8b  :    0 - 0x0
    "00000000", -- 3468 - 0xd8c  :    0 - 0x0
    "00000000", -- 3469 - 0xd8d  :    0 - 0x0
    "00000000", -- 3470 - 0xd8e  :    0 - 0x0
    "00000000", -- 3471 - 0xd8f  :    0 - 0x0
    "00000000", -- 3472 - 0xd90  :    0 - 0x0 -- Sprite 0xd9
    "00000000", -- 3473 - 0xd91  :    0 - 0x0
    "00000000", -- 3474 - 0xd92  :    0 - 0x0
    "00000000", -- 3475 - 0xd93  :    0 - 0x0
    "00000000", -- 3476 - 0xd94  :    0 - 0x0
    "00000000", -- 3477 - 0xd95  :    0 - 0x0
    "00000000", -- 3478 - 0xd96  :    0 - 0x0
    "00000000", -- 3479 - 0xd97  :    0 - 0x0
    "00000000", -- 3480 - 0xd98  :    0 - 0x0
    "00000000", -- 3481 - 0xd99  :    0 - 0x0
    "00000000", -- 3482 - 0xd9a  :    0 - 0x0
    "00000000", -- 3483 - 0xd9b  :    0 - 0x0
    "00000000", -- 3484 - 0xd9c  :    0 - 0x0
    "00000000", -- 3485 - 0xd9d  :    0 - 0x0
    "00000000", -- 3486 - 0xd9e  :    0 - 0x0
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "00000000", -- 3488 - 0xda0  :    0 - 0x0 -- Sprite 0xda
    "00000000", -- 3489 - 0xda1  :    0 - 0x0
    "00000000", -- 3490 - 0xda2  :    0 - 0x0
    "00000000", -- 3491 - 0xda3  :    0 - 0x0
    "00000000", -- 3492 - 0xda4  :    0 - 0x0
    "00000000", -- 3493 - 0xda5  :    0 - 0x0
    "00000000", -- 3494 - 0xda6  :    0 - 0x0
    "00000000", -- 3495 - 0xda7  :    0 - 0x0
    "00000000", -- 3496 - 0xda8  :    0 - 0x0
    "00000000", -- 3497 - 0xda9  :    0 - 0x0
    "00000000", -- 3498 - 0xdaa  :    0 - 0x0
    "00000000", -- 3499 - 0xdab  :    0 - 0x0
    "00000000", -- 3500 - 0xdac  :    0 - 0x0
    "00000000", -- 3501 - 0xdad  :    0 - 0x0
    "00000000", -- 3502 - 0xdae  :    0 - 0x0
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00000000", -- 3504 - 0xdb0  :    0 - 0x0 -- Sprite 0xdb
    "00000000", -- 3505 - 0xdb1  :    0 - 0x0
    "00000000", -- 3506 - 0xdb2  :    0 - 0x0
    "00000000", -- 3507 - 0xdb3  :    0 - 0x0
    "00000000", -- 3508 - 0xdb4  :    0 - 0x0
    "00000000", -- 3509 - 0xdb5  :    0 - 0x0
    "00000000", -- 3510 - 0xdb6  :    0 - 0x0
    "00000000", -- 3511 - 0xdb7  :    0 - 0x0
    "00000000", -- 3512 - 0xdb8  :    0 - 0x0
    "00000000", -- 3513 - 0xdb9  :    0 - 0x0
    "00000000", -- 3514 - 0xdba  :    0 - 0x0
    "00000000", -- 3515 - 0xdbb  :    0 - 0x0
    "00000000", -- 3516 - 0xdbc  :    0 - 0x0
    "00000000", -- 3517 - 0xdbd  :    0 - 0x0
    "00000000", -- 3518 - 0xdbe  :    0 - 0x0
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0 -- Sprite 0xdc
    "00000000", -- 3521 - 0xdc1  :    0 - 0x0
    "00000000", -- 3522 - 0xdc2  :    0 - 0x0
    "00000000", -- 3523 - 0xdc3  :    0 - 0x0
    "00000000", -- 3524 - 0xdc4  :    0 - 0x0
    "00000000", -- 3525 - 0xdc5  :    0 - 0x0
    "00000000", -- 3526 - 0xdc6  :    0 - 0x0
    "00000000", -- 3527 - 0xdc7  :    0 - 0x0
    "00000000", -- 3528 - 0xdc8  :    0 - 0x0
    "00000000", -- 3529 - 0xdc9  :    0 - 0x0
    "00000000", -- 3530 - 0xdca  :    0 - 0x0
    "00000000", -- 3531 - 0xdcb  :    0 - 0x0
    "00000000", -- 3532 - 0xdcc  :    0 - 0x0
    "00000000", -- 3533 - 0xdcd  :    0 - 0x0
    "00000000", -- 3534 - 0xdce  :    0 - 0x0
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "00000000", -- 3536 - 0xdd0  :    0 - 0x0 -- Sprite 0xdd
    "00000000", -- 3537 - 0xdd1  :    0 - 0x0
    "00000000", -- 3538 - 0xdd2  :    0 - 0x0
    "00000000", -- 3539 - 0xdd3  :    0 - 0x0
    "00000000", -- 3540 - 0xdd4  :    0 - 0x0
    "00000000", -- 3541 - 0xdd5  :    0 - 0x0
    "00000000", -- 3542 - 0xdd6  :    0 - 0x0
    "00000000", -- 3543 - 0xdd7  :    0 - 0x0
    "00000000", -- 3544 - 0xdd8  :    0 - 0x0
    "00000000", -- 3545 - 0xdd9  :    0 - 0x0
    "00000000", -- 3546 - 0xdda  :    0 - 0x0
    "00000000", -- 3547 - 0xddb  :    0 - 0x0
    "00000000", -- 3548 - 0xddc  :    0 - 0x0
    "00000000", -- 3549 - 0xddd  :    0 - 0x0
    "00000000", -- 3550 - 0xdde  :    0 - 0x0
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "00000000", -- 3552 - 0xde0  :    0 - 0x0 -- Sprite 0xde
    "00000000", -- 3553 - 0xde1  :    0 - 0x0
    "00000000", -- 3554 - 0xde2  :    0 - 0x0
    "00000000", -- 3555 - 0xde3  :    0 - 0x0
    "00000000", -- 3556 - 0xde4  :    0 - 0x0
    "00000000", -- 3557 - 0xde5  :    0 - 0x0
    "00000000", -- 3558 - 0xde6  :    0 - 0x0
    "00000000", -- 3559 - 0xde7  :    0 - 0x0
    "00000000", -- 3560 - 0xde8  :    0 - 0x0
    "00000000", -- 3561 - 0xde9  :    0 - 0x0
    "00000000", -- 3562 - 0xdea  :    0 - 0x0
    "00000000", -- 3563 - 0xdeb  :    0 - 0x0
    "00000000", -- 3564 - 0xdec  :    0 - 0x0
    "00000000", -- 3565 - 0xded  :    0 - 0x0
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "00000000", -- 3568 - 0xdf0  :    0 - 0x0 -- Sprite 0xdf
    "00000000", -- 3569 - 0xdf1  :    0 - 0x0
    "00000000", -- 3570 - 0xdf2  :    0 - 0x0
    "00000000", -- 3571 - 0xdf3  :    0 - 0x0
    "00000000", -- 3572 - 0xdf4  :    0 - 0x0
    "00000000", -- 3573 - 0xdf5  :    0 - 0x0
    "00000000", -- 3574 - 0xdf6  :    0 - 0x0
    "00000000", -- 3575 - 0xdf7  :    0 - 0x0
    "00000000", -- 3576 - 0xdf8  :    0 - 0x0
    "00000000", -- 3577 - 0xdf9  :    0 - 0x0
    "00000000", -- 3578 - 0xdfa  :    0 - 0x0
    "00000000", -- 3579 - 0xdfb  :    0 - 0x0
    "00000000", -- 3580 - 0xdfc  :    0 - 0x0
    "00000000", -- 3581 - 0xdfd  :    0 - 0x0
    "00000000", -- 3582 - 0xdfe  :    0 - 0x0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "00000000", -- 3584 - 0xe00  :    0 - 0x0 -- Sprite 0xe0
    "00000000", -- 3585 - 0xe01  :    0 - 0x0
    "00000000", -- 3586 - 0xe02  :    0 - 0x0
    "00000000", -- 3587 - 0xe03  :    0 - 0x0
    "00000000", -- 3588 - 0xe04  :    0 - 0x0
    "00000000", -- 3589 - 0xe05  :    0 - 0x0
    "00000000", -- 3590 - 0xe06  :    0 - 0x0
    "00000000", -- 3591 - 0xe07  :    0 - 0x0
    "00000000", -- 3592 - 0xe08  :    0 - 0x0
    "00000000", -- 3593 - 0xe09  :    0 - 0x0
    "00000000", -- 3594 - 0xe0a  :    0 - 0x0
    "00000000", -- 3595 - 0xe0b  :    0 - 0x0
    "00000000", -- 3596 - 0xe0c  :    0 - 0x0
    "00000000", -- 3597 - 0xe0d  :    0 - 0x0
    "00000000", -- 3598 - 0xe0e  :    0 - 0x0
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "00000000", -- 3600 - 0xe10  :    0 - 0x0 -- Sprite 0xe1
    "00000000", -- 3601 - 0xe11  :    0 - 0x0
    "00000000", -- 3602 - 0xe12  :    0 - 0x0
    "00000000", -- 3603 - 0xe13  :    0 - 0x0
    "00000000", -- 3604 - 0xe14  :    0 - 0x0
    "00000000", -- 3605 - 0xe15  :    0 - 0x0
    "00000000", -- 3606 - 0xe16  :    0 - 0x0
    "00000000", -- 3607 - 0xe17  :    0 - 0x0
    "00000000", -- 3608 - 0xe18  :    0 - 0x0
    "00000000", -- 3609 - 0xe19  :    0 - 0x0
    "00000000", -- 3610 - 0xe1a  :    0 - 0x0
    "00000000", -- 3611 - 0xe1b  :    0 - 0x0
    "00000000", -- 3612 - 0xe1c  :    0 - 0x0
    "00000000", -- 3613 - 0xe1d  :    0 - 0x0
    "00000000", -- 3614 - 0xe1e  :    0 - 0x0
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "00000000", -- 3616 - 0xe20  :    0 - 0x0 -- Sprite 0xe2
    "00000000", -- 3617 - 0xe21  :    0 - 0x0
    "00000000", -- 3618 - 0xe22  :    0 - 0x0
    "00000000", -- 3619 - 0xe23  :    0 - 0x0
    "00000000", -- 3620 - 0xe24  :    0 - 0x0
    "00000000", -- 3621 - 0xe25  :    0 - 0x0
    "00000000", -- 3622 - 0xe26  :    0 - 0x0
    "00000000", -- 3623 - 0xe27  :    0 - 0x0
    "00000000", -- 3624 - 0xe28  :    0 - 0x0
    "00000000", -- 3625 - 0xe29  :    0 - 0x0
    "00000000", -- 3626 - 0xe2a  :    0 - 0x0
    "00000000", -- 3627 - 0xe2b  :    0 - 0x0
    "00000000", -- 3628 - 0xe2c  :    0 - 0x0
    "00000000", -- 3629 - 0xe2d  :    0 - 0x0
    "00000000", -- 3630 - 0xe2e  :    0 - 0x0
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "00000000", -- 3632 - 0xe30  :    0 - 0x0 -- Sprite 0xe3
    "00000000", -- 3633 - 0xe31  :    0 - 0x0
    "00000000", -- 3634 - 0xe32  :    0 - 0x0
    "00000000", -- 3635 - 0xe33  :    0 - 0x0
    "00000000", -- 3636 - 0xe34  :    0 - 0x0
    "00000000", -- 3637 - 0xe35  :    0 - 0x0
    "00000000", -- 3638 - 0xe36  :    0 - 0x0
    "00000000", -- 3639 - 0xe37  :    0 - 0x0
    "00000000", -- 3640 - 0xe38  :    0 - 0x0
    "00000000", -- 3641 - 0xe39  :    0 - 0x0
    "00000000", -- 3642 - 0xe3a  :    0 - 0x0
    "00000000", -- 3643 - 0xe3b  :    0 - 0x0
    "00000000", -- 3644 - 0xe3c  :    0 - 0x0
    "00000000", -- 3645 - 0xe3d  :    0 - 0x0
    "00000000", -- 3646 - 0xe3e  :    0 - 0x0
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "00000000", -- 3648 - 0xe40  :    0 - 0x0 -- Sprite 0xe4
    "00000000", -- 3649 - 0xe41  :    0 - 0x0
    "00000000", -- 3650 - 0xe42  :    0 - 0x0
    "00000000", -- 3651 - 0xe43  :    0 - 0x0
    "00000000", -- 3652 - 0xe44  :    0 - 0x0
    "00000000", -- 3653 - 0xe45  :    0 - 0x0
    "00000000", -- 3654 - 0xe46  :    0 - 0x0
    "00000000", -- 3655 - 0xe47  :    0 - 0x0
    "00000000", -- 3656 - 0xe48  :    0 - 0x0
    "00000000", -- 3657 - 0xe49  :    0 - 0x0
    "00000000", -- 3658 - 0xe4a  :    0 - 0x0
    "00000000", -- 3659 - 0xe4b  :    0 - 0x0
    "00000000", -- 3660 - 0xe4c  :    0 - 0x0
    "00000000", -- 3661 - 0xe4d  :    0 - 0x0
    "00000000", -- 3662 - 0xe4e  :    0 - 0x0
    "00000000", -- 3663 - 0xe4f  :    0 - 0x0
    "00000000", -- 3664 - 0xe50  :    0 - 0x0 -- Sprite 0xe5
    "00000000", -- 3665 - 0xe51  :    0 - 0x0
    "00000000", -- 3666 - 0xe52  :    0 - 0x0
    "00000000", -- 3667 - 0xe53  :    0 - 0x0
    "00000000", -- 3668 - 0xe54  :    0 - 0x0
    "00000000", -- 3669 - 0xe55  :    0 - 0x0
    "00000000", -- 3670 - 0xe56  :    0 - 0x0
    "00000000", -- 3671 - 0xe57  :    0 - 0x0
    "00000000", -- 3672 - 0xe58  :    0 - 0x0
    "00000000", -- 3673 - 0xe59  :    0 - 0x0
    "00000000", -- 3674 - 0xe5a  :    0 - 0x0
    "00000000", -- 3675 - 0xe5b  :    0 - 0x0
    "00000000", -- 3676 - 0xe5c  :    0 - 0x0
    "00000000", -- 3677 - 0xe5d  :    0 - 0x0
    "00000000", -- 3678 - 0xe5e  :    0 - 0x0
    "00000000", -- 3679 - 0xe5f  :    0 - 0x0
    "00000000", -- 3680 - 0xe60  :    0 - 0x0 -- Sprite 0xe6
    "00000000", -- 3681 - 0xe61  :    0 - 0x0
    "00000000", -- 3682 - 0xe62  :    0 - 0x0
    "00000000", -- 3683 - 0xe63  :    0 - 0x0
    "00000000", -- 3684 - 0xe64  :    0 - 0x0
    "00000000", -- 3685 - 0xe65  :    0 - 0x0
    "00000000", -- 3686 - 0xe66  :    0 - 0x0
    "00000000", -- 3687 - 0xe67  :    0 - 0x0
    "00000000", -- 3688 - 0xe68  :    0 - 0x0
    "00000000", -- 3689 - 0xe69  :    0 - 0x0
    "00000000", -- 3690 - 0xe6a  :    0 - 0x0
    "00000000", -- 3691 - 0xe6b  :    0 - 0x0
    "00000000", -- 3692 - 0xe6c  :    0 - 0x0
    "00000000", -- 3693 - 0xe6d  :    0 - 0x0
    "00000000", -- 3694 - 0xe6e  :    0 - 0x0
    "00000000", -- 3695 - 0xe6f  :    0 - 0x0
    "00000000", -- 3696 - 0xe70  :    0 - 0x0 -- Sprite 0xe7
    "00000000", -- 3697 - 0xe71  :    0 - 0x0
    "00000000", -- 3698 - 0xe72  :    0 - 0x0
    "00000000", -- 3699 - 0xe73  :    0 - 0x0
    "00000000", -- 3700 - 0xe74  :    0 - 0x0
    "00000000", -- 3701 - 0xe75  :    0 - 0x0
    "00000000", -- 3702 - 0xe76  :    0 - 0x0
    "00000000", -- 3703 - 0xe77  :    0 - 0x0
    "00000000", -- 3704 - 0xe78  :    0 - 0x0
    "00000000", -- 3705 - 0xe79  :    0 - 0x0
    "00000000", -- 3706 - 0xe7a  :    0 - 0x0
    "00000000", -- 3707 - 0xe7b  :    0 - 0x0
    "00000000", -- 3708 - 0xe7c  :    0 - 0x0
    "00000000", -- 3709 - 0xe7d  :    0 - 0x0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "00000000", -- 3712 - 0xe80  :    0 - 0x0 -- Sprite 0xe8
    "00000000", -- 3713 - 0xe81  :    0 - 0x0
    "00000000", -- 3714 - 0xe82  :    0 - 0x0
    "00000000", -- 3715 - 0xe83  :    0 - 0x0
    "00000000", -- 3716 - 0xe84  :    0 - 0x0
    "00000000", -- 3717 - 0xe85  :    0 - 0x0
    "00000000", -- 3718 - 0xe86  :    0 - 0x0
    "00000000", -- 3719 - 0xe87  :    0 - 0x0
    "00000000", -- 3720 - 0xe88  :    0 - 0x0
    "00000000", -- 3721 - 0xe89  :    0 - 0x0
    "00000000", -- 3722 - 0xe8a  :    0 - 0x0
    "00000000", -- 3723 - 0xe8b  :    0 - 0x0
    "00000000", -- 3724 - 0xe8c  :    0 - 0x0
    "00000000", -- 3725 - 0xe8d  :    0 - 0x0
    "00000000", -- 3726 - 0xe8e  :    0 - 0x0
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "00000000", -- 3728 - 0xe90  :    0 - 0x0 -- Sprite 0xe9
    "00000000", -- 3729 - 0xe91  :    0 - 0x0
    "00000000", -- 3730 - 0xe92  :    0 - 0x0
    "00000000", -- 3731 - 0xe93  :    0 - 0x0
    "00000000", -- 3732 - 0xe94  :    0 - 0x0
    "00000000", -- 3733 - 0xe95  :    0 - 0x0
    "00000000", -- 3734 - 0xe96  :    0 - 0x0
    "00000000", -- 3735 - 0xe97  :    0 - 0x0
    "00000000", -- 3736 - 0xe98  :    0 - 0x0
    "00000000", -- 3737 - 0xe99  :    0 - 0x0
    "00000000", -- 3738 - 0xe9a  :    0 - 0x0
    "00000000", -- 3739 - 0xe9b  :    0 - 0x0
    "00000000", -- 3740 - 0xe9c  :    0 - 0x0
    "00000000", -- 3741 - 0xe9d  :    0 - 0x0
    "00000000", -- 3742 - 0xe9e  :    0 - 0x0
    "00000000", -- 3743 - 0xe9f  :    0 - 0x0
    "00000000", -- 3744 - 0xea0  :    0 - 0x0 -- Sprite 0xea
    "00000000", -- 3745 - 0xea1  :    0 - 0x0
    "00000000", -- 3746 - 0xea2  :    0 - 0x0
    "00000000", -- 3747 - 0xea3  :    0 - 0x0
    "00000000", -- 3748 - 0xea4  :    0 - 0x0
    "00000000", -- 3749 - 0xea5  :    0 - 0x0
    "00000000", -- 3750 - 0xea6  :    0 - 0x0
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "00000000", -- 3752 - 0xea8  :    0 - 0x0
    "00000000", -- 3753 - 0xea9  :    0 - 0x0
    "00000000", -- 3754 - 0xeaa  :    0 - 0x0
    "00000000", -- 3755 - 0xeab  :    0 - 0x0
    "00000000", -- 3756 - 0xeac  :    0 - 0x0
    "00000000", -- 3757 - 0xead  :    0 - 0x0
    "00000000", -- 3758 - 0xeae  :    0 - 0x0
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0 -- Sprite 0xeb
    "00000000", -- 3761 - 0xeb1  :    0 - 0x0
    "00000000", -- 3762 - 0xeb2  :    0 - 0x0
    "00000000", -- 3763 - 0xeb3  :    0 - 0x0
    "00000000", -- 3764 - 0xeb4  :    0 - 0x0
    "00000000", -- 3765 - 0xeb5  :    0 - 0x0
    "00000000", -- 3766 - 0xeb6  :    0 - 0x0
    "00000000", -- 3767 - 0xeb7  :    0 - 0x0
    "00000000", -- 3768 - 0xeb8  :    0 - 0x0
    "00000000", -- 3769 - 0xeb9  :    0 - 0x0
    "00000000", -- 3770 - 0xeba  :    0 - 0x0
    "00000000", -- 3771 - 0xebb  :    0 - 0x0
    "00000000", -- 3772 - 0xebc  :    0 - 0x0
    "00000000", -- 3773 - 0xebd  :    0 - 0x0
    "00000000", -- 3774 - 0xebe  :    0 - 0x0
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Sprite 0xec
    "00000000", -- 3777 - 0xec1  :    0 - 0x0
    "00000000", -- 3778 - 0xec2  :    0 - 0x0
    "00000000", -- 3779 - 0xec3  :    0 - 0x0
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00000000", -- 3781 - 0xec5  :    0 - 0x0
    "00000000", -- 3782 - 0xec6  :    0 - 0x0
    "00000000", -- 3783 - 0xec7  :    0 - 0x0
    "00000000", -- 3784 - 0xec8  :    0 - 0x0
    "00000000", -- 3785 - 0xec9  :    0 - 0x0
    "00000000", -- 3786 - 0xeca  :    0 - 0x0
    "00000000", -- 3787 - 0xecb  :    0 - 0x0
    "00000000", -- 3788 - 0xecc  :    0 - 0x0
    "00000000", -- 3789 - 0xecd  :    0 - 0x0
    "00000000", -- 3790 - 0xece  :    0 - 0x0
    "00000000", -- 3791 - 0xecf  :    0 - 0x0
    "00000000", -- 3792 - 0xed0  :    0 - 0x0 -- Sprite 0xed
    "00000000", -- 3793 - 0xed1  :    0 - 0x0
    "00000000", -- 3794 - 0xed2  :    0 - 0x0
    "00000000", -- 3795 - 0xed3  :    0 - 0x0
    "00000000", -- 3796 - 0xed4  :    0 - 0x0
    "00000000", -- 3797 - 0xed5  :    0 - 0x0
    "00000000", -- 3798 - 0xed6  :    0 - 0x0
    "00000000", -- 3799 - 0xed7  :    0 - 0x0
    "00000000", -- 3800 - 0xed8  :    0 - 0x0
    "00000000", -- 3801 - 0xed9  :    0 - 0x0
    "00000000", -- 3802 - 0xeda  :    0 - 0x0
    "00000000", -- 3803 - 0xedb  :    0 - 0x0
    "00000000", -- 3804 - 0xedc  :    0 - 0x0
    "00000000", -- 3805 - 0xedd  :    0 - 0x0
    "00000000", -- 3806 - 0xede  :    0 - 0x0
    "00000000", -- 3807 - 0xedf  :    0 - 0x0
    "00000000", -- 3808 - 0xee0  :    0 - 0x0 -- Sprite 0xee
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000000", -- 3811 - 0xee3  :    0 - 0x0
    "00000000", -- 3812 - 0xee4  :    0 - 0x0
    "00000000", -- 3813 - 0xee5  :    0 - 0x0
    "00000000", -- 3814 - 0xee6  :    0 - 0x0
    "00000000", -- 3815 - 0xee7  :    0 - 0x0
    "00000000", -- 3816 - 0xee8  :    0 - 0x0
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "00000000", -- 3818 - 0xeea  :    0 - 0x0
    "00000000", -- 3819 - 0xeeb  :    0 - 0x0
    "00000000", -- 3820 - 0xeec  :    0 - 0x0
    "00000000", -- 3821 - 0xeed  :    0 - 0x0
    "00000000", -- 3822 - 0xeee  :    0 - 0x0
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "00000000", -- 3824 - 0xef0  :    0 - 0x0 -- Sprite 0xef
    "00000000", -- 3825 - 0xef1  :    0 - 0x0
    "00000000", -- 3826 - 0xef2  :    0 - 0x0
    "00000000", -- 3827 - 0xef3  :    0 - 0x0
    "00000000", -- 3828 - 0xef4  :    0 - 0x0
    "00000000", -- 3829 - 0xef5  :    0 - 0x0
    "00000000", -- 3830 - 0xef6  :    0 - 0x0
    "00000000", -- 3831 - 0xef7  :    0 - 0x0
    "00000000", -- 3832 - 0xef8  :    0 - 0x0
    "00000000", -- 3833 - 0xef9  :    0 - 0x0
    "00000000", -- 3834 - 0xefa  :    0 - 0x0
    "00000000", -- 3835 - 0xefb  :    0 - 0x0
    "00000000", -- 3836 - 0xefc  :    0 - 0x0
    "00000000", -- 3837 - 0xefd  :    0 - 0x0
    "00000000", -- 3838 - 0xefe  :    0 - 0x0
    "00000000", -- 3839 - 0xeff  :    0 - 0x0
    "00000000", -- 3840 - 0xf00  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 3841 - 0xf01  :    0 - 0x0
    "00000000", -- 3842 - 0xf02  :    0 - 0x0
    "00000000", -- 3843 - 0xf03  :    0 - 0x0
    "00000000", -- 3844 - 0xf04  :    0 - 0x0
    "00000000", -- 3845 - 0xf05  :    0 - 0x0
    "00000000", -- 3846 - 0xf06  :    0 - 0x0
    "00000000", -- 3847 - 0xf07  :    0 - 0x0
    "00000000", -- 3848 - 0xf08  :    0 - 0x0
    "00000000", -- 3849 - 0xf09  :    0 - 0x0
    "00000000", -- 3850 - 0xf0a  :    0 - 0x0
    "00000000", -- 3851 - 0xf0b  :    0 - 0x0
    "00000000", -- 3852 - 0xf0c  :    0 - 0x0
    "00000000", -- 3853 - 0xf0d  :    0 - 0x0
    "00000000", -- 3854 - 0xf0e  :    0 - 0x0
    "00000000", -- 3855 - 0xf0f  :    0 - 0x0
    "00000000", -- 3856 - 0xf10  :    0 - 0x0 -- Sprite 0xf1
    "00000000", -- 3857 - 0xf11  :    0 - 0x0
    "00000000", -- 3858 - 0xf12  :    0 - 0x0
    "00000000", -- 3859 - 0xf13  :    0 - 0x0
    "00000000", -- 3860 - 0xf14  :    0 - 0x0
    "00000000", -- 3861 - 0xf15  :    0 - 0x0
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "00000000", -- 3864 - 0xf18  :    0 - 0x0
    "00000000", -- 3865 - 0xf19  :    0 - 0x0
    "00000000", -- 3866 - 0xf1a  :    0 - 0x0
    "00000000", -- 3867 - 0xf1b  :    0 - 0x0
    "00000000", -- 3868 - 0xf1c  :    0 - 0x0
    "00000000", -- 3869 - 0xf1d  :    0 - 0x0
    "00000000", -- 3870 - 0xf1e  :    0 - 0x0
    "00000000", -- 3871 - 0xf1f  :    0 - 0x0
    "00000000", -- 3872 - 0xf20  :    0 - 0x0 -- Sprite 0xf2
    "00000000", -- 3873 - 0xf21  :    0 - 0x0
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000000", -- 3876 - 0xf24  :    0 - 0x0
    "00000000", -- 3877 - 0xf25  :    0 - 0x0
    "00000000", -- 3878 - 0xf26  :    0 - 0x0
    "00000000", -- 3879 - 0xf27  :    0 - 0x0
    "00000000", -- 3880 - 0xf28  :    0 - 0x0
    "00000000", -- 3881 - 0xf29  :    0 - 0x0
    "00000000", -- 3882 - 0xf2a  :    0 - 0x0
    "00000000", -- 3883 - 0xf2b  :    0 - 0x0
    "00000000", -- 3884 - 0xf2c  :    0 - 0x0
    "00000000", -- 3885 - 0xf2d  :    0 - 0x0
    "00000000", -- 3886 - 0xf2e  :    0 - 0x0
    "00000000", -- 3887 - 0xf2f  :    0 - 0x0
    "00000000", -- 3888 - 0xf30  :    0 - 0x0 -- Sprite 0xf3
    "00000000", -- 3889 - 0xf31  :    0 - 0x0
    "00000000", -- 3890 - 0xf32  :    0 - 0x0
    "00000000", -- 3891 - 0xf33  :    0 - 0x0
    "00000000", -- 3892 - 0xf34  :    0 - 0x0
    "00000000", -- 3893 - 0xf35  :    0 - 0x0
    "00000000", -- 3894 - 0xf36  :    0 - 0x0
    "00000000", -- 3895 - 0xf37  :    0 - 0x0
    "00000000", -- 3896 - 0xf38  :    0 - 0x0
    "00000000", -- 3897 - 0xf39  :    0 - 0x0
    "00000000", -- 3898 - 0xf3a  :    0 - 0x0
    "00000000", -- 3899 - 0xf3b  :    0 - 0x0
    "00000000", -- 3900 - 0xf3c  :    0 - 0x0
    "00000000", -- 3901 - 0xf3d  :    0 - 0x0
    "00000000", -- 3902 - 0xf3e  :    0 - 0x0
    "00000000", -- 3903 - 0xf3f  :    0 - 0x0
    "00000000", -- 3904 - 0xf40  :    0 - 0x0 -- Sprite 0xf4
    "00000000", -- 3905 - 0xf41  :    0 - 0x0
    "00000000", -- 3906 - 0xf42  :    0 - 0x0
    "00000000", -- 3907 - 0xf43  :    0 - 0x0
    "00000000", -- 3908 - 0xf44  :    0 - 0x0
    "00000000", -- 3909 - 0xf45  :    0 - 0x0
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "00000000", -- 3911 - 0xf47  :    0 - 0x0
    "00000000", -- 3912 - 0xf48  :    0 - 0x0
    "00000000", -- 3913 - 0xf49  :    0 - 0x0
    "00000000", -- 3914 - 0xf4a  :    0 - 0x0
    "00000000", -- 3915 - 0xf4b  :    0 - 0x0
    "00000000", -- 3916 - 0xf4c  :    0 - 0x0
    "00000000", -- 3917 - 0xf4d  :    0 - 0x0
    "00000000", -- 3918 - 0xf4e  :    0 - 0x0
    "00000000", -- 3919 - 0xf4f  :    0 - 0x0
    "00000000", -- 3920 - 0xf50  :    0 - 0x0 -- Sprite 0xf5
    "00000000", -- 3921 - 0xf51  :    0 - 0x0
    "00000000", -- 3922 - 0xf52  :    0 - 0x0
    "00000000", -- 3923 - 0xf53  :    0 - 0x0
    "00000000", -- 3924 - 0xf54  :    0 - 0x0
    "00000000", -- 3925 - 0xf55  :    0 - 0x0
    "00000000", -- 3926 - 0xf56  :    0 - 0x0
    "00000000", -- 3927 - 0xf57  :    0 - 0x0
    "00000000", -- 3928 - 0xf58  :    0 - 0x0
    "00000000", -- 3929 - 0xf59  :    0 - 0x0
    "00000000", -- 3930 - 0xf5a  :    0 - 0x0
    "00000000", -- 3931 - 0xf5b  :    0 - 0x0
    "00000000", -- 3932 - 0xf5c  :    0 - 0x0
    "00000000", -- 3933 - 0xf5d  :    0 - 0x0
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Sprite 0xf6
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00000000", -- 3941 - 0xf65  :    0 - 0x0
    "00000000", -- 3942 - 0xf66  :    0 - 0x0
    "00000000", -- 3943 - 0xf67  :    0 - 0x0
    "00000000", -- 3944 - 0xf68  :    0 - 0x0
    "00000000", -- 3945 - 0xf69  :    0 - 0x0
    "00000000", -- 3946 - 0xf6a  :    0 - 0x0
    "00000000", -- 3947 - 0xf6b  :    0 - 0x0
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "00000000", -- 3949 - 0xf6d  :    0 - 0x0
    "00000000", -- 3950 - 0xf6e  :    0 - 0x0
    "00000000", -- 3951 - 0xf6f  :    0 - 0x0
    "00000000", -- 3952 - 0xf70  :    0 - 0x0 -- Sprite 0xf7
    "00000000", -- 3953 - 0xf71  :    0 - 0x0
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00000000", -- 3958 - 0xf76  :    0 - 0x0
    "00000000", -- 3959 - 0xf77  :    0 - 0x0
    "00000000", -- 3960 - 0xf78  :    0 - 0x0
    "00000000", -- 3961 - 0xf79  :    0 - 0x0
    "00000000", -- 3962 - 0xf7a  :    0 - 0x0
    "00000000", -- 3963 - 0xf7b  :    0 - 0x0
    "00000000", -- 3964 - 0xf7c  :    0 - 0x0
    "00000000", -- 3965 - 0xf7d  :    0 - 0x0
    "00000000", -- 3966 - 0xf7e  :    0 - 0x0
    "00000000", -- 3967 - 0xf7f  :    0 - 0x0
    "00000000", -- 3968 - 0xf80  :    0 - 0x0 -- Sprite 0xf8
    "00000000", -- 3969 - 0xf81  :    0 - 0x0
    "00000000", -- 3970 - 0xf82  :    0 - 0x0
    "00000000", -- 3971 - 0xf83  :    0 - 0x0
    "00000000", -- 3972 - 0xf84  :    0 - 0x0
    "00000000", -- 3973 - 0xf85  :    0 - 0x0
    "00000000", -- 3974 - 0xf86  :    0 - 0x0
    "00000000", -- 3975 - 0xf87  :    0 - 0x0
    "00000000", -- 3976 - 0xf88  :    0 - 0x0
    "00000000", -- 3977 - 0xf89  :    0 - 0x0
    "00000000", -- 3978 - 0xf8a  :    0 - 0x0
    "00000000", -- 3979 - 0xf8b  :    0 - 0x0
    "00000000", -- 3980 - 0xf8c  :    0 - 0x0
    "00000000", -- 3981 - 0xf8d  :    0 - 0x0
    "00000000", -- 3982 - 0xf8e  :    0 - 0x0
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "00000000", -- 3984 - 0xf90  :    0 - 0x0 -- Sprite 0xf9
    "00000000", -- 3985 - 0xf91  :    0 - 0x0
    "00000000", -- 3986 - 0xf92  :    0 - 0x0
    "00000000", -- 3987 - 0xf93  :    0 - 0x0
    "00000000", -- 3988 - 0xf94  :    0 - 0x0
    "00000000", -- 3989 - 0xf95  :    0 - 0x0
    "00000000", -- 3990 - 0xf96  :    0 - 0x0
    "00000000", -- 3991 - 0xf97  :    0 - 0x0
    "00000000", -- 3992 - 0xf98  :    0 - 0x0
    "00000000", -- 3993 - 0xf99  :    0 - 0x0
    "00000000", -- 3994 - 0xf9a  :    0 - 0x0
    "00000000", -- 3995 - 0xf9b  :    0 - 0x0
    "00000000", -- 3996 - 0xf9c  :    0 - 0x0
    "00000000", -- 3997 - 0xf9d  :    0 - 0x0
    "00000000", -- 3998 - 0xf9e  :    0 - 0x0
    "00000000", -- 3999 - 0xf9f  :    0 - 0x0
    "00000000", -- 4000 - 0xfa0  :    0 - 0x0 -- Sprite 0xfa
    "00000000", -- 4001 - 0xfa1  :    0 - 0x0
    "00000000", -- 4002 - 0xfa2  :    0 - 0x0
    "00000000", -- 4003 - 0xfa3  :    0 - 0x0
    "00000000", -- 4004 - 0xfa4  :    0 - 0x0
    "00000000", -- 4005 - 0xfa5  :    0 - 0x0
    "00000000", -- 4006 - 0xfa6  :    0 - 0x0
    "00000000", -- 4007 - 0xfa7  :    0 - 0x0
    "00000000", -- 4008 - 0xfa8  :    0 - 0x0
    "00000000", -- 4009 - 0xfa9  :    0 - 0x0
    "00000000", -- 4010 - 0xfaa  :    0 - 0x0
    "00000000", -- 4011 - 0xfab  :    0 - 0x0
    "00000000", -- 4012 - 0xfac  :    0 - 0x0
    "00000000", -- 4013 - 0xfad  :    0 - 0x0
    "00000000", -- 4014 - 0xfae  :    0 - 0x0
    "00000000", -- 4015 - 0xfaf  :    0 - 0x0
    "00000000", -- 4016 - 0xfb0  :    0 - 0x0 -- Sprite 0xfb
    "00000000", -- 4017 - 0xfb1  :    0 - 0x0
    "00000000", -- 4018 - 0xfb2  :    0 - 0x0
    "00000000", -- 4019 - 0xfb3  :    0 - 0x0
    "00000000", -- 4020 - 0xfb4  :    0 - 0x0
    "00000000", -- 4021 - 0xfb5  :    0 - 0x0
    "00000000", -- 4022 - 0xfb6  :    0 - 0x0
    "00000000", -- 4023 - 0xfb7  :    0 - 0x0
    "00000000", -- 4024 - 0xfb8  :    0 - 0x0
    "00000000", -- 4025 - 0xfb9  :    0 - 0x0
    "00000000", -- 4026 - 0xfba  :    0 - 0x0
    "00000000", -- 4027 - 0xfbb  :    0 - 0x0
    "00000000", -- 4028 - 0xfbc  :    0 - 0x0
    "00000000", -- 4029 - 0xfbd  :    0 - 0x0
    "00000000", -- 4030 - 0xfbe  :    0 - 0x0
    "00000000", -- 4031 - 0xfbf  :    0 - 0x0
    "00000000", -- 4032 - 0xfc0  :    0 - 0x0 -- Sprite 0xfc
    "00000000", -- 4033 - 0xfc1  :    0 - 0x0
    "00000000", -- 4034 - 0xfc2  :    0 - 0x0
    "00000000", -- 4035 - 0xfc3  :    0 - 0x0
    "00000000", -- 4036 - 0xfc4  :    0 - 0x0
    "00000000", -- 4037 - 0xfc5  :    0 - 0x0
    "00000000", -- 4038 - 0xfc6  :    0 - 0x0
    "00000000", -- 4039 - 0xfc7  :    0 - 0x0
    "00000000", -- 4040 - 0xfc8  :    0 - 0x0
    "00000000", -- 4041 - 0xfc9  :    0 - 0x0
    "00000000", -- 4042 - 0xfca  :    0 - 0x0
    "00000000", -- 4043 - 0xfcb  :    0 - 0x0
    "00000000", -- 4044 - 0xfcc  :    0 - 0x0
    "00000000", -- 4045 - 0xfcd  :    0 - 0x0
    "00000000", -- 4046 - 0xfce  :    0 - 0x0
    "00000000", -- 4047 - 0xfcf  :    0 - 0x0
    "00000000", -- 4048 - 0xfd0  :    0 - 0x0 -- Sprite 0xfd
    "00000000", -- 4049 - 0xfd1  :    0 - 0x0
    "00000000", -- 4050 - 0xfd2  :    0 - 0x0
    "00000000", -- 4051 - 0xfd3  :    0 - 0x0
    "00000000", -- 4052 - 0xfd4  :    0 - 0x0
    "00000000", -- 4053 - 0xfd5  :    0 - 0x0
    "00000000", -- 4054 - 0xfd6  :    0 - 0x0
    "00000000", -- 4055 - 0xfd7  :    0 - 0x0
    "00000000", -- 4056 - 0xfd8  :    0 - 0x0
    "00000000", -- 4057 - 0xfd9  :    0 - 0x0
    "00000000", -- 4058 - 0xfda  :    0 - 0x0
    "00000000", -- 4059 - 0xfdb  :    0 - 0x0
    "00000000", -- 4060 - 0xfdc  :    0 - 0x0
    "00000000", -- 4061 - 0xfdd  :    0 - 0x0
    "00000000", -- 4062 - 0xfde  :    0 - 0x0
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00000000", -- 4064 - 0xfe0  :    0 - 0x0 -- Sprite 0xfe
    "00000000", -- 4065 - 0xfe1  :    0 - 0x0
    "00000000", -- 4066 - 0xfe2  :    0 - 0x0
    "00000000", -- 4067 - 0xfe3  :    0 - 0x0
    "00000000", -- 4068 - 0xfe4  :    0 - 0x0
    "00000000", -- 4069 - 0xfe5  :    0 - 0x0
    "00000000", -- 4070 - 0xfe6  :    0 - 0x0
    "00000000", -- 4071 - 0xfe7  :    0 - 0x0
    "00000000", -- 4072 - 0xfe8  :    0 - 0x0
    "00000000", -- 4073 - 0xfe9  :    0 - 0x0
    "00000000", -- 4074 - 0xfea  :    0 - 0x0
    "00000000", -- 4075 - 0xfeb  :    0 - 0x0
    "00000000", -- 4076 - 0xfec  :    0 - 0x0
    "00000000", -- 4077 - 0xfed  :    0 - 0x0
    "00000000", -- 4078 - 0xfee  :    0 - 0x0
    "00000000", -- 4079 - 0xfef  :    0 - 0x0
    "00000000", -- 4080 - 0xff0  :    0 - 0x0 -- Sprite 0xff
    "00000000", -- 4081 - 0xff1  :    0 - 0x0
    "00000000", -- 4082 - 0xff2  :    0 - 0x0
    "00000000", -- 4083 - 0xff3  :    0 - 0x0
    "00000000", -- 4084 - 0xff4  :    0 - 0x0
    "00000000", -- 4085 - 0xff5  :    0 - 0x0
    "00000000", -- 4086 - 0xff6  :    0 - 0x0
    "00000000", -- 4087 - 0xff7  :    0 - 0x0
    "00000000", -- 4088 - 0xff8  :    0 - 0x0
    "00000000", -- 4089 - 0xff9  :    0 - 0x0
    "00000000", -- 4090 - 0xffa  :    0 - 0x0
    "00000000", -- 4091 - 0xffb  :    0 - 0x0
    "00000000", -- 4092 - 0xffc  :    0 - 0x0
    "00000000", -- 4093 - 0xffd  :    0 - 0x0
    "00000000", -- 4094 - 0xffe  :    0 - 0x0
    "00000000", -- 4095 - 0xfff  :    0 - 0x0
          -- Pattern Table 1---------
    "00111110", -- 4096 - 0x1000  :   62 - 0x3e -- Background 0x0
    "01111111", -- 4097 - 0x1001  :  127 - 0x7f
    "01110111", -- 4098 - 0x1002  :  119 - 0x77
    "01111111", -- 4099 - 0x1003  :  127 - 0x7f
    "01111111", -- 4100 - 0x1004  :  127 - 0x7f
    "01110111", -- 4101 - 0x1005  :  119 - 0x77
    "01111111", -- 4102 - 0x1006  :  127 - 0x7f
    "00111110", -- 4103 - 0x1007  :   62 - 0x3e
    "11000011", -- 4104 - 0x1008  :  195 - 0xc3
    "10000001", -- 4105 - 0x1009  :  129 - 0x81
    "10011001", -- 4106 - 0x100a  :  153 - 0x99
    "10010001", -- 4107 - 0x100b  :  145 - 0x91
    "10001001", -- 4108 - 0x100c  :  137 - 0x89
    "10011001", -- 4109 - 0x100d  :  153 - 0x99
    "10000001", -- 4110 - 0x100e  :  129 - 0x81
    "11000011", -- 4111 - 0x100f  :  195 - 0xc3
    "00011100", -- 4112 - 0x1010  :   28 - 0x1c -- Background 0x1
    "00111100", -- 4113 - 0x1011  :   60 - 0x3c
    "01111100", -- 4114 - 0x1012  :  124 - 0x7c
    "00011100", -- 4115 - 0x1013  :   28 - 0x1c
    "00011100", -- 4116 - 0x1014  :   28 - 0x1c
    "00011100", -- 4117 - 0x1015  :   28 - 0x1c
    "01111111", -- 4118 - 0x1016  :  127 - 0x7f
    "01111111", -- 4119 - 0x1017  :  127 - 0x7f
    "11100111", -- 4120 - 0x1018  :  231 - 0xe7
    "11000111", -- 4121 - 0x1019  :  199 - 0xc7
    "10000111", -- 4122 - 0x101a  :  135 - 0x87
    "11100111", -- 4123 - 0x101b  :  231 - 0xe7
    "11100111", -- 4124 - 0x101c  :  231 - 0xe7
    "11100111", -- 4125 - 0x101d  :  231 - 0xe7
    "10000001", -- 4126 - 0x101e  :  129 - 0x81
    "10000001", -- 4127 - 0x101f  :  129 - 0x81
    "00111110", -- 4128 - 0x1020  :   62 - 0x3e -- Background 0x2
    "01111111", -- 4129 - 0x1021  :  127 - 0x7f
    "00000111", -- 4130 - 0x1022  :    7 - 0x7
    "00111111", -- 4131 - 0x1023  :   63 - 0x3f
    "01111111", -- 4132 - 0x1024  :  127 - 0x7f
    "01110000", -- 4133 - 0x1025  :  112 - 0x70
    "01111111", -- 4134 - 0x1026  :  127 - 0x7f
    "01111111", -- 4135 - 0x1027  :  127 - 0x7f
    "11000011", -- 4136 - 0x1028  :  195 - 0xc3
    "10000001", -- 4137 - 0x1029  :  129 - 0x81
    "11111001", -- 4138 - 0x102a  :  249 - 0xf9
    "11000001", -- 4139 - 0x102b  :  193 - 0xc1
    "10000001", -- 4140 - 0x102c  :  129 - 0x81
    "10011111", -- 4141 - 0x102d  :  159 - 0x9f
    "10000001", -- 4142 - 0x102e  :  129 - 0x81
    "10000001", -- 4143 - 0x102f  :  129 - 0x81
    "00111110", -- 4144 - 0x1030  :   62 - 0x3e -- Background 0x3
    "01111111", -- 4145 - 0x1031  :  127 - 0x7f
    "00000111", -- 4146 - 0x1032  :    7 - 0x7
    "00011111", -- 4147 - 0x1033  :   31 - 0x1f
    "00011111", -- 4148 - 0x1034  :   31 - 0x1f
    "00000111", -- 4149 - 0x1035  :    7 - 0x7
    "01111111", -- 4150 - 0x1036  :  127 - 0x7f
    "00111110", -- 4151 - 0x1037  :   62 - 0x3e
    "11000011", -- 4152 - 0x1038  :  195 - 0xc3
    "10000001", -- 4153 - 0x1039  :  129 - 0x81
    "11111001", -- 4154 - 0x103a  :  249 - 0xf9
    "11100001", -- 4155 - 0x103b  :  225 - 0xe1
    "11100001", -- 4156 - 0x103c  :  225 - 0xe1
    "11111001", -- 4157 - 0x103d  :  249 - 0xf9
    "10000001", -- 4158 - 0x103e  :  129 - 0x81
    "11000011", -- 4159 - 0x103f  :  195 - 0xc3
    "00110000", -- 4160 - 0x1040  :   48 - 0x30 -- Background 0x4
    "01110000", -- 4161 - 0x1041  :  112 - 0x70
    "01110111", -- 4162 - 0x1042  :  119 - 0x77
    "01110111", -- 4163 - 0x1043  :  119 - 0x77
    "01111111", -- 4164 - 0x1044  :  127 - 0x7f
    "01111111", -- 4165 - 0x1045  :  127 - 0x7f
    "00000111", -- 4166 - 0x1046  :    7 - 0x7
    "00000111", -- 4167 - 0x1047  :    7 - 0x7
    "11011111", -- 4168 - 0x1048  :  223 - 0xdf
    "10011111", -- 4169 - 0x1049  :  159 - 0x9f
    "10011001", -- 4170 - 0x104a  :  153 - 0x99
    "10011001", -- 4171 - 0x104b  :  153 - 0x99
    "10000000", -- 4172 - 0x104c  :  128 - 0x80
    "10000000", -- 4173 - 0x104d  :  128 - 0x80
    "11111001", -- 4174 - 0x104e  :  249 - 0xf9
    "11111001", -- 4175 - 0x104f  :  249 - 0xf9
    "01111111", -- 4176 - 0x1050  :  127 - 0x7f -- Background 0x5
    "01111111", -- 4177 - 0x1051  :  127 - 0x7f
    "01110000", -- 4178 - 0x1052  :  112 - 0x70
    "01111110", -- 4179 - 0x1053  :  126 - 0x7e
    "01111111", -- 4180 - 0x1054  :  127 - 0x7f
    "00000111", -- 4181 - 0x1055  :    7 - 0x7
    "01111111", -- 4182 - 0x1056  :  127 - 0x7f
    "00111110", -- 4183 - 0x1057  :   62 - 0x3e
    "10000001", -- 4184 - 0x1058  :  129 - 0x81
    "10000001", -- 4185 - 0x1059  :  129 - 0x81
    "10011111", -- 4186 - 0x105a  :  159 - 0x9f
    "10000011", -- 4187 - 0x105b  :  131 - 0x83
    "10000001", -- 4188 - 0x105c  :  129 - 0x81
    "11111001", -- 4189 - 0x105d  :  249 - 0xf9
    "10000001", -- 4190 - 0x105e  :  129 - 0x81
    "11000011", -- 4191 - 0x105f  :  195 - 0xc3
    "00111110", -- 4192 - 0x1060  :   62 - 0x3e -- Background 0x6
    "01111111", -- 4193 - 0x1061  :  127 - 0x7f
    "01110000", -- 4194 - 0x1062  :  112 - 0x70
    "01111110", -- 4195 - 0x1063  :  126 - 0x7e
    "01111111", -- 4196 - 0x1064  :  127 - 0x7f
    "01110111", -- 4197 - 0x1065  :  119 - 0x77
    "01111111", -- 4198 - 0x1066  :  127 - 0x7f
    "00111110", -- 4199 - 0x1067  :   62 - 0x3e
    "11000011", -- 4200 - 0x1068  :  195 - 0xc3
    "10000001", -- 4201 - 0x1069  :  129 - 0x81
    "10011111", -- 4202 - 0x106a  :  159 - 0x9f
    "10000011", -- 4203 - 0x106b  :  131 - 0x83
    "10000001", -- 4204 - 0x106c  :  129 - 0x81
    "10011001", -- 4205 - 0x106d  :  153 - 0x99
    "10000001", -- 4206 - 0x106e  :  129 - 0x81
    "11000011", -- 4207 - 0x106f  :  195 - 0xc3
    "01111111", -- 4208 - 0x1070  :  127 - 0x7f -- Background 0x7
    "01111111", -- 4209 - 0x1071  :  127 - 0x7f
    "00000111", -- 4210 - 0x1072  :    7 - 0x7
    "00001110", -- 4211 - 0x1073  :   14 - 0xe
    "00001110", -- 4212 - 0x1074  :   14 - 0xe
    "00011100", -- 4213 - 0x1075  :   28 - 0x1c
    "00011100", -- 4214 - 0x1076  :   28 - 0x1c
    "00011100", -- 4215 - 0x1077  :   28 - 0x1c
    "10000001", -- 4216 - 0x1078  :  129 - 0x81
    "10000001", -- 4217 - 0x1079  :  129 - 0x81
    "11111001", -- 4218 - 0x107a  :  249 - 0xf9
    "11110011", -- 4219 - 0x107b  :  243 - 0xf3
    "11110011", -- 4220 - 0x107c  :  243 - 0xf3
    "11100111", -- 4221 - 0x107d  :  231 - 0xe7
    "11100111", -- 4222 - 0x107e  :  231 - 0xe7
    "11100111", -- 4223 - 0x107f  :  231 - 0xe7
    "00111110", -- 4224 - 0x1080  :   62 - 0x3e -- Background 0x8
    "01111111", -- 4225 - 0x1081  :  127 - 0x7f
    "01110111", -- 4226 - 0x1082  :  119 - 0x77
    "00111110", -- 4227 - 0x1083  :   62 - 0x3e
    "01111111", -- 4228 - 0x1084  :  127 - 0x7f
    "01110111", -- 4229 - 0x1085  :  119 - 0x77
    "01111111", -- 4230 - 0x1086  :  127 - 0x7f
    "00111110", -- 4231 - 0x1087  :   62 - 0x3e
    "11000011", -- 4232 - 0x1088  :  195 - 0xc3
    "10000001", -- 4233 - 0x1089  :  129 - 0x81
    "10011001", -- 4234 - 0x108a  :  153 - 0x99
    "11000011", -- 4235 - 0x108b  :  195 - 0xc3
    "10000001", -- 4236 - 0x108c  :  129 - 0x81
    "10011001", -- 4237 - 0x108d  :  153 - 0x99
    "10000001", -- 4238 - 0x108e  :  129 - 0x81
    "11000011", -- 4239 - 0x108f  :  195 - 0xc3
    "00111110", -- 4240 - 0x1090  :   62 - 0x3e -- Background 0x9
    "01111111", -- 4241 - 0x1091  :  127 - 0x7f
    "01110111", -- 4242 - 0x1092  :  119 - 0x77
    "01111111", -- 4243 - 0x1093  :  127 - 0x7f
    "00111111", -- 4244 - 0x1094  :   63 - 0x3f
    "00000111", -- 4245 - 0x1095  :    7 - 0x7
    "01111111", -- 4246 - 0x1096  :  127 - 0x7f
    "00111110", -- 4247 - 0x1097  :   62 - 0x3e
    "11000011", -- 4248 - 0x1098  :  195 - 0xc3
    "10000001", -- 4249 - 0x1099  :  129 - 0x81
    "10011001", -- 4250 - 0x109a  :  153 - 0x99
    "10000001", -- 4251 - 0x109b  :  129 - 0x81
    "11000001", -- 4252 - 0x109c  :  193 - 0xc1
    "11111001", -- 4253 - 0x109d  :  249 - 0xf9
    "10000001", -- 4254 - 0x109e  :  129 - 0x81
    "11000011", -- 4255 - 0x109f  :  195 - 0xc3
    "00000000", -- 4256 - 0x10a0  :    0 - 0x0 -- Background 0xa
    "00000000", -- 4257 - 0x10a1  :    0 - 0x0
    "00000000", -- 4258 - 0x10a2  :    0 - 0x0
    "00000000", -- 4259 - 0x10a3  :    0 - 0x0
    "00000000", -- 4260 - 0x10a4  :    0 - 0x0
    "00110000", -- 4261 - 0x10a5  :   48 - 0x30
    "01111000", -- 4262 - 0x10a6  :  120 - 0x78
    "00110000", -- 4263 - 0x10a7  :   48 - 0x30
    "11111111", -- 4264 - 0x10a8  :  255 - 0xff
    "11111111", -- 4265 - 0x10a9  :  255 - 0xff
    "11111111", -- 4266 - 0x10aa  :  255 - 0xff
    "11111111", -- 4267 - 0x10ab  :  255 - 0xff
    "11111111", -- 4268 - 0x10ac  :  255 - 0xff
    "11011111", -- 4269 - 0x10ad  :  223 - 0xdf
    "10001111", -- 4270 - 0x10ae  :  143 - 0x8f
    "11011111", -- 4271 - 0x10af  :  223 - 0xdf
    "01110000", -- 4272 - 0x10b0  :  112 - 0x70 -- Background 0xb
    "11111000", -- 4273 - 0x10b1  :  248 - 0xf8
    "11111000", -- 4274 - 0x10b2  :  248 - 0xf8
    "11111000", -- 4275 - 0x10b3  :  248 - 0xf8
    "01110000", -- 4276 - 0x10b4  :  112 - 0x70
    "00000000", -- 4277 - 0x10b5  :    0 - 0x0
    "01110000", -- 4278 - 0x10b6  :  112 - 0x70
    "01110000", -- 4279 - 0x10b7  :  112 - 0x70
    "10011111", -- 4280 - 0x10b8  :  159 - 0x9f
    "00001111", -- 4281 - 0x10b9  :   15 - 0xf
    "00001111", -- 4282 - 0x10ba  :   15 - 0xf
    "00001111", -- 4283 - 0x10bb  :   15 - 0xf
    "10011111", -- 4284 - 0x10bc  :  159 - 0x9f
    "11111111", -- 4285 - 0x10bd  :  255 - 0xff
    "10011111", -- 4286 - 0x10be  :  159 - 0x9f
    "10011111", -- 4287 - 0x10bf  :  159 - 0x9f
    "01111000", -- 4288 - 0x10c0  :  120 - 0x78 -- Background 0xc
    "11111100", -- 4289 - 0x10c1  :  252 - 0xfc
    "00011100", -- 4290 - 0x10c2  :   28 - 0x1c
    "00111000", -- 4291 - 0x10c3  :   56 - 0x38
    "00110000", -- 4292 - 0x10c4  :   48 - 0x30
    "00000000", -- 4293 - 0x10c5  :    0 - 0x0
    "01110000", -- 4294 - 0x10c6  :  112 - 0x70
    "01110000", -- 4295 - 0x10c7  :  112 - 0x70
    "10001111", -- 4296 - 0x10c8  :  143 - 0x8f
    "00100111", -- 4297 - 0x10c9  :   39 - 0x27
    "11100111", -- 4298 - 0x10ca  :  231 - 0xe7
    "11001111", -- 4299 - 0x10cb  :  207 - 0xcf
    "11011111", -- 4300 - 0x10cc  :  223 - 0xdf
    "11111111", -- 4301 - 0x10cd  :  255 - 0xff
    "10011111", -- 4302 - 0x10ce  :  159 - 0x9f
    "10011111", -- 4303 - 0x10cf  :  159 - 0x9f
    "00111100", -- 4304 - 0x10d0  :   60 - 0x3c -- Background 0xd
    "01111110", -- 4305 - 0x10d1  :  126 - 0x7e
    "11011011", -- 4306 - 0x10d2  :  219 - 0xdb
    "11011111", -- 4307 - 0x10d3  :  223 - 0xdf
    "11000011", -- 4308 - 0x10d4  :  195 - 0xc3
    "01100110", -- 4309 - 0x10d5  :  102 - 0x66
    "00111100", -- 4310 - 0x10d6  :   60 - 0x3c
    "00000000", -- 4311 - 0x10d7  :    0 - 0x0
    "11000111", -- 4312 - 0x10d8  :  199 - 0xc7
    "10101011", -- 4313 - 0x10d9  :  171 - 0xab
    "01101101", -- 4314 - 0x10da  :  109 - 0x6d
    "01100101", -- 4315 - 0x10db  :  101 - 0x65
    "01111101", -- 4316 - 0x10dc  :  125 - 0x7d
    "10111011", -- 4317 - 0x10dd  :  187 - 0xbb
    "11000111", -- 4318 - 0x10de  :  199 - 0xc7
    "11111111", -- 4319 - 0x10df  :  255 - 0xff
    "00000000", -- 4320 - 0x10e0  :    0 - 0x0 -- Background 0xe
    "00000000", -- 4321 - 0x10e1  :    0 - 0x0
    "00000000", -- 4322 - 0x10e2  :    0 - 0x0
    "00111100", -- 4323 - 0x10e3  :   60 - 0x3c
    "00111110", -- 4324 - 0x10e4  :   62 - 0x3e
    "00011110", -- 4325 - 0x10e5  :   30 - 0x1e
    "00000000", -- 4326 - 0x10e6  :    0 - 0x0
    "00000000", -- 4327 - 0x10e7  :    0 - 0x0
    "11111111", -- 4328 - 0x10e8  :  255 - 0xff
    "11111111", -- 4329 - 0x10e9  :  255 - 0xff
    "11111111", -- 4330 - 0x10ea  :  255 - 0xff
    "11000011", -- 4331 - 0x10eb  :  195 - 0xc3
    "11000011", -- 4332 - 0x10ec  :  195 - 0xc3
    "11111111", -- 4333 - 0x10ed  :  255 - 0xff
    "11111111", -- 4334 - 0x10ee  :  255 - 0xff
    "11111111", -- 4335 - 0x10ef  :  255 - 0xff
    "11111111", -- 4336 - 0x10f0  :  255 - 0xff -- Background 0xf
    "11111111", -- 4337 - 0x10f1  :  255 - 0xff
    "11111111", -- 4338 - 0x10f2  :  255 - 0xff
    "11111111", -- 4339 - 0x10f3  :  255 - 0xff
    "11111111", -- 4340 - 0x10f4  :  255 - 0xff
    "11111111", -- 4341 - 0x10f5  :  255 - 0xff
    "11100000", -- 4342 - 0x10f6  :  224 - 0xe0
    "11100000", -- 4343 - 0x10f7  :  224 - 0xe0
    "00000001", -- 4344 - 0x10f8  :    1 - 0x1
    "00101001", -- 4345 - 0x10f9  :   41 - 0x29
    "01010101", -- 4346 - 0x10fa  :   85 - 0x55
    "00101001", -- 4347 - 0x10fb  :   41 - 0x29
    "01010101", -- 4348 - 0x10fc  :   85 - 0x55
    "00000001", -- 4349 - 0x10fd  :    1 - 0x1
    "00111111", -- 4350 - 0x10fe  :   63 - 0x3f
    "00111111", -- 4351 - 0x10ff  :   63 - 0x3f
    "00001110", -- 4352 - 0x1100  :   14 - 0xe -- Background 0x10
    "00001110", -- 4353 - 0x1101  :   14 - 0xe
    "00011100", -- 4354 - 0x1102  :   28 - 0x1c
    "00011100", -- 4355 - 0x1103  :   28 - 0x1c
    "00011100", -- 4356 - 0x1104  :   28 - 0x1c
    "00011100", -- 4357 - 0x1105  :   28 - 0x1c
    "00111000", -- 4358 - 0x1106  :   56 - 0x38
    "00111000", -- 4359 - 0x1107  :   56 - 0x38
    "11110011", -- 4360 - 0x1108  :  243 - 0xf3
    "11110011", -- 4361 - 0x1109  :  243 - 0xf3
    "11100111", -- 4362 - 0x110a  :  231 - 0xe7
    "11100111", -- 4363 - 0x110b  :  231 - 0xe7
    "11100111", -- 4364 - 0x110c  :  231 - 0xe7
    "11100111", -- 4365 - 0x110d  :  231 - 0xe7
    "11001111", -- 4366 - 0x110e  :  207 - 0xcf
    "11001111", -- 4367 - 0x110f  :  207 - 0xcf
    "00011100", -- 4368 - 0x1110  :   28 - 0x1c -- Background 0x11
    "00111110", -- 4369 - 0x1111  :   62 - 0x3e
    "01110111", -- 4370 - 0x1112  :  119 - 0x77
    "01110111", -- 4371 - 0x1113  :  119 - 0x77
    "01111111", -- 4372 - 0x1114  :  127 - 0x7f
    "01111111", -- 4373 - 0x1115  :  127 - 0x7f
    "01110111", -- 4374 - 0x1116  :  119 - 0x77
    "01110111", -- 4375 - 0x1117  :  119 - 0x77
    "11100111", -- 4376 - 0x1118  :  231 - 0xe7
    "11000011", -- 4377 - 0x1119  :  195 - 0xc3
    "10011001", -- 4378 - 0x111a  :  153 - 0x99
    "10011001", -- 4379 - 0x111b  :  153 - 0x99
    "10000001", -- 4380 - 0x111c  :  129 - 0x81
    "10000001", -- 4381 - 0x111d  :  129 - 0x81
    "10011001", -- 4382 - 0x111e  :  153 - 0x99
    "10011001", -- 4383 - 0x111f  :  153 - 0x99
    "01111110", -- 4384 - 0x1120  :  126 - 0x7e -- Background 0x12
    "01110111", -- 4385 - 0x1121  :  119 - 0x77
    "01110111", -- 4386 - 0x1122  :  119 - 0x77
    "01111110", -- 4387 - 0x1123  :  126 - 0x7e
    "01111110", -- 4388 - 0x1124  :  126 - 0x7e
    "01110111", -- 4389 - 0x1125  :  119 - 0x77
    "01110111", -- 4390 - 0x1126  :  119 - 0x77
    "01111110", -- 4391 - 0x1127  :  126 - 0x7e
    "10000011", -- 4392 - 0x1128  :  131 - 0x83
    "10011001", -- 4393 - 0x1129  :  153 - 0x99
    "10011001", -- 4394 - 0x112a  :  153 - 0x99
    "10000011", -- 4395 - 0x112b  :  131 - 0x83
    "10000011", -- 4396 - 0x112c  :  131 - 0x83
    "10011001", -- 4397 - 0x112d  :  153 - 0x99
    "10011001", -- 4398 - 0x112e  :  153 - 0x99
    "10000011", -- 4399 - 0x112f  :  131 - 0x83
    "00111110", -- 4400 - 0x1130  :   62 - 0x3e -- Background 0x13
    "01111111", -- 4401 - 0x1131  :  127 - 0x7f
    "01110111", -- 4402 - 0x1132  :  119 - 0x77
    "01110000", -- 4403 - 0x1133  :  112 - 0x70
    "01110000", -- 4404 - 0x1134  :  112 - 0x70
    "01110111", -- 4405 - 0x1135  :  119 - 0x77
    "01111111", -- 4406 - 0x1136  :  127 - 0x7f
    "00111110", -- 4407 - 0x1137  :   62 - 0x3e
    "11000011", -- 4408 - 0x1138  :  195 - 0xc3
    "10000001", -- 4409 - 0x1139  :  129 - 0x81
    "10011001", -- 4410 - 0x113a  :  153 - 0x99
    "10011111", -- 4411 - 0x113b  :  159 - 0x9f
    "10011111", -- 4412 - 0x113c  :  159 - 0x9f
    "10011001", -- 4413 - 0x113d  :  153 - 0x99
    "10000001", -- 4414 - 0x113e  :  129 - 0x81
    "11000011", -- 4415 - 0x113f  :  195 - 0xc3
    "01111110", -- 4416 - 0x1140  :  126 - 0x7e -- Background 0x14
    "01111111", -- 4417 - 0x1141  :  127 - 0x7f
    "01110111", -- 4418 - 0x1142  :  119 - 0x77
    "01110111", -- 4419 - 0x1143  :  119 - 0x77
    "01110111", -- 4420 - 0x1144  :  119 - 0x77
    "01110111", -- 4421 - 0x1145  :  119 - 0x77
    "01111111", -- 4422 - 0x1146  :  127 - 0x7f
    "01111110", -- 4423 - 0x1147  :  126 - 0x7e
    "10000011", -- 4424 - 0x1148  :  131 - 0x83
    "10000001", -- 4425 - 0x1149  :  129 - 0x81
    "10011001", -- 4426 - 0x114a  :  153 - 0x99
    "10011001", -- 4427 - 0x114b  :  153 - 0x99
    "10011001", -- 4428 - 0x114c  :  153 - 0x99
    "10011001", -- 4429 - 0x114d  :  153 - 0x99
    "10000001", -- 4430 - 0x114e  :  129 - 0x81
    "10000011", -- 4431 - 0x114f  :  131 - 0x83
    "01111111", -- 4432 - 0x1150  :  127 - 0x7f -- Background 0x15
    "01111111", -- 4433 - 0x1151  :  127 - 0x7f
    "01110000", -- 4434 - 0x1152  :  112 - 0x70
    "01111100", -- 4435 - 0x1153  :  124 - 0x7c
    "01111100", -- 4436 - 0x1154  :  124 - 0x7c
    "01110000", -- 4437 - 0x1155  :  112 - 0x70
    "01111111", -- 4438 - 0x1156  :  127 - 0x7f
    "01111111", -- 4439 - 0x1157  :  127 - 0x7f
    "10000001", -- 4440 - 0x1158  :  129 - 0x81
    "10000001", -- 4441 - 0x1159  :  129 - 0x81
    "10011111", -- 4442 - 0x115a  :  159 - 0x9f
    "10000111", -- 4443 - 0x115b  :  135 - 0x87
    "10000111", -- 4444 - 0x115c  :  135 - 0x87
    "10011111", -- 4445 - 0x115d  :  159 - 0x9f
    "10000001", -- 4446 - 0x115e  :  129 - 0x81
    "10000001", -- 4447 - 0x115f  :  129 - 0x81
    "01111111", -- 4448 - 0x1160  :  127 - 0x7f -- Background 0x16
    "01111111", -- 4449 - 0x1161  :  127 - 0x7f
    "01110000", -- 4450 - 0x1162  :  112 - 0x70
    "01111100", -- 4451 - 0x1163  :  124 - 0x7c
    "01111100", -- 4452 - 0x1164  :  124 - 0x7c
    "01110000", -- 4453 - 0x1165  :  112 - 0x70
    "01110000", -- 4454 - 0x1166  :  112 - 0x70
    "01110000", -- 4455 - 0x1167  :  112 - 0x70
    "10000001", -- 4456 - 0x1168  :  129 - 0x81
    "10000001", -- 4457 - 0x1169  :  129 - 0x81
    "10011111", -- 4458 - 0x116a  :  159 - 0x9f
    "10000111", -- 4459 - 0x116b  :  135 - 0x87
    "10000111", -- 4460 - 0x116c  :  135 - 0x87
    "10011111", -- 4461 - 0x116d  :  159 - 0x9f
    "10011111", -- 4462 - 0x116e  :  159 - 0x9f
    "10011111", -- 4463 - 0x116f  :  159 - 0x9f
    "00111110", -- 4464 - 0x1170  :   62 - 0x3e -- Background 0x17
    "01111111", -- 4465 - 0x1171  :  127 - 0x7f
    "01110111", -- 4466 - 0x1172  :  119 - 0x77
    "01110000", -- 4467 - 0x1173  :  112 - 0x70
    "01111111", -- 4468 - 0x1174  :  127 - 0x7f
    "01110111", -- 4469 - 0x1175  :  119 - 0x77
    "01111111", -- 4470 - 0x1176  :  127 - 0x7f
    "00111110", -- 4471 - 0x1177  :   62 - 0x3e
    "11000011", -- 4472 - 0x1178  :  195 - 0xc3
    "10000001", -- 4473 - 0x1179  :  129 - 0x81
    "10011001", -- 4474 - 0x117a  :  153 - 0x99
    "10011111", -- 4475 - 0x117b  :  159 - 0x9f
    "10010001", -- 4476 - 0x117c  :  145 - 0x91
    "10011001", -- 4477 - 0x117d  :  153 - 0x99
    "10000001", -- 4478 - 0x117e  :  129 - 0x81
    "11000011", -- 4479 - 0x117f  :  195 - 0xc3
    "01110111", -- 4480 - 0x1180  :  119 - 0x77 -- Background 0x18
    "01110111", -- 4481 - 0x1181  :  119 - 0x77
    "01110111", -- 4482 - 0x1182  :  119 - 0x77
    "01111111", -- 4483 - 0x1183  :  127 - 0x7f
    "01111111", -- 4484 - 0x1184  :  127 - 0x7f
    "01110111", -- 4485 - 0x1185  :  119 - 0x77
    "01110111", -- 4486 - 0x1186  :  119 - 0x77
    "01110111", -- 4487 - 0x1187  :  119 - 0x77
    "10011001", -- 4488 - 0x1188  :  153 - 0x99
    "10011001", -- 4489 - 0x1189  :  153 - 0x99
    "10011001", -- 4490 - 0x118a  :  153 - 0x99
    "10000001", -- 4491 - 0x118b  :  129 - 0x81
    "10000001", -- 4492 - 0x118c  :  129 - 0x81
    "10011001", -- 4493 - 0x118d  :  153 - 0x99
    "10011001", -- 4494 - 0x118e  :  153 - 0x99
    "10011001", -- 4495 - 0x118f  :  153 - 0x99
    "00111110", -- 4496 - 0x1190  :   62 - 0x3e -- Background 0x19
    "00111110", -- 4497 - 0x1191  :   62 - 0x3e
    "00011100", -- 4498 - 0x1192  :   28 - 0x1c
    "00011100", -- 4499 - 0x1193  :   28 - 0x1c
    "00011100", -- 4500 - 0x1194  :   28 - 0x1c
    "00011100", -- 4501 - 0x1195  :   28 - 0x1c
    "00111110", -- 4502 - 0x1196  :   62 - 0x3e
    "00111110", -- 4503 - 0x1197  :   62 - 0x3e
    "11000011", -- 4504 - 0x1198  :  195 - 0xc3
    "11000011", -- 4505 - 0x1199  :  195 - 0xc3
    "11100111", -- 4506 - 0x119a  :  231 - 0xe7
    "11100111", -- 4507 - 0x119b  :  231 - 0xe7
    "11100111", -- 4508 - 0x119c  :  231 - 0xe7
    "11100111", -- 4509 - 0x119d  :  231 - 0xe7
    "11000011", -- 4510 - 0x119e  :  195 - 0xc3
    "11000011", -- 4511 - 0x119f  :  195 - 0xc3
    "00000111", -- 4512 - 0x11a0  :    7 - 0x7 -- Background 0x1a
    "00000111", -- 4513 - 0x11a1  :    7 - 0x7
    "00000111", -- 4514 - 0x11a2  :    7 - 0x7
    "00000111", -- 4515 - 0x11a3  :    7 - 0x7
    "00000111", -- 4516 - 0x11a4  :    7 - 0x7
    "01110111", -- 4517 - 0x11a5  :  119 - 0x77
    "01111111", -- 4518 - 0x11a6  :  127 - 0x7f
    "00111110", -- 4519 - 0x11a7  :   62 - 0x3e
    "11111001", -- 4520 - 0x11a8  :  249 - 0xf9
    "11111001", -- 4521 - 0x11a9  :  249 - 0xf9
    "11111001", -- 4522 - 0x11aa  :  249 - 0xf9
    "11111001", -- 4523 - 0x11ab  :  249 - 0xf9
    "11111001", -- 4524 - 0x11ac  :  249 - 0xf9
    "10011001", -- 4525 - 0x11ad  :  153 - 0x99
    "10000001", -- 4526 - 0x11ae  :  129 - 0x81
    "11000011", -- 4527 - 0x11af  :  195 - 0xc3
    "01110011", -- 4528 - 0x11b0  :  115 - 0x73 -- Background 0x1b
    "01110111", -- 4529 - 0x11b1  :  119 - 0x77
    "01111110", -- 4530 - 0x11b2  :  126 - 0x7e
    "01111100", -- 4531 - 0x11b3  :  124 - 0x7c
    "01111110", -- 4532 - 0x11b4  :  126 - 0x7e
    "01110111", -- 4533 - 0x11b5  :  119 - 0x77
    "01110111", -- 4534 - 0x11b6  :  119 - 0x77
    "01110111", -- 4535 - 0x11b7  :  119 - 0x77
    "10011101", -- 4536 - 0x11b8  :  157 - 0x9d
    "10011001", -- 4537 - 0x11b9  :  153 - 0x99
    "10010011", -- 4538 - 0x11ba  :  147 - 0x93
    "10000111", -- 4539 - 0x11bb  :  135 - 0x87
    "10000011", -- 4540 - 0x11bc  :  131 - 0x83
    "10011001", -- 4541 - 0x11bd  :  153 - 0x99
    "10011001", -- 4542 - 0x11be  :  153 - 0x99
    "10011001", -- 4543 - 0x11bf  :  153 - 0x99
    "01110000", -- 4544 - 0x11c0  :  112 - 0x70 -- Background 0x1c
    "01110000", -- 4545 - 0x11c1  :  112 - 0x70
    "01110000", -- 4546 - 0x11c2  :  112 - 0x70
    "01110000", -- 4547 - 0x11c3  :  112 - 0x70
    "01110000", -- 4548 - 0x11c4  :  112 - 0x70
    "01110000", -- 4549 - 0x11c5  :  112 - 0x70
    "01111111", -- 4550 - 0x11c6  :  127 - 0x7f
    "01111111", -- 4551 - 0x11c7  :  127 - 0x7f
    "10011111", -- 4552 - 0x11c8  :  159 - 0x9f
    "10011111", -- 4553 - 0x11c9  :  159 - 0x9f
    "10011111", -- 4554 - 0x11ca  :  159 - 0x9f
    "10011111", -- 4555 - 0x11cb  :  159 - 0x9f
    "10011111", -- 4556 - 0x11cc  :  159 - 0x9f
    "10011111", -- 4557 - 0x11cd  :  159 - 0x9f
    "10000001", -- 4558 - 0x11ce  :  129 - 0x81
    "10000001", -- 4559 - 0x11cf  :  129 - 0x81
    "11100111", -- 4560 - 0x11d0  :  231 - 0xe7 -- Background 0x1d
    "11111111", -- 4561 - 0x11d1  :  255 - 0xff
    "11111111", -- 4562 - 0x11d2  :  255 - 0xff
    "11111111", -- 4563 - 0x11d3  :  255 - 0xff
    "11111111", -- 4564 - 0x11d4  :  255 - 0xff
    "11100111", -- 4565 - 0x11d5  :  231 - 0xe7
    "11100111", -- 4566 - 0x11d6  :  231 - 0xe7
    "11100111", -- 4567 - 0x11d7  :  231 - 0xe7
    "00111001", -- 4568 - 0x11d8  :   57 - 0x39
    "00010001", -- 4569 - 0x11d9  :   17 - 0x11
    "00000001", -- 4570 - 0x11da  :    1 - 0x1
    "00000001", -- 4571 - 0x11db  :    1 - 0x1
    "00101001", -- 4572 - 0x11dc  :   41 - 0x29
    "00111001", -- 4573 - 0x11dd  :   57 - 0x39
    "00111001", -- 4574 - 0x11de  :   57 - 0x39
    "00111001", -- 4575 - 0x11df  :   57 - 0x39
    "01110111", -- 4576 - 0x11e0  :  119 - 0x77 -- Background 0x1e
    "01110111", -- 4577 - 0x11e1  :  119 - 0x77
    "01111111", -- 4578 - 0x11e2  :  127 - 0x7f
    "01111111", -- 4579 - 0x11e3  :  127 - 0x7f
    "01111111", -- 4580 - 0x11e4  :  127 - 0x7f
    "01111111", -- 4581 - 0x11e5  :  127 - 0x7f
    "01110111", -- 4582 - 0x11e6  :  119 - 0x77
    "01110111", -- 4583 - 0x11e7  :  119 - 0x77
    "10011001", -- 4584 - 0x11e8  :  153 - 0x99
    "10011001", -- 4585 - 0x11e9  :  153 - 0x99
    "10001001", -- 4586 - 0x11ea  :  137 - 0x89
    "10000001", -- 4587 - 0x11eb  :  129 - 0x81
    "10000001", -- 4588 - 0x11ec  :  129 - 0x81
    "10010001", -- 4589 - 0x11ed  :  145 - 0x91
    "10011001", -- 4590 - 0x11ee  :  153 - 0x99
    "10011001", -- 4591 - 0x11ef  :  153 - 0x99
    "00111100", -- 4592 - 0x11f0  :   60 - 0x3c -- Background 0x1f
    "01111110", -- 4593 - 0x11f1  :  126 - 0x7e
    "11100111", -- 4594 - 0x11f2  :  231 - 0xe7
    "11100111", -- 4595 - 0x11f3  :  231 - 0xe7
    "11100111", -- 4596 - 0x11f4  :  231 - 0xe7
    "11100111", -- 4597 - 0x11f5  :  231 - 0xe7
    "01111110", -- 4598 - 0x11f6  :  126 - 0x7e
    "00111100", -- 4599 - 0x11f7  :   60 - 0x3c
    "11000111", -- 4600 - 0x11f8  :  199 - 0xc7
    "10000011", -- 4601 - 0x11f9  :  131 - 0x83
    "00111001", -- 4602 - 0x11fa  :   57 - 0x39
    "00111001", -- 4603 - 0x11fb  :   57 - 0x39
    "00111001", -- 4604 - 0x11fc  :   57 - 0x39
    "00111001", -- 4605 - 0x11fd  :   57 - 0x39
    "10000011", -- 4606 - 0x11fe  :  131 - 0x83
    "11000111", -- 4607 - 0x11ff  :  199 - 0xc7
    "01111110", -- 4608 - 0x1200  :  126 - 0x7e -- Background 0x20
    "01111111", -- 4609 - 0x1201  :  127 - 0x7f
    "01110111", -- 4610 - 0x1202  :  119 - 0x77
    "01110111", -- 4611 - 0x1203  :  119 - 0x77
    "01111111", -- 4612 - 0x1204  :  127 - 0x7f
    "01111110", -- 4613 - 0x1205  :  126 - 0x7e
    "01110000", -- 4614 - 0x1206  :  112 - 0x70
    "01110000", -- 4615 - 0x1207  :  112 - 0x70
    "10000011", -- 4616 - 0x1208  :  131 - 0x83
    "10000001", -- 4617 - 0x1209  :  129 - 0x81
    "10011001", -- 4618 - 0x120a  :  153 - 0x99
    "10011001", -- 4619 - 0x120b  :  153 - 0x99
    "10000001", -- 4620 - 0x120c  :  129 - 0x81
    "10000011", -- 4621 - 0x120d  :  131 - 0x83
    "10011111", -- 4622 - 0x120e  :  159 - 0x9f
    "10011111", -- 4623 - 0x120f  :  159 - 0x9f
    "00111100", -- 4624 - 0x1210  :   60 - 0x3c -- Background 0x21
    "01111110", -- 4625 - 0x1211  :  126 - 0x7e
    "11100111", -- 4626 - 0x1212  :  231 - 0xe7
    "11100111", -- 4627 - 0x1213  :  231 - 0xe7
    "11100111", -- 4628 - 0x1214  :  231 - 0xe7
    "11101110", -- 4629 - 0x1215  :  238 - 0xee
    "01111111", -- 4630 - 0x1216  :  127 - 0x7f
    "00111111", -- 4631 - 0x1217  :   63 - 0x3f
    "11000111", -- 4632 - 0x1218  :  199 - 0xc7
    "10000011", -- 4633 - 0x1219  :  131 - 0x83
    "00111001", -- 4634 - 0x121a  :   57 - 0x39
    "00111001", -- 4635 - 0x121b  :   57 - 0x39
    "00111001", -- 4636 - 0x121c  :   57 - 0x39
    "00110011", -- 4637 - 0x121d  :   51 - 0x33
    "10000001", -- 4638 - 0x121e  :  129 - 0x81
    "11001001", -- 4639 - 0x121f  :  201 - 0xc9
    "01111110", -- 4640 - 0x1220  :  126 - 0x7e -- Background 0x22
    "01111111", -- 4641 - 0x1221  :  127 - 0x7f
    "01110111", -- 4642 - 0x1222  :  119 - 0x77
    "01110111", -- 4643 - 0x1223  :  119 - 0x77
    "01111111", -- 4644 - 0x1224  :  127 - 0x7f
    "01111110", -- 4645 - 0x1225  :  126 - 0x7e
    "01110111", -- 4646 - 0x1226  :  119 - 0x77
    "01110111", -- 4647 - 0x1227  :  119 - 0x77
    "10000011", -- 4648 - 0x1228  :  131 - 0x83
    "10000001", -- 4649 - 0x1229  :  129 - 0x81
    "10011001", -- 4650 - 0x122a  :  153 - 0x99
    "10011001", -- 4651 - 0x122b  :  153 - 0x99
    "10000001", -- 4652 - 0x122c  :  129 - 0x81
    "10000011", -- 4653 - 0x122d  :  131 - 0x83
    "10011001", -- 4654 - 0x122e  :  153 - 0x99
    "10011001", -- 4655 - 0x122f  :  153 - 0x99
    "00111110", -- 4656 - 0x1230  :   62 - 0x3e -- Background 0x23
    "01111111", -- 4657 - 0x1231  :  127 - 0x7f
    "01110000", -- 4658 - 0x1232  :  112 - 0x70
    "01111110", -- 4659 - 0x1233  :  126 - 0x7e
    "00111111", -- 4660 - 0x1234  :   63 - 0x3f
    "00000111", -- 4661 - 0x1235  :    7 - 0x7
    "01111111", -- 4662 - 0x1236  :  127 - 0x7f
    "00111110", -- 4663 - 0x1237  :   62 - 0x3e
    "11000011", -- 4664 - 0x1238  :  195 - 0xc3
    "10000001", -- 4665 - 0x1239  :  129 - 0x81
    "10011111", -- 4666 - 0x123a  :  159 - 0x9f
    "10000011", -- 4667 - 0x123b  :  131 - 0x83
    "11000001", -- 4668 - 0x123c  :  193 - 0xc1
    "11111001", -- 4669 - 0x123d  :  249 - 0xf9
    "10000001", -- 4670 - 0x123e  :  129 - 0x81
    "11000011", -- 4671 - 0x123f  :  195 - 0xc3
    "01111111", -- 4672 - 0x1240  :  127 - 0x7f -- Background 0x24
    "01111111", -- 4673 - 0x1241  :  127 - 0x7f
    "00011100", -- 4674 - 0x1242  :   28 - 0x1c
    "00011100", -- 4675 - 0x1243  :   28 - 0x1c
    "00011100", -- 4676 - 0x1244  :   28 - 0x1c
    "00011100", -- 4677 - 0x1245  :   28 - 0x1c
    "00011100", -- 4678 - 0x1246  :   28 - 0x1c
    "00011100", -- 4679 - 0x1247  :   28 - 0x1c
    "10000001", -- 4680 - 0x1248  :  129 - 0x81
    "10000001", -- 4681 - 0x1249  :  129 - 0x81
    "11100111", -- 4682 - 0x124a  :  231 - 0xe7
    "11100111", -- 4683 - 0x124b  :  231 - 0xe7
    "11100111", -- 4684 - 0x124c  :  231 - 0xe7
    "11100111", -- 4685 - 0x124d  :  231 - 0xe7
    "11100111", -- 4686 - 0x124e  :  231 - 0xe7
    "11100111", -- 4687 - 0x124f  :  231 - 0xe7
    "01110111", -- 4688 - 0x1250  :  119 - 0x77 -- Background 0x25
    "01110111", -- 4689 - 0x1251  :  119 - 0x77
    "01110111", -- 4690 - 0x1252  :  119 - 0x77
    "01110111", -- 4691 - 0x1253  :  119 - 0x77
    "01110111", -- 4692 - 0x1254  :  119 - 0x77
    "01110111", -- 4693 - 0x1255  :  119 - 0x77
    "01111111", -- 4694 - 0x1256  :  127 - 0x7f
    "00111110", -- 4695 - 0x1257  :   62 - 0x3e
    "10011001", -- 4696 - 0x1258  :  153 - 0x99
    "10011001", -- 4697 - 0x1259  :  153 - 0x99
    "10011001", -- 4698 - 0x125a  :  153 - 0x99
    "10011001", -- 4699 - 0x125b  :  153 - 0x99
    "10011001", -- 4700 - 0x125c  :  153 - 0x99
    "10011001", -- 4701 - 0x125d  :  153 - 0x99
    "10000001", -- 4702 - 0x125e  :  129 - 0x81
    "11000011", -- 4703 - 0x125f  :  195 - 0xc3
    "01110111", -- 4704 - 0x1260  :  119 - 0x77 -- Background 0x26
    "01110111", -- 4705 - 0x1261  :  119 - 0x77
    "01110111", -- 4706 - 0x1262  :  119 - 0x77
    "01110111", -- 4707 - 0x1263  :  119 - 0x77
    "01110111", -- 4708 - 0x1264  :  119 - 0x77
    "01110111", -- 4709 - 0x1265  :  119 - 0x77
    "00111110", -- 4710 - 0x1266  :   62 - 0x3e
    "00011100", -- 4711 - 0x1267  :   28 - 0x1c
    "10011001", -- 4712 - 0x1268  :  153 - 0x99
    "10011001", -- 4713 - 0x1269  :  153 - 0x99
    "10011001", -- 4714 - 0x126a  :  153 - 0x99
    "10011001", -- 4715 - 0x126b  :  153 - 0x99
    "10011001", -- 4716 - 0x126c  :  153 - 0x99
    "10011001", -- 4717 - 0x126d  :  153 - 0x99
    "11000011", -- 4718 - 0x126e  :  195 - 0xc3
    "11100111", -- 4719 - 0x126f  :  231 - 0xe7
    "11100111", -- 4720 - 0x1270  :  231 - 0xe7 -- Background 0x27
    "11100111", -- 4721 - 0x1271  :  231 - 0xe7
    "11100111", -- 4722 - 0x1272  :  231 - 0xe7
    "11100111", -- 4723 - 0x1273  :  231 - 0xe7
    "11110111", -- 4724 - 0x1274  :  247 - 0xf7
    "11111111", -- 4725 - 0x1275  :  255 - 0xff
    "11111111", -- 4726 - 0x1276  :  255 - 0xff
    "01111110", -- 4727 - 0x1277  :  126 - 0x7e
    "00111001", -- 4728 - 0x1278  :   57 - 0x39
    "00111001", -- 4729 - 0x1279  :   57 - 0x39
    "00111001", -- 4730 - 0x127a  :   57 - 0x39
    "00111001", -- 4731 - 0x127b  :   57 - 0x39
    "00101001", -- 4732 - 0x127c  :   41 - 0x29
    "00000001", -- 4733 - 0x127d  :    1 - 0x1
    "00000001", -- 4734 - 0x127e  :    1 - 0x1
    "10010011", -- 4735 - 0x127f  :  147 - 0x93
    "01110111", -- 4736 - 0x1280  :  119 - 0x77 -- Background 0x28
    "01110111", -- 4737 - 0x1281  :  119 - 0x77
    "01110111", -- 4738 - 0x1282  :  119 - 0x77
    "00111110", -- 4739 - 0x1283  :   62 - 0x3e
    "00111110", -- 4740 - 0x1284  :   62 - 0x3e
    "01110111", -- 4741 - 0x1285  :  119 - 0x77
    "01110111", -- 4742 - 0x1286  :  119 - 0x77
    "01110111", -- 4743 - 0x1287  :  119 - 0x77
    "10011001", -- 4744 - 0x1288  :  153 - 0x99
    "10011001", -- 4745 - 0x1289  :  153 - 0x99
    "10011001", -- 4746 - 0x128a  :  153 - 0x99
    "11000011", -- 4747 - 0x128b  :  195 - 0xc3
    "11000011", -- 4748 - 0x128c  :  195 - 0xc3
    "10011001", -- 4749 - 0x128d  :  153 - 0x99
    "10011001", -- 4750 - 0x128e  :  153 - 0x99
    "10011001", -- 4751 - 0x128f  :  153 - 0x99
    "01110111", -- 4752 - 0x1290  :  119 - 0x77 -- Background 0x29
    "01110111", -- 4753 - 0x1291  :  119 - 0x77
    "01110111", -- 4754 - 0x1292  :  119 - 0x77
    "01111111", -- 4755 - 0x1293  :  127 - 0x7f
    "00111110", -- 4756 - 0x1294  :   62 - 0x3e
    "00011100", -- 4757 - 0x1295  :   28 - 0x1c
    "00011100", -- 4758 - 0x1296  :   28 - 0x1c
    "00011100", -- 4759 - 0x1297  :   28 - 0x1c
    "10011001", -- 4760 - 0x1298  :  153 - 0x99
    "10011001", -- 4761 - 0x1299  :  153 - 0x99
    "10011001", -- 4762 - 0x129a  :  153 - 0x99
    "10000001", -- 4763 - 0x129b  :  129 - 0x81
    "11000011", -- 4764 - 0x129c  :  195 - 0xc3
    "11100111", -- 4765 - 0x129d  :  231 - 0xe7
    "11100111", -- 4766 - 0x129e  :  231 - 0xe7
    "11100111", -- 4767 - 0x129f  :  231 - 0xe7
    "01111111", -- 4768 - 0x12a0  :  127 - 0x7f -- Background 0x2a
    "01111111", -- 4769 - 0x12a1  :  127 - 0x7f
    "00001110", -- 4770 - 0x12a2  :   14 - 0xe
    "00011100", -- 4771 - 0x12a3  :   28 - 0x1c
    "00011100", -- 4772 - 0x12a4  :   28 - 0x1c
    "00111000", -- 4773 - 0x12a5  :   56 - 0x38
    "01111111", -- 4774 - 0x12a6  :  127 - 0x7f
    "01111111", -- 4775 - 0x12a7  :  127 - 0x7f
    "10000001", -- 4776 - 0x12a8  :  129 - 0x81
    "10000001", -- 4777 - 0x12a9  :  129 - 0x81
    "11110011", -- 4778 - 0x12aa  :  243 - 0xf3
    "11100111", -- 4779 - 0x12ab  :  231 - 0xe7
    "11100111", -- 4780 - 0x12ac  :  231 - 0xe7
    "11001111", -- 4781 - 0x12ad  :  207 - 0xcf
    "10000001", -- 4782 - 0x12ae  :  129 - 0x81
    "10000001", -- 4783 - 0x12af  :  129 - 0x81
    "00111110", -- 4784 - 0x12b0  :   62 - 0x3e -- Background 0x2b
    "01100011", -- 4785 - 0x12b1  :   99 - 0x63
    "01101111", -- 4786 - 0x12b2  :  111 - 0x6f
    "01111111", -- 4787 - 0x12b3  :  127 - 0x7f
    "01111111", -- 4788 - 0x12b4  :  127 - 0x7f
    "01111110", -- 4789 - 0x12b5  :  126 - 0x7e
    "01100000", -- 4790 - 0x12b6  :   96 - 0x60
    "00111111", -- 4791 - 0x12b7  :   63 - 0x3f
    "11000011", -- 4792 - 0x12b8  :  195 - 0xc3
    "10111101", -- 4793 - 0x12b9  :  189 - 0xbd
    "10110101", -- 4794 - 0x12ba  :  181 - 0xb5
    "10101001", -- 4795 - 0x12bb  :  169 - 0xa9
    "10101001", -- 4796 - 0x12bc  :  169 - 0xa9
    "10100011", -- 4797 - 0x12bd  :  163 - 0xa3
    "10111111", -- 4798 - 0x12be  :  191 - 0xbf
    "11000001", -- 4799 - 0x12bf  :  193 - 0xc1
    "00000000", -- 4800 - 0x12c0  :    0 - 0x0 -- Background 0x2c
    "01110000", -- 4801 - 0x12c1  :  112 - 0x70
    "01111100", -- 4802 - 0x12c2  :  124 - 0x7c
    "01111111", -- 4803 - 0x12c3  :  127 - 0x7f
    "01111111", -- 4804 - 0x12c4  :  127 - 0x7f
    "01111100", -- 4805 - 0x12c5  :  124 - 0x7c
    "01110000", -- 4806 - 0x12c6  :  112 - 0x70
    "00000000", -- 4807 - 0x12c7  :    0 - 0x0
    "11111111", -- 4808 - 0x12c8  :  255 - 0xff
    "10011111", -- 4809 - 0x12c9  :  159 - 0x9f
    "10000111", -- 4810 - 0x12ca  :  135 - 0x87
    "10000001", -- 4811 - 0x12cb  :  129 - 0x81
    "10000001", -- 4812 - 0x12cc  :  129 - 0x81
    "10000111", -- 4813 - 0x12cd  :  135 - 0x87
    "10011111", -- 4814 - 0x12ce  :  159 - 0x9f
    "11111111", -- 4815 - 0x12cf  :  255 - 0xff
    "00000000", -- 4816 - 0x12d0  :    0 - 0x0 -- Background 0x2d
    "01110000", -- 4817 - 0x12d1  :  112 - 0x70
    "01110000", -- 4818 - 0x12d2  :  112 - 0x70
    "00000000", -- 4819 - 0x12d3  :    0 - 0x0
    "00000000", -- 4820 - 0x12d4  :    0 - 0x0
    "01110000", -- 4821 - 0x12d5  :  112 - 0x70
    "01110000", -- 4822 - 0x12d6  :  112 - 0x70
    "00000000", -- 4823 - 0x12d7  :    0 - 0x0
    "11111111", -- 4824 - 0x12d8  :  255 - 0xff
    "10011111", -- 4825 - 0x12d9  :  159 - 0x9f
    "10011111", -- 4826 - 0x12da  :  159 - 0x9f
    "11111111", -- 4827 - 0x12db  :  255 - 0xff
    "11111111", -- 4828 - 0x12dc  :  255 - 0xff
    "10011111", -- 4829 - 0x12dd  :  159 - 0x9f
    "10011111", -- 4830 - 0x12de  :  159 - 0x9f
    "11111111", -- 4831 - 0x12df  :  255 - 0xff
    "00000000", -- 4832 - 0x12e0  :    0 - 0x0 -- Background 0x2e
    "00000000", -- 4833 - 0x12e1  :    0 - 0x0
    "00000000", -- 4834 - 0x12e2  :    0 - 0x0
    "00000000", -- 4835 - 0x12e3  :    0 - 0x0
    "00000000", -- 4836 - 0x12e4  :    0 - 0x0
    "00000000", -- 4837 - 0x12e5  :    0 - 0x0
    "00000000", -- 4838 - 0x12e6  :    0 - 0x0
    "00000000", -- 4839 - 0x12e7  :    0 - 0x0
    "00000000", -- 4840 - 0x12e8  :    0 - 0x0
    "00000000", -- 4841 - 0x12e9  :    0 - 0x0
    "00000000", -- 4842 - 0x12ea  :    0 - 0x0
    "00000000", -- 4843 - 0x12eb  :    0 - 0x0
    "00000000", -- 4844 - 0x12ec  :    0 - 0x0
    "00000000", -- 4845 - 0x12ed  :    0 - 0x0
    "00000000", -- 4846 - 0x12ee  :    0 - 0x0
    "00000000", -- 4847 - 0x12ef  :    0 - 0x0
    "00000000", -- 4848 - 0x12f0  :    0 - 0x0 -- Background 0x2f
    "00000000", -- 4849 - 0x12f1  :    0 - 0x0
    "00000000", -- 4850 - 0x12f2  :    0 - 0x0
    "00000000", -- 4851 - 0x12f3  :    0 - 0x0
    "00000000", -- 4852 - 0x12f4  :    0 - 0x0
    "00000000", -- 4853 - 0x12f5  :    0 - 0x0
    "00000000", -- 4854 - 0x12f6  :    0 - 0x0
    "00000000", -- 4855 - 0x12f7  :    0 - 0x0
    "00000000", -- 4856 - 0x12f8  :    0 - 0x0
    "00000000", -- 4857 - 0x12f9  :    0 - 0x0
    "00000000", -- 4858 - 0x12fa  :    0 - 0x0
    "00000000", -- 4859 - 0x12fb  :    0 - 0x0
    "00000000", -- 4860 - 0x12fc  :    0 - 0x0
    "00000000", -- 4861 - 0x12fd  :    0 - 0x0
    "00000000", -- 4862 - 0x12fe  :    0 - 0x0
    "00000000", -- 4863 - 0x12ff  :    0 - 0x0
    "00000000", -- 4864 - 0x1300  :    0 - 0x0 -- Background 0x30
    "00000000", -- 4865 - 0x1301  :    0 - 0x0
    "00000000", -- 4866 - 0x1302  :    0 - 0x0
    "00000000", -- 4867 - 0x1303  :    0 - 0x0
    "00000000", -- 4868 - 0x1304  :    0 - 0x0
    "00000000", -- 4869 - 0x1305  :    0 - 0x0
    "00000000", -- 4870 - 0x1306  :    0 - 0x0
    "00000000", -- 4871 - 0x1307  :    0 - 0x0
    "00000000", -- 4872 - 0x1308  :    0 - 0x0
    "00000000", -- 4873 - 0x1309  :    0 - 0x0
    "00000000", -- 4874 - 0x130a  :    0 - 0x0
    "00000000", -- 4875 - 0x130b  :    0 - 0x0
    "00000000", -- 4876 - 0x130c  :    0 - 0x0
    "00000000", -- 4877 - 0x130d  :    0 - 0x0
    "00000000", -- 4878 - 0x130e  :    0 - 0x0
    "00000000", -- 4879 - 0x130f  :    0 - 0x0
    "00000000", -- 4880 - 0x1310  :    0 - 0x0 -- Background 0x31
    "00000000", -- 4881 - 0x1311  :    0 - 0x0
    "00000000", -- 4882 - 0x1312  :    0 - 0x0
    "00000000", -- 4883 - 0x1313  :    0 - 0x0
    "00000000", -- 4884 - 0x1314  :    0 - 0x0
    "00000000", -- 4885 - 0x1315  :    0 - 0x0
    "00000000", -- 4886 - 0x1316  :    0 - 0x0
    "00000000", -- 4887 - 0x1317  :    0 - 0x0
    "00000000", -- 4888 - 0x1318  :    0 - 0x0
    "00000000", -- 4889 - 0x1319  :    0 - 0x0
    "00000000", -- 4890 - 0x131a  :    0 - 0x0
    "00000000", -- 4891 - 0x131b  :    0 - 0x0
    "00000000", -- 4892 - 0x131c  :    0 - 0x0
    "00000000", -- 4893 - 0x131d  :    0 - 0x0
    "00000000", -- 4894 - 0x131e  :    0 - 0x0
    "00000000", -- 4895 - 0x131f  :    0 - 0x0
    "00000000", -- 4896 - 0x1320  :    0 - 0x0 -- Background 0x32
    "00000000", -- 4897 - 0x1321  :    0 - 0x0
    "00000000", -- 4898 - 0x1322  :    0 - 0x0
    "00000000", -- 4899 - 0x1323  :    0 - 0x0
    "00000000", -- 4900 - 0x1324  :    0 - 0x0
    "00000000", -- 4901 - 0x1325  :    0 - 0x0
    "00000000", -- 4902 - 0x1326  :    0 - 0x0
    "00000000", -- 4903 - 0x1327  :    0 - 0x0
    "00000000", -- 4904 - 0x1328  :    0 - 0x0
    "00000000", -- 4905 - 0x1329  :    0 - 0x0
    "00000000", -- 4906 - 0x132a  :    0 - 0x0
    "00000000", -- 4907 - 0x132b  :    0 - 0x0
    "00000000", -- 4908 - 0x132c  :    0 - 0x0
    "00000000", -- 4909 - 0x132d  :    0 - 0x0
    "00000000", -- 4910 - 0x132e  :    0 - 0x0
    "00000000", -- 4911 - 0x132f  :    0 - 0x0
    "00000000", -- 4912 - 0x1330  :    0 - 0x0 -- Background 0x33
    "00000000", -- 4913 - 0x1331  :    0 - 0x0
    "00000000", -- 4914 - 0x1332  :    0 - 0x0
    "00000000", -- 4915 - 0x1333  :    0 - 0x0
    "00000000", -- 4916 - 0x1334  :    0 - 0x0
    "00000000", -- 4917 - 0x1335  :    0 - 0x0
    "00000000", -- 4918 - 0x1336  :    0 - 0x0
    "00000000", -- 4919 - 0x1337  :    0 - 0x0
    "00000000", -- 4920 - 0x1338  :    0 - 0x0
    "00000000", -- 4921 - 0x1339  :    0 - 0x0
    "00000000", -- 4922 - 0x133a  :    0 - 0x0
    "00000000", -- 4923 - 0x133b  :    0 - 0x0
    "00000000", -- 4924 - 0x133c  :    0 - 0x0
    "00000000", -- 4925 - 0x133d  :    0 - 0x0
    "00000000", -- 4926 - 0x133e  :    0 - 0x0
    "00000000", -- 4927 - 0x133f  :    0 - 0x0
    "00000000", -- 4928 - 0x1340  :    0 - 0x0 -- Background 0x34
    "00000000", -- 4929 - 0x1341  :    0 - 0x0
    "00000000", -- 4930 - 0x1342  :    0 - 0x0
    "00000000", -- 4931 - 0x1343  :    0 - 0x0
    "00000000", -- 4932 - 0x1344  :    0 - 0x0
    "00000000", -- 4933 - 0x1345  :    0 - 0x0
    "00000000", -- 4934 - 0x1346  :    0 - 0x0
    "00000000", -- 4935 - 0x1347  :    0 - 0x0
    "00000000", -- 4936 - 0x1348  :    0 - 0x0
    "00000000", -- 4937 - 0x1349  :    0 - 0x0
    "00000000", -- 4938 - 0x134a  :    0 - 0x0
    "00000000", -- 4939 - 0x134b  :    0 - 0x0
    "00000000", -- 4940 - 0x134c  :    0 - 0x0
    "00000000", -- 4941 - 0x134d  :    0 - 0x0
    "00000000", -- 4942 - 0x134e  :    0 - 0x0
    "00000000", -- 4943 - 0x134f  :    0 - 0x0
    "00000000", -- 4944 - 0x1350  :    0 - 0x0 -- Background 0x35
    "00000000", -- 4945 - 0x1351  :    0 - 0x0
    "00000000", -- 4946 - 0x1352  :    0 - 0x0
    "00000000", -- 4947 - 0x1353  :    0 - 0x0
    "00000000", -- 4948 - 0x1354  :    0 - 0x0
    "00000000", -- 4949 - 0x1355  :    0 - 0x0
    "00000000", -- 4950 - 0x1356  :    0 - 0x0
    "00000000", -- 4951 - 0x1357  :    0 - 0x0
    "00000000", -- 4952 - 0x1358  :    0 - 0x0
    "00000000", -- 4953 - 0x1359  :    0 - 0x0
    "00000000", -- 4954 - 0x135a  :    0 - 0x0
    "00000000", -- 4955 - 0x135b  :    0 - 0x0
    "00000000", -- 4956 - 0x135c  :    0 - 0x0
    "00000000", -- 4957 - 0x135d  :    0 - 0x0
    "00000000", -- 4958 - 0x135e  :    0 - 0x0
    "00000000", -- 4959 - 0x135f  :    0 - 0x0
    "00000000", -- 4960 - 0x1360  :    0 - 0x0 -- Background 0x36
    "00000000", -- 4961 - 0x1361  :    0 - 0x0
    "00000000", -- 4962 - 0x1362  :    0 - 0x0
    "00000000", -- 4963 - 0x1363  :    0 - 0x0
    "00000000", -- 4964 - 0x1364  :    0 - 0x0
    "00000000", -- 4965 - 0x1365  :    0 - 0x0
    "00000000", -- 4966 - 0x1366  :    0 - 0x0
    "00000000", -- 4967 - 0x1367  :    0 - 0x0
    "00000000", -- 4968 - 0x1368  :    0 - 0x0
    "00000000", -- 4969 - 0x1369  :    0 - 0x0
    "00000000", -- 4970 - 0x136a  :    0 - 0x0
    "00000000", -- 4971 - 0x136b  :    0 - 0x0
    "00000000", -- 4972 - 0x136c  :    0 - 0x0
    "00000000", -- 4973 - 0x136d  :    0 - 0x0
    "00000000", -- 4974 - 0x136e  :    0 - 0x0
    "00000000", -- 4975 - 0x136f  :    0 - 0x0
    "00000000", -- 4976 - 0x1370  :    0 - 0x0 -- Background 0x37
    "00000000", -- 4977 - 0x1371  :    0 - 0x0
    "00000000", -- 4978 - 0x1372  :    0 - 0x0
    "00000000", -- 4979 - 0x1373  :    0 - 0x0
    "00000000", -- 4980 - 0x1374  :    0 - 0x0
    "00000000", -- 4981 - 0x1375  :    0 - 0x0
    "00000000", -- 4982 - 0x1376  :    0 - 0x0
    "00000000", -- 4983 - 0x1377  :    0 - 0x0
    "00000000", -- 4984 - 0x1378  :    0 - 0x0
    "00000000", -- 4985 - 0x1379  :    0 - 0x0
    "00000000", -- 4986 - 0x137a  :    0 - 0x0
    "00000000", -- 4987 - 0x137b  :    0 - 0x0
    "00000000", -- 4988 - 0x137c  :    0 - 0x0
    "00000000", -- 4989 - 0x137d  :    0 - 0x0
    "00000000", -- 4990 - 0x137e  :    0 - 0x0
    "00000000", -- 4991 - 0x137f  :    0 - 0x0
    "00000000", -- 4992 - 0x1380  :    0 - 0x0 -- Background 0x38
    "00000000", -- 4993 - 0x1381  :    0 - 0x0
    "00000000", -- 4994 - 0x1382  :    0 - 0x0
    "00000000", -- 4995 - 0x1383  :    0 - 0x0
    "00000000", -- 4996 - 0x1384  :    0 - 0x0
    "00000000", -- 4997 - 0x1385  :    0 - 0x0
    "00000000", -- 4998 - 0x1386  :    0 - 0x0
    "00000000", -- 4999 - 0x1387  :    0 - 0x0
    "00000000", -- 5000 - 0x1388  :    0 - 0x0
    "00000000", -- 5001 - 0x1389  :    0 - 0x0
    "00000000", -- 5002 - 0x138a  :    0 - 0x0
    "00000000", -- 5003 - 0x138b  :    0 - 0x0
    "00000000", -- 5004 - 0x138c  :    0 - 0x0
    "00000000", -- 5005 - 0x138d  :    0 - 0x0
    "00000000", -- 5006 - 0x138e  :    0 - 0x0
    "00000000", -- 5007 - 0x138f  :    0 - 0x0
    "00000000", -- 5008 - 0x1390  :    0 - 0x0 -- Background 0x39
    "00000000", -- 5009 - 0x1391  :    0 - 0x0
    "00000000", -- 5010 - 0x1392  :    0 - 0x0
    "00000000", -- 5011 - 0x1393  :    0 - 0x0
    "00000000", -- 5012 - 0x1394  :    0 - 0x0
    "00000000", -- 5013 - 0x1395  :    0 - 0x0
    "00000000", -- 5014 - 0x1396  :    0 - 0x0
    "00000000", -- 5015 - 0x1397  :    0 - 0x0
    "00000000", -- 5016 - 0x1398  :    0 - 0x0
    "00000000", -- 5017 - 0x1399  :    0 - 0x0
    "00000000", -- 5018 - 0x139a  :    0 - 0x0
    "00000000", -- 5019 - 0x139b  :    0 - 0x0
    "00000000", -- 5020 - 0x139c  :    0 - 0x0
    "00000000", -- 5021 - 0x139d  :    0 - 0x0
    "00000000", -- 5022 - 0x139e  :    0 - 0x0
    "00000000", -- 5023 - 0x139f  :    0 - 0x0
    "00000000", -- 5024 - 0x13a0  :    0 - 0x0 -- Background 0x3a
    "00000000", -- 5025 - 0x13a1  :    0 - 0x0
    "00000000", -- 5026 - 0x13a2  :    0 - 0x0
    "00000000", -- 5027 - 0x13a3  :    0 - 0x0
    "00000000", -- 5028 - 0x13a4  :    0 - 0x0
    "00000000", -- 5029 - 0x13a5  :    0 - 0x0
    "00000000", -- 5030 - 0x13a6  :    0 - 0x0
    "00000000", -- 5031 - 0x13a7  :    0 - 0x0
    "00000000", -- 5032 - 0x13a8  :    0 - 0x0
    "00000000", -- 5033 - 0x13a9  :    0 - 0x0
    "00000000", -- 5034 - 0x13aa  :    0 - 0x0
    "00000000", -- 5035 - 0x13ab  :    0 - 0x0
    "00000000", -- 5036 - 0x13ac  :    0 - 0x0
    "00000000", -- 5037 - 0x13ad  :    0 - 0x0
    "00000000", -- 5038 - 0x13ae  :    0 - 0x0
    "00000000", -- 5039 - 0x13af  :    0 - 0x0
    "00000000", -- 5040 - 0x13b0  :    0 - 0x0 -- Background 0x3b
    "00000000", -- 5041 - 0x13b1  :    0 - 0x0
    "00000000", -- 5042 - 0x13b2  :    0 - 0x0
    "00000000", -- 5043 - 0x13b3  :    0 - 0x0
    "00000000", -- 5044 - 0x13b4  :    0 - 0x0
    "00000000", -- 5045 - 0x13b5  :    0 - 0x0
    "00000000", -- 5046 - 0x13b6  :    0 - 0x0
    "00000000", -- 5047 - 0x13b7  :    0 - 0x0
    "00000000", -- 5048 - 0x13b8  :    0 - 0x0
    "00000000", -- 5049 - 0x13b9  :    0 - 0x0
    "00000000", -- 5050 - 0x13ba  :    0 - 0x0
    "00000000", -- 5051 - 0x13bb  :    0 - 0x0
    "00000000", -- 5052 - 0x13bc  :    0 - 0x0
    "00000000", -- 5053 - 0x13bd  :    0 - 0x0
    "00000000", -- 5054 - 0x13be  :    0 - 0x0
    "00000000", -- 5055 - 0x13bf  :    0 - 0x0
    "00000000", -- 5056 - 0x13c0  :    0 - 0x0 -- Background 0x3c
    "00000000", -- 5057 - 0x13c1  :    0 - 0x0
    "00000000", -- 5058 - 0x13c2  :    0 - 0x0
    "00000000", -- 5059 - 0x13c3  :    0 - 0x0
    "00000000", -- 5060 - 0x13c4  :    0 - 0x0
    "00000000", -- 5061 - 0x13c5  :    0 - 0x0
    "00000000", -- 5062 - 0x13c6  :    0 - 0x0
    "00000000", -- 5063 - 0x13c7  :    0 - 0x0
    "00000000", -- 5064 - 0x13c8  :    0 - 0x0
    "00000000", -- 5065 - 0x13c9  :    0 - 0x0
    "00000000", -- 5066 - 0x13ca  :    0 - 0x0
    "00000000", -- 5067 - 0x13cb  :    0 - 0x0
    "00000000", -- 5068 - 0x13cc  :    0 - 0x0
    "00000000", -- 5069 - 0x13cd  :    0 - 0x0
    "00000000", -- 5070 - 0x13ce  :    0 - 0x0
    "00000000", -- 5071 - 0x13cf  :    0 - 0x0
    "00000000", -- 5072 - 0x13d0  :    0 - 0x0 -- Background 0x3d
    "00000000", -- 5073 - 0x13d1  :    0 - 0x0
    "00000000", -- 5074 - 0x13d2  :    0 - 0x0
    "00000000", -- 5075 - 0x13d3  :    0 - 0x0
    "00000000", -- 5076 - 0x13d4  :    0 - 0x0
    "00000000", -- 5077 - 0x13d5  :    0 - 0x0
    "00000000", -- 5078 - 0x13d6  :    0 - 0x0
    "00000000", -- 5079 - 0x13d7  :    0 - 0x0
    "00000000", -- 5080 - 0x13d8  :    0 - 0x0
    "00000000", -- 5081 - 0x13d9  :    0 - 0x0
    "00000000", -- 5082 - 0x13da  :    0 - 0x0
    "00000000", -- 5083 - 0x13db  :    0 - 0x0
    "00000000", -- 5084 - 0x13dc  :    0 - 0x0
    "00000000", -- 5085 - 0x13dd  :    0 - 0x0
    "00000000", -- 5086 - 0x13de  :    0 - 0x0
    "00000000", -- 5087 - 0x13df  :    0 - 0x0
    "00000000", -- 5088 - 0x13e0  :    0 - 0x0 -- Background 0x3e
    "00000000", -- 5089 - 0x13e1  :    0 - 0x0
    "00000000", -- 5090 - 0x13e2  :    0 - 0x0
    "00000000", -- 5091 - 0x13e3  :    0 - 0x0
    "00000000", -- 5092 - 0x13e4  :    0 - 0x0
    "00000000", -- 5093 - 0x13e5  :    0 - 0x0
    "00000000", -- 5094 - 0x13e6  :    0 - 0x0
    "00000000", -- 5095 - 0x13e7  :    0 - 0x0
    "00000000", -- 5096 - 0x13e8  :    0 - 0x0
    "00000000", -- 5097 - 0x13e9  :    0 - 0x0
    "00000000", -- 5098 - 0x13ea  :    0 - 0x0
    "00000000", -- 5099 - 0x13eb  :    0 - 0x0
    "00000000", -- 5100 - 0x13ec  :    0 - 0x0
    "00000000", -- 5101 - 0x13ed  :    0 - 0x0
    "00000000", -- 5102 - 0x13ee  :    0 - 0x0
    "00000000", -- 5103 - 0x13ef  :    0 - 0x0
    "00000000", -- 5104 - 0x13f0  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 5105 - 0x13f1  :    0 - 0x0
    "00000000", -- 5106 - 0x13f2  :    0 - 0x0
    "00000000", -- 5107 - 0x13f3  :    0 - 0x0
    "00000000", -- 5108 - 0x13f4  :    0 - 0x0
    "00000000", -- 5109 - 0x13f5  :    0 - 0x0
    "00000000", -- 5110 - 0x13f6  :    0 - 0x0
    "00000000", -- 5111 - 0x13f7  :    0 - 0x0
    "00000000", -- 5112 - 0x13f8  :    0 - 0x0
    "00000000", -- 5113 - 0x13f9  :    0 - 0x0
    "00000000", -- 5114 - 0x13fa  :    0 - 0x0
    "00000000", -- 5115 - 0x13fb  :    0 - 0x0
    "00000000", -- 5116 - 0x13fc  :    0 - 0x0
    "00000000", -- 5117 - 0x13fd  :    0 - 0x0
    "00000000", -- 5118 - 0x13fe  :    0 - 0x0
    "00000000", -- 5119 - 0x13ff  :    0 - 0x0
    "00000000", -- 5120 - 0x1400  :    0 - 0x0 -- Background 0x40
    "00000000", -- 5121 - 0x1401  :    0 - 0x0
    "00000000", -- 5122 - 0x1402  :    0 - 0x0
    "00000000", -- 5123 - 0x1403  :    0 - 0x0
    "00000000", -- 5124 - 0x1404  :    0 - 0x0
    "00000000", -- 5125 - 0x1405  :    0 - 0x0
    "00000000", -- 5126 - 0x1406  :    0 - 0x0
    "00000000", -- 5127 - 0x1407  :    0 - 0x0
    "00000000", -- 5128 - 0x1408  :    0 - 0x0
    "00000000", -- 5129 - 0x1409  :    0 - 0x0
    "00000000", -- 5130 - 0x140a  :    0 - 0x0
    "00000000", -- 5131 - 0x140b  :    0 - 0x0
    "00000000", -- 5132 - 0x140c  :    0 - 0x0
    "00000000", -- 5133 - 0x140d  :    0 - 0x0
    "00000000", -- 5134 - 0x140e  :    0 - 0x0
    "00000000", -- 5135 - 0x140f  :    0 - 0x0
    "00000000", -- 5136 - 0x1410  :    0 - 0x0 -- Background 0x41
    "00000000", -- 5137 - 0x1411  :    0 - 0x0
    "00000000", -- 5138 - 0x1412  :    0 - 0x0
    "00000000", -- 5139 - 0x1413  :    0 - 0x0
    "00000000", -- 5140 - 0x1414  :    0 - 0x0
    "00000000", -- 5141 - 0x1415  :    0 - 0x0
    "00000000", -- 5142 - 0x1416  :    0 - 0x0
    "00000000", -- 5143 - 0x1417  :    0 - 0x0
    "00000000", -- 5144 - 0x1418  :    0 - 0x0
    "00000000", -- 5145 - 0x1419  :    0 - 0x0
    "00000000", -- 5146 - 0x141a  :    0 - 0x0
    "00000000", -- 5147 - 0x141b  :    0 - 0x0
    "00000000", -- 5148 - 0x141c  :    0 - 0x0
    "00000000", -- 5149 - 0x141d  :    0 - 0x0
    "00000000", -- 5150 - 0x141e  :    0 - 0x0
    "00000000", -- 5151 - 0x141f  :    0 - 0x0
    "00000000", -- 5152 - 0x1420  :    0 - 0x0 -- Background 0x42
    "00000000", -- 5153 - 0x1421  :    0 - 0x0
    "00000000", -- 5154 - 0x1422  :    0 - 0x0
    "00000000", -- 5155 - 0x1423  :    0 - 0x0
    "00000000", -- 5156 - 0x1424  :    0 - 0x0
    "00000000", -- 5157 - 0x1425  :    0 - 0x0
    "00000000", -- 5158 - 0x1426  :    0 - 0x0
    "00000000", -- 5159 - 0x1427  :    0 - 0x0
    "00000000", -- 5160 - 0x1428  :    0 - 0x0
    "00000000", -- 5161 - 0x1429  :    0 - 0x0
    "00000000", -- 5162 - 0x142a  :    0 - 0x0
    "00000000", -- 5163 - 0x142b  :    0 - 0x0
    "00000000", -- 5164 - 0x142c  :    0 - 0x0
    "00000000", -- 5165 - 0x142d  :    0 - 0x0
    "00000000", -- 5166 - 0x142e  :    0 - 0x0
    "00000000", -- 5167 - 0x142f  :    0 - 0x0
    "00000000", -- 5168 - 0x1430  :    0 - 0x0 -- Background 0x43
    "00000000", -- 5169 - 0x1431  :    0 - 0x0
    "00000000", -- 5170 - 0x1432  :    0 - 0x0
    "00000000", -- 5171 - 0x1433  :    0 - 0x0
    "00000000", -- 5172 - 0x1434  :    0 - 0x0
    "00000000", -- 5173 - 0x1435  :    0 - 0x0
    "00000000", -- 5174 - 0x1436  :    0 - 0x0
    "00000000", -- 5175 - 0x1437  :    0 - 0x0
    "00000000", -- 5176 - 0x1438  :    0 - 0x0
    "00000000", -- 5177 - 0x1439  :    0 - 0x0
    "00000000", -- 5178 - 0x143a  :    0 - 0x0
    "00000000", -- 5179 - 0x143b  :    0 - 0x0
    "00000000", -- 5180 - 0x143c  :    0 - 0x0
    "00000000", -- 5181 - 0x143d  :    0 - 0x0
    "00000000", -- 5182 - 0x143e  :    0 - 0x0
    "00000000", -- 5183 - 0x143f  :    0 - 0x0
    "00000000", -- 5184 - 0x1440  :    0 - 0x0 -- Background 0x44
    "00000000", -- 5185 - 0x1441  :    0 - 0x0
    "00000000", -- 5186 - 0x1442  :    0 - 0x0
    "00000000", -- 5187 - 0x1443  :    0 - 0x0
    "00000000", -- 5188 - 0x1444  :    0 - 0x0
    "00000000", -- 5189 - 0x1445  :    0 - 0x0
    "00000000", -- 5190 - 0x1446  :    0 - 0x0
    "00000000", -- 5191 - 0x1447  :    0 - 0x0
    "00000000", -- 5192 - 0x1448  :    0 - 0x0
    "00000000", -- 5193 - 0x1449  :    0 - 0x0
    "00000000", -- 5194 - 0x144a  :    0 - 0x0
    "00000000", -- 5195 - 0x144b  :    0 - 0x0
    "00000000", -- 5196 - 0x144c  :    0 - 0x0
    "00000000", -- 5197 - 0x144d  :    0 - 0x0
    "00000000", -- 5198 - 0x144e  :    0 - 0x0
    "00000000", -- 5199 - 0x144f  :    0 - 0x0
    "00000000", -- 5200 - 0x1450  :    0 - 0x0 -- Background 0x45
    "00000000", -- 5201 - 0x1451  :    0 - 0x0
    "00000000", -- 5202 - 0x1452  :    0 - 0x0
    "00000000", -- 5203 - 0x1453  :    0 - 0x0
    "00000000", -- 5204 - 0x1454  :    0 - 0x0
    "00000000", -- 5205 - 0x1455  :    0 - 0x0
    "00000000", -- 5206 - 0x1456  :    0 - 0x0
    "00000000", -- 5207 - 0x1457  :    0 - 0x0
    "00000000", -- 5208 - 0x1458  :    0 - 0x0
    "00000000", -- 5209 - 0x1459  :    0 - 0x0
    "00000000", -- 5210 - 0x145a  :    0 - 0x0
    "00000000", -- 5211 - 0x145b  :    0 - 0x0
    "00000000", -- 5212 - 0x145c  :    0 - 0x0
    "00000000", -- 5213 - 0x145d  :    0 - 0x0
    "00000000", -- 5214 - 0x145e  :    0 - 0x0
    "00000000", -- 5215 - 0x145f  :    0 - 0x0
    "00000000", -- 5216 - 0x1460  :    0 - 0x0 -- Background 0x46
    "00000000", -- 5217 - 0x1461  :    0 - 0x0
    "00000000", -- 5218 - 0x1462  :    0 - 0x0
    "00000000", -- 5219 - 0x1463  :    0 - 0x0
    "00000000", -- 5220 - 0x1464  :    0 - 0x0
    "00000000", -- 5221 - 0x1465  :    0 - 0x0
    "00000000", -- 5222 - 0x1466  :    0 - 0x0
    "00000000", -- 5223 - 0x1467  :    0 - 0x0
    "00000000", -- 5224 - 0x1468  :    0 - 0x0
    "00000000", -- 5225 - 0x1469  :    0 - 0x0
    "00000000", -- 5226 - 0x146a  :    0 - 0x0
    "00000000", -- 5227 - 0x146b  :    0 - 0x0
    "00000000", -- 5228 - 0x146c  :    0 - 0x0
    "00000000", -- 5229 - 0x146d  :    0 - 0x0
    "00000000", -- 5230 - 0x146e  :    0 - 0x0
    "00000000", -- 5231 - 0x146f  :    0 - 0x0
    "00000000", -- 5232 - 0x1470  :    0 - 0x0 -- Background 0x47
    "00000000", -- 5233 - 0x1471  :    0 - 0x0
    "00000000", -- 5234 - 0x1472  :    0 - 0x0
    "00000000", -- 5235 - 0x1473  :    0 - 0x0
    "00000000", -- 5236 - 0x1474  :    0 - 0x0
    "00000000", -- 5237 - 0x1475  :    0 - 0x0
    "00000000", -- 5238 - 0x1476  :    0 - 0x0
    "00000000", -- 5239 - 0x1477  :    0 - 0x0
    "00000000", -- 5240 - 0x1478  :    0 - 0x0
    "00000000", -- 5241 - 0x1479  :    0 - 0x0
    "00000000", -- 5242 - 0x147a  :    0 - 0x0
    "00000000", -- 5243 - 0x147b  :    0 - 0x0
    "00000000", -- 5244 - 0x147c  :    0 - 0x0
    "00000000", -- 5245 - 0x147d  :    0 - 0x0
    "00000000", -- 5246 - 0x147e  :    0 - 0x0
    "00000000", -- 5247 - 0x147f  :    0 - 0x0
    "00000000", -- 5248 - 0x1480  :    0 - 0x0 -- Background 0x48
    "00000000", -- 5249 - 0x1481  :    0 - 0x0
    "00000000", -- 5250 - 0x1482  :    0 - 0x0
    "00000000", -- 5251 - 0x1483  :    0 - 0x0
    "00000000", -- 5252 - 0x1484  :    0 - 0x0
    "00000000", -- 5253 - 0x1485  :    0 - 0x0
    "00000000", -- 5254 - 0x1486  :    0 - 0x0
    "00000000", -- 5255 - 0x1487  :    0 - 0x0
    "00000000", -- 5256 - 0x1488  :    0 - 0x0
    "00000000", -- 5257 - 0x1489  :    0 - 0x0
    "00000000", -- 5258 - 0x148a  :    0 - 0x0
    "00000000", -- 5259 - 0x148b  :    0 - 0x0
    "00000000", -- 5260 - 0x148c  :    0 - 0x0
    "00000000", -- 5261 - 0x148d  :    0 - 0x0
    "00000000", -- 5262 - 0x148e  :    0 - 0x0
    "00000000", -- 5263 - 0x148f  :    0 - 0x0
    "00000000", -- 5264 - 0x1490  :    0 - 0x0 -- Background 0x49
    "00000000", -- 5265 - 0x1491  :    0 - 0x0
    "00000000", -- 5266 - 0x1492  :    0 - 0x0
    "00000000", -- 5267 - 0x1493  :    0 - 0x0
    "00000000", -- 5268 - 0x1494  :    0 - 0x0
    "00000000", -- 5269 - 0x1495  :    0 - 0x0
    "00000000", -- 5270 - 0x1496  :    0 - 0x0
    "00000000", -- 5271 - 0x1497  :    0 - 0x0
    "00000000", -- 5272 - 0x1498  :    0 - 0x0
    "00000000", -- 5273 - 0x1499  :    0 - 0x0
    "00000000", -- 5274 - 0x149a  :    0 - 0x0
    "00000000", -- 5275 - 0x149b  :    0 - 0x0
    "00000000", -- 5276 - 0x149c  :    0 - 0x0
    "00000000", -- 5277 - 0x149d  :    0 - 0x0
    "00000000", -- 5278 - 0x149e  :    0 - 0x0
    "00000000", -- 5279 - 0x149f  :    0 - 0x0
    "00000000", -- 5280 - 0x14a0  :    0 - 0x0 -- Background 0x4a
    "00000000", -- 5281 - 0x14a1  :    0 - 0x0
    "00000000", -- 5282 - 0x14a2  :    0 - 0x0
    "00000000", -- 5283 - 0x14a3  :    0 - 0x0
    "00000000", -- 5284 - 0x14a4  :    0 - 0x0
    "00000000", -- 5285 - 0x14a5  :    0 - 0x0
    "00000000", -- 5286 - 0x14a6  :    0 - 0x0
    "00000000", -- 5287 - 0x14a7  :    0 - 0x0
    "00000000", -- 5288 - 0x14a8  :    0 - 0x0
    "00000000", -- 5289 - 0x14a9  :    0 - 0x0
    "00000000", -- 5290 - 0x14aa  :    0 - 0x0
    "00000000", -- 5291 - 0x14ab  :    0 - 0x0
    "00000000", -- 5292 - 0x14ac  :    0 - 0x0
    "00000000", -- 5293 - 0x14ad  :    0 - 0x0
    "00000000", -- 5294 - 0x14ae  :    0 - 0x0
    "00000000", -- 5295 - 0x14af  :    0 - 0x0
    "00000000", -- 5296 - 0x14b0  :    0 - 0x0 -- Background 0x4b
    "00000000", -- 5297 - 0x14b1  :    0 - 0x0
    "00000000", -- 5298 - 0x14b2  :    0 - 0x0
    "00000000", -- 5299 - 0x14b3  :    0 - 0x0
    "00000000", -- 5300 - 0x14b4  :    0 - 0x0
    "00000000", -- 5301 - 0x14b5  :    0 - 0x0
    "00000000", -- 5302 - 0x14b6  :    0 - 0x0
    "00000000", -- 5303 - 0x14b7  :    0 - 0x0
    "00000000", -- 5304 - 0x14b8  :    0 - 0x0
    "00000000", -- 5305 - 0x14b9  :    0 - 0x0
    "00000000", -- 5306 - 0x14ba  :    0 - 0x0
    "00000000", -- 5307 - 0x14bb  :    0 - 0x0
    "00000000", -- 5308 - 0x14bc  :    0 - 0x0
    "00000000", -- 5309 - 0x14bd  :    0 - 0x0
    "00000000", -- 5310 - 0x14be  :    0 - 0x0
    "00000000", -- 5311 - 0x14bf  :    0 - 0x0
    "00000000", -- 5312 - 0x14c0  :    0 - 0x0 -- Background 0x4c
    "00000000", -- 5313 - 0x14c1  :    0 - 0x0
    "00000000", -- 5314 - 0x14c2  :    0 - 0x0
    "00000000", -- 5315 - 0x14c3  :    0 - 0x0
    "00000000", -- 5316 - 0x14c4  :    0 - 0x0
    "00000000", -- 5317 - 0x14c5  :    0 - 0x0
    "00000000", -- 5318 - 0x14c6  :    0 - 0x0
    "00000000", -- 5319 - 0x14c7  :    0 - 0x0
    "00000000", -- 5320 - 0x14c8  :    0 - 0x0
    "00000000", -- 5321 - 0x14c9  :    0 - 0x0
    "00000000", -- 5322 - 0x14ca  :    0 - 0x0
    "00000000", -- 5323 - 0x14cb  :    0 - 0x0
    "00000000", -- 5324 - 0x14cc  :    0 - 0x0
    "00000000", -- 5325 - 0x14cd  :    0 - 0x0
    "00000000", -- 5326 - 0x14ce  :    0 - 0x0
    "00000000", -- 5327 - 0x14cf  :    0 - 0x0
    "00000000", -- 5328 - 0x14d0  :    0 - 0x0 -- Background 0x4d
    "00000000", -- 5329 - 0x14d1  :    0 - 0x0
    "00000000", -- 5330 - 0x14d2  :    0 - 0x0
    "00000000", -- 5331 - 0x14d3  :    0 - 0x0
    "00000000", -- 5332 - 0x14d4  :    0 - 0x0
    "00000000", -- 5333 - 0x14d5  :    0 - 0x0
    "00000000", -- 5334 - 0x14d6  :    0 - 0x0
    "00000000", -- 5335 - 0x14d7  :    0 - 0x0
    "00000000", -- 5336 - 0x14d8  :    0 - 0x0
    "00000000", -- 5337 - 0x14d9  :    0 - 0x0
    "00000000", -- 5338 - 0x14da  :    0 - 0x0
    "00000000", -- 5339 - 0x14db  :    0 - 0x0
    "00000000", -- 5340 - 0x14dc  :    0 - 0x0
    "00000000", -- 5341 - 0x14dd  :    0 - 0x0
    "00000000", -- 5342 - 0x14de  :    0 - 0x0
    "00000000", -- 5343 - 0x14df  :    0 - 0x0
    "00000000", -- 5344 - 0x14e0  :    0 - 0x0 -- Background 0x4e
    "00000000", -- 5345 - 0x14e1  :    0 - 0x0
    "00000000", -- 5346 - 0x14e2  :    0 - 0x0
    "00000000", -- 5347 - 0x14e3  :    0 - 0x0
    "00000000", -- 5348 - 0x14e4  :    0 - 0x0
    "00000000", -- 5349 - 0x14e5  :    0 - 0x0
    "00000000", -- 5350 - 0x14e6  :    0 - 0x0
    "00000000", -- 5351 - 0x14e7  :    0 - 0x0
    "00000000", -- 5352 - 0x14e8  :    0 - 0x0
    "00000000", -- 5353 - 0x14e9  :    0 - 0x0
    "00000000", -- 5354 - 0x14ea  :    0 - 0x0
    "00000000", -- 5355 - 0x14eb  :    0 - 0x0
    "00000000", -- 5356 - 0x14ec  :    0 - 0x0
    "00000000", -- 5357 - 0x14ed  :    0 - 0x0
    "00000000", -- 5358 - 0x14ee  :    0 - 0x0
    "00000000", -- 5359 - 0x14ef  :    0 - 0x0
    "00000000", -- 5360 - 0x14f0  :    0 - 0x0 -- Background 0x4f
    "00000000", -- 5361 - 0x14f1  :    0 - 0x0
    "00000000", -- 5362 - 0x14f2  :    0 - 0x0
    "00000000", -- 5363 - 0x14f3  :    0 - 0x0
    "00000000", -- 5364 - 0x14f4  :    0 - 0x0
    "00000000", -- 5365 - 0x14f5  :    0 - 0x0
    "00000000", -- 5366 - 0x14f6  :    0 - 0x0
    "00000000", -- 5367 - 0x14f7  :    0 - 0x0
    "00000000", -- 5368 - 0x14f8  :    0 - 0x0
    "00000000", -- 5369 - 0x14f9  :    0 - 0x0
    "00000000", -- 5370 - 0x14fa  :    0 - 0x0
    "00000000", -- 5371 - 0x14fb  :    0 - 0x0
    "00000000", -- 5372 - 0x14fc  :    0 - 0x0
    "00000000", -- 5373 - 0x14fd  :    0 - 0x0
    "00000000", -- 5374 - 0x14fe  :    0 - 0x0
    "00000000", -- 5375 - 0x14ff  :    0 - 0x0
    "00000000", -- 5376 - 0x1500  :    0 - 0x0 -- Background 0x50
    "00000000", -- 5377 - 0x1501  :    0 - 0x0
    "00000000", -- 5378 - 0x1502  :    0 - 0x0
    "00000000", -- 5379 - 0x1503  :    0 - 0x0
    "00000000", -- 5380 - 0x1504  :    0 - 0x0
    "00000000", -- 5381 - 0x1505  :    0 - 0x0
    "00000000", -- 5382 - 0x1506  :    0 - 0x0
    "00000000", -- 5383 - 0x1507  :    0 - 0x0
    "00000000", -- 5384 - 0x1508  :    0 - 0x0
    "00000000", -- 5385 - 0x1509  :    0 - 0x0
    "00000000", -- 5386 - 0x150a  :    0 - 0x0
    "00000000", -- 5387 - 0x150b  :    0 - 0x0
    "00000000", -- 5388 - 0x150c  :    0 - 0x0
    "00000000", -- 5389 - 0x150d  :    0 - 0x0
    "00000000", -- 5390 - 0x150e  :    0 - 0x0
    "00000000", -- 5391 - 0x150f  :    0 - 0x0
    "00000000", -- 5392 - 0x1510  :    0 - 0x0 -- Background 0x51
    "00000000", -- 5393 - 0x1511  :    0 - 0x0
    "00000000", -- 5394 - 0x1512  :    0 - 0x0
    "00000000", -- 5395 - 0x1513  :    0 - 0x0
    "00000000", -- 5396 - 0x1514  :    0 - 0x0
    "00000000", -- 5397 - 0x1515  :    0 - 0x0
    "00000000", -- 5398 - 0x1516  :    0 - 0x0
    "00000000", -- 5399 - 0x1517  :    0 - 0x0
    "00000000", -- 5400 - 0x1518  :    0 - 0x0
    "00000000", -- 5401 - 0x1519  :    0 - 0x0
    "00000000", -- 5402 - 0x151a  :    0 - 0x0
    "00000000", -- 5403 - 0x151b  :    0 - 0x0
    "00000000", -- 5404 - 0x151c  :    0 - 0x0
    "00000000", -- 5405 - 0x151d  :    0 - 0x0
    "00000000", -- 5406 - 0x151e  :    0 - 0x0
    "00000000", -- 5407 - 0x151f  :    0 - 0x0
    "00000000", -- 5408 - 0x1520  :    0 - 0x0 -- Background 0x52
    "00000000", -- 5409 - 0x1521  :    0 - 0x0
    "00000000", -- 5410 - 0x1522  :    0 - 0x0
    "00000000", -- 5411 - 0x1523  :    0 - 0x0
    "00000000", -- 5412 - 0x1524  :    0 - 0x0
    "00000000", -- 5413 - 0x1525  :    0 - 0x0
    "00000000", -- 5414 - 0x1526  :    0 - 0x0
    "00000000", -- 5415 - 0x1527  :    0 - 0x0
    "00000000", -- 5416 - 0x1528  :    0 - 0x0
    "00000000", -- 5417 - 0x1529  :    0 - 0x0
    "00000000", -- 5418 - 0x152a  :    0 - 0x0
    "00000000", -- 5419 - 0x152b  :    0 - 0x0
    "00000000", -- 5420 - 0x152c  :    0 - 0x0
    "00000000", -- 5421 - 0x152d  :    0 - 0x0
    "00000000", -- 5422 - 0x152e  :    0 - 0x0
    "00000000", -- 5423 - 0x152f  :    0 - 0x0
    "00000000", -- 5424 - 0x1530  :    0 - 0x0 -- Background 0x53
    "00000000", -- 5425 - 0x1531  :    0 - 0x0
    "00000000", -- 5426 - 0x1532  :    0 - 0x0
    "00000000", -- 5427 - 0x1533  :    0 - 0x0
    "00000000", -- 5428 - 0x1534  :    0 - 0x0
    "00000000", -- 5429 - 0x1535  :    0 - 0x0
    "00000000", -- 5430 - 0x1536  :    0 - 0x0
    "00000000", -- 5431 - 0x1537  :    0 - 0x0
    "00000000", -- 5432 - 0x1538  :    0 - 0x0
    "00000000", -- 5433 - 0x1539  :    0 - 0x0
    "00000000", -- 5434 - 0x153a  :    0 - 0x0
    "00000000", -- 5435 - 0x153b  :    0 - 0x0
    "00000000", -- 5436 - 0x153c  :    0 - 0x0
    "00000000", -- 5437 - 0x153d  :    0 - 0x0
    "00000000", -- 5438 - 0x153e  :    0 - 0x0
    "00000000", -- 5439 - 0x153f  :    0 - 0x0
    "00000000", -- 5440 - 0x1540  :    0 - 0x0 -- Background 0x54
    "00000000", -- 5441 - 0x1541  :    0 - 0x0
    "00000000", -- 5442 - 0x1542  :    0 - 0x0
    "00000000", -- 5443 - 0x1543  :    0 - 0x0
    "00000000", -- 5444 - 0x1544  :    0 - 0x0
    "00000000", -- 5445 - 0x1545  :    0 - 0x0
    "00000000", -- 5446 - 0x1546  :    0 - 0x0
    "00000000", -- 5447 - 0x1547  :    0 - 0x0
    "00000000", -- 5448 - 0x1548  :    0 - 0x0
    "00000000", -- 5449 - 0x1549  :    0 - 0x0
    "00000000", -- 5450 - 0x154a  :    0 - 0x0
    "00000000", -- 5451 - 0x154b  :    0 - 0x0
    "00000000", -- 5452 - 0x154c  :    0 - 0x0
    "00000000", -- 5453 - 0x154d  :    0 - 0x0
    "00000000", -- 5454 - 0x154e  :    0 - 0x0
    "00000000", -- 5455 - 0x154f  :    0 - 0x0
    "00000000", -- 5456 - 0x1550  :    0 - 0x0 -- Background 0x55
    "00000000", -- 5457 - 0x1551  :    0 - 0x0
    "00000000", -- 5458 - 0x1552  :    0 - 0x0
    "00000000", -- 5459 - 0x1553  :    0 - 0x0
    "00000000", -- 5460 - 0x1554  :    0 - 0x0
    "00000000", -- 5461 - 0x1555  :    0 - 0x0
    "00000000", -- 5462 - 0x1556  :    0 - 0x0
    "00000000", -- 5463 - 0x1557  :    0 - 0x0
    "00000000", -- 5464 - 0x1558  :    0 - 0x0
    "00000000", -- 5465 - 0x1559  :    0 - 0x0
    "00000000", -- 5466 - 0x155a  :    0 - 0x0
    "00000000", -- 5467 - 0x155b  :    0 - 0x0
    "00000000", -- 5468 - 0x155c  :    0 - 0x0
    "00000000", -- 5469 - 0x155d  :    0 - 0x0
    "00000000", -- 5470 - 0x155e  :    0 - 0x0
    "00000000", -- 5471 - 0x155f  :    0 - 0x0
    "00000000", -- 5472 - 0x1560  :    0 - 0x0 -- Background 0x56
    "00000000", -- 5473 - 0x1561  :    0 - 0x0
    "00000000", -- 5474 - 0x1562  :    0 - 0x0
    "00000000", -- 5475 - 0x1563  :    0 - 0x0
    "00000000", -- 5476 - 0x1564  :    0 - 0x0
    "00000000", -- 5477 - 0x1565  :    0 - 0x0
    "00000000", -- 5478 - 0x1566  :    0 - 0x0
    "00000000", -- 5479 - 0x1567  :    0 - 0x0
    "00000000", -- 5480 - 0x1568  :    0 - 0x0
    "00000000", -- 5481 - 0x1569  :    0 - 0x0
    "00000000", -- 5482 - 0x156a  :    0 - 0x0
    "00000000", -- 5483 - 0x156b  :    0 - 0x0
    "00000000", -- 5484 - 0x156c  :    0 - 0x0
    "00000000", -- 5485 - 0x156d  :    0 - 0x0
    "00000000", -- 5486 - 0x156e  :    0 - 0x0
    "00000000", -- 5487 - 0x156f  :    0 - 0x0
    "00000000", -- 5488 - 0x1570  :    0 - 0x0 -- Background 0x57
    "00000000", -- 5489 - 0x1571  :    0 - 0x0
    "00000000", -- 5490 - 0x1572  :    0 - 0x0
    "00000000", -- 5491 - 0x1573  :    0 - 0x0
    "00000000", -- 5492 - 0x1574  :    0 - 0x0
    "00000000", -- 5493 - 0x1575  :    0 - 0x0
    "00000000", -- 5494 - 0x1576  :    0 - 0x0
    "00000000", -- 5495 - 0x1577  :    0 - 0x0
    "00000000", -- 5496 - 0x1578  :    0 - 0x0
    "00000000", -- 5497 - 0x1579  :    0 - 0x0
    "00000000", -- 5498 - 0x157a  :    0 - 0x0
    "00000000", -- 5499 - 0x157b  :    0 - 0x0
    "00000000", -- 5500 - 0x157c  :    0 - 0x0
    "00000000", -- 5501 - 0x157d  :    0 - 0x0
    "00000000", -- 5502 - 0x157e  :    0 - 0x0
    "00000000", -- 5503 - 0x157f  :    0 - 0x0
    "00000000", -- 5504 - 0x1580  :    0 - 0x0 -- Background 0x58
    "00000000", -- 5505 - 0x1581  :    0 - 0x0
    "00000000", -- 5506 - 0x1582  :    0 - 0x0
    "00000000", -- 5507 - 0x1583  :    0 - 0x0
    "00000000", -- 5508 - 0x1584  :    0 - 0x0
    "00000000", -- 5509 - 0x1585  :    0 - 0x0
    "00000000", -- 5510 - 0x1586  :    0 - 0x0
    "00000000", -- 5511 - 0x1587  :    0 - 0x0
    "00000000", -- 5512 - 0x1588  :    0 - 0x0
    "00000000", -- 5513 - 0x1589  :    0 - 0x0
    "00000000", -- 5514 - 0x158a  :    0 - 0x0
    "00000000", -- 5515 - 0x158b  :    0 - 0x0
    "00000000", -- 5516 - 0x158c  :    0 - 0x0
    "00000000", -- 5517 - 0x158d  :    0 - 0x0
    "00000000", -- 5518 - 0x158e  :    0 - 0x0
    "00000000", -- 5519 - 0x158f  :    0 - 0x0
    "00000000", -- 5520 - 0x1590  :    0 - 0x0 -- Background 0x59
    "00000000", -- 5521 - 0x1591  :    0 - 0x0
    "00000000", -- 5522 - 0x1592  :    0 - 0x0
    "00000000", -- 5523 - 0x1593  :    0 - 0x0
    "00000000", -- 5524 - 0x1594  :    0 - 0x0
    "00000000", -- 5525 - 0x1595  :    0 - 0x0
    "00000000", -- 5526 - 0x1596  :    0 - 0x0
    "00000000", -- 5527 - 0x1597  :    0 - 0x0
    "00000000", -- 5528 - 0x1598  :    0 - 0x0
    "00000000", -- 5529 - 0x1599  :    0 - 0x0
    "00000000", -- 5530 - 0x159a  :    0 - 0x0
    "00000000", -- 5531 - 0x159b  :    0 - 0x0
    "00000000", -- 5532 - 0x159c  :    0 - 0x0
    "00000000", -- 5533 - 0x159d  :    0 - 0x0
    "00000000", -- 5534 - 0x159e  :    0 - 0x0
    "00000000", -- 5535 - 0x159f  :    0 - 0x0
    "00000000", -- 5536 - 0x15a0  :    0 - 0x0 -- Background 0x5a
    "00000000", -- 5537 - 0x15a1  :    0 - 0x0
    "00000000", -- 5538 - 0x15a2  :    0 - 0x0
    "00000000", -- 5539 - 0x15a3  :    0 - 0x0
    "00000000", -- 5540 - 0x15a4  :    0 - 0x0
    "00000000", -- 5541 - 0x15a5  :    0 - 0x0
    "00000000", -- 5542 - 0x15a6  :    0 - 0x0
    "00000000", -- 5543 - 0x15a7  :    0 - 0x0
    "00000000", -- 5544 - 0x15a8  :    0 - 0x0
    "00000000", -- 5545 - 0x15a9  :    0 - 0x0
    "00000000", -- 5546 - 0x15aa  :    0 - 0x0
    "00000000", -- 5547 - 0x15ab  :    0 - 0x0
    "00000000", -- 5548 - 0x15ac  :    0 - 0x0
    "00000000", -- 5549 - 0x15ad  :    0 - 0x0
    "00000000", -- 5550 - 0x15ae  :    0 - 0x0
    "00000000", -- 5551 - 0x15af  :    0 - 0x0
    "00000000", -- 5552 - 0x15b0  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 5553 - 0x15b1  :    0 - 0x0
    "00000000", -- 5554 - 0x15b2  :    0 - 0x0
    "00000000", -- 5555 - 0x15b3  :    0 - 0x0
    "00000000", -- 5556 - 0x15b4  :    0 - 0x0
    "00000000", -- 5557 - 0x15b5  :    0 - 0x0
    "00000000", -- 5558 - 0x15b6  :    0 - 0x0
    "00000000", -- 5559 - 0x15b7  :    0 - 0x0
    "00000000", -- 5560 - 0x15b8  :    0 - 0x0
    "00000000", -- 5561 - 0x15b9  :    0 - 0x0
    "00000000", -- 5562 - 0x15ba  :    0 - 0x0
    "00000000", -- 5563 - 0x15bb  :    0 - 0x0
    "00000000", -- 5564 - 0x15bc  :    0 - 0x0
    "00000000", -- 5565 - 0x15bd  :    0 - 0x0
    "00000000", -- 5566 - 0x15be  :    0 - 0x0
    "00000000", -- 5567 - 0x15bf  :    0 - 0x0
    "00000000", -- 5568 - 0x15c0  :    0 - 0x0 -- Background 0x5c
    "00000000", -- 5569 - 0x15c1  :    0 - 0x0
    "00000000", -- 5570 - 0x15c2  :    0 - 0x0
    "00000000", -- 5571 - 0x15c3  :    0 - 0x0
    "00000000", -- 5572 - 0x15c4  :    0 - 0x0
    "00000000", -- 5573 - 0x15c5  :    0 - 0x0
    "00000000", -- 5574 - 0x15c6  :    0 - 0x0
    "00000000", -- 5575 - 0x15c7  :    0 - 0x0
    "00000000", -- 5576 - 0x15c8  :    0 - 0x0
    "00000000", -- 5577 - 0x15c9  :    0 - 0x0
    "00000000", -- 5578 - 0x15ca  :    0 - 0x0
    "00000000", -- 5579 - 0x15cb  :    0 - 0x0
    "00000000", -- 5580 - 0x15cc  :    0 - 0x0
    "00000000", -- 5581 - 0x15cd  :    0 - 0x0
    "00000000", -- 5582 - 0x15ce  :    0 - 0x0
    "00000000", -- 5583 - 0x15cf  :    0 - 0x0
    "00000000", -- 5584 - 0x15d0  :    0 - 0x0 -- Background 0x5d
    "00000000", -- 5585 - 0x15d1  :    0 - 0x0
    "00000000", -- 5586 - 0x15d2  :    0 - 0x0
    "00000000", -- 5587 - 0x15d3  :    0 - 0x0
    "00000000", -- 5588 - 0x15d4  :    0 - 0x0
    "00000000", -- 5589 - 0x15d5  :    0 - 0x0
    "00000000", -- 5590 - 0x15d6  :    0 - 0x0
    "00000000", -- 5591 - 0x15d7  :    0 - 0x0
    "00000000", -- 5592 - 0x15d8  :    0 - 0x0
    "00000000", -- 5593 - 0x15d9  :    0 - 0x0
    "00000000", -- 5594 - 0x15da  :    0 - 0x0
    "00000000", -- 5595 - 0x15db  :    0 - 0x0
    "00000000", -- 5596 - 0x15dc  :    0 - 0x0
    "00000000", -- 5597 - 0x15dd  :    0 - 0x0
    "00000000", -- 5598 - 0x15de  :    0 - 0x0
    "00000000", -- 5599 - 0x15df  :    0 - 0x0
    "00000000", -- 5600 - 0x15e0  :    0 - 0x0 -- Background 0x5e
    "00000000", -- 5601 - 0x15e1  :    0 - 0x0
    "00000000", -- 5602 - 0x15e2  :    0 - 0x0
    "00000000", -- 5603 - 0x15e3  :    0 - 0x0
    "00000000", -- 5604 - 0x15e4  :    0 - 0x0
    "00000000", -- 5605 - 0x15e5  :    0 - 0x0
    "00000000", -- 5606 - 0x15e6  :    0 - 0x0
    "00000000", -- 5607 - 0x15e7  :    0 - 0x0
    "00000000", -- 5608 - 0x15e8  :    0 - 0x0
    "00000000", -- 5609 - 0x15e9  :    0 - 0x0
    "00000000", -- 5610 - 0x15ea  :    0 - 0x0
    "00000000", -- 5611 - 0x15eb  :    0 - 0x0
    "00000000", -- 5612 - 0x15ec  :    0 - 0x0
    "00000000", -- 5613 - 0x15ed  :    0 - 0x0
    "00000000", -- 5614 - 0x15ee  :    0 - 0x0
    "00000000", -- 5615 - 0x15ef  :    0 - 0x0
    "00000000", -- 5616 - 0x15f0  :    0 - 0x0 -- Background 0x5f
    "00000000", -- 5617 - 0x15f1  :    0 - 0x0
    "00000000", -- 5618 - 0x15f2  :    0 - 0x0
    "00000000", -- 5619 - 0x15f3  :    0 - 0x0
    "00000000", -- 5620 - 0x15f4  :    0 - 0x0
    "00000000", -- 5621 - 0x15f5  :    0 - 0x0
    "00000000", -- 5622 - 0x15f6  :    0 - 0x0
    "00000000", -- 5623 - 0x15f7  :    0 - 0x0
    "00000000", -- 5624 - 0x15f8  :    0 - 0x0
    "00000000", -- 5625 - 0x15f9  :    0 - 0x0
    "00000000", -- 5626 - 0x15fa  :    0 - 0x0
    "00000000", -- 5627 - 0x15fb  :    0 - 0x0
    "00000000", -- 5628 - 0x15fc  :    0 - 0x0
    "00000000", -- 5629 - 0x15fd  :    0 - 0x0
    "00000000", -- 5630 - 0x15fe  :    0 - 0x0
    "00000000", -- 5631 - 0x15ff  :    0 - 0x0
    "00000000", -- 5632 - 0x1600  :    0 - 0x0 -- Background 0x60
    "00000000", -- 5633 - 0x1601  :    0 - 0x0
    "00000000", -- 5634 - 0x1602  :    0 - 0x0
    "00000000", -- 5635 - 0x1603  :    0 - 0x0
    "00000000", -- 5636 - 0x1604  :    0 - 0x0
    "00000000", -- 5637 - 0x1605  :    0 - 0x0
    "00000000", -- 5638 - 0x1606  :    0 - 0x0
    "00000000", -- 5639 - 0x1607  :    0 - 0x0
    "00000000", -- 5640 - 0x1608  :    0 - 0x0
    "00000000", -- 5641 - 0x1609  :    0 - 0x0
    "00000000", -- 5642 - 0x160a  :    0 - 0x0
    "00000000", -- 5643 - 0x160b  :    0 - 0x0
    "00000000", -- 5644 - 0x160c  :    0 - 0x0
    "00000000", -- 5645 - 0x160d  :    0 - 0x0
    "00000000", -- 5646 - 0x160e  :    0 - 0x0
    "00000000", -- 5647 - 0x160f  :    0 - 0x0
    "00000000", -- 5648 - 0x1610  :    0 - 0x0 -- Background 0x61
    "00000000", -- 5649 - 0x1611  :    0 - 0x0
    "00000000", -- 5650 - 0x1612  :    0 - 0x0
    "00000000", -- 5651 - 0x1613  :    0 - 0x0
    "00000000", -- 5652 - 0x1614  :    0 - 0x0
    "00000000", -- 5653 - 0x1615  :    0 - 0x0
    "00000000", -- 5654 - 0x1616  :    0 - 0x0
    "00000000", -- 5655 - 0x1617  :    0 - 0x0
    "00000000", -- 5656 - 0x1618  :    0 - 0x0
    "00000000", -- 5657 - 0x1619  :    0 - 0x0
    "00000000", -- 5658 - 0x161a  :    0 - 0x0
    "00000000", -- 5659 - 0x161b  :    0 - 0x0
    "00000000", -- 5660 - 0x161c  :    0 - 0x0
    "00000000", -- 5661 - 0x161d  :    0 - 0x0
    "00000000", -- 5662 - 0x161e  :    0 - 0x0
    "00000000", -- 5663 - 0x161f  :    0 - 0x0
    "00000000", -- 5664 - 0x1620  :    0 - 0x0 -- Background 0x62
    "00000000", -- 5665 - 0x1621  :    0 - 0x0
    "00000000", -- 5666 - 0x1622  :    0 - 0x0
    "00000000", -- 5667 - 0x1623  :    0 - 0x0
    "00000000", -- 5668 - 0x1624  :    0 - 0x0
    "00000000", -- 5669 - 0x1625  :    0 - 0x0
    "00000000", -- 5670 - 0x1626  :    0 - 0x0
    "00000000", -- 5671 - 0x1627  :    0 - 0x0
    "00000000", -- 5672 - 0x1628  :    0 - 0x0
    "00000000", -- 5673 - 0x1629  :    0 - 0x0
    "00000000", -- 5674 - 0x162a  :    0 - 0x0
    "00000000", -- 5675 - 0x162b  :    0 - 0x0
    "00000000", -- 5676 - 0x162c  :    0 - 0x0
    "00000000", -- 5677 - 0x162d  :    0 - 0x0
    "00000000", -- 5678 - 0x162e  :    0 - 0x0
    "00000000", -- 5679 - 0x162f  :    0 - 0x0
    "00000000", -- 5680 - 0x1630  :    0 - 0x0 -- Background 0x63
    "00000000", -- 5681 - 0x1631  :    0 - 0x0
    "00000000", -- 5682 - 0x1632  :    0 - 0x0
    "00000000", -- 5683 - 0x1633  :    0 - 0x0
    "00000000", -- 5684 - 0x1634  :    0 - 0x0
    "00000000", -- 5685 - 0x1635  :    0 - 0x0
    "00000000", -- 5686 - 0x1636  :    0 - 0x0
    "00000000", -- 5687 - 0x1637  :    0 - 0x0
    "00000000", -- 5688 - 0x1638  :    0 - 0x0
    "00000000", -- 5689 - 0x1639  :    0 - 0x0
    "00000000", -- 5690 - 0x163a  :    0 - 0x0
    "00000000", -- 5691 - 0x163b  :    0 - 0x0
    "00000000", -- 5692 - 0x163c  :    0 - 0x0
    "00000000", -- 5693 - 0x163d  :    0 - 0x0
    "00000000", -- 5694 - 0x163e  :    0 - 0x0
    "00000000", -- 5695 - 0x163f  :    0 - 0x0
    "00000000", -- 5696 - 0x1640  :    0 - 0x0 -- Background 0x64
    "00000000", -- 5697 - 0x1641  :    0 - 0x0
    "00000000", -- 5698 - 0x1642  :    0 - 0x0
    "00000000", -- 5699 - 0x1643  :    0 - 0x0
    "00000000", -- 5700 - 0x1644  :    0 - 0x0
    "00000000", -- 5701 - 0x1645  :    0 - 0x0
    "00000000", -- 5702 - 0x1646  :    0 - 0x0
    "00000000", -- 5703 - 0x1647  :    0 - 0x0
    "00000000", -- 5704 - 0x1648  :    0 - 0x0
    "00000000", -- 5705 - 0x1649  :    0 - 0x0
    "00000000", -- 5706 - 0x164a  :    0 - 0x0
    "00000000", -- 5707 - 0x164b  :    0 - 0x0
    "00000000", -- 5708 - 0x164c  :    0 - 0x0
    "00000000", -- 5709 - 0x164d  :    0 - 0x0
    "00000000", -- 5710 - 0x164e  :    0 - 0x0
    "00000000", -- 5711 - 0x164f  :    0 - 0x0
    "00000000", -- 5712 - 0x1650  :    0 - 0x0 -- Background 0x65
    "00000000", -- 5713 - 0x1651  :    0 - 0x0
    "00000000", -- 5714 - 0x1652  :    0 - 0x0
    "00000000", -- 5715 - 0x1653  :    0 - 0x0
    "00000000", -- 5716 - 0x1654  :    0 - 0x0
    "00000000", -- 5717 - 0x1655  :    0 - 0x0
    "00000000", -- 5718 - 0x1656  :    0 - 0x0
    "00000000", -- 5719 - 0x1657  :    0 - 0x0
    "00000000", -- 5720 - 0x1658  :    0 - 0x0
    "00000000", -- 5721 - 0x1659  :    0 - 0x0
    "00000000", -- 5722 - 0x165a  :    0 - 0x0
    "00000000", -- 5723 - 0x165b  :    0 - 0x0
    "00000000", -- 5724 - 0x165c  :    0 - 0x0
    "00000000", -- 5725 - 0x165d  :    0 - 0x0
    "00000000", -- 5726 - 0x165e  :    0 - 0x0
    "00000000", -- 5727 - 0x165f  :    0 - 0x0
    "00000000", -- 5728 - 0x1660  :    0 - 0x0 -- Background 0x66
    "00000000", -- 5729 - 0x1661  :    0 - 0x0
    "00000000", -- 5730 - 0x1662  :    0 - 0x0
    "00000000", -- 5731 - 0x1663  :    0 - 0x0
    "00000000", -- 5732 - 0x1664  :    0 - 0x0
    "00000000", -- 5733 - 0x1665  :    0 - 0x0
    "00000000", -- 5734 - 0x1666  :    0 - 0x0
    "00000000", -- 5735 - 0x1667  :    0 - 0x0
    "00000000", -- 5736 - 0x1668  :    0 - 0x0
    "00000000", -- 5737 - 0x1669  :    0 - 0x0
    "00000000", -- 5738 - 0x166a  :    0 - 0x0
    "00000000", -- 5739 - 0x166b  :    0 - 0x0
    "00000000", -- 5740 - 0x166c  :    0 - 0x0
    "00000000", -- 5741 - 0x166d  :    0 - 0x0
    "00000000", -- 5742 - 0x166e  :    0 - 0x0
    "00000000", -- 5743 - 0x166f  :    0 - 0x0
    "00000000", -- 5744 - 0x1670  :    0 - 0x0 -- Background 0x67
    "00000000", -- 5745 - 0x1671  :    0 - 0x0
    "00000000", -- 5746 - 0x1672  :    0 - 0x0
    "00000000", -- 5747 - 0x1673  :    0 - 0x0
    "00000000", -- 5748 - 0x1674  :    0 - 0x0
    "00000000", -- 5749 - 0x1675  :    0 - 0x0
    "00000000", -- 5750 - 0x1676  :    0 - 0x0
    "00000000", -- 5751 - 0x1677  :    0 - 0x0
    "00000000", -- 5752 - 0x1678  :    0 - 0x0
    "00000000", -- 5753 - 0x1679  :    0 - 0x0
    "00000000", -- 5754 - 0x167a  :    0 - 0x0
    "00000000", -- 5755 - 0x167b  :    0 - 0x0
    "00000000", -- 5756 - 0x167c  :    0 - 0x0
    "00000000", -- 5757 - 0x167d  :    0 - 0x0
    "00000000", -- 5758 - 0x167e  :    0 - 0x0
    "00000000", -- 5759 - 0x167f  :    0 - 0x0
    "00000000", -- 5760 - 0x1680  :    0 - 0x0 -- Background 0x68
    "00000000", -- 5761 - 0x1681  :    0 - 0x0
    "00000000", -- 5762 - 0x1682  :    0 - 0x0
    "00000000", -- 5763 - 0x1683  :    0 - 0x0
    "00000000", -- 5764 - 0x1684  :    0 - 0x0
    "00000000", -- 5765 - 0x1685  :    0 - 0x0
    "00000000", -- 5766 - 0x1686  :    0 - 0x0
    "00000000", -- 5767 - 0x1687  :    0 - 0x0
    "00000000", -- 5768 - 0x1688  :    0 - 0x0
    "00000000", -- 5769 - 0x1689  :    0 - 0x0
    "00000000", -- 5770 - 0x168a  :    0 - 0x0
    "00000000", -- 5771 - 0x168b  :    0 - 0x0
    "00000000", -- 5772 - 0x168c  :    0 - 0x0
    "00000000", -- 5773 - 0x168d  :    0 - 0x0
    "00000000", -- 5774 - 0x168e  :    0 - 0x0
    "00000000", -- 5775 - 0x168f  :    0 - 0x0
    "00000000", -- 5776 - 0x1690  :    0 - 0x0 -- Background 0x69
    "00000000", -- 5777 - 0x1691  :    0 - 0x0
    "00000000", -- 5778 - 0x1692  :    0 - 0x0
    "00000000", -- 5779 - 0x1693  :    0 - 0x0
    "00000000", -- 5780 - 0x1694  :    0 - 0x0
    "00000000", -- 5781 - 0x1695  :    0 - 0x0
    "00000000", -- 5782 - 0x1696  :    0 - 0x0
    "00000000", -- 5783 - 0x1697  :    0 - 0x0
    "00000000", -- 5784 - 0x1698  :    0 - 0x0
    "00000000", -- 5785 - 0x1699  :    0 - 0x0
    "00000000", -- 5786 - 0x169a  :    0 - 0x0
    "00000000", -- 5787 - 0x169b  :    0 - 0x0
    "00000000", -- 5788 - 0x169c  :    0 - 0x0
    "00000000", -- 5789 - 0x169d  :    0 - 0x0
    "00000000", -- 5790 - 0x169e  :    0 - 0x0
    "00000000", -- 5791 - 0x169f  :    0 - 0x0
    "00000000", -- 5792 - 0x16a0  :    0 - 0x0 -- Background 0x6a
    "00000000", -- 5793 - 0x16a1  :    0 - 0x0
    "00000000", -- 5794 - 0x16a2  :    0 - 0x0
    "00000000", -- 5795 - 0x16a3  :    0 - 0x0
    "00000000", -- 5796 - 0x16a4  :    0 - 0x0
    "00000000", -- 5797 - 0x16a5  :    0 - 0x0
    "00000000", -- 5798 - 0x16a6  :    0 - 0x0
    "00000000", -- 5799 - 0x16a7  :    0 - 0x0
    "00000000", -- 5800 - 0x16a8  :    0 - 0x0
    "00000000", -- 5801 - 0x16a9  :    0 - 0x0
    "00000000", -- 5802 - 0x16aa  :    0 - 0x0
    "00000000", -- 5803 - 0x16ab  :    0 - 0x0
    "00000000", -- 5804 - 0x16ac  :    0 - 0x0
    "00000000", -- 5805 - 0x16ad  :    0 - 0x0
    "00000000", -- 5806 - 0x16ae  :    0 - 0x0
    "00000000", -- 5807 - 0x16af  :    0 - 0x0
    "00000000", -- 5808 - 0x16b0  :    0 - 0x0 -- Background 0x6b
    "00000000", -- 5809 - 0x16b1  :    0 - 0x0
    "00000000", -- 5810 - 0x16b2  :    0 - 0x0
    "00000000", -- 5811 - 0x16b3  :    0 - 0x0
    "00000000", -- 5812 - 0x16b4  :    0 - 0x0
    "00000000", -- 5813 - 0x16b5  :    0 - 0x0
    "00000000", -- 5814 - 0x16b6  :    0 - 0x0
    "00000000", -- 5815 - 0x16b7  :    0 - 0x0
    "00000000", -- 5816 - 0x16b8  :    0 - 0x0
    "00000000", -- 5817 - 0x16b9  :    0 - 0x0
    "00000000", -- 5818 - 0x16ba  :    0 - 0x0
    "00000000", -- 5819 - 0x16bb  :    0 - 0x0
    "00000000", -- 5820 - 0x16bc  :    0 - 0x0
    "00000000", -- 5821 - 0x16bd  :    0 - 0x0
    "00000000", -- 5822 - 0x16be  :    0 - 0x0
    "00000000", -- 5823 - 0x16bf  :    0 - 0x0
    "00000000", -- 5824 - 0x16c0  :    0 - 0x0 -- Background 0x6c
    "00000000", -- 5825 - 0x16c1  :    0 - 0x0
    "00000000", -- 5826 - 0x16c2  :    0 - 0x0
    "00000000", -- 5827 - 0x16c3  :    0 - 0x0
    "00000000", -- 5828 - 0x16c4  :    0 - 0x0
    "00000000", -- 5829 - 0x16c5  :    0 - 0x0
    "00000000", -- 5830 - 0x16c6  :    0 - 0x0
    "00000000", -- 5831 - 0x16c7  :    0 - 0x0
    "00000000", -- 5832 - 0x16c8  :    0 - 0x0
    "00000000", -- 5833 - 0x16c9  :    0 - 0x0
    "00000000", -- 5834 - 0x16ca  :    0 - 0x0
    "00000000", -- 5835 - 0x16cb  :    0 - 0x0
    "00000000", -- 5836 - 0x16cc  :    0 - 0x0
    "00000000", -- 5837 - 0x16cd  :    0 - 0x0
    "00000000", -- 5838 - 0x16ce  :    0 - 0x0
    "00000000", -- 5839 - 0x16cf  :    0 - 0x0
    "00000000", -- 5840 - 0x16d0  :    0 - 0x0 -- Background 0x6d
    "00000000", -- 5841 - 0x16d1  :    0 - 0x0
    "00000000", -- 5842 - 0x16d2  :    0 - 0x0
    "00000000", -- 5843 - 0x16d3  :    0 - 0x0
    "00000000", -- 5844 - 0x16d4  :    0 - 0x0
    "00000000", -- 5845 - 0x16d5  :    0 - 0x0
    "00000000", -- 5846 - 0x16d6  :    0 - 0x0
    "00000000", -- 5847 - 0x16d7  :    0 - 0x0
    "00000000", -- 5848 - 0x16d8  :    0 - 0x0
    "00000000", -- 5849 - 0x16d9  :    0 - 0x0
    "00000000", -- 5850 - 0x16da  :    0 - 0x0
    "00000000", -- 5851 - 0x16db  :    0 - 0x0
    "00000000", -- 5852 - 0x16dc  :    0 - 0x0
    "00000000", -- 5853 - 0x16dd  :    0 - 0x0
    "00000000", -- 5854 - 0x16de  :    0 - 0x0
    "00000000", -- 5855 - 0x16df  :    0 - 0x0
    "00000000", -- 5856 - 0x16e0  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 5857 - 0x16e1  :    0 - 0x0
    "00000000", -- 5858 - 0x16e2  :    0 - 0x0
    "00000000", -- 5859 - 0x16e3  :    0 - 0x0
    "00000000", -- 5860 - 0x16e4  :    0 - 0x0
    "00000000", -- 5861 - 0x16e5  :    0 - 0x0
    "00000000", -- 5862 - 0x16e6  :    0 - 0x0
    "00000000", -- 5863 - 0x16e7  :    0 - 0x0
    "00000000", -- 5864 - 0x16e8  :    0 - 0x0
    "00000000", -- 5865 - 0x16e9  :    0 - 0x0
    "00000000", -- 5866 - 0x16ea  :    0 - 0x0
    "00000000", -- 5867 - 0x16eb  :    0 - 0x0
    "00000000", -- 5868 - 0x16ec  :    0 - 0x0
    "00000000", -- 5869 - 0x16ed  :    0 - 0x0
    "00000000", -- 5870 - 0x16ee  :    0 - 0x0
    "00000000", -- 5871 - 0x16ef  :    0 - 0x0
    "00000000", -- 5872 - 0x16f0  :    0 - 0x0 -- Background 0x6f
    "00000000", -- 5873 - 0x16f1  :    0 - 0x0
    "00000000", -- 5874 - 0x16f2  :    0 - 0x0
    "00000000", -- 5875 - 0x16f3  :    0 - 0x0
    "00000000", -- 5876 - 0x16f4  :    0 - 0x0
    "00000000", -- 5877 - 0x16f5  :    0 - 0x0
    "00000000", -- 5878 - 0x16f6  :    0 - 0x0
    "00000000", -- 5879 - 0x16f7  :    0 - 0x0
    "00000000", -- 5880 - 0x16f8  :    0 - 0x0
    "00000000", -- 5881 - 0x16f9  :    0 - 0x0
    "00000000", -- 5882 - 0x16fa  :    0 - 0x0
    "00000000", -- 5883 - 0x16fb  :    0 - 0x0
    "00000000", -- 5884 - 0x16fc  :    0 - 0x0
    "00000000", -- 5885 - 0x16fd  :    0 - 0x0
    "00000000", -- 5886 - 0x16fe  :    0 - 0x0
    "00000000", -- 5887 - 0x16ff  :    0 - 0x0
    "00000000", -- 5888 - 0x1700  :    0 - 0x0 -- Background 0x70
    "00000000", -- 5889 - 0x1701  :    0 - 0x0
    "00000000", -- 5890 - 0x1702  :    0 - 0x0
    "00000000", -- 5891 - 0x1703  :    0 - 0x0
    "00000000", -- 5892 - 0x1704  :    0 - 0x0
    "00000000", -- 5893 - 0x1705  :    0 - 0x0
    "00000000", -- 5894 - 0x1706  :    0 - 0x0
    "00000000", -- 5895 - 0x1707  :    0 - 0x0
    "00000000", -- 5896 - 0x1708  :    0 - 0x0
    "00000000", -- 5897 - 0x1709  :    0 - 0x0
    "00000000", -- 5898 - 0x170a  :    0 - 0x0
    "00000000", -- 5899 - 0x170b  :    0 - 0x0
    "00000000", -- 5900 - 0x170c  :    0 - 0x0
    "00000000", -- 5901 - 0x170d  :    0 - 0x0
    "00000000", -- 5902 - 0x170e  :    0 - 0x0
    "00000000", -- 5903 - 0x170f  :    0 - 0x0
    "00000000", -- 5904 - 0x1710  :    0 - 0x0 -- Background 0x71
    "00000000", -- 5905 - 0x1711  :    0 - 0x0
    "00000000", -- 5906 - 0x1712  :    0 - 0x0
    "00000000", -- 5907 - 0x1713  :    0 - 0x0
    "00000000", -- 5908 - 0x1714  :    0 - 0x0
    "00000000", -- 5909 - 0x1715  :    0 - 0x0
    "00000000", -- 5910 - 0x1716  :    0 - 0x0
    "00000000", -- 5911 - 0x1717  :    0 - 0x0
    "00000000", -- 5912 - 0x1718  :    0 - 0x0
    "00000000", -- 5913 - 0x1719  :    0 - 0x0
    "00000000", -- 5914 - 0x171a  :    0 - 0x0
    "00000000", -- 5915 - 0x171b  :    0 - 0x0
    "00000000", -- 5916 - 0x171c  :    0 - 0x0
    "00000000", -- 5917 - 0x171d  :    0 - 0x0
    "00000000", -- 5918 - 0x171e  :    0 - 0x0
    "00000000", -- 5919 - 0x171f  :    0 - 0x0
    "00000000", -- 5920 - 0x1720  :    0 - 0x0 -- Background 0x72
    "00000000", -- 5921 - 0x1721  :    0 - 0x0
    "00000000", -- 5922 - 0x1722  :    0 - 0x0
    "00000000", -- 5923 - 0x1723  :    0 - 0x0
    "00000000", -- 5924 - 0x1724  :    0 - 0x0
    "00000000", -- 5925 - 0x1725  :    0 - 0x0
    "00000000", -- 5926 - 0x1726  :    0 - 0x0
    "00000000", -- 5927 - 0x1727  :    0 - 0x0
    "00000000", -- 5928 - 0x1728  :    0 - 0x0
    "00000000", -- 5929 - 0x1729  :    0 - 0x0
    "00000000", -- 5930 - 0x172a  :    0 - 0x0
    "00000000", -- 5931 - 0x172b  :    0 - 0x0
    "00000000", -- 5932 - 0x172c  :    0 - 0x0
    "00000000", -- 5933 - 0x172d  :    0 - 0x0
    "00000000", -- 5934 - 0x172e  :    0 - 0x0
    "00000000", -- 5935 - 0x172f  :    0 - 0x0
    "00000000", -- 5936 - 0x1730  :    0 - 0x0 -- Background 0x73
    "00000000", -- 5937 - 0x1731  :    0 - 0x0
    "00000000", -- 5938 - 0x1732  :    0 - 0x0
    "00000000", -- 5939 - 0x1733  :    0 - 0x0
    "00000000", -- 5940 - 0x1734  :    0 - 0x0
    "00000000", -- 5941 - 0x1735  :    0 - 0x0
    "00000000", -- 5942 - 0x1736  :    0 - 0x0
    "00000000", -- 5943 - 0x1737  :    0 - 0x0
    "00000000", -- 5944 - 0x1738  :    0 - 0x0
    "00000000", -- 5945 - 0x1739  :    0 - 0x0
    "00000000", -- 5946 - 0x173a  :    0 - 0x0
    "00000000", -- 5947 - 0x173b  :    0 - 0x0
    "00000000", -- 5948 - 0x173c  :    0 - 0x0
    "00000000", -- 5949 - 0x173d  :    0 - 0x0
    "00000000", -- 5950 - 0x173e  :    0 - 0x0
    "00000000", -- 5951 - 0x173f  :    0 - 0x0
    "00000000", -- 5952 - 0x1740  :    0 - 0x0 -- Background 0x74
    "00000000", -- 5953 - 0x1741  :    0 - 0x0
    "00000000", -- 5954 - 0x1742  :    0 - 0x0
    "00000000", -- 5955 - 0x1743  :    0 - 0x0
    "00000000", -- 5956 - 0x1744  :    0 - 0x0
    "00000000", -- 5957 - 0x1745  :    0 - 0x0
    "00000000", -- 5958 - 0x1746  :    0 - 0x0
    "00000000", -- 5959 - 0x1747  :    0 - 0x0
    "00000000", -- 5960 - 0x1748  :    0 - 0x0
    "00000000", -- 5961 - 0x1749  :    0 - 0x0
    "00000000", -- 5962 - 0x174a  :    0 - 0x0
    "00000000", -- 5963 - 0x174b  :    0 - 0x0
    "00000000", -- 5964 - 0x174c  :    0 - 0x0
    "00000000", -- 5965 - 0x174d  :    0 - 0x0
    "00000000", -- 5966 - 0x174e  :    0 - 0x0
    "00000000", -- 5967 - 0x174f  :    0 - 0x0
    "00000000", -- 5968 - 0x1750  :    0 - 0x0 -- Background 0x75
    "00000000", -- 5969 - 0x1751  :    0 - 0x0
    "00000000", -- 5970 - 0x1752  :    0 - 0x0
    "00000000", -- 5971 - 0x1753  :    0 - 0x0
    "00000000", -- 5972 - 0x1754  :    0 - 0x0
    "00000000", -- 5973 - 0x1755  :    0 - 0x0
    "00000000", -- 5974 - 0x1756  :    0 - 0x0
    "00000000", -- 5975 - 0x1757  :    0 - 0x0
    "00000000", -- 5976 - 0x1758  :    0 - 0x0
    "00000000", -- 5977 - 0x1759  :    0 - 0x0
    "00000000", -- 5978 - 0x175a  :    0 - 0x0
    "00000000", -- 5979 - 0x175b  :    0 - 0x0
    "00000000", -- 5980 - 0x175c  :    0 - 0x0
    "00000000", -- 5981 - 0x175d  :    0 - 0x0
    "00000000", -- 5982 - 0x175e  :    0 - 0x0
    "00000000", -- 5983 - 0x175f  :    0 - 0x0
    "00000000", -- 5984 - 0x1760  :    0 - 0x0 -- Background 0x76
    "00000000", -- 5985 - 0x1761  :    0 - 0x0
    "00000000", -- 5986 - 0x1762  :    0 - 0x0
    "00000000", -- 5987 - 0x1763  :    0 - 0x0
    "00000000", -- 5988 - 0x1764  :    0 - 0x0
    "00000000", -- 5989 - 0x1765  :    0 - 0x0
    "00000000", -- 5990 - 0x1766  :    0 - 0x0
    "00000000", -- 5991 - 0x1767  :    0 - 0x0
    "00000000", -- 5992 - 0x1768  :    0 - 0x0
    "00000000", -- 5993 - 0x1769  :    0 - 0x0
    "00000000", -- 5994 - 0x176a  :    0 - 0x0
    "00000000", -- 5995 - 0x176b  :    0 - 0x0
    "00000000", -- 5996 - 0x176c  :    0 - 0x0
    "00000000", -- 5997 - 0x176d  :    0 - 0x0
    "00000000", -- 5998 - 0x176e  :    0 - 0x0
    "00000000", -- 5999 - 0x176f  :    0 - 0x0
    "00000000", -- 6000 - 0x1770  :    0 - 0x0 -- Background 0x77
    "00000000", -- 6001 - 0x1771  :    0 - 0x0
    "00000000", -- 6002 - 0x1772  :    0 - 0x0
    "00000000", -- 6003 - 0x1773  :    0 - 0x0
    "00000000", -- 6004 - 0x1774  :    0 - 0x0
    "00000000", -- 6005 - 0x1775  :    0 - 0x0
    "00000000", -- 6006 - 0x1776  :    0 - 0x0
    "00000000", -- 6007 - 0x1777  :    0 - 0x0
    "00000000", -- 6008 - 0x1778  :    0 - 0x0
    "00000000", -- 6009 - 0x1779  :    0 - 0x0
    "00000000", -- 6010 - 0x177a  :    0 - 0x0
    "00000000", -- 6011 - 0x177b  :    0 - 0x0
    "00000000", -- 6012 - 0x177c  :    0 - 0x0
    "00000000", -- 6013 - 0x177d  :    0 - 0x0
    "00000000", -- 6014 - 0x177e  :    0 - 0x0
    "00000000", -- 6015 - 0x177f  :    0 - 0x0
    "00000000", -- 6016 - 0x1780  :    0 - 0x0 -- Background 0x78
    "00000000", -- 6017 - 0x1781  :    0 - 0x0
    "00000000", -- 6018 - 0x1782  :    0 - 0x0
    "00000000", -- 6019 - 0x1783  :    0 - 0x0
    "00000000", -- 6020 - 0x1784  :    0 - 0x0
    "00000000", -- 6021 - 0x1785  :    0 - 0x0
    "00000000", -- 6022 - 0x1786  :    0 - 0x0
    "00000000", -- 6023 - 0x1787  :    0 - 0x0
    "00000000", -- 6024 - 0x1788  :    0 - 0x0
    "00000000", -- 6025 - 0x1789  :    0 - 0x0
    "00000000", -- 6026 - 0x178a  :    0 - 0x0
    "00000000", -- 6027 - 0x178b  :    0 - 0x0
    "00000000", -- 6028 - 0x178c  :    0 - 0x0
    "00000000", -- 6029 - 0x178d  :    0 - 0x0
    "00000000", -- 6030 - 0x178e  :    0 - 0x0
    "00000000", -- 6031 - 0x178f  :    0 - 0x0
    "00000000", -- 6032 - 0x1790  :    0 - 0x0 -- Background 0x79
    "00000000", -- 6033 - 0x1791  :    0 - 0x0
    "00000000", -- 6034 - 0x1792  :    0 - 0x0
    "00000000", -- 6035 - 0x1793  :    0 - 0x0
    "00000000", -- 6036 - 0x1794  :    0 - 0x0
    "00000000", -- 6037 - 0x1795  :    0 - 0x0
    "00000000", -- 6038 - 0x1796  :    0 - 0x0
    "00000000", -- 6039 - 0x1797  :    0 - 0x0
    "00000000", -- 6040 - 0x1798  :    0 - 0x0
    "00000000", -- 6041 - 0x1799  :    0 - 0x0
    "00000000", -- 6042 - 0x179a  :    0 - 0x0
    "00000000", -- 6043 - 0x179b  :    0 - 0x0
    "00000000", -- 6044 - 0x179c  :    0 - 0x0
    "00000000", -- 6045 - 0x179d  :    0 - 0x0
    "00000000", -- 6046 - 0x179e  :    0 - 0x0
    "00000000", -- 6047 - 0x179f  :    0 - 0x0
    "00000000", -- 6048 - 0x17a0  :    0 - 0x0 -- Background 0x7a
    "00000000", -- 6049 - 0x17a1  :    0 - 0x0
    "00000000", -- 6050 - 0x17a2  :    0 - 0x0
    "00000000", -- 6051 - 0x17a3  :    0 - 0x0
    "00000000", -- 6052 - 0x17a4  :    0 - 0x0
    "00000000", -- 6053 - 0x17a5  :    0 - 0x0
    "00000000", -- 6054 - 0x17a6  :    0 - 0x0
    "00000000", -- 6055 - 0x17a7  :    0 - 0x0
    "00000000", -- 6056 - 0x17a8  :    0 - 0x0
    "00000000", -- 6057 - 0x17a9  :    0 - 0x0
    "00000000", -- 6058 - 0x17aa  :    0 - 0x0
    "00000000", -- 6059 - 0x17ab  :    0 - 0x0
    "00000000", -- 6060 - 0x17ac  :    0 - 0x0
    "00000000", -- 6061 - 0x17ad  :    0 - 0x0
    "00000000", -- 6062 - 0x17ae  :    0 - 0x0
    "00000000", -- 6063 - 0x17af  :    0 - 0x0
    "00000000", -- 6064 - 0x17b0  :    0 - 0x0 -- Background 0x7b
    "00000000", -- 6065 - 0x17b1  :    0 - 0x0
    "00000000", -- 6066 - 0x17b2  :    0 - 0x0
    "00000000", -- 6067 - 0x17b3  :    0 - 0x0
    "00000000", -- 6068 - 0x17b4  :    0 - 0x0
    "00000000", -- 6069 - 0x17b5  :    0 - 0x0
    "00000000", -- 6070 - 0x17b6  :    0 - 0x0
    "00000000", -- 6071 - 0x17b7  :    0 - 0x0
    "00000000", -- 6072 - 0x17b8  :    0 - 0x0
    "00000000", -- 6073 - 0x17b9  :    0 - 0x0
    "00000000", -- 6074 - 0x17ba  :    0 - 0x0
    "00000000", -- 6075 - 0x17bb  :    0 - 0x0
    "00000000", -- 6076 - 0x17bc  :    0 - 0x0
    "00000000", -- 6077 - 0x17bd  :    0 - 0x0
    "00000000", -- 6078 - 0x17be  :    0 - 0x0
    "00000000", -- 6079 - 0x17bf  :    0 - 0x0
    "00000000", -- 6080 - 0x17c0  :    0 - 0x0 -- Background 0x7c
    "00000000", -- 6081 - 0x17c1  :    0 - 0x0
    "00000000", -- 6082 - 0x17c2  :    0 - 0x0
    "00000000", -- 6083 - 0x17c3  :    0 - 0x0
    "00000000", -- 6084 - 0x17c4  :    0 - 0x0
    "00000000", -- 6085 - 0x17c5  :    0 - 0x0
    "00000000", -- 6086 - 0x17c6  :    0 - 0x0
    "00000000", -- 6087 - 0x17c7  :    0 - 0x0
    "00000000", -- 6088 - 0x17c8  :    0 - 0x0
    "00000000", -- 6089 - 0x17c9  :    0 - 0x0
    "00000000", -- 6090 - 0x17ca  :    0 - 0x0
    "00000000", -- 6091 - 0x17cb  :    0 - 0x0
    "00000000", -- 6092 - 0x17cc  :    0 - 0x0
    "00000000", -- 6093 - 0x17cd  :    0 - 0x0
    "00000000", -- 6094 - 0x17ce  :    0 - 0x0
    "00000000", -- 6095 - 0x17cf  :    0 - 0x0
    "00000000", -- 6096 - 0x17d0  :    0 - 0x0 -- Background 0x7d
    "00000000", -- 6097 - 0x17d1  :    0 - 0x0
    "00000000", -- 6098 - 0x17d2  :    0 - 0x0
    "00000000", -- 6099 - 0x17d3  :    0 - 0x0
    "00000000", -- 6100 - 0x17d4  :    0 - 0x0
    "00000000", -- 6101 - 0x17d5  :    0 - 0x0
    "00000000", -- 6102 - 0x17d6  :    0 - 0x0
    "00000000", -- 6103 - 0x17d7  :    0 - 0x0
    "00000000", -- 6104 - 0x17d8  :    0 - 0x0
    "00000000", -- 6105 - 0x17d9  :    0 - 0x0
    "00000000", -- 6106 - 0x17da  :    0 - 0x0
    "00000000", -- 6107 - 0x17db  :    0 - 0x0
    "00000000", -- 6108 - 0x17dc  :    0 - 0x0
    "00000000", -- 6109 - 0x17dd  :    0 - 0x0
    "00000000", -- 6110 - 0x17de  :    0 - 0x0
    "00000000", -- 6111 - 0x17df  :    0 - 0x0
    "00000000", -- 6112 - 0x17e0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 6113 - 0x17e1  :    0 - 0x0
    "00000000", -- 6114 - 0x17e2  :    0 - 0x0
    "00000000", -- 6115 - 0x17e3  :    0 - 0x0
    "00000000", -- 6116 - 0x17e4  :    0 - 0x0
    "00000000", -- 6117 - 0x17e5  :    0 - 0x0
    "00000000", -- 6118 - 0x17e6  :    0 - 0x0
    "00000000", -- 6119 - 0x17e7  :    0 - 0x0
    "00000000", -- 6120 - 0x17e8  :    0 - 0x0
    "00000000", -- 6121 - 0x17e9  :    0 - 0x0
    "00000000", -- 6122 - 0x17ea  :    0 - 0x0
    "00000000", -- 6123 - 0x17eb  :    0 - 0x0
    "00000000", -- 6124 - 0x17ec  :    0 - 0x0
    "00000000", -- 6125 - 0x17ed  :    0 - 0x0
    "00000000", -- 6126 - 0x17ee  :    0 - 0x0
    "00000000", -- 6127 - 0x17ef  :    0 - 0x0
    "00000000", -- 6128 - 0x17f0  :    0 - 0x0 -- Background 0x7f
    "00000000", -- 6129 - 0x17f1  :    0 - 0x0
    "00000000", -- 6130 - 0x17f2  :    0 - 0x0
    "00000000", -- 6131 - 0x17f3  :    0 - 0x0
    "00000000", -- 6132 - 0x17f4  :    0 - 0x0
    "00000000", -- 6133 - 0x17f5  :    0 - 0x0
    "00000000", -- 6134 - 0x17f6  :    0 - 0x0
    "00000000", -- 6135 - 0x17f7  :    0 - 0x0
    "00000000", -- 6136 - 0x17f8  :    0 - 0x0
    "00000000", -- 6137 - 0x17f9  :    0 - 0x0
    "00000000", -- 6138 - 0x17fa  :    0 - 0x0
    "00000000", -- 6139 - 0x17fb  :    0 - 0x0
    "00000000", -- 6140 - 0x17fc  :    0 - 0x0
    "00000000", -- 6141 - 0x17fd  :    0 - 0x0
    "00000000", -- 6142 - 0x17fe  :    0 - 0x0
    "00000000", -- 6143 - 0x17ff  :    0 - 0x0
    "00000000", -- 6144 - 0x1800  :    0 - 0x0 -- Background 0x80
    "00000000", -- 6145 - 0x1801  :    0 - 0x0
    "00000000", -- 6146 - 0x1802  :    0 - 0x0
    "00000000", -- 6147 - 0x1803  :    0 - 0x0
    "00000000", -- 6148 - 0x1804  :    0 - 0x0
    "00000000", -- 6149 - 0x1805  :    0 - 0x0
    "00000000", -- 6150 - 0x1806  :    0 - 0x0
    "00000000", -- 6151 - 0x1807  :    0 - 0x0
    "00000000", -- 6152 - 0x1808  :    0 - 0x0
    "00000000", -- 6153 - 0x1809  :    0 - 0x0
    "00000000", -- 6154 - 0x180a  :    0 - 0x0
    "00000000", -- 6155 - 0x180b  :    0 - 0x0
    "00000000", -- 6156 - 0x180c  :    0 - 0x0
    "00000000", -- 6157 - 0x180d  :    0 - 0x0
    "00000000", -- 6158 - 0x180e  :    0 - 0x0
    "00000000", -- 6159 - 0x180f  :    0 - 0x0
    "00000000", -- 6160 - 0x1810  :    0 - 0x0 -- Background 0x81
    "00000000", -- 6161 - 0x1811  :    0 - 0x0
    "00000000", -- 6162 - 0x1812  :    0 - 0x0
    "00000000", -- 6163 - 0x1813  :    0 - 0x0
    "00000000", -- 6164 - 0x1814  :    0 - 0x0
    "00000000", -- 6165 - 0x1815  :    0 - 0x0
    "00000000", -- 6166 - 0x1816  :    0 - 0x0
    "00000000", -- 6167 - 0x1817  :    0 - 0x0
    "00000000", -- 6168 - 0x1818  :    0 - 0x0
    "00000000", -- 6169 - 0x1819  :    0 - 0x0
    "00000000", -- 6170 - 0x181a  :    0 - 0x0
    "00000000", -- 6171 - 0x181b  :    0 - 0x0
    "00000000", -- 6172 - 0x181c  :    0 - 0x0
    "00000000", -- 6173 - 0x181d  :    0 - 0x0
    "00000000", -- 6174 - 0x181e  :    0 - 0x0
    "00000000", -- 6175 - 0x181f  :    0 - 0x0
    "00000000", -- 6176 - 0x1820  :    0 - 0x0 -- Background 0x82
    "00000000", -- 6177 - 0x1821  :    0 - 0x0
    "00000000", -- 6178 - 0x1822  :    0 - 0x0
    "00000000", -- 6179 - 0x1823  :    0 - 0x0
    "00000000", -- 6180 - 0x1824  :    0 - 0x0
    "00000000", -- 6181 - 0x1825  :    0 - 0x0
    "00000000", -- 6182 - 0x1826  :    0 - 0x0
    "00000000", -- 6183 - 0x1827  :    0 - 0x0
    "00000000", -- 6184 - 0x1828  :    0 - 0x0
    "00000000", -- 6185 - 0x1829  :    0 - 0x0
    "00000000", -- 6186 - 0x182a  :    0 - 0x0
    "00000000", -- 6187 - 0x182b  :    0 - 0x0
    "00000000", -- 6188 - 0x182c  :    0 - 0x0
    "00000000", -- 6189 - 0x182d  :    0 - 0x0
    "00000000", -- 6190 - 0x182e  :    0 - 0x0
    "00000000", -- 6191 - 0x182f  :    0 - 0x0
    "00000000", -- 6192 - 0x1830  :    0 - 0x0 -- Background 0x83
    "00000000", -- 6193 - 0x1831  :    0 - 0x0
    "00000000", -- 6194 - 0x1832  :    0 - 0x0
    "00000000", -- 6195 - 0x1833  :    0 - 0x0
    "00000000", -- 6196 - 0x1834  :    0 - 0x0
    "00000000", -- 6197 - 0x1835  :    0 - 0x0
    "00000000", -- 6198 - 0x1836  :    0 - 0x0
    "00000000", -- 6199 - 0x1837  :    0 - 0x0
    "00000000", -- 6200 - 0x1838  :    0 - 0x0
    "00000000", -- 6201 - 0x1839  :    0 - 0x0
    "00000000", -- 6202 - 0x183a  :    0 - 0x0
    "00000000", -- 6203 - 0x183b  :    0 - 0x0
    "00000000", -- 6204 - 0x183c  :    0 - 0x0
    "00000000", -- 6205 - 0x183d  :    0 - 0x0
    "00000000", -- 6206 - 0x183e  :    0 - 0x0
    "00000000", -- 6207 - 0x183f  :    0 - 0x0
    "00000000", -- 6208 - 0x1840  :    0 - 0x0 -- Background 0x84
    "00000000", -- 6209 - 0x1841  :    0 - 0x0
    "00000000", -- 6210 - 0x1842  :    0 - 0x0
    "00000000", -- 6211 - 0x1843  :    0 - 0x0
    "00000000", -- 6212 - 0x1844  :    0 - 0x0
    "00000000", -- 6213 - 0x1845  :    0 - 0x0
    "00000000", -- 6214 - 0x1846  :    0 - 0x0
    "00000000", -- 6215 - 0x1847  :    0 - 0x0
    "00000000", -- 6216 - 0x1848  :    0 - 0x0
    "00000000", -- 6217 - 0x1849  :    0 - 0x0
    "00000000", -- 6218 - 0x184a  :    0 - 0x0
    "00000000", -- 6219 - 0x184b  :    0 - 0x0
    "00000000", -- 6220 - 0x184c  :    0 - 0x0
    "00000000", -- 6221 - 0x184d  :    0 - 0x0
    "00000000", -- 6222 - 0x184e  :    0 - 0x0
    "00000000", -- 6223 - 0x184f  :    0 - 0x0
    "00000000", -- 6224 - 0x1850  :    0 - 0x0 -- Background 0x85
    "00000000", -- 6225 - 0x1851  :    0 - 0x0
    "00000000", -- 6226 - 0x1852  :    0 - 0x0
    "00000000", -- 6227 - 0x1853  :    0 - 0x0
    "00000000", -- 6228 - 0x1854  :    0 - 0x0
    "00000000", -- 6229 - 0x1855  :    0 - 0x0
    "00000000", -- 6230 - 0x1856  :    0 - 0x0
    "00000000", -- 6231 - 0x1857  :    0 - 0x0
    "00000000", -- 6232 - 0x1858  :    0 - 0x0
    "00000000", -- 6233 - 0x1859  :    0 - 0x0
    "00000000", -- 6234 - 0x185a  :    0 - 0x0
    "00000000", -- 6235 - 0x185b  :    0 - 0x0
    "00000000", -- 6236 - 0x185c  :    0 - 0x0
    "00000000", -- 6237 - 0x185d  :    0 - 0x0
    "00000000", -- 6238 - 0x185e  :    0 - 0x0
    "00000000", -- 6239 - 0x185f  :    0 - 0x0
    "00000000", -- 6240 - 0x1860  :    0 - 0x0 -- Background 0x86
    "00000000", -- 6241 - 0x1861  :    0 - 0x0
    "00000000", -- 6242 - 0x1862  :    0 - 0x0
    "00000000", -- 6243 - 0x1863  :    0 - 0x0
    "00000000", -- 6244 - 0x1864  :    0 - 0x0
    "00000000", -- 6245 - 0x1865  :    0 - 0x0
    "00000000", -- 6246 - 0x1866  :    0 - 0x0
    "00000000", -- 6247 - 0x1867  :    0 - 0x0
    "00000000", -- 6248 - 0x1868  :    0 - 0x0
    "00000000", -- 6249 - 0x1869  :    0 - 0x0
    "00000000", -- 6250 - 0x186a  :    0 - 0x0
    "00000000", -- 6251 - 0x186b  :    0 - 0x0
    "00000000", -- 6252 - 0x186c  :    0 - 0x0
    "00000000", -- 6253 - 0x186d  :    0 - 0x0
    "00000000", -- 6254 - 0x186e  :    0 - 0x0
    "00000000", -- 6255 - 0x186f  :    0 - 0x0
    "00000000", -- 6256 - 0x1870  :    0 - 0x0 -- Background 0x87
    "00000000", -- 6257 - 0x1871  :    0 - 0x0
    "00000000", -- 6258 - 0x1872  :    0 - 0x0
    "00000000", -- 6259 - 0x1873  :    0 - 0x0
    "00000000", -- 6260 - 0x1874  :    0 - 0x0
    "00000000", -- 6261 - 0x1875  :    0 - 0x0
    "00000000", -- 6262 - 0x1876  :    0 - 0x0
    "00000000", -- 6263 - 0x1877  :    0 - 0x0
    "00000000", -- 6264 - 0x1878  :    0 - 0x0
    "00000000", -- 6265 - 0x1879  :    0 - 0x0
    "00000000", -- 6266 - 0x187a  :    0 - 0x0
    "00000000", -- 6267 - 0x187b  :    0 - 0x0
    "00000000", -- 6268 - 0x187c  :    0 - 0x0
    "00000000", -- 6269 - 0x187d  :    0 - 0x0
    "00000000", -- 6270 - 0x187e  :    0 - 0x0
    "00000000", -- 6271 - 0x187f  :    0 - 0x0
    "00000000", -- 6272 - 0x1880  :    0 - 0x0 -- Background 0x88
    "00000000", -- 6273 - 0x1881  :    0 - 0x0
    "00000000", -- 6274 - 0x1882  :    0 - 0x0
    "00000000", -- 6275 - 0x1883  :    0 - 0x0
    "00000000", -- 6276 - 0x1884  :    0 - 0x0
    "00000000", -- 6277 - 0x1885  :    0 - 0x0
    "00000000", -- 6278 - 0x1886  :    0 - 0x0
    "00000000", -- 6279 - 0x1887  :    0 - 0x0
    "00000000", -- 6280 - 0x1888  :    0 - 0x0
    "00000000", -- 6281 - 0x1889  :    0 - 0x0
    "00000000", -- 6282 - 0x188a  :    0 - 0x0
    "00000000", -- 6283 - 0x188b  :    0 - 0x0
    "00000000", -- 6284 - 0x188c  :    0 - 0x0
    "00000000", -- 6285 - 0x188d  :    0 - 0x0
    "00000000", -- 6286 - 0x188e  :    0 - 0x0
    "00000000", -- 6287 - 0x188f  :    0 - 0x0
    "00000000", -- 6288 - 0x1890  :    0 - 0x0 -- Background 0x89
    "00000000", -- 6289 - 0x1891  :    0 - 0x0
    "00000000", -- 6290 - 0x1892  :    0 - 0x0
    "00000000", -- 6291 - 0x1893  :    0 - 0x0
    "00000000", -- 6292 - 0x1894  :    0 - 0x0
    "00000000", -- 6293 - 0x1895  :    0 - 0x0
    "00000000", -- 6294 - 0x1896  :    0 - 0x0
    "00000000", -- 6295 - 0x1897  :    0 - 0x0
    "00000000", -- 6296 - 0x1898  :    0 - 0x0
    "00000000", -- 6297 - 0x1899  :    0 - 0x0
    "00000000", -- 6298 - 0x189a  :    0 - 0x0
    "00000000", -- 6299 - 0x189b  :    0 - 0x0
    "00000000", -- 6300 - 0x189c  :    0 - 0x0
    "00000000", -- 6301 - 0x189d  :    0 - 0x0
    "00000000", -- 6302 - 0x189e  :    0 - 0x0
    "00000000", -- 6303 - 0x189f  :    0 - 0x0
    "00000000", -- 6304 - 0x18a0  :    0 - 0x0 -- Background 0x8a
    "00000000", -- 6305 - 0x18a1  :    0 - 0x0
    "00000000", -- 6306 - 0x18a2  :    0 - 0x0
    "00000000", -- 6307 - 0x18a3  :    0 - 0x0
    "00000000", -- 6308 - 0x18a4  :    0 - 0x0
    "00000000", -- 6309 - 0x18a5  :    0 - 0x0
    "00000000", -- 6310 - 0x18a6  :    0 - 0x0
    "00000000", -- 6311 - 0x18a7  :    0 - 0x0
    "00000000", -- 6312 - 0x18a8  :    0 - 0x0
    "00000000", -- 6313 - 0x18a9  :    0 - 0x0
    "00000000", -- 6314 - 0x18aa  :    0 - 0x0
    "00000000", -- 6315 - 0x18ab  :    0 - 0x0
    "00000000", -- 6316 - 0x18ac  :    0 - 0x0
    "00000000", -- 6317 - 0x18ad  :    0 - 0x0
    "00000000", -- 6318 - 0x18ae  :    0 - 0x0
    "00000000", -- 6319 - 0x18af  :    0 - 0x0
    "00000000", -- 6320 - 0x18b0  :    0 - 0x0 -- Background 0x8b
    "00000000", -- 6321 - 0x18b1  :    0 - 0x0
    "00000000", -- 6322 - 0x18b2  :    0 - 0x0
    "00000000", -- 6323 - 0x18b3  :    0 - 0x0
    "00000000", -- 6324 - 0x18b4  :    0 - 0x0
    "00000000", -- 6325 - 0x18b5  :    0 - 0x0
    "00000000", -- 6326 - 0x18b6  :    0 - 0x0
    "00000000", -- 6327 - 0x18b7  :    0 - 0x0
    "00000000", -- 6328 - 0x18b8  :    0 - 0x0
    "00000000", -- 6329 - 0x18b9  :    0 - 0x0
    "00000000", -- 6330 - 0x18ba  :    0 - 0x0
    "00000000", -- 6331 - 0x18bb  :    0 - 0x0
    "00000000", -- 6332 - 0x18bc  :    0 - 0x0
    "00000000", -- 6333 - 0x18bd  :    0 - 0x0
    "00000000", -- 6334 - 0x18be  :    0 - 0x0
    "00000000", -- 6335 - 0x18bf  :    0 - 0x0
    "00000000", -- 6336 - 0x18c0  :    0 - 0x0 -- Background 0x8c
    "00000000", -- 6337 - 0x18c1  :    0 - 0x0
    "00000000", -- 6338 - 0x18c2  :    0 - 0x0
    "00000000", -- 6339 - 0x18c3  :    0 - 0x0
    "00000000", -- 6340 - 0x18c4  :    0 - 0x0
    "00000000", -- 6341 - 0x18c5  :    0 - 0x0
    "00000000", -- 6342 - 0x18c6  :    0 - 0x0
    "00000000", -- 6343 - 0x18c7  :    0 - 0x0
    "00000000", -- 6344 - 0x18c8  :    0 - 0x0
    "00000000", -- 6345 - 0x18c9  :    0 - 0x0
    "00000000", -- 6346 - 0x18ca  :    0 - 0x0
    "00000000", -- 6347 - 0x18cb  :    0 - 0x0
    "00000000", -- 6348 - 0x18cc  :    0 - 0x0
    "00000000", -- 6349 - 0x18cd  :    0 - 0x0
    "00000000", -- 6350 - 0x18ce  :    0 - 0x0
    "00000000", -- 6351 - 0x18cf  :    0 - 0x0
    "00000000", -- 6352 - 0x18d0  :    0 - 0x0 -- Background 0x8d
    "00000000", -- 6353 - 0x18d1  :    0 - 0x0
    "00000000", -- 6354 - 0x18d2  :    0 - 0x0
    "00000000", -- 6355 - 0x18d3  :    0 - 0x0
    "00000000", -- 6356 - 0x18d4  :    0 - 0x0
    "00000000", -- 6357 - 0x18d5  :    0 - 0x0
    "00000000", -- 6358 - 0x18d6  :    0 - 0x0
    "00000000", -- 6359 - 0x18d7  :    0 - 0x0
    "00000000", -- 6360 - 0x18d8  :    0 - 0x0
    "00000000", -- 6361 - 0x18d9  :    0 - 0x0
    "00000000", -- 6362 - 0x18da  :    0 - 0x0
    "00000000", -- 6363 - 0x18db  :    0 - 0x0
    "00000000", -- 6364 - 0x18dc  :    0 - 0x0
    "00000000", -- 6365 - 0x18dd  :    0 - 0x0
    "00000000", -- 6366 - 0x18de  :    0 - 0x0
    "00000000", -- 6367 - 0x18df  :    0 - 0x0
    "00000000", -- 6368 - 0x18e0  :    0 - 0x0 -- Background 0x8e
    "00000000", -- 6369 - 0x18e1  :    0 - 0x0
    "00000000", -- 6370 - 0x18e2  :    0 - 0x0
    "00000000", -- 6371 - 0x18e3  :    0 - 0x0
    "00000000", -- 6372 - 0x18e4  :    0 - 0x0
    "00000000", -- 6373 - 0x18e5  :    0 - 0x0
    "00000000", -- 6374 - 0x18e6  :    0 - 0x0
    "00000000", -- 6375 - 0x18e7  :    0 - 0x0
    "00000000", -- 6376 - 0x18e8  :    0 - 0x0
    "00000000", -- 6377 - 0x18e9  :    0 - 0x0
    "00000000", -- 6378 - 0x18ea  :    0 - 0x0
    "00000000", -- 6379 - 0x18eb  :    0 - 0x0
    "00000000", -- 6380 - 0x18ec  :    0 - 0x0
    "00000000", -- 6381 - 0x18ed  :    0 - 0x0
    "00000000", -- 6382 - 0x18ee  :    0 - 0x0
    "00000000", -- 6383 - 0x18ef  :    0 - 0x0
    "00000000", -- 6384 - 0x18f0  :    0 - 0x0 -- Background 0x8f
    "00000000", -- 6385 - 0x18f1  :    0 - 0x0
    "00000000", -- 6386 - 0x18f2  :    0 - 0x0
    "00000000", -- 6387 - 0x18f3  :    0 - 0x0
    "00000000", -- 6388 - 0x18f4  :    0 - 0x0
    "00000000", -- 6389 - 0x18f5  :    0 - 0x0
    "00000000", -- 6390 - 0x18f6  :    0 - 0x0
    "00000000", -- 6391 - 0x18f7  :    0 - 0x0
    "00000000", -- 6392 - 0x18f8  :    0 - 0x0
    "00000000", -- 6393 - 0x18f9  :    0 - 0x0
    "00000000", -- 6394 - 0x18fa  :    0 - 0x0
    "00000000", -- 6395 - 0x18fb  :    0 - 0x0
    "00000000", -- 6396 - 0x18fc  :    0 - 0x0
    "00000000", -- 6397 - 0x18fd  :    0 - 0x0
    "00000000", -- 6398 - 0x18fe  :    0 - 0x0
    "00000000", -- 6399 - 0x18ff  :    0 - 0x0
    "00000000", -- 6400 - 0x1900  :    0 - 0x0 -- Background 0x90
    "00000000", -- 6401 - 0x1901  :    0 - 0x0
    "00000000", -- 6402 - 0x1902  :    0 - 0x0
    "00000000", -- 6403 - 0x1903  :    0 - 0x0
    "00000000", -- 6404 - 0x1904  :    0 - 0x0
    "00000000", -- 6405 - 0x1905  :    0 - 0x0
    "00000000", -- 6406 - 0x1906  :    0 - 0x0
    "00000000", -- 6407 - 0x1907  :    0 - 0x0
    "00000000", -- 6408 - 0x1908  :    0 - 0x0
    "00000000", -- 6409 - 0x1909  :    0 - 0x0
    "00000000", -- 6410 - 0x190a  :    0 - 0x0
    "00000000", -- 6411 - 0x190b  :    0 - 0x0
    "00000000", -- 6412 - 0x190c  :    0 - 0x0
    "00000000", -- 6413 - 0x190d  :    0 - 0x0
    "00000000", -- 6414 - 0x190e  :    0 - 0x0
    "00000000", -- 6415 - 0x190f  :    0 - 0x0
    "00000000", -- 6416 - 0x1910  :    0 - 0x0 -- Background 0x91
    "00000000", -- 6417 - 0x1911  :    0 - 0x0
    "00000000", -- 6418 - 0x1912  :    0 - 0x0
    "00000000", -- 6419 - 0x1913  :    0 - 0x0
    "00000000", -- 6420 - 0x1914  :    0 - 0x0
    "00000000", -- 6421 - 0x1915  :    0 - 0x0
    "00000000", -- 6422 - 0x1916  :    0 - 0x0
    "00000000", -- 6423 - 0x1917  :    0 - 0x0
    "00000000", -- 6424 - 0x1918  :    0 - 0x0
    "00000000", -- 6425 - 0x1919  :    0 - 0x0
    "00000000", -- 6426 - 0x191a  :    0 - 0x0
    "00000000", -- 6427 - 0x191b  :    0 - 0x0
    "00000000", -- 6428 - 0x191c  :    0 - 0x0
    "00000000", -- 6429 - 0x191d  :    0 - 0x0
    "00000000", -- 6430 - 0x191e  :    0 - 0x0
    "00000000", -- 6431 - 0x191f  :    0 - 0x0
    "00000000", -- 6432 - 0x1920  :    0 - 0x0 -- Background 0x92
    "00000000", -- 6433 - 0x1921  :    0 - 0x0
    "00000000", -- 6434 - 0x1922  :    0 - 0x0
    "00000000", -- 6435 - 0x1923  :    0 - 0x0
    "00000000", -- 6436 - 0x1924  :    0 - 0x0
    "00000000", -- 6437 - 0x1925  :    0 - 0x0
    "00000000", -- 6438 - 0x1926  :    0 - 0x0
    "00000000", -- 6439 - 0x1927  :    0 - 0x0
    "00000000", -- 6440 - 0x1928  :    0 - 0x0
    "00000000", -- 6441 - 0x1929  :    0 - 0x0
    "00000000", -- 6442 - 0x192a  :    0 - 0x0
    "00000000", -- 6443 - 0x192b  :    0 - 0x0
    "00000000", -- 6444 - 0x192c  :    0 - 0x0
    "00000000", -- 6445 - 0x192d  :    0 - 0x0
    "00000000", -- 6446 - 0x192e  :    0 - 0x0
    "00000000", -- 6447 - 0x192f  :    0 - 0x0
    "00000000", -- 6448 - 0x1930  :    0 - 0x0 -- Background 0x93
    "00000000", -- 6449 - 0x1931  :    0 - 0x0
    "00000000", -- 6450 - 0x1932  :    0 - 0x0
    "00000000", -- 6451 - 0x1933  :    0 - 0x0
    "00000000", -- 6452 - 0x1934  :    0 - 0x0
    "00000000", -- 6453 - 0x1935  :    0 - 0x0
    "00000000", -- 6454 - 0x1936  :    0 - 0x0
    "00000000", -- 6455 - 0x1937  :    0 - 0x0
    "00000000", -- 6456 - 0x1938  :    0 - 0x0
    "00000000", -- 6457 - 0x1939  :    0 - 0x0
    "00000000", -- 6458 - 0x193a  :    0 - 0x0
    "00000000", -- 6459 - 0x193b  :    0 - 0x0
    "00000000", -- 6460 - 0x193c  :    0 - 0x0
    "00000000", -- 6461 - 0x193d  :    0 - 0x0
    "00000000", -- 6462 - 0x193e  :    0 - 0x0
    "00000000", -- 6463 - 0x193f  :    0 - 0x0
    "00000000", -- 6464 - 0x1940  :    0 - 0x0 -- Background 0x94
    "00000000", -- 6465 - 0x1941  :    0 - 0x0
    "00000000", -- 6466 - 0x1942  :    0 - 0x0
    "00000000", -- 6467 - 0x1943  :    0 - 0x0
    "00000000", -- 6468 - 0x1944  :    0 - 0x0
    "00000000", -- 6469 - 0x1945  :    0 - 0x0
    "00000000", -- 6470 - 0x1946  :    0 - 0x0
    "00000000", -- 6471 - 0x1947  :    0 - 0x0
    "00000000", -- 6472 - 0x1948  :    0 - 0x0
    "00000000", -- 6473 - 0x1949  :    0 - 0x0
    "00000000", -- 6474 - 0x194a  :    0 - 0x0
    "00000000", -- 6475 - 0x194b  :    0 - 0x0
    "00000000", -- 6476 - 0x194c  :    0 - 0x0
    "00000000", -- 6477 - 0x194d  :    0 - 0x0
    "00000000", -- 6478 - 0x194e  :    0 - 0x0
    "00000000", -- 6479 - 0x194f  :    0 - 0x0
    "00000000", -- 6480 - 0x1950  :    0 - 0x0 -- Background 0x95
    "00000000", -- 6481 - 0x1951  :    0 - 0x0
    "00000000", -- 6482 - 0x1952  :    0 - 0x0
    "00000000", -- 6483 - 0x1953  :    0 - 0x0
    "00000000", -- 6484 - 0x1954  :    0 - 0x0
    "00000000", -- 6485 - 0x1955  :    0 - 0x0
    "00000000", -- 6486 - 0x1956  :    0 - 0x0
    "00000000", -- 6487 - 0x1957  :    0 - 0x0
    "00000000", -- 6488 - 0x1958  :    0 - 0x0
    "00000000", -- 6489 - 0x1959  :    0 - 0x0
    "00000000", -- 6490 - 0x195a  :    0 - 0x0
    "00000000", -- 6491 - 0x195b  :    0 - 0x0
    "00000000", -- 6492 - 0x195c  :    0 - 0x0
    "00000000", -- 6493 - 0x195d  :    0 - 0x0
    "00000000", -- 6494 - 0x195e  :    0 - 0x0
    "00000000", -- 6495 - 0x195f  :    0 - 0x0
    "00000000", -- 6496 - 0x1960  :    0 - 0x0 -- Background 0x96
    "00000000", -- 6497 - 0x1961  :    0 - 0x0
    "00000000", -- 6498 - 0x1962  :    0 - 0x0
    "00000000", -- 6499 - 0x1963  :    0 - 0x0
    "00000000", -- 6500 - 0x1964  :    0 - 0x0
    "00000000", -- 6501 - 0x1965  :    0 - 0x0
    "00000000", -- 6502 - 0x1966  :    0 - 0x0
    "00000000", -- 6503 - 0x1967  :    0 - 0x0
    "00000000", -- 6504 - 0x1968  :    0 - 0x0
    "00000000", -- 6505 - 0x1969  :    0 - 0x0
    "00000000", -- 6506 - 0x196a  :    0 - 0x0
    "00000000", -- 6507 - 0x196b  :    0 - 0x0
    "00000000", -- 6508 - 0x196c  :    0 - 0x0
    "00000000", -- 6509 - 0x196d  :    0 - 0x0
    "00000000", -- 6510 - 0x196e  :    0 - 0x0
    "00000000", -- 6511 - 0x196f  :    0 - 0x0
    "00000000", -- 6512 - 0x1970  :    0 - 0x0 -- Background 0x97
    "00000000", -- 6513 - 0x1971  :    0 - 0x0
    "00000000", -- 6514 - 0x1972  :    0 - 0x0
    "00000000", -- 6515 - 0x1973  :    0 - 0x0
    "00000000", -- 6516 - 0x1974  :    0 - 0x0
    "00000000", -- 6517 - 0x1975  :    0 - 0x0
    "00000000", -- 6518 - 0x1976  :    0 - 0x0
    "00000000", -- 6519 - 0x1977  :    0 - 0x0
    "00000000", -- 6520 - 0x1978  :    0 - 0x0
    "00000000", -- 6521 - 0x1979  :    0 - 0x0
    "00000000", -- 6522 - 0x197a  :    0 - 0x0
    "00000000", -- 6523 - 0x197b  :    0 - 0x0
    "00000000", -- 6524 - 0x197c  :    0 - 0x0
    "00000000", -- 6525 - 0x197d  :    0 - 0x0
    "00000000", -- 6526 - 0x197e  :    0 - 0x0
    "00000000", -- 6527 - 0x197f  :    0 - 0x0
    "00000000", -- 6528 - 0x1980  :    0 - 0x0 -- Background 0x98
    "00000000", -- 6529 - 0x1981  :    0 - 0x0
    "00000000", -- 6530 - 0x1982  :    0 - 0x0
    "00000000", -- 6531 - 0x1983  :    0 - 0x0
    "00000000", -- 6532 - 0x1984  :    0 - 0x0
    "00000000", -- 6533 - 0x1985  :    0 - 0x0
    "00000000", -- 6534 - 0x1986  :    0 - 0x0
    "00000000", -- 6535 - 0x1987  :    0 - 0x0
    "00000000", -- 6536 - 0x1988  :    0 - 0x0
    "00000000", -- 6537 - 0x1989  :    0 - 0x0
    "00000000", -- 6538 - 0x198a  :    0 - 0x0
    "00000000", -- 6539 - 0x198b  :    0 - 0x0
    "00000000", -- 6540 - 0x198c  :    0 - 0x0
    "00000000", -- 6541 - 0x198d  :    0 - 0x0
    "00000000", -- 6542 - 0x198e  :    0 - 0x0
    "00000000", -- 6543 - 0x198f  :    0 - 0x0
    "00000000", -- 6544 - 0x1990  :    0 - 0x0 -- Background 0x99
    "00000000", -- 6545 - 0x1991  :    0 - 0x0
    "00000000", -- 6546 - 0x1992  :    0 - 0x0
    "00000000", -- 6547 - 0x1993  :    0 - 0x0
    "00000000", -- 6548 - 0x1994  :    0 - 0x0
    "00000000", -- 6549 - 0x1995  :    0 - 0x0
    "00000000", -- 6550 - 0x1996  :    0 - 0x0
    "00000000", -- 6551 - 0x1997  :    0 - 0x0
    "00000000", -- 6552 - 0x1998  :    0 - 0x0
    "00000000", -- 6553 - 0x1999  :    0 - 0x0
    "00000000", -- 6554 - 0x199a  :    0 - 0x0
    "00000000", -- 6555 - 0x199b  :    0 - 0x0
    "00000000", -- 6556 - 0x199c  :    0 - 0x0
    "00000000", -- 6557 - 0x199d  :    0 - 0x0
    "00000000", -- 6558 - 0x199e  :    0 - 0x0
    "00000000", -- 6559 - 0x199f  :    0 - 0x0
    "00000000", -- 6560 - 0x19a0  :    0 - 0x0 -- Background 0x9a
    "00000000", -- 6561 - 0x19a1  :    0 - 0x0
    "00000000", -- 6562 - 0x19a2  :    0 - 0x0
    "00000000", -- 6563 - 0x19a3  :    0 - 0x0
    "00000000", -- 6564 - 0x19a4  :    0 - 0x0
    "00000000", -- 6565 - 0x19a5  :    0 - 0x0
    "00000000", -- 6566 - 0x19a6  :    0 - 0x0
    "00000000", -- 6567 - 0x19a7  :    0 - 0x0
    "00000000", -- 6568 - 0x19a8  :    0 - 0x0
    "00000000", -- 6569 - 0x19a9  :    0 - 0x0
    "00000000", -- 6570 - 0x19aa  :    0 - 0x0
    "00000000", -- 6571 - 0x19ab  :    0 - 0x0
    "00000000", -- 6572 - 0x19ac  :    0 - 0x0
    "00000000", -- 6573 - 0x19ad  :    0 - 0x0
    "00000000", -- 6574 - 0x19ae  :    0 - 0x0
    "00000000", -- 6575 - 0x19af  :    0 - 0x0
    "00000000", -- 6576 - 0x19b0  :    0 - 0x0 -- Background 0x9b
    "00000000", -- 6577 - 0x19b1  :    0 - 0x0
    "00000000", -- 6578 - 0x19b2  :    0 - 0x0
    "00000000", -- 6579 - 0x19b3  :    0 - 0x0
    "00000000", -- 6580 - 0x19b4  :    0 - 0x0
    "00000000", -- 6581 - 0x19b5  :    0 - 0x0
    "00000000", -- 6582 - 0x19b6  :    0 - 0x0
    "00000000", -- 6583 - 0x19b7  :    0 - 0x0
    "00000000", -- 6584 - 0x19b8  :    0 - 0x0
    "00000000", -- 6585 - 0x19b9  :    0 - 0x0
    "00000000", -- 6586 - 0x19ba  :    0 - 0x0
    "00000000", -- 6587 - 0x19bb  :    0 - 0x0
    "00000000", -- 6588 - 0x19bc  :    0 - 0x0
    "00000000", -- 6589 - 0x19bd  :    0 - 0x0
    "00000000", -- 6590 - 0x19be  :    0 - 0x0
    "00000000", -- 6591 - 0x19bf  :    0 - 0x0
    "00000000", -- 6592 - 0x19c0  :    0 - 0x0 -- Background 0x9c
    "00000000", -- 6593 - 0x19c1  :    0 - 0x0
    "00000000", -- 6594 - 0x19c2  :    0 - 0x0
    "00000000", -- 6595 - 0x19c3  :    0 - 0x0
    "00000000", -- 6596 - 0x19c4  :    0 - 0x0
    "00000000", -- 6597 - 0x19c5  :    0 - 0x0
    "00000000", -- 6598 - 0x19c6  :    0 - 0x0
    "00000000", -- 6599 - 0x19c7  :    0 - 0x0
    "00000000", -- 6600 - 0x19c8  :    0 - 0x0
    "00000000", -- 6601 - 0x19c9  :    0 - 0x0
    "00000000", -- 6602 - 0x19ca  :    0 - 0x0
    "00000000", -- 6603 - 0x19cb  :    0 - 0x0
    "00000000", -- 6604 - 0x19cc  :    0 - 0x0
    "00000000", -- 6605 - 0x19cd  :    0 - 0x0
    "00000000", -- 6606 - 0x19ce  :    0 - 0x0
    "00000000", -- 6607 - 0x19cf  :    0 - 0x0
    "00000000", -- 6608 - 0x19d0  :    0 - 0x0 -- Background 0x9d
    "00000000", -- 6609 - 0x19d1  :    0 - 0x0
    "00000000", -- 6610 - 0x19d2  :    0 - 0x0
    "00000000", -- 6611 - 0x19d3  :    0 - 0x0
    "00000000", -- 6612 - 0x19d4  :    0 - 0x0
    "00000000", -- 6613 - 0x19d5  :    0 - 0x0
    "00000000", -- 6614 - 0x19d6  :    0 - 0x0
    "00000000", -- 6615 - 0x19d7  :    0 - 0x0
    "00000000", -- 6616 - 0x19d8  :    0 - 0x0
    "00000000", -- 6617 - 0x19d9  :    0 - 0x0
    "00000000", -- 6618 - 0x19da  :    0 - 0x0
    "00000000", -- 6619 - 0x19db  :    0 - 0x0
    "00000000", -- 6620 - 0x19dc  :    0 - 0x0
    "00000000", -- 6621 - 0x19dd  :    0 - 0x0
    "00000000", -- 6622 - 0x19de  :    0 - 0x0
    "00000000", -- 6623 - 0x19df  :    0 - 0x0
    "00000000", -- 6624 - 0x19e0  :    0 - 0x0 -- Background 0x9e
    "00000000", -- 6625 - 0x19e1  :    0 - 0x0
    "00000000", -- 6626 - 0x19e2  :    0 - 0x0
    "00000000", -- 6627 - 0x19e3  :    0 - 0x0
    "00000000", -- 6628 - 0x19e4  :    0 - 0x0
    "00000000", -- 6629 - 0x19e5  :    0 - 0x0
    "00000000", -- 6630 - 0x19e6  :    0 - 0x0
    "00000000", -- 6631 - 0x19e7  :    0 - 0x0
    "00000000", -- 6632 - 0x19e8  :    0 - 0x0
    "00000000", -- 6633 - 0x19e9  :    0 - 0x0
    "00000000", -- 6634 - 0x19ea  :    0 - 0x0
    "00000000", -- 6635 - 0x19eb  :    0 - 0x0
    "00000000", -- 6636 - 0x19ec  :    0 - 0x0
    "00000000", -- 6637 - 0x19ed  :    0 - 0x0
    "00000000", -- 6638 - 0x19ee  :    0 - 0x0
    "00000000", -- 6639 - 0x19ef  :    0 - 0x0
    "00000000", -- 6640 - 0x19f0  :    0 - 0x0 -- Background 0x9f
    "00000000", -- 6641 - 0x19f1  :    0 - 0x0
    "00000000", -- 6642 - 0x19f2  :    0 - 0x0
    "00000000", -- 6643 - 0x19f3  :    0 - 0x0
    "00000000", -- 6644 - 0x19f4  :    0 - 0x0
    "00000000", -- 6645 - 0x19f5  :    0 - 0x0
    "00000000", -- 6646 - 0x19f6  :    0 - 0x0
    "00000000", -- 6647 - 0x19f7  :    0 - 0x0
    "00000000", -- 6648 - 0x19f8  :    0 - 0x0
    "00000000", -- 6649 - 0x19f9  :    0 - 0x0
    "00000000", -- 6650 - 0x19fa  :    0 - 0x0
    "00000000", -- 6651 - 0x19fb  :    0 - 0x0
    "00000000", -- 6652 - 0x19fc  :    0 - 0x0
    "00000000", -- 6653 - 0x19fd  :    0 - 0x0
    "00000000", -- 6654 - 0x19fe  :    0 - 0x0
    "00000000", -- 6655 - 0x19ff  :    0 - 0x0
    "00000000", -- 6656 - 0x1a00  :    0 - 0x0 -- Background 0xa0
    "00000000", -- 6657 - 0x1a01  :    0 - 0x0
    "00000000", -- 6658 - 0x1a02  :    0 - 0x0
    "00000000", -- 6659 - 0x1a03  :    0 - 0x0
    "00000000", -- 6660 - 0x1a04  :    0 - 0x0
    "00000000", -- 6661 - 0x1a05  :    0 - 0x0
    "00000000", -- 6662 - 0x1a06  :    0 - 0x0
    "00000000", -- 6663 - 0x1a07  :    0 - 0x0
    "00000000", -- 6664 - 0x1a08  :    0 - 0x0
    "00000000", -- 6665 - 0x1a09  :    0 - 0x0
    "00000000", -- 6666 - 0x1a0a  :    0 - 0x0
    "00000000", -- 6667 - 0x1a0b  :    0 - 0x0
    "00000000", -- 6668 - 0x1a0c  :    0 - 0x0
    "00000000", -- 6669 - 0x1a0d  :    0 - 0x0
    "00000000", -- 6670 - 0x1a0e  :    0 - 0x0
    "00000000", -- 6671 - 0x1a0f  :    0 - 0x0
    "00000000", -- 6672 - 0x1a10  :    0 - 0x0 -- Background 0xa1
    "00000000", -- 6673 - 0x1a11  :    0 - 0x0
    "00000000", -- 6674 - 0x1a12  :    0 - 0x0
    "00000000", -- 6675 - 0x1a13  :    0 - 0x0
    "00000000", -- 6676 - 0x1a14  :    0 - 0x0
    "00000000", -- 6677 - 0x1a15  :    0 - 0x0
    "00000000", -- 6678 - 0x1a16  :    0 - 0x0
    "00000000", -- 6679 - 0x1a17  :    0 - 0x0
    "00000000", -- 6680 - 0x1a18  :    0 - 0x0
    "00000000", -- 6681 - 0x1a19  :    0 - 0x0
    "00000000", -- 6682 - 0x1a1a  :    0 - 0x0
    "00000000", -- 6683 - 0x1a1b  :    0 - 0x0
    "00000000", -- 6684 - 0x1a1c  :    0 - 0x0
    "00000000", -- 6685 - 0x1a1d  :    0 - 0x0
    "00000000", -- 6686 - 0x1a1e  :    0 - 0x0
    "00000000", -- 6687 - 0x1a1f  :    0 - 0x0
    "00000000", -- 6688 - 0x1a20  :    0 - 0x0 -- Background 0xa2
    "00000000", -- 6689 - 0x1a21  :    0 - 0x0
    "00000000", -- 6690 - 0x1a22  :    0 - 0x0
    "00000000", -- 6691 - 0x1a23  :    0 - 0x0
    "00000000", -- 6692 - 0x1a24  :    0 - 0x0
    "00000000", -- 6693 - 0x1a25  :    0 - 0x0
    "00000000", -- 6694 - 0x1a26  :    0 - 0x0
    "00000000", -- 6695 - 0x1a27  :    0 - 0x0
    "00000000", -- 6696 - 0x1a28  :    0 - 0x0
    "00000000", -- 6697 - 0x1a29  :    0 - 0x0
    "00000000", -- 6698 - 0x1a2a  :    0 - 0x0
    "00000000", -- 6699 - 0x1a2b  :    0 - 0x0
    "00000000", -- 6700 - 0x1a2c  :    0 - 0x0
    "00000000", -- 6701 - 0x1a2d  :    0 - 0x0
    "00000000", -- 6702 - 0x1a2e  :    0 - 0x0
    "00000000", -- 6703 - 0x1a2f  :    0 - 0x0
    "00000000", -- 6704 - 0x1a30  :    0 - 0x0 -- Background 0xa3
    "00000000", -- 6705 - 0x1a31  :    0 - 0x0
    "00000000", -- 6706 - 0x1a32  :    0 - 0x0
    "00000000", -- 6707 - 0x1a33  :    0 - 0x0
    "00000000", -- 6708 - 0x1a34  :    0 - 0x0
    "00000000", -- 6709 - 0x1a35  :    0 - 0x0
    "00000000", -- 6710 - 0x1a36  :    0 - 0x0
    "00000000", -- 6711 - 0x1a37  :    0 - 0x0
    "00000000", -- 6712 - 0x1a38  :    0 - 0x0
    "00000000", -- 6713 - 0x1a39  :    0 - 0x0
    "00000000", -- 6714 - 0x1a3a  :    0 - 0x0
    "00000000", -- 6715 - 0x1a3b  :    0 - 0x0
    "00000000", -- 6716 - 0x1a3c  :    0 - 0x0
    "00000000", -- 6717 - 0x1a3d  :    0 - 0x0
    "00000000", -- 6718 - 0x1a3e  :    0 - 0x0
    "00000000", -- 6719 - 0x1a3f  :    0 - 0x0
    "00000000", -- 6720 - 0x1a40  :    0 - 0x0 -- Background 0xa4
    "00000000", -- 6721 - 0x1a41  :    0 - 0x0
    "00000000", -- 6722 - 0x1a42  :    0 - 0x0
    "00000000", -- 6723 - 0x1a43  :    0 - 0x0
    "00000000", -- 6724 - 0x1a44  :    0 - 0x0
    "00000000", -- 6725 - 0x1a45  :    0 - 0x0
    "00000000", -- 6726 - 0x1a46  :    0 - 0x0
    "00000000", -- 6727 - 0x1a47  :    0 - 0x0
    "00000000", -- 6728 - 0x1a48  :    0 - 0x0
    "00000000", -- 6729 - 0x1a49  :    0 - 0x0
    "00000000", -- 6730 - 0x1a4a  :    0 - 0x0
    "00000000", -- 6731 - 0x1a4b  :    0 - 0x0
    "00000000", -- 6732 - 0x1a4c  :    0 - 0x0
    "00000000", -- 6733 - 0x1a4d  :    0 - 0x0
    "00000000", -- 6734 - 0x1a4e  :    0 - 0x0
    "00000000", -- 6735 - 0x1a4f  :    0 - 0x0
    "00000000", -- 6736 - 0x1a50  :    0 - 0x0 -- Background 0xa5
    "00000000", -- 6737 - 0x1a51  :    0 - 0x0
    "00000000", -- 6738 - 0x1a52  :    0 - 0x0
    "00000000", -- 6739 - 0x1a53  :    0 - 0x0
    "00000000", -- 6740 - 0x1a54  :    0 - 0x0
    "00000000", -- 6741 - 0x1a55  :    0 - 0x0
    "00000000", -- 6742 - 0x1a56  :    0 - 0x0
    "00000000", -- 6743 - 0x1a57  :    0 - 0x0
    "00000000", -- 6744 - 0x1a58  :    0 - 0x0
    "00000000", -- 6745 - 0x1a59  :    0 - 0x0
    "00000000", -- 6746 - 0x1a5a  :    0 - 0x0
    "00000000", -- 6747 - 0x1a5b  :    0 - 0x0
    "00000000", -- 6748 - 0x1a5c  :    0 - 0x0
    "00000000", -- 6749 - 0x1a5d  :    0 - 0x0
    "00000000", -- 6750 - 0x1a5e  :    0 - 0x0
    "00000000", -- 6751 - 0x1a5f  :    0 - 0x0
    "00000000", -- 6752 - 0x1a60  :    0 - 0x0 -- Background 0xa6
    "00000000", -- 6753 - 0x1a61  :    0 - 0x0
    "00000000", -- 6754 - 0x1a62  :    0 - 0x0
    "00000000", -- 6755 - 0x1a63  :    0 - 0x0
    "00000000", -- 6756 - 0x1a64  :    0 - 0x0
    "00000000", -- 6757 - 0x1a65  :    0 - 0x0
    "00000000", -- 6758 - 0x1a66  :    0 - 0x0
    "00000000", -- 6759 - 0x1a67  :    0 - 0x0
    "00000000", -- 6760 - 0x1a68  :    0 - 0x0
    "00000000", -- 6761 - 0x1a69  :    0 - 0x0
    "00000000", -- 6762 - 0x1a6a  :    0 - 0x0
    "00000000", -- 6763 - 0x1a6b  :    0 - 0x0
    "00000000", -- 6764 - 0x1a6c  :    0 - 0x0
    "00000000", -- 6765 - 0x1a6d  :    0 - 0x0
    "00000000", -- 6766 - 0x1a6e  :    0 - 0x0
    "00000000", -- 6767 - 0x1a6f  :    0 - 0x0
    "00000000", -- 6768 - 0x1a70  :    0 - 0x0 -- Background 0xa7
    "00000000", -- 6769 - 0x1a71  :    0 - 0x0
    "00000000", -- 6770 - 0x1a72  :    0 - 0x0
    "00000000", -- 6771 - 0x1a73  :    0 - 0x0
    "00000000", -- 6772 - 0x1a74  :    0 - 0x0
    "00000000", -- 6773 - 0x1a75  :    0 - 0x0
    "00000000", -- 6774 - 0x1a76  :    0 - 0x0
    "00000000", -- 6775 - 0x1a77  :    0 - 0x0
    "00000000", -- 6776 - 0x1a78  :    0 - 0x0
    "00000000", -- 6777 - 0x1a79  :    0 - 0x0
    "00000000", -- 6778 - 0x1a7a  :    0 - 0x0
    "00000000", -- 6779 - 0x1a7b  :    0 - 0x0
    "00000000", -- 6780 - 0x1a7c  :    0 - 0x0
    "00000000", -- 6781 - 0x1a7d  :    0 - 0x0
    "00000000", -- 6782 - 0x1a7e  :    0 - 0x0
    "00000000", -- 6783 - 0x1a7f  :    0 - 0x0
    "00000000", -- 6784 - 0x1a80  :    0 - 0x0 -- Background 0xa8
    "00000000", -- 6785 - 0x1a81  :    0 - 0x0
    "00000000", -- 6786 - 0x1a82  :    0 - 0x0
    "00000000", -- 6787 - 0x1a83  :    0 - 0x0
    "00000000", -- 6788 - 0x1a84  :    0 - 0x0
    "00000000", -- 6789 - 0x1a85  :    0 - 0x0
    "00000000", -- 6790 - 0x1a86  :    0 - 0x0
    "00000000", -- 6791 - 0x1a87  :    0 - 0x0
    "00000000", -- 6792 - 0x1a88  :    0 - 0x0
    "00000000", -- 6793 - 0x1a89  :    0 - 0x0
    "00000000", -- 6794 - 0x1a8a  :    0 - 0x0
    "00000000", -- 6795 - 0x1a8b  :    0 - 0x0
    "00000000", -- 6796 - 0x1a8c  :    0 - 0x0
    "00000000", -- 6797 - 0x1a8d  :    0 - 0x0
    "00000000", -- 6798 - 0x1a8e  :    0 - 0x0
    "00000000", -- 6799 - 0x1a8f  :    0 - 0x0
    "00000000", -- 6800 - 0x1a90  :    0 - 0x0 -- Background 0xa9
    "00000000", -- 6801 - 0x1a91  :    0 - 0x0
    "00000000", -- 6802 - 0x1a92  :    0 - 0x0
    "00000000", -- 6803 - 0x1a93  :    0 - 0x0
    "00000000", -- 6804 - 0x1a94  :    0 - 0x0
    "00000000", -- 6805 - 0x1a95  :    0 - 0x0
    "00000000", -- 6806 - 0x1a96  :    0 - 0x0
    "00000000", -- 6807 - 0x1a97  :    0 - 0x0
    "00000000", -- 6808 - 0x1a98  :    0 - 0x0
    "00000000", -- 6809 - 0x1a99  :    0 - 0x0
    "00000000", -- 6810 - 0x1a9a  :    0 - 0x0
    "00000000", -- 6811 - 0x1a9b  :    0 - 0x0
    "00000000", -- 6812 - 0x1a9c  :    0 - 0x0
    "00000000", -- 6813 - 0x1a9d  :    0 - 0x0
    "00000000", -- 6814 - 0x1a9e  :    0 - 0x0
    "00000000", -- 6815 - 0x1a9f  :    0 - 0x0
    "00000000", -- 6816 - 0x1aa0  :    0 - 0x0 -- Background 0xaa
    "00000000", -- 6817 - 0x1aa1  :    0 - 0x0
    "00000000", -- 6818 - 0x1aa2  :    0 - 0x0
    "00000000", -- 6819 - 0x1aa3  :    0 - 0x0
    "00000000", -- 6820 - 0x1aa4  :    0 - 0x0
    "00000000", -- 6821 - 0x1aa5  :    0 - 0x0
    "00000000", -- 6822 - 0x1aa6  :    0 - 0x0
    "00000000", -- 6823 - 0x1aa7  :    0 - 0x0
    "00000000", -- 6824 - 0x1aa8  :    0 - 0x0
    "00000000", -- 6825 - 0x1aa9  :    0 - 0x0
    "00000000", -- 6826 - 0x1aaa  :    0 - 0x0
    "00000000", -- 6827 - 0x1aab  :    0 - 0x0
    "00000000", -- 6828 - 0x1aac  :    0 - 0x0
    "00000000", -- 6829 - 0x1aad  :    0 - 0x0
    "00000000", -- 6830 - 0x1aae  :    0 - 0x0
    "00000000", -- 6831 - 0x1aaf  :    0 - 0x0
    "00000000", -- 6832 - 0x1ab0  :    0 - 0x0 -- Background 0xab
    "00000000", -- 6833 - 0x1ab1  :    0 - 0x0
    "00000000", -- 6834 - 0x1ab2  :    0 - 0x0
    "00000000", -- 6835 - 0x1ab3  :    0 - 0x0
    "00000000", -- 6836 - 0x1ab4  :    0 - 0x0
    "00000000", -- 6837 - 0x1ab5  :    0 - 0x0
    "00000000", -- 6838 - 0x1ab6  :    0 - 0x0
    "00000000", -- 6839 - 0x1ab7  :    0 - 0x0
    "00000000", -- 6840 - 0x1ab8  :    0 - 0x0
    "00000000", -- 6841 - 0x1ab9  :    0 - 0x0
    "00000000", -- 6842 - 0x1aba  :    0 - 0x0
    "00000000", -- 6843 - 0x1abb  :    0 - 0x0
    "00000000", -- 6844 - 0x1abc  :    0 - 0x0
    "00000000", -- 6845 - 0x1abd  :    0 - 0x0
    "00000000", -- 6846 - 0x1abe  :    0 - 0x0
    "00000000", -- 6847 - 0x1abf  :    0 - 0x0
    "00000000", -- 6848 - 0x1ac0  :    0 - 0x0 -- Background 0xac
    "00000000", -- 6849 - 0x1ac1  :    0 - 0x0
    "00000000", -- 6850 - 0x1ac2  :    0 - 0x0
    "00000000", -- 6851 - 0x1ac3  :    0 - 0x0
    "00000000", -- 6852 - 0x1ac4  :    0 - 0x0
    "00000000", -- 6853 - 0x1ac5  :    0 - 0x0
    "00000000", -- 6854 - 0x1ac6  :    0 - 0x0
    "00000000", -- 6855 - 0x1ac7  :    0 - 0x0
    "00000000", -- 6856 - 0x1ac8  :    0 - 0x0
    "00000000", -- 6857 - 0x1ac9  :    0 - 0x0
    "00000000", -- 6858 - 0x1aca  :    0 - 0x0
    "00000000", -- 6859 - 0x1acb  :    0 - 0x0
    "00000000", -- 6860 - 0x1acc  :    0 - 0x0
    "00000000", -- 6861 - 0x1acd  :    0 - 0x0
    "00000000", -- 6862 - 0x1ace  :    0 - 0x0
    "00000000", -- 6863 - 0x1acf  :    0 - 0x0
    "00000000", -- 6864 - 0x1ad0  :    0 - 0x0 -- Background 0xad
    "00000000", -- 6865 - 0x1ad1  :    0 - 0x0
    "00000000", -- 6866 - 0x1ad2  :    0 - 0x0
    "00000000", -- 6867 - 0x1ad3  :    0 - 0x0
    "00000000", -- 6868 - 0x1ad4  :    0 - 0x0
    "00000000", -- 6869 - 0x1ad5  :    0 - 0x0
    "00000000", -- 6870 - 0x1ad6  :    0 - 0x0
    "00000000", -- 6871 - 0x1ad7  :    0 - 0x0
    "00000000", -- 6872 - 0x1ad8  :    0 - 0x0
    "00000000", -- 6873 - 0x1ad9  :    0 - 0x0
    "00000000", -- 6874 - 0x1ada  :    0 - 0x0
    "00000000", -- 6875 - 0x1adb  :    0 - 0x0
    "00000000", -- 6876 - 0x1adc  :    0 - 0x0
    "00000000", -- 6877 - 0x1add  :    0 - 0x0
    "00000000", -- 6878 - 0x1ade  :    0 - 0x0
    "00000000", -- 6879 - 0x1adf  :    0 - 0x0
    "00000000", -- 6880 - 0x1ae0  :    0 - 0x0 -- Background 0xae
    "00000000", -- 6881 - 0x1ae1  :    0 - 0x0
    "00000000", -- 6882 - 0x1ae2  :    0 - 0x0
    "00000000", -- 6883 - 0x1ae3  :    0 - 0x0
    "00000000", -- 6884 - 0x1ae4  :    0 - 0x0
    "00000000", -- 6885 - 0x1ae5  :    0 - 0x0
    "00000000", -- 6886 - 0x1ae6  :    0 - 0x0
    "00000000", -- 6887 - 0x1ae7  :    0 - 0x0
    "00000000", -- 6888 - 0x1ae8  :    0 - 0x0
    "00000000", -- 6889 - 0x1ae9  :    0 - 0x0
    "00000000", -- 6890 - 0x1aea  :    0 - 0x0
    "00000000", -- 6891 - 0x1aeb  :    0 - 0x0
    "00000000", -- 6892 - 0x1aec  :    0 - 0x0
    "00000000", -- 6893 - 0x1aed  :    0 - 0x0
    "00000000", -- 6894 - 0x1aee  :    0 - 0x0
    "00000000", -- 6895 - 0x1aef  :    0 - 0x0
    "00000000", -- 6896 - 0x1af0  :    0 - 0x0 -- Background 0xaf
    "00000000", -- 6897 - 0x1af1  :    0 - 0x0
    "00000000", -- 6898 - 0x1af2  :    0 - 0x0
    "00000000", -- 6899 - 0x1af3  :    0 - 0x0
    "00000000", -- 6900 - 0x1af4  :    0 - 0x0
    "00000000", -- 6901 - 0x1af5  :    0 - 0x0
    "00000000", -- 6902 - 0x1af6  :    0 - 0x0
    "00000000", -- 6903 - 0x1af7  :    0 - 0x0
    "00000000", -- 6904 - 0x1af8  :    0 - 0x0
    "00000000", -- 6905 - 0x1af9  :    0 - 0x0
    "00000000", -- 6906 - 0x1afa  :    0 - 0x0
    "00000000", -- 6907 - 0x1afb  :    0 - 0x0
    "00000000", -- 6908 - 0x1afc  :    0 - 0x0
    "00000000", -- 6909 - 0x1afd  :    0 - 0x0
    "00000000", -- 6910 - 0x1afe  :    0 - 0x0
    "00000000", -- 6911 - 0x1aff  :    0 - 0x0
    "00000000", -- 6912 - 0x1b00  :    0 - 0x0 -- Background 0xb0
    "00000000", -- 6913 - 0x1b01  :    0 - 0x0
    "00000000", -- 6914 - 0x1b02  :    0 - 0x0
    "00000000", -- 6915 - 0x1b03  :    0 - 0x0
    "00000000", -- 6916 - 0x1b04  :    0 - 0x0
    "00000000", -- 6917 - 0x1b05  :    0 - 0x0
    "00000000", -- 6918 - 0x1b06  :    0 - 0x0
    "00000000", -- 6919 - 0x1b07  :    0 - 0x0
    "00000000", -- 6920 - 0x1b08  :    0 - 0x0
    "00000000", -- 6921 - 0x1b09  :    0 - 0x0
    "00000000", -- 6922 - 0x1b0a  :    0 - 0x0
    "00000000", -- 6923 - 0x1b0b  :    0 - 0x0
    "00000000", -- 6924 - 0x1b0c  :    0 - 0x0
    "00000000", -- 6925 - 0x1b0d  :    0 - 0x0
    "00000000", -- 6926 - 0x1b0e  :    0 - 0x0
    "00000000", -- 6927 - 0x1b0f  :    0 - 0x0
    "00000000", -- 6928 - 0x1b10  :    0 - 0x0 -- Background 0xb1
    "00000000", -- 6929 - 0x1b11  :    0 - 0x0
    "00000000", -- 6930 - 0x1b12  :    0 - 0x0
    "00000000", -- 6931 - 0x1b13  :    0 - 0x0
    "00000000", -- 6932 - 0x1b14  :    0 - 0x0
    "00000000", -- 6933 - 0x1b15  :    0 - 0x0
    "00000000", -- 6934 - 0x1b16  :    0 - 0x0
    "00000000", -- 6935 - 0x1b17  :    0 - 0x0
    "00000000", -- 6936 - 0x1b18  :    0 - 0x0
    "00000000", -- 6937 - 0x1b19  :    0 - 0x0
    "00000000", -- 6938 - 0x1b1a  :    0 - 0x0
    "00000000", -- 6939 - 0x1b1b  :    0 - 0x0
    "00000000", -- 6940 - 0x1b1c  :    0 - 0x0
    "00000000", -- 6941 - 0x1b1d  :    0 - 0x0
    "00000000", -- 6942 - 0x1b1e  :    0 - 0x0
    "00000000", -- 6943 - 0x1b1f  :    0 - 0x0
    "00000000", -- 6944 - 0x1b20  :    0 - 0x0 -- Background 0xb2
    "00000000", -- 6945 - 0x1b21  :    0 - 0x0
    "00000000", -- 6946 - 0x1b22  :    0 - 0x0
    "00000000", -- 6947 - 0x1b23  :    0 - 0x0
    "00000000", -- 6948 - 0x1b24  :    0 - 0x0
    "00000000", -- 6949 - 0x1b25  :    0 - 0x0
    "00000000", -- 6950 - 0x1b26  :    0 - 0x0
    "00000000", -- 6951 - 0x1b27  :    0 - 0x0
    "00000000", -- 6952 - 0x1b28  :    0 - 0x0
    "00000000", -- 6953 - 0x1b29  :    0 - 0x0
    "00000000", -- 6954 - 0x1b2a  :    0 - 0x0
    "00000000", -- 6955 - 0x1b2b  :    0 - 0x0
    "00000000", -- 6956 - 0x1b2c  :    0 - 0x0
    "00000000", -- 6957 - 0x1b2d  :    0 - 0x0
    "00000000", -- 6958 - 0x1b2e  :    0 - 0x0
    "00000000", -- 6959 - 0x1b2f  :    0 - 0x0
    "00000000", -- 6960 - 0x1b30  :    0 - 0x0 -- Background 0xb3
    "00000000", -- 6961 - 0x1b31  :    0 - 0x0
    "00000000", -- 6962 - 0x1b32  :    0 - 0x0
    "00000000", -- 6963 - 0x1b33  :    0 - 0x0
    "00000000", -- 6964 - 0x1b34  :    0 - 0x0
    "00000000", -- 6965 - 0x1b35  :    0 - 0x0
    "00000000", -- 6966 - 0x1b36  :    0 - 0x0
    "00000000", -- 6967 - 0x1b37  :    0 - 0x0
    "00000000", -- 6968 - 0x1b38  :    0 - 0x0
    "00000000", -- 6969 - 0x1b39  :    0 - 0x0
    "00000000", -- 6970 - 0x1b3a  :    0 - 0x0
    "00000000", -- 6971 - 0x1b3b  :    0 - 0x0
    "00000000", -- 6972 - 0x1b3c  :    0 - 0x0
    "00000000", -- 6973 - 0x1b3d  :    0 - 0x0
    "00000000", -- 6974 - 0x1b3e  :    0 - 0x0
    "00000000", -- 6975 - 0x1b3f  :    0 - 0x0
    "00000000", -- 6976 - 0x1b40  :    0 - 0x0 -- Background 0xb4
    "00000000", -- 6977 - 0x1b41  :    0 - 0x0
    "00000000", -- 6978 - 0x1b42  :    0 - 0x0
    "00000000", -- 6979 - 0x1b43  :    0 - 0x0
    "00000000", -- 6980 - 0x1b44  :    0 - 0x0
    "00000000", -- 6981 - 0x1b45  :    0 - 0x0
    "00000000", -- 6982 - 0x1b46  :    0 - 0x0
    "00000000", -- 6983 - 0x1b47  :    0 - 0x0
    "00000000", -- 6984 - 0x1b48  :    0 - 0x0
    "00000000", -- 6985 - 0x1b49  :    0 - 0x0
    "00000000", -- 6986 - 0x1b4a  :    0 - 0x0
    "00000000", -- 6987 - 0x1b4b  :    0 - 0x0
    "00000000", -- 6988 - 0x1b4c  :    0 - 0x0
    "00000000", -- 6989 - 0x1b4d  :    0 - 0x0
    "00000000", -- 6990 - 0x1b4e  :    0 - 0x0
    "00000000", -- 6991 - 0x1b4f  :    0 - 0x0
    "00000000", -- 6992 - 0x1b50  :    0 - 0x0 -- Background 0xb5
    "00000000", -- 6993 - 0x1b51  :    0 - 0x0
    "00000000", -- 6994 - 0x1b52  :    0 - 0x0
    "00000000", -- 6995 - 0x1b53  :    0 - 0x0
    "00000000", -- 6996 - 0x1b54  :    0 - 0x0
    "00000000", -- 6997 - 0x1b55  :    0 - 0x0
    "00000000", -- 6998 - 0x1b56  :    0 - 0x0
    "00000000", -- 6999 - 0x1b57  :    0 - 0x0
    "00000000", -- 7000 - 0x1b58  :    0 - 0x0
    "00000000", -- 7001 - 0x1b59  :    0 - 0x0
    "00000000", -- 7002 - 0x1b5a  :    0 - 0x0
    "00000000", -- 7003 - 0x1b5b  :    0 - 0x0
    "00000000", -- 7004 - 0x1b5c  :    0 - 0x0
    "00000000", -- 7005 - 0x1b5d  :    0 - 0x0
    "00000000", -- 7006 - 0x1b5e  :    0 - 0x0
    "00000000", -- 7007 - 0x1b5f  :    0 - 0x0
    "00000000", -- 7008 - 0x1b60  :    0 - 0x0 -- Background 0xb6
    "00000000", -- 7009 - 0x1b61  :    0 - 0x0
    "00000000", -- 7010 - 0x1b62  :    0 - 0x0
    "00000000", -- 7011 - 0x1b63  :    0 - 0x0
    "00000000", -- 7012 - 0x1b64  :    0 - 0x0
    "00000000", -- 7013 - 0x1b65  :    0 - 0x0
    "00000000", -- 7014 - 0x1b66  :    0 - 0x0
    "00000000", -- 7015 - 0x1b67  :    0 - 0x0
    "00000000", -- 7016 - 0x1b68  :    0 - 0x0
    "00000000", -- 7017 - 0x1b69  :    0 - 0x0
    "00000000", -- 7018 - 0x1b6a  :    0 - 0x0
    "00000000", -- 7019 - 0x1b6b  :    0 - 0x0
    "00000000", -- 7020 - 0x1b6c  :    0 - 0x0
    "00000000", -- 7021 - 0x1b6d  :    0 - 0x0
    "00000000", -- 7022 - 0x1b6e  :    0 - 0x0
    "00000000", -- 7023 - 0x1b6f  :    0 - 0x0
    "00000000", -- 7024 - 0x1b70  :    0 - 0x0 -- Background 0xb7
    "00000000", -- 7025 - 0x1b71  :    0 - 0x0
    "00000000", -- 7026 - 0x1b72  :    0 - 0x0
    "00000000", -- 7027 - 0x1b73  :    0 - 0x0
    "00000000", -- 7028 - 0x1b74  :    0 - 0x0
    "00000000", -- 7029 - 0x1b75  :    0 - 0x0
    "00000000", -- 7030 - 0x1b76  :    0 - 0x0
    "00000000", -- 7031 - 0x1b77  :    0 - 0x0
    "00000000", -- 7032 - 0x1b78  :    0 - 0x0
    "00000000", -- 7033 - 0x1b79  :    0 - 0x0
    "00000000", -- 7034 - 0x1b7a  :    0 - 0x0
    "00000000", -- 7035 - 0x1b7b  :    0 - 0x0
    "00000000", -- 7036 - 0x1b7c  :    0 - 0x0
    "00000000", -- 7037 - 0x1b7d  :    0 - 0x0
    "00000000", -- 7038 - 0x1b7e  :    0 - 0x0
    "00000000", -- 7039 - 0x1b7f  :    0 - 0x0
    "00000000", -- 7040 - 0x1b80  :    0 - 0x0 -- Background 0xb8
    "00000000", -- 7041 - 0x1b81  :    0 - 0x0
    "00000000", -- 7042 - 0x1b82  :    0 - 0x0
    "00000000", -- 7043 - 0x1b83  :    0 - 0x0
    "00000000", -- 7044 - 0x1b84  :    0 - 0x0
    "00000000", -- 7045 - 0x1b85  :    0 - 0x0
    "00000000", -- 7046 - 0x1b86  :    0 - 0x0
    "00000000", -- 7047 - 0x1b87  :    0 - 0x0
    "00000000", -- 7048 - 0x1b88  :    0 - 0x0
    "00000000", -- 7049 - 0x1b89  :    0 - 0x0
    "00000000", -- 7050 - 0x1b8a  :    0 - 0x0
    "00000000", -- 7051 - 0x1b8b  :    0 - 0x0
    "00000000", -- 7052 - 0x1b8c  :    0 - 0x0
    "00000000", -- 7053 - 0x1b8d  :    0 - 0x0
    "00000000", -- 7054 - 0x1b8e  :    0 - 0x0
    "00000000", -- 7055 - 0x1b8f  :    0 - 0x0
    "00000000", -- 7056 - 0x1b90  :    0 - 0x0 -- Background 0xb9
    "00000000", -- 7057 - 0x1b91  :    0 - 0x0
    "00000000", -- 7058 - 0x1b92  :    0 - 0x0
    "00000000", -- 7059 - 0x1b93  :    0 - 0x0
    "00000000", -- 7060 - 0x1b94  :    0 - 0x0
    "00000000", -- 7061 - 0x1b95  :    0 - 0x0
    "00000000", -- 7062 - 0x1b96  :    0 - 0x0
    "00000000", -- 7063 - 0x1b97  :    0 - 0x0
    "00000000", -- 7064 - 0x1b98  :    0 - 0x0
    "00000000", -- 7065 - 0x1b99  :    0 - 0x0
    "00000000", -- 7066 - 0x1b9a  :    0 - 0x0
    "00000000", -- 7067 - 0x1b9b  :    0 - 0x0
    "00000000", -- 7068 - 0x1b9c  :    0 - 0x0
    "00000000", -- 7069 - 0x1b9d  :    0 - 0x0
    "00000000", -- 7070 - 0x1b9e  :    0 - 0x0
    "00000000", -- 7071 - 0x1b9f  :    0 - 0x0
    "00000000", -- 7072 - 0x1ba0  :    0 - 0x0 -- Background 0xba
    "00000000", -- 7073 - 0x1ba1  :    0 - 0x0
    "00000000", -- 7074 - 0x1ba2  :    0 - 0x0
    "00000000", -- 7075 - 0x1ba3  :    0 - 0x0
    "00000000", -- 7076 - 0x1ba4  :    0 - 0x0
    "00000000", -- 7077 - 0x1ba5  :    0 - 0x0
    "00000000", -- 7078 - 0x1ba6  :    0 - 0x0
    "00000000", -- 7079 - 0x1ba7  :    0 - 0x0
    "00000000", -- 7080 - 0x1ba8  :    0 - 0x0
    "00000000", -- 7081 - 0x1ba9  :    0 - 0x0
    "00000000", -- 7082 - 0x1baa  :    0 - 0x0
    "00000000", -- 7083 - 0x1bab  :    0 - 0x0
    "00000000", -- 7084 - 0x1bac  :    0 - 0x0
    "00000000", -- 7085 - 0x1bad  :    0 - 0x0
    "00000000", -- 7086 - 0x1bae  :    0 - 0x0
    "00000000", -- 7087 - 0x1baf  :    0 - 0x0
    "00000000", -- 7088 - 0x1bb0  :    0 - 0x0 -- Background 0xbb
    "00000000", -- 7089 - 0x1bb1  :    0 - 0x0
    "00000000", -- 7090 - 0x1bb2  :    0 - 0x0
    "00000000", -- 7091 - 0x1bb3  :    0 - 0x0
    "00000000", -- 7092 - 0x1bb4  :    0 - 0x0
    "00000000", -- 7093 - 0x1bb5  :    0 - 0x0
    "00000000", -- 7094 - 0x1bb6  :    0 - 0x0
    "00000000", -- 7095 - 0x1bb7  :    0 - 0x0
    "00000000", -- 7096 - 0x1bb8  :    0 - 0x0
    "00000000", -- 7097 - 0x1bb9  :    0 - 0x0
    "00000000", -- 7098 - 0x1bba  :    0 - 0x0
    "00000000", -- 7099 - 0x1bbb  :    0 - 0x0
    "00000000", -- 7100 - 0x1bbc  :    0 - 0x0
    "00000000", -- 7101 - 0x1bbd  :    0 - 0x0
    "00000000", -- 7102 - 0x1bbe  :    0 - 0x0
    "00000000", -- 7103 - 0x1bbf  :    0 - 0x0
    "00000000", -- 7104 - 0x1bc0  :    0 - 0x0 -- Background 0xbc
    "00000000", -- 7105 - 0x1bc1  :    0 - 0x0
    "00000000", -- 7106 - 0x1bc2  :    0 - 0x0
    "00000000", -- 7107 - 0x1bc3  :    0 - 0x0
    "00000000", -- 7108 - 0x1bc4  :    0 - 0x0
    "00000000", -- 7109 - 0x1bc5  :    0 - 0x0
    "00000000", -- 7110 - 0x1bc6  :    0 - 0x0
    "00000000", -- 7111 - 0x1bc7  :    0 - 0x0
    "00000000", -- 7112 - 0x1bc8  :    0 - 0x0
    "00000000", -- 7113 - 0x1bc9  :    0 - 0x0
    "00000000", -- 7114 - 0x1bca  :    0 - 0x0
    "00000000", -- 7115 - 0x1bcb  :    0 - 0x0
    "00000000", -- 7116 - 0x1bcc  :    0 - 0x0
    "00000000", -- 7117 - 0x1bcd  :    0 - 0x0
    "00000000", -- 7118 - 0x1bce  :    0 - 0x0
    "00000000", -- 7119 - 0x1bcf  :    0 - 0x0
    "00000000", -- 7120 - 0x1bd0  :    0 - 0x0 -- Background 0xbd
    "00000000", -- 7121 - 0x1bd1  :    0 - 0x0
    "00000000", -- 7122 - 0x1bd2  :    0 - 0x0
    "00000000", -- 7123 - 0x1bd3  :    0 - 0x0
    "00000000", -- 7124 - 0x1bd4  :    0 - 0x0
    "00000000", -- 7125 - 0x1bd5  :    0 - 0x0
    "00000000", -- 7126 - 0x1bd6  :    0 - 0x0
    "00000000", -- 7127 - 0x1bd7  :    0 - 0x0
    "00000000", -- 7128 - 0x1bd8  :    0 - 0x0
    "00000000", -- 7129 - 0x1bd9  :    0 - 0x0
    "00000000", -- 7130 - 0x1bda  :    0 - 0x0
    "00000000", -- 7131 - 0x1bdb  :    0 - 0x0
    "00000000", -- 7132 - 0x1bdc  :    0 - 0x0
    "00000000", -- 7133 - 0x1bdd  :    0 - 0x0
    "00000000", -- 7134 - 0x1bde  :    0 - 0x0
    "00000000", -- 7135 - 0x1bdf  :    0 - 0x0
    "00000000", -- 7136 - 0x1be0  :    0 - 0x0 -- Background 0xbe
    "00000000", -- 7137 - 0x1be1  :    0 - 0x0
    "00000000", -- 7138 - 0x1be2  :    0 - 0x0
    "00000000", -- 7139 - 0x1be3  :    0 - 0x0
    "00000000", -- 7140 - 0x1be4  :    0 - 0x0
    "00000000", -- 7141 - 0x1be5  :    0 - 0x0
    "00000000", -- 7142 - 0x1be6  :    0 - 0x0
    "00000000", -- 7143 - 0x1be7  :    0 - 0x0
    "00000000", -- 7144 - 0x1be8  :    0 - 0x0
    "00000000", -- 7145 - 0x1be9  :    0 - 0x0
    "00000000", -- 7146 - 0x1bea  :    0 - 0x0
    "00000000", -- 7147 - 0x1beb  :    0 - 0x0
    "00000000", -- 7148 - 0x1bec  :    0 - 0x0
    "00000000", -- 7149 - 0x1bed  :    0 - 0x0
    "00000000", -- 7150 - 0x1bee  :    0 - 0x0
    "00000000", -- 7151 - 0x1bef  :    0 - 0x0
    "00000000", -- 7152 - 0x1bf0  :    0 - 0x0 -- Background 0xbf
    "00000000", -- 7153 - 0x1bf1  :    0 - 0x0
    "00000000", -- 7154 - 0x1bf2  :    0 - 0x0
    "00000000", -- 7155 - 0x1bf3  :    0 - 0x0
    "00000000", -- 7156 - 0x1bf4  :    0 - 0x0
    "00000000", -- 7157 - 0x1bf5  :    0 - 0x0
    "00000000", -- 7158 - 0x1bf6  :    0 - 0x0
    "00000000", -- 7159 - 0x1bf7  :    0 - 0x0
    "00000000", -- 7160 - 0x1bf8  :    0 - 0x0
    "00000000", -- 7161 - 0x1bf9  :    0 - 0x0
    "00000000", -- 7162 - 0x1bfa  :    0 - 0x0
    "00000000", -- 7163 - 0x1bfb  :    0 - 0x0
    "00000000", -- 7164 - 0x1bfc  :    0 - 0x0
    "00000000", -- 7165 - 0x1bfd  :    0 - 0x0
    "00000000", -- 7166 - 0x1bfe  :    0 - 0x0
    "00000000", -- 7167 - 0x1bff  :    0 - 0x0
    "00000000", -- 7168 - 0x1c00  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 7169 - 0x1c01  :    0 - 0x0
    "00000000", -- 7170 - 0x1c02  :    0 - 0x0
    "00000000", -- 7171 - 0x1c03  :    0 - 0x0
    "00000000", -- 7172 - 0x1c04  :    0 - 0x0
    "00000000", -- 7173 - 0x1c05  :    0 - 0x0
    "00000000", -- 7174 - 0x1c06  :    0 - 0x0
    "00000000", -- 7175 - 0x1c07  :    0 - 0x0
    "00000000", -- 7176 - 0x1c08  :    0 - 0x0
    "00000000", -- 7177 - 0x1c09  :    0 - 0x0
    "00000000", -- 7178 - 0x1c0a  :    0 - 0x0
    "00000000", -- 7179 - 0x1c0b  :    0 - 0x0
    "00000000", -- 7180 - 0x1c0c  :    0 - 0x0
    "00000000", -- 7181 - 0x1c0d  :    0 - 0x0
    "00000000", -- 7182 - 0x1c0e  :    0 - 0x0
    "00000000", -- 7183 - 0x1c0f  :    0 - 0x0
    "00000000", -- 7184 - 0x1c10  :    0 - 0x0 -- Background 0xc1
    "00000000", -- 7185 - 0x1c11  :    0 - 0x0
    "00000000", -- 7186 - 0x1c12  :    0 - 0x0
    "00000000", -- 7187 - 0x1c13  :    0 - 0x0
    "00000000", -- 7188 - 0x1c14  :    0 - 0x0
    "00000000", -- 7189 - 0x1c15  :    0 - 0x0
    "00000000", -- 7190 - 0x1c16  :    0 - 0x0
    "00000000", -- 7191 - 0x1c17  :    0 - 0x0
    "00000000", -- 7192 - 0x1c18  :    0 - 0x0
    "00000000", -- 7193 - 0x1c19  :    0 - 0x0
    "00000000", -- 7194 - 0x1c1a  :    0 - 0x0
    "00000000", -- 7195 - 0x1c1b  :    0 - 0x0
    "00000000", -- 7196 - 0x1c1c  :    0 - 0x0
    "00000000", -- 7197 - 0x1c1d  :    0 - 0x0
    "00000000", -- 7198 - 0x1c1e  :    0 - 0x0
    "00000000", -- 7199 - 0x1c1f  :    0 - 0x0
    "00000000", -- 7200 - 0x1c20  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 7201 - 0x1c21  :    0 - 0x0
    "00000000", -- 7202 - 0x1c22  :    0 - 0x0
    "00000000", -- 7203 - 0x1c23  :    0 - 0x0
    "00000000", -- 7204 - 0x1c24  :    0 - 0x0
    "00000000", -- 7205 - 0x1c25  :    0 - 0x0
    "00000000", -- 7206 - 0x1c26  :    0 - 0x0
    "00000000", -- 7207 - 0x1c27  :    0 - 0x0
    "00000000", -- 7208 - 0x1c28  :    0 - 0x0
    "00000000", -- 7209 - 0x1c29  :    0 - 0x0
    "00000000", -- 7210 - 0x1c2a  :    0 - 0x0
    "00000000", -- 7211 - 0x1c2b  :    0 - 0x0
    "00000000", -- 7212 - 0x1c2c  :    0 - 0x0
    "00000000", -- 7213 - 0x1c2d  :    0 - 0x0
    "00000000", -- 7214 - 0x1c2e  :    0 - 0x0
    "00000000", -- 7215 - 0x1c2f  :    0 - 0x0
    "00000000", -- 7216 - 0x1c30  :    0 - 0x0 -- Background 0xc3
    "00000000", -- 7217 - 0x1c31  :    0 - 0x0
    "00000000", -- 7218 - 0x1c32  :    0 - 0x0
    "00000000", -- 7219 - 0x1c33  :    0 - 0x0
    "00000000", -- 7220 - 0x1c34  :    0 - 0x0
    "00000000", -- 7221 - 0x1c35  :    0 - 0x0
    "00000000", -- 7222 - 0x1c36  :    0 - 0x0
    "00000000", -- 7223 - 0x1c37  :    0 - 0x0
    "00000000", -- 7224 - 0x1c38  :    0 - 0x0
    "00000000", -- 7225 - 0x1c39  :    0 - 0x0
    "00000000", -- 7226 - 0x1c3a  :    0 - 0x0
    "00000000", -- 7227 - 0x1c3b  :    0 - 0x0
    "00000000", -- 7228 - 0x1c3c  :    0 - 0x0
    "00000000", -- 7229 - 0x1c3d  :    0 - 0x0
    "00000000", -- 7230 - 0x1c3e  :    0 - 0x0
    "00000000", -- 7231 - 0x1c3f  :    0 - 0x0
    "00000000", -- 7232 - 0x1c40  :    0 - 0x0 -- Background 0xc4
    "00000000", -- 7233 - 0x1c41  :    0 - 0x0
    "00000000", -- 7234 - 0x1c42  :    0 - 0x0
    "00000000", -- 7235 - 0x1c43  :    0 - 0x0
    "00000000", -- 7236 - 0x1c44  :    0 - 0x0
    "00000000", -- 7237 - 0x1c45  :    0 - 0x0
    "00000000", -- 7238 - 0x1c46  :    0 - 0x0
    "00000000", -- 7239 - 0x1c47  :    0 - 0x0
    "00000000", -- 7240 - 0x1c48  :    0 - 0x0
    "00000000", -- 7241 - 0x1c49  :    0 - 0x0
    "00000000", -- 7242 - 0x1c4a  :    0 - 0x0
    "00000000", -- 7243 - 0x1c4b  :    0 - 0x0
    "00000000", -- 7244 - 0x1c4c  :    0 - 0x0
    "00000000", -- 7245 - 0x1c4d  :    0 - 0x0
    "00000000", -- 7246 - 0x1c4e  :    0 - 0x0
    "00000000", -- 7247 - 0x1c4f  :    0 - 0x0
    "00000000", -- 7248 - 0x1c50  :    0 - 0x0 -- Background 0xc5
    "00000000", -- 7249 - 0x1c51  :    0 - 0x0
    "00000000", -- 7250 - 0x1c52  :    0 - 0x0
    "00000000", -- 7251 - 0x1c53  :    0 - 0x0
    "00000000", -- 7252 - 0x1c54  :    0 - 0x0
    "00000000", -- 7253 - 0x1c55  :    0 - 0x0
    "00000000", -- 7254 - 0x1c56  :    0 - 0x0
    "00000000", -- 7255 - 0x1c57  :    0 - 0x0
    "00000000", -- 7256 - 0x1c58  :    0 - 0x0
    "00000000", -- 7257 - 0x1c59  :    0 - 0x0
    "00000000", -- 7258 - 0x1c5a  :    0 - 0x0
    "00000000", -- 7259 - 0x1c5b  :    0 - 0x0
    "00000000", -- 7260 - 0x1c5c  :    0 - 0x0
    "00000000", -- 7261 - 0x1c5d  :    0 - 0x0
    "00000000", -- 7262 - 0x1c5e  :    0 - 0x0
    "00000000", -- 7263 - 0x1c5f  :    0 - 0x0
    "00000000", -- 7264 - 0x1c60  :    0 - 0x0 -- Background 0xc6
    "00000000", -- 7265 - 0x1c61  :    0 - 0x0
    "00000000", -- 7266 - 0x1c62  :    0 - 0x0
    "00000000", -- 7267 - 0x1c63  :    0 - 0x0
    "00000000", -- 7268 - 0x1c64  :    0 - 0x0
    "00000000", -- 7269 - 0x1c65  :    0 - 0x0
    "00000000", -- 7270 - 0x1c66  :    0 - 0x0
    "00000000", -- 7271 - 0x1c67  :    0 - 0x0
    "00000000", -- 7272 - 0x1c68  :    0 - 0x0
    "00000000", -- 7273 - 0x1c69  :    0 - 0x0
    "00000000", -- 7274 - 0x1c6a  :    0 - 0x0
    "00000000", -- 7275 - 0x1c6b  :    0 - 0x0
    "00000000", -- 7276 - 0x1c6c  :    0 - 0x0
    "00000000", -- 7277 - 0x1c6d  :    0 - 0x0
    "00000000", -- 7278 - 0x1c6e  :    0 - 0x0
    "00000000", -- 7279 - 0x1c6f  :    0 - 0x0
    "00000000", -- 7280 - 0x1c70  :    0 - 0x0 -- Background 0xc7
    "00000000", -- 7281 - 0x1c71  :    0 - 0x0
    "00000000", -- 7282 - 0x1c72  :    0 - 0x0
    "00000000", -- 7283 - 0x1c73  :    0 - 0x0
    "00000000", -- 7284 - 0x1c74  :    0 - 0x0
    "00000000", -- 7285 - 0x1c75  :    0 - 0x0
    "00000000", -- 7286 - 0x1c76  :    0 - 0x0
    "00000000", -- 7287 - 0x1c77  :    0 - 0x0
    "00000000", -- 7288 - 0x1c78  :    0 - 0x0
    "00000000", -- 7289 - 0x1c79  :    0 - 0x0
    "00000000", -- 7290 - 0x1c7a  :    0 - 0x0
    "00000000", -- 7291 - 0x1c7b  :    0 - 0x0
    "00000000", -- 7292 - 0x1c7c  :    0 - 0x0
    "00000000", -- 7293 - 0x1c7d  :    0 - 0x0
    "00000000", -- 7294 - 0x1c7e  :    0 - 0x0
    "00000000", -- 7295 - 0x1c7f  :    0 - 0x0
    "00000000", -- 7296 - 0x1c80  :    0 - 0x0 -- Background 0xc8
    "00000000", -- 7297 - 0x1c81  :    0 - 0x0
    "00000000", -- 7298 - 0x1c82  :    0 - 0x0
    "00000000", -- 7299 - 0x1c83  :    0 - 0x0
    "00000000", -- 7300 - 0x1c84  :    0 - 0x0
    "00000000", -- 7301 - 0x1c85  :    0 - 0x0
    "00000000", -- 7302 - 0x1c86  :    0 - 0x0
    "00000000", -- 7303 - 0x1c87  :    0 - 0x0
    "00000000", -- 7304 - 0x1c88  :    0 - 0x0
    "00000000", -- 7305 - 0x1c89  :    0 - 0x0
    "00000000", -- 7306 - 0x1c8a  :    0 - 0x0
    "00000000", -- 7307 - 0x1c8b  :    0 - 0x0
    "00000000", -- 7308 - 0x1c8c  :    0 - 0x0
    "00000000", -- 7309 - 0x1c8d  :    0 - 0x0
    "00000000", -- 7310 - 0x1c8e  :    0 - 0x0
    "00000000", -- 7311 - 0x1c8f  :    0 - 0x0
    "00000000", -- 7312 - 0x1c90  :    0 - 0x0 -- Background 0xc9
    "00000000", -- 7313 - 0x1c91  :    0 - 0x0
    "00000000", -- 7314 - 0x1c92  :    0 - 0x0
    "00000000", -- 7315 - 0x1c93  :    0 - 0x0
    "00000000", -- 7316 - 0x1c94  :    0 - 0x0
    "00000000", -- 7317 - 0x1c95  :    0 - 0x0
    "00000000", -- 7318 - 0x1c96  :    0 - 0x0
    "00000000", -- 7319 - 0x1c97  :    0 - 0x0
    "00000000", -- 7320 - 0x1c98  :    0 - 0x0
    "00000000", -- 7321 - 0x1c99  :    0 - 0x0
    "00000000", -- 7322 - 0x1c9a  :    0 - 0x0
    "00000000", -- 7323 - 0x1c9b  :    0 - 0x0
    "00000000", -- 7324 - 0x1c9c  :    0 - 0x0
    "00000000", -- 7325 - 0x1c9d  :    0 - 0x0
    "00000000", -- 7326 - 0x1c9e  :    0 - 0x0
    "00000000", -- 7327 - 0x1c9f  :    0 - 0x0
    "00000000", -- 7328 - 0x1ca0  :    0 - 0x0 -- Background 0xca
    "00000000", -- 7329 - 0x1ca1  :    0 - 0x0
    "00000000", -- 7330 - 0x1ca2  :    0 - 0x0
    "00000000", -- 7331 - 0x1ca3  :    0 - 0x0
    "00000000", -- 7332 - 0x1ca4  :    0 - 0x0
    "00000000", -- 7333 - 0x1ca5  :    0 - 0x0
    "00000000", -- 7334 - 0x1ca6  :    0 - 0x0
    "00000000", -- 7335 - 0x1ca7  :    0 - 0x0
    "00000000", -- 7336 - 0x1ca8  :    0 - 0x0
    "00000000", -- 7337 - 0x1ca9  :    0 - 0x0
    "00000000", -- 7338 - 0x1caa  :    0 - 0x0
    "00000000", -- 7339 - 0x1cab  :    0 - 0x0
    "00000000", -- 7340 - 0x1cac  :    0 - 0x0
    "00000000", -- 7341 - 0x1cad  :    0 - 0x0
    "00000000", -- 7342 - 0x1cae  :    0 - 0x0
    "00000000", -- 7343 - 0x1caf  :    0 - 0x0
    "00000000", -- 7344 - 0x1cb0  :    0 - 0x0 -- Background 0xcb
    "00000000", -- 7345 - 0x1cb1  :    0 - 0x0
    "00000000", -- 7346 - 0x1cb2  :    0 - 0x0
    "00000000", -- 7347 - 0x1cb3  :    0 - 0x0
    "00000000", -- 7348 - 0x1cb4  :    0 - 0x0
    "00000000", -- 7349 - 0x1cb5  :    0 - 0x0
    "00000000", -- 7350 - 0x1cb6  :    0 - 0x0
    "00000000", -- 7351 - 0x1cb7  :    0 - 0x0
    "00000000", -- 7352 - 0x1cb8  :    0 - 0x0
    "00000000", -- 7353 - 0x1cb9  :    0 - 0x0
    "00000000", -- 7354 - 0x1cba  :    0 - 0x0
    "00000000", -- 7355 - 0x1cbb  :    0 - 0x0
    "00000000", -- 7356 - 0x1cbc  :    0 - 0x0
    "00000000", -- 7357 - 0x1cbd  :    0 - 0x0
    "00000000", -- 7358 - 0x1cbe  :    0 - 0x0
    "00000000", -- 7359 - 0x1cbf  :    0 - 0x0
    "00000000", -- 7360 - 0x1cc0  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 7361 - 0x1cc1  :    0 - 0x0
    "00000000", -- 7362 - 0x1cc2  :    0 - 0x0
    "00000000", -- 7363 - 0x1cc3  :    0 - 0x0
    "00000000", -- 7364 - 0x1cc4  :    0 - 0x0
    "00000000", -- 7365 - 0x1cc5  :    0 - 0x0
    "00000000", -- 7366 - 0x1cc6  :    0 - 0x0
    "00000000", -- 7367 - 0x1cc7  :    0 - 0x0
    "00000000", -- 7368 - 0x1cc8  :    0 - 0x0
    "00000000", -- 7369 - 0x1cc9  :    0 - 0x0
    "00000000", -- 7370 - 0x1cca  :    0 - 0x0
    "00000000", -- 7371 - 0x1ccb  :    0 - 0x0
    "00000000", -- 7372 - 0x1ccc  :    0 - 0x0
    "00000000", -- 7373 - 0x1ccd  :    0 - 0x0
    "00000000", -- 7374 - 0x1cce  :    0 - 0x0
    "00000000", -- 7375 - 0x1ccf  :    0 - 0x0
    "00111111", -- 7376 - 0x1cd0  :   63 - 0x3f -- Background 0xcd
    "01111111", -- 7377 - 0x1cd1  :  127 - 0x7f
    "11111111", -- 7378 - 0x1cd2  :  255 - 0xff
    "11110000", -- 7379 - 0x1cd3  :  240 - 0xf0
    "11100000", -- 7380 - 0x1cd4  :  224 - 0xe0
    "11100011", -- 7381 - 0x1cd5  :  227 - 0xe3
    "11100111", -- 7382 - 0x1cd6  :  231 - 0xe7
    "11100111", -- 7383 - 0x1cd7  :  231 - 0xe7
    "11000000", -- 7384 - 0x1cd8  :  192 - 0xc0
    "10000000", -- 7385 - 0x1cd9  :  128 - 0x80
    "00000000", -- 7386 - 0x1cda  :    0 - 0x0
    "00001111", -- 7387 - 0x1cdb  :   15 - 0xf
    "00011111", -- 7388 - 0x1cdc  :   31 - 0x1f
    "00011100", -- 7389 - 0x1cdd  :   28 - 0x1c
    "00011000", -- 7390 - 0x1cde  :   24 - 0x18
    "00011000", -- 7391 - 0x1cdf  :   24 - 0x18
    "11111100", -- 7392 - 0x1ce0  :  252 - 0xfc -- Background 0xce
    "11111110", -- 7393 - 0x1ce1  :  254 - 0xfe
    "11111111", -- 7394 - 0x1ce2  :  255 - 0xff
    "00001111", -- 7395 - 0x1ce3  :   15 - 0xf
    "00000111", -- 7396 - 0x1ce4  :    7 - 0x7
    "11000111", -- 7397 - 0x1ce5  :  199 - 0xc7
    "11100111", -- 7398 - 0x1ce6  :  231 - 0xe7
    "11100111", -- 7399 - 0x1ce7  :  231 - 0xe7
    "00000011", -- 7400 - 0x1ce8  :    3 - 0x3
    "00000001", -- 7401 - 0x1ce9  :    1 - 0x1
    "00000000", -- 7402 - 0x1cea  :    0 - 0x0
    "11110000", -- 7403 - 0x1ceb  :  240 - 0xf0
    "11111000", -- 7404 - 0x1cec  :  248 - 0xf8
    "00111000", -- 7405 - 0x1ced  :   56 - 0x38
    "00011000", -- 7406 - 0x1cee  :   24 - 0x18
    "00011000", -- 7407 - 0x1cef  :   24 - 0x18
    "00000000", -- 7408 - 0x1cf0  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 7409 - 0x1cf1  :    0 - 0x0
    "00000000", -- 7410 - 0x1cf2  :    0 - 0x0
    "00000000", -- 7411 - 0x1cf3  :    0 - 0x0
    "00000000", -- 7412 - 0x1cf4  :    0 - 0x0
    "00000000", -- 7413 - 0x1cf5  :    0 - 0x0
    "00000000", -- 7414 - 0x1cf6  :    0 - 0x0
    "00000000", -- 7415 - 0x1cf7  :    0 - 0x0
    "00000000", -- 7416 - 0x1cf8  :    0 - 0x0
    "00000000", -- 7417 - 0x1cf9  :    0 - 0x0
    "00000000", -- 7418 - 0x1cfa  :    0 - 0x0
    "00000000", -- 7419 - 0x1cfb  :    0 - 0x0
    "00000000", -- 7420 - 0x1cfc  :    0 - 0x0
    "00000000", -- 7421 - 0x1cfd  :    0 - 0x0
    "00000000", -- 7422 - 0x1cfe  :    0 - 0x0
    "00000000", -- 7423 - 0x1cff  :    0 - 0x0
    "00000000", -- 7424 - 0x1d00  :    0 - 0x0 -- Background 0xd0
    "00000000", -- 7425 - 0x1d01  :    0 - 0x0
    "00000000", -- 7426 - 0x1d02  :    0 - 0x0
    "00000000", -- 7427 - 0x1d03  :    0 - 0x0
    "00000000", -- 7428 - 0x1d04  :    0 - 0x0
    "00000000", -- 7429 - 0x1d05  :    0 - 0x0
    "00000000", -- 7430 - 0x1d06  :    0 - 0x0
    "00000000", -- 7431 - 0x1d07  :    0 - 0x0
    "00000000", -- 7432 - 0x1d08  :    0 - 0x0
    "00000000", -- 7433 - 0x1d09  :    0 - 0x0
    "00000000", -- 7434 - 0x1d0a  :    0 - 0x0
    "00000000", -- 7435 - 0x1d0b  :    0 - 0x0
    "00000000", -- 7436 - 0x1d0c  :    0 - 0x0
    "00000000", -- 7437 - 0x1d0d  :    0 - 0x0
    "00000000", -- 7438 - 0x1d0e  :    0 - 0x0
    "00000000", -- 7439 - 0x1d0f  :    0 - 0x0
    "00000000", -- 7440 - 0x1d10  :    0 - 0x0 -- Background 0xd1
    "00000000", -- 7441 - 0x1d11  :    0 - 0x0
    "00000000", -- 7442 - 0x1d12  :    0 - 0x0
    "00000000", -- 7443 - 0x1d13  :    0 - 0x0
    "00000000", -- 7444 - 0x1d14  :    0 - 0x0
    "00000000", -- 7445 - 0x1d15  :    0 - 0x0
    "00000000", -- 7446 - 0x1d16  :    0 - 0x0
    "00000000", -- 7447 - 0x1d17  :    0 - 0x0
    "00000000", -- 7448 - 0x1d18  :    0 - 0x0
    "00000000", -- 7449 - 0x1d19  :    0 - 0x0
    "00000000", -- 7450 - 0x1d1a  :    0 - 0x0
    "00000000", -- 7451 - 0x1d1b  :    0 - 0x0
    "00000000", -- 7452 - 0x1d1c  :    0 - 0x0
    "00000000", -- 7453 - 0x1d1d  :    0 - 0x0
    "00000000", -- 7454 - 0x1d1e  :    0 - 0x0
    "00000000", -- 7455 - 0x1d1f  :    0 - 0x0
    "00000000", -- 7456 - 0x1d20  :    0 - 0x0 -- Background 0xd2
    "00000000", -- 7457 - 0x1d21  :    0 - 0x0
    "00000000", -- 7458 - 0x1d22  :    0 - 0x0
    "00000000", -- 7459 - 0x1d23  :    0 - 0x0
    "00000000", -- 7460 - 0x1d24  :    0 - 0x0
    "00000000", -- 7461 - 0x1d25  :    0 - 0x0
    "00000000", -- 7462 - 0x1d26  :    0 - 0x0
    "00000000", -- 7463 - 0x1d27  :    0 - 0x0
    "00000000", -- 7464 - 0x1d28  :    0 - 0x0
    "00000000", -- 7465 - 0x1d29  :    0 - 0x0
    "00000000", -- 7466 - 0x1d2a  :    0 - 0x0
    "00000000", -- 7467 - 0x1d2b  :    0 - 0x0
    "00000000", -- 7468 - 0x1d2c  :    0 - 0x0
    "00000000", -- 7469 - 0x1d2d  :    0 - 0x0
    "00000000", -- 7470 - 0x1d2e  :    0 - 0x0
    "00000000", -- 7471 - 0x1d2f  :    0 - 0x0
    "00000000", -- 7472 - 0x1d30  :    0 - 0x0 -- Background 0xd3
    "00000000", -- 7473 - 0x1d31  :    0 - 0x0
    "00000000", -- 7474 - 0x1d32  :    0 - 0x0
    "00000000", -- 7475 - 0x1d33  :    0 - 0x0
    "00000000", -- 7476 - 0x1d34  :    0 - 0x0
    "00000000", -- 7477 - 0x1d35  :    0 - 0x0
    "00000000", -- 7478 - 0x1d36  :    0 - 0x0
    "00000000", -- 7479 - 0x1d37  :    0 - 0x0
    "00000000", -- 7480 - 0x1d38  :    0 - 0x0
    "00000000", -- 7481 - 0x1d39  :    0 - 0x0
    "00000000", -- 7482 - 0x1d3a  :    0 - 0x0
    "00000000", -- 7483 - 0x1d3b  :    0 - 0x0
    "00000000", -- 7484 - 0x1d3c  :    0 - 0x0
    "00000000", -- 7485 - 0x1d3d  :    0 - 0x0
    "00000000", -- 7486 - 0x1d3e  :    0 - 0x0
    "00000000", -- 7487 - 0x1d3f  :    0 - 0x0
    "00000000", -- 7488 - 0x1d40  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 7489 - 0x1d41  :    0 - 0x0
    "00000000", -- 7490 - 0x1d42  :    0 - 0x0
    "00000000", -- 7491 - 0x1d43  :    0 - 0x0
    "00000000", -- 7492 - 0x1d44  :    0 - 0x0
    "00000000", -- 7493 - 0x1d45  :    0 - 0x0
    "00000000", -- 7494 - 0x1d46  :    0 - 0x0
    "00000000", -- 7495 - 0x1d47  :    0 - 0x0
    "00000000", -- 7496 - 0x1d48  :    0 - 0x0
    "00000000", -- 7497 - 0x1d49  :    0 - 0x0
    "00000000", -- 7498 - 0x1d4a  :    0 - 0x0
    "00000000", -- 7499 - 0x1d4b  :    0 - 0x0
    "00000000", -- 7500 - 0x1d4c  :    0 - 0x0
    "00000000", -- 7501 - 0x1d4d  :    0 - 0x0
    "00000000", -- 7502 - 0x1d4e  :    0 - 0x0
    "00000000", -- 7503 - 0x1d4f  :    0 - 0x0
    "00000000", -- 7504 - 0x1d50  :    0 - 0x0 -- Background 0xd5
    "00000000", -- 7505 - 0x1d51  :    0 - 0x0
    "00000000", -- 7506 - 0x1d52  :    0 - 0x0
    "00000000", -- 7507 - 0x1d53  :    0 - 0x0
    "00000000", -- 7508 - 0x1d54  :    0 - 0x0
    "00000000", -- 7509 - 0x1d55  :    0 - 0x0
    "00000000", -- 7510 - 0x1d56  :    0 - 0x0
    "00000000", -- 7511 - 0x1d57  :    0 - 0x0
    "00000000", -- 7512 - 0x1d58  :    0 - 0x0
    "00000000", -- 7513 - 0x1d59  :    0 - 0x0
    "00000000", -- 7514 - 0x1d5a  :    0 - 0x0
    "00000000", -- 7515 - 0x1d5b  :    0 - 0x0
    "00000000", -- 7516 - 0x1d5c  :    0 - 0x0
    "00000000", -- 7517 - 0x1d5d  :    0 - 0x0
    "00000000", -- 7518 - 0x1d5e  :    0 - 0x0
    "00000000", -- 7519 - 0x1d5f  :    0 - 0x0
    "00000000", -- 7520 - 0x1d60  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 7521 - 0x1d61  :    0 - 0x0
    "00000000", -- 7522 - 0x1d62  :    0 - 0x0
    "00000000", -- 7523 - 0x1d63  :    0 - 0x0
    "00000000", -- 7524 - 0x1d64  :    0 - 0x0
    "00000000", -- 7525 - 0x1d65  :    0 - 0x0
    "00000000", -- 7526 - 0x1d66  :    0 - 0x0
    "00000000", -- 7527 - 0x1d67  :    0 - 0x0
    "00000000", -- 7528 - 0x1d68  :    0 - 0x0
    "00000000", -- 7529 - 0x1d69  :    0 - 0x0
    "00000000", -- 7530 - 0x1d6a  :    0 - 0x0
    "00000000", -- 7531 - 0x1d6b  :    0 - 0x0
    "00000000", -- 7532 - 0x1d6c  :    0 - 0x0
    "00000000", -- 7533 - 0x1d6d  :    0 - 0x0
    "00000000", -- 7534 - 0x1d6e  :    0 - 0x0
    "00000000", -- 7535 - 0x1d6f  :    0 - 0x0
    "00000000", -- 7536 - 0x1d70  :    0 - 0x0 -- Background 0xd7
    "00000000", -- 7537 - 0x1d71  :    0 - 0x0
    "00000000", -- 7538 - 0x1d72  :    0 - 0x0
    "00000000", -- 7539 - 0x1d73  :    0 - 0x0
    "00000000", -- 7540 - 0x1d74  :    0 - 0x0
    "00000000", -- 7541 - 0x1d75  :    0 - 0x0
    "00000000", -- 7542 - 0x1d76  :    0 - 0x0
    "00000000", -- 7543 - 0x1d77  :    0 - 0x0
    "00000000", -- 7544 - 0x1d78  :    0 - 0x0
    "00000000", -- 7545 - 0x1d79  :    0 - 0x0
    "00000000", -- 7546 - 0x1d7a  :    0 - 0x0
    "00000000", -- 7547 - 0x1d7b  :    0 - 0x0
    "00000000", -- 7548 - 0x1d7c  :    0 - 0x0
    "00000000", -- 7549 - 0x1d7d  :    0 - 0x0
    "00000000", -- 7550 - 0x1d7e  :    0 - 0x0
    "00000000", -- 7551 - 0x1d7f  :    0 - 0x0
    "00000000", -- 7552 - 0x1d80  :    0 - 0x0 -- Background 0xd8
    "00000000", -- 7553 - 0x1d81  :    0 - 0x0
    "00000000", -- 7554 - 0x1d82  :    0 - 0x0
    "00000000", -- 7555 - 0x1d83  :    0 - 0x0
    "00000000", -- 7556 - 0x1d84  :    0 - 0x0
    "00000000", -- 7557 - 0x1d85  :    0 - 0x0
    "00000000", -- 7558 - 0x1d86  :    0 - 0x0
    "00000000", -- 7559 - 0x1d87  :    0 - 0x0
    "00000000", -- 7560 - 0x1d88  :    0 - 0x0
    "00000000", -- 7561 - 0x1d89  :    0 - 0x0
    "00000000", -- 7562 - 0x1d8a  :    0 - 0x0
    "00000000", -- 7563 - 0x1d8b  :    0 - 0x0
    "00000000", -- 7564 - 0x1d8c  :    0 - 0x0
    "00000000", -- 7565 - 0x1d8d  :    0 - 0x0
    "00000000", -- 7566 - 0x1d8e  :    0 - 0x0
    "00000000", -- 7567 - 0x1d8f  :    0 - 0x0
    "00000000", -- 7568 - 0x1d90  :    0 - 0x0 -- Background 0xd9
    "00000000", -- 7569 - 0x1d91  :    0 - 0x0
    "00000000", -- 7570 - 0x1d92  :    0 - 0x0
    "00000000", -- 7571 - 0x1d93  :    0 - 0x0
    "00000000", -- 7572 - 0x1d94  :    0 - 0x0
    "00000000", -- 7573 - 0x1d95  :    0 - 0x0
    "00000000", -- 7574 - 0x1d96  :    0 - 0x0
    "00000000", -- 7575 - 0x1d97  :    0 - 0x0
    "00000000", -- 7576 - 0x1d98  :    0 - 0x0
    "00000000", -- 7577 - 0x1d99  :    0 - 0x0
    "00000000", -- 7578 - 0x1d9a  :    0 - 0x0
    "00000000", -- 7579 - 0x1d9b  :    0 - 0x0
    "00000000", -- 7580 - 0x1d9c  :    0 - 0x0
    "00000000", -- 7581 - 0x1d9d  :    0 - 0x0
    "00000000", -- 7582 - 0x1d9e  :    0 - 0x0
    "00000000", -- 7583 - 0x1d9f  :    0 - 0x0
    "00000000", -- 7584 - 0x1da0  :    0 - 0x0 -- Background 0xda
    "00000000", -- 7585 - 0x1da1  :    0 - 0x0
    "00000000", -- 7586 - 0x1da2  :    0 - 0x0
    "00000000", -- 7587 - 0x1da3  :    0 - 0x0
    "00000000", -- 7588 - 0x1da4  :    0 - 0x0
    "00000000", -- 7589 - 0x1da5  :    0 - 0x0
    "00000000", -- 7590 - 0x1da6  :    0 - 0x0
    "00000000", -- 7591 - 0x1da7  :    0 - 0x0
    "00000000", -- 7592 - 0x1da8  :    0 - 0x0
    "00000000", -- 7593 - 0x1da9  :    0 - 0x0
    "00000000", -- 7594 - 0x1daa  :    0 - 0x0
    "00000000", -- 7595 - 0x1dab  :    0 - 0x0
    "00000000", -- 7596 - 0x1dac  :    0 - 0x0
    "00000000", -- 7597 - 0x1dad  :    0 - 0x0
    "00000000", -- 7598 - 0x1dae  :    0 - 0x0
    "00000000", -- 7599 - 0x1daf  :    0 - 0x0
    "00000000", -- 7600 - 0x1db0  :    0 - 0x0 -- Background 0xdb
    "00000000", -- 7601 - 0x1db1  :    0 - 0x0
    "00000000", -- 7602 - 0x1db2  :    0 - 0x0
    "00000000", -- 7603 - 0x1db3  :    0 - 0x0
    "00000000", -- 7604 - 0x1db4  :    0 - 0x0
    "00000000", -- 7605 - 0x1db5  :    0 - 0x0
    "00000000", -- 7606 - 0x1db6  :    0 - 0x0
    "00000000", -- 7607 - 0x1db7  :    0 - 0x0
    "00000000", -- 7608 - 0x1db8  :    0 - 0x0
    "00000000", -- 7609 - 0x1db9  :    0 - 0x0
    "00000000", -- 7610 - 0x1dba  :    0 - 0x0
    "00000000", -- 7611 - 0x1dbb  :    0 - 0x0
    "00000000", -- 7612 - 0x1dbc  :    0 - 0x0
    "00000000", -- 7613 - 0x1dbd  :    0 - 0x0
    "00000000", -- 7614 - 0x1dbe  :    0 - 0x0
    "00000000", -- 7615 - 0x1dbf  :    0 - 0x0
    "00000000", -- 7616 - 0x1dc0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 7617 - 0x1dc1  :    0 - 0x0
    "00000000", -- 7618 - 0x1dc2  :    0 - 0x0
    "00000000", -- 7619 - 0x1dc3  :    0 - 0x0
    "00000000", -- 7620 - 0x1dc4  :    0 - 0x0
    "00000000", -- 7621 - 0x1dc5  :    0 - 0x0
    "00000000", -- 7622 - 0x1dc6  :    0 - 0x0
    "00000000", -- 7623 - 0x1dc7  :    0 - 0x0
    "00000000", -- 7624 - 0x1dc8  :    0 - 0x0
    "00000000", -- 7625 - 0x1dc9  :    0 - 0x0
    "00000000", -- 7626 - 0x1dca  :    0 - 0x0
    "00000000", -- 7627 - 0x1dcb  :    0 - 0x0
    "00000000", -- 7628 - 0x1dcc  :    0 - 0x0
    "00000000", -- 7629 - 0x1dcd  :    0 - 0x0
    "00000000", -- 7630 - 0x1dce  :    0 - 0x0
    "00000000", -- 7631 - 0x1dcf  :    0 - 0x0
    "11100111", -- 7632 - 0x1dd0  :  231 - 0xe7 -- Background 0xdd
    "11100111", -- 7633 - 0x1dd1  :  231 - 0xe7
    "11100011", -- 7634 - 0x1dd2  :  227 - 0xe3
    "11100000", -- 7635 - 0x1dd3  :  224 - 0xe0
    "11110000", -- 7636 - 0x1dd4  :  240 - 0xf0
    "11111111", -- 7637 - 0x1dd5  :  255 - 0xff
    "01111111", -- 7638 - 0x1dd6  :  127 - 0x7f
    "00111111", -- 7639 - 0x1dd7  :   63 - 0x3f
    "00011000", -- 7640 - 0x1dd8  :   24 - 0x18
    "00011000", -- 7641 - 0x1dd9  :   24 - 0x18
    "00011100", -- 7642 - 0x1dda  :   28 - 0x1c
    "00011111", -- 7643 - 0x1ddb  :   31 - 0x1f
    "00001111", -- 7644 - 0x1ddc  :   15 - 0xf
    "00000000", -- 7645 - 0x1ddd  :    0 - 0x0
    "10000000", -- 7646 - 0x1dde  :  128 - 0x80
    "11000000", -- 7647 - 0x1ddf  :  192 - 0xc0
    "11100111", -- 7648 - 0x1de0  :  231 - 0xe7 -- Background 0xde
    "11100111", -- 7649 - 0x1de1  :  231 - 0xe7
    "11000111", -- 7650 - 0x1de2  :  199 - 0xc7
    "00000111", -- 7651 - 0x1de3  :    7 - 0x7
    "00001111", -- 7652 - 0x1de4  :   15 - 0xf
    "11111111", -- 7653 - 0x1de5  :  255 - 0xff
    "11111110", -- 7654 - 0x1de6  :  254 - 0xfe
    "11111100", -- 7655 - 0x1de7  :  252 - 0xfc
    "00011000", -- 7656 - 0x1de8  :   24 - 0x18
    "00011000", -- 7657 - 0x1de9  :   24 - 0x18
    "00111000", -- 7658 - 0x1dea  :   56 - 0x38
    "11111000", -- 7659 - 0x1deb  :  248 - 0xf8
    "11110000", -- 7660 - 0x1dec  :  240 - 0xf0
    "00000000", -- 7661 - 0x1ded  :    0 - 0x0
    "00000001", -- 7662 - 0x1dee  :    1 - 0x1
    "00000011", -- 7663 - 0x1def  :    3 - 0x3
    "00000000", -- 7664 - 0x1df0  :    0 - 0x0 -- Background 0xdf
    "00000000", -- 7665 - 0x1df1  :    0 - 0x0
    "00000000", -- 7666 - 0x1df2  :    0 - 0x0
    "00000000", -- 7667 - 0x1df3  :    0 - 0x0
    "00000000", -- 7668 - 0x1df4  :    0 - 0x0
    "00000000", -- 7669 - 0x1df5  :    0 - 0x0
    "00000000", -- 7670 - 0x1df6  :    0 - 0x0
    "00000000", -- 7671 - 0x1df7  :    0 - 0x0
    "00000000", -- 7672 - 0x1df8  :    0 - 0x0
    "00000000", -- 7673 - 0x1df9  :    0 - 0x0
    "00000000", -- 7674 - 0x1dfa  :    0 - 0x0
    "00000000", -- 7675 - 0x1dfb  :    0 - 0x0
    "00000000", -- 7676 - 0x1dfc  :    0 - 0x0
    "00000000", -- 7677 - 0x1dfd  :    0 - 0x0
    "00000000", -- 7678 - 0x1dfe  :    0 - 0x0
    "00000000", -- 7679 - 0x1dff  :    0 - 0x0
    "00000000", -- 7680 - 0x1e00  :    0 - 0x0 -- Background 0xe0
    "00000000", -- 7681 - 0x1e01  :    0 - 0x0
    "00000000", -- 7682 - 0x1e02  :    0 - 0x0
    "00000000", -- 7683 - 0x1e03  :    0 - 0x0
    "00000000", -- 7684 - 0x1e04  :    0 - 0x0
    "00000000", -- 7685 - 0x1e05  :    0 - 0x0
    "00000000", -- 7686 - 0x1e06  :    0 - 0x0
    "00000000", -- 7687 - 0x1e07  :    0 - 0x0
    "00000000", -- 7688 - 0x1e08  :    0 - 0x0
    "00000000", -- 7689 - 0x1e09  :    0 - 0x0
    "00000000", -- 7690 - 0x1e0a  :    0 - 0x0
    "00000000", -- 7691 - 0x1e0b  :    0 - 0x0
    "00000000", -- 7692 - 0x1e0c  :    0 - 0x0
    "00000000", -- 7693 - 0x1e0d  :    0 - 0x0
    "00000000", -- 7694 - 0x1e0e  :    0 - 0x0
    "00000000", -- 7695 - 0x1e0f  :    0 - 0x0
    "00000000", -- 7696 - 0x1e10  :    0 - 0x0 -- Background 0xe1
    "00000000", -- 7697 - 0x1e11  :    0 - 0x0
    "00000000", -- 7698 - 0x1e12  :    0 - 0x0
    "00000000", -- 7699 - 0x1e13  :    0 - 0x0
    "00000000", -- 7700 - 0x1e14  :    0 - 0x0
    "00000000", -- 7701 - 0x1e15  :    0 - 0x0
    "00000000", -- 7702 - 0x1e16  :    0 - 0x0
    "00000000", -- 7703 - 0x1e17  :    0 - 0x0
    "00000000", -- 7704 - 0x1e18  :    0 - 0x0
    "00000000", -- 7705 - 0x1e19  :    0 - 0x0
    "00000000", -- 7706 - 0x1e1a  :    0 - 0x0
    "00000000", -- 7707 - 0x1e1b  :    0 - 0x0
    "00000000", -- 7708 - 0x1e1c  :    0 - 0x0
    "00000000", -- 7709 - 0x1e1d  :    0 - 0x0
    "00000000", -- 7710 - 0x1e1e  :    0 - 0x0
    "00000000", -- 7711 - 0x1e1f  :    0 - 0x0
    "00000000", -- 7712 - 0x1e20  :    0 - 0x0 -- Background 0xe2
    "00000000", -- 7713 - 0x1e21  :    0 - 0x0
    "00000000", -- 7714 - 0x1e22  :    0 - 0x0
    "00000000", -- 7715 - 0x1e23  :    0 - 0x0
    "00000000", -- 7716 - 0x1e24  :    0 - 0x0
    "00000000", -- 7717 - 0x1e25  :    0 - 0x0
    "00000000", -- 7718 - 0x1e26  :    0 - 0x0
    "00000000", -- 7719 - 0x1e27  :    0 - 0x0
    "00000000", -- 7720 - 0x1e28  :    0 - 0x0
    "00000000", -- 7721 - 0x1e29  :    0 - 0x0
    "00000000", -- 7722 - 0x1e2a  :    0 - 0x0
    "00000000", -- 7723 - 0x1e2b  :    0 - 0x0
    "00000000", -- 7724 - 0x1e2c  :    0 - 0x0
    "00000000", -- 7725 - 0x1e2d  :    0 - 0x0
    "00000000", -- 7726 - 0x1e2e  :    0 - 0x0
    "00000000", -- 7727 - 0x1e2f  :    0 - 0x0
    "00000000", -- 7728 - 0x1e30  :    0 - 0x0 -- Background 0xe3
    "00000000", -- 7729 - 0x1e31  :    0 - 0x0
    "00000000", -- 7730 - 0x1e32  :    0 - 0x0
    "00000000", -- 7731 - 0x1e33  :    0 - 0x0
    "00000000", -- 7732 - 0x1e34  :    0 - 0x0
    "00000000", -- 7733 - 0x1e35  :    0 - 0x0
    "00000000", -- 7734 - 0x1e36  :    0 - 0x0
    "00000000", -- 7735 - 0x1e37  :    0 - 0x0
    "00000000", -- 7736 - 0x1e38  :    0 - 0x0
    "00000000", -- 7737 - 0x1e39  :    0 - 0x0
    "00000000", -- 7738 - 0x1e3a  :    0 - 0x0
    "00000000", -- 7739 - 0x1e3b  :    0 - 0x0
    "00000000", -- 7740 - 0x1e3c  :    0 - 0x0
    "00000000", -- 7741 - 0x1e3d  :    0 - 0x0
    "00000000", -- 7742 - 0x1e3e  :    0 - 0x0
    "00000000", -- 7743 - 0x1e3f  :    0 - 0x0
    "00000000", -- 7744 - 0x1e40  :    0 - 0x0 -- Background 0xe4
    "00000000", -- 7745 - 0x1e41  :    0 - 0x0
    "00000000", -- 7746 - 0x1e42  :    0 - 0x0
    "00000000", -- 7747 - 0x1e43  :    0 - 0x0
    "00000000", -- 7748 - 0x1e44  :    0 - 0x0
    "00000000", -- 7749 - 0x1e45  :    0 - 0x0
    "00000000", -- 7750 - 0x1e46  :    0 - 0x0
    "00000000", -- 7751 - 0x1e47  :    0 - 0x0
    "00000000", -- 7752 - 0x1e48  :    0 - 0x0
    "00000000", -- 7753 - 0x1e49  :    0 - 0x0
    "00000000", -- 7754 - 0x1e4a  :    0 - 0x0
    "00000000", -- 7755 - 0x1e4b  :    0 - 0x0
    "00000000", -- 7756 - 0x1e4c  :    0 - 0x0
    "00000000", -- 7757 - 0x1e4d  :    0 - 0x0
    "00000000", -- 7758 - 0x1e4e  :    0 - 0x0
    "00000000", -- 7759 - 0x1e4f  :    0 - 0x0
    "01111111", -- 7760 - 0x1e50  :  127 - 0x7f -- Background 0xe5
    "11111111", -- 7761 - 0x1e51  :  255 - 0xff
    "11111111", -- 7762 - 0x1e52  :  255 - 0xff
    "11100000", -- 7763 - 0x1e53  :  224 - 0xe0
    "11100000", -- 7764 - 0x1e54  :  224 - 0xe0
    "11100000", -- 7765 - 0x1e55  :  224 - 0xe0
    "11100000", -- 7766 - 0x1e56  :  224 - 0xe0
    "11100001", -- 7767 - 0x1e57  :  225 - 0xe1
    "00000000", -- 7768 - 0x1e58  :    0 - 0x0
    "00000000", -- 7769 - 0x1e59  :    0 - 0x0
    "00000000", -- 7770 - 0x1e5a  :    0 - 0x0
    "00000000", -- 7771 - 0x1e5b  :    0 - 0x0
    "00000000", -- 7772 - 0x1e5c  :    0 - 0x0
    "00000000", -- 7773 - 0x1e5d  :    0 - 0x0
    "00000000", -- 7774 - 0x1e5e  :    0 - 0x0
    "00000000", -- 7775 - 0x1e5f  :    0 - 0x0
    "11111110", -- 7776 - 0x1e60  :  254 - 0xfe -- Background 0xe6
    "11111111", -- 7777 - 0x1e61  :  255 - 0xff
    "11111111", -- 7778 - 0x1e62  :  255 - 0xff
    "00000111", -- 7779 - 0x1e63  :    7 - 0x7
    "00000111", -- 7780 - 0x1e64  :    7 - 0x7
    "00000111", -- 7781 - 0x1e65  :    7 - 0x7
    "00000111", -- 7782 - 0x1e66  :    7 - 0x7
    "10000111", -- 7783 - 0x1e67  :  135 - 0x87
    "00000000", -- 7784 - 0x1e68  :    0 - 0x0
    "00000000", -- 7785 - 0x1e69  :    0 - 0x0
    "00000000", -- 7786 - 0x1e6a  :    0 - 0x0
    "00000000", -- 7787 - 0x1e6b  :    0 - 0x0
    "00000000", -- 7788 - 0x1e6c  :    0 - 0x0
    "00000000", -- 7789 - 0x1e6d  :    0 - 0x0
    "00000000", -- 7790 - 0x1e6e  :    0 - 0x0
    "00000000", -- 7791 - 0x1e6f  :    0 - 0x0
    "00011111", -- 7792 - 0x1e70  :   31 - 0x1f -- Background 0xe7
    "00100000", -- 7793 - 0x1e71  :   32 - 0x20
    "01000000", -- 7794 - 0x1e72  :   64 - 0x40
    "10000000", -- 7795 - 0x1e73  :  128 - 0x80
    "10000000", -- 7796 - 0x1e74  :  128 - 0x80
    "10000011", -- 7797 - 0x1e75  :  131 - 0x83
    "10000111", -- 7798 - 0x1e76  :  135 - 0x87
    "10000111", -- 7799 - 0x1e77  :  135 - 0x87
    "11100000", -- 7800 - 0x1e78  :  224 - 0xe0
    "11000000", -- 7801 - 0x1e79  :  192 - 0xc0
    "10000000", -- 7802 - 0x1e7a  :  128 - 0x80
    "00000000", -- 7803 - 0x1e7b  :    0 - 0x0
    "00000000", -- 7804 - 0x1e7c  :    0 - 0x0
    "00000000", -- 7805 - 0x1e7d  :    0 - 0x0
    "00000000", -- 7806 - 0x1e7e  :    0 - 0x0
    "00000000", -- 7807 - 0x1e7f  :    0 - 0x0
    "11111000", -- 7808 - 0x1e80  :  248 - 0xf8 -- Background 0xe8
    "00000100", -- 7809 - 0x1e81  :    4 - 0x4
    "00000010", -- 7810 - 0x1e82  :    2 - 0x2
    "00000001", -- 7811 - 0x1e83  :    1 - 0x1
    "00000001", -- 7812 - 0x1e84  :    1 - 0x1
    "11000001", -- 7813 - 0x1e85  :  193 - 0xc1
    "11100001", -- 7814 - 0x1e86  :  225 - 0xe1
    "11100001", -- 7815 - 0x1e87  :  225 - 0xe1
    "00000111", -- 7816 - 0x1e88  :    7 - 0x7
    "00000011", -- 7817 - 0x1e89  :    3 - 0x3
    "00000001", -- 7818 - 0x1e8a  :    1 - 0x1
    "00000000", -- 7819 - 0x1e8b  :    0 - 0x0
    "00000000", -- 7820 - 0x1e8c  :    0 - 0x0
    "00000000", -- 7821 - 0x1e8d  :    0 - 0x0
    "00000000", -- 7822 - 0x1e8e  :    0 - 0x0
    "00000000", -- 7823 - 0x1e8f  :    0 - 0x0
    "00000000", -- 7824 - 0x1e90  :    0 - 0x0 -- Background 0xe9
    "00000000", -- 7825 - 0x1e91  :    0 - 0x0
    "00001000", -- 7826 - 0x1e92  :    8 - 0x8
    "00010100", -- 7827 - 0x1e93  :   20 - 0x14
    "00000000", -- 7828 - 0x1e94  :    0 - 0x0
    "00000000", -- 7829 - 0x1e95  :    0 - 0x0
    "01000000", -- 7830 - 0x1e96  :   64 - 0x40
    "10100000", -- 7831 - 0x1e97  :  160 - 0xa0
    "11111111", -- 7832 - 0x1e98  :  255 - 0xff
    "11111111", -- 7833 - 0x1e99  :  255 - 0xff
    "11111111", -- 7834 - 0x1e9a  :  255 - 0xff
    "11111111", -- 7835 - 0x1e9b  :  255 - 0xff
    "11111111", -- 7836 - 0x1e9c  :  255 - 0xff
    "11111111", -- 7837 - 0x1e9d  :  255 - 0xff
    "11111111", -- 7838 - 0x1e9e  :  255 - 0xff
    "11111111", -- 7839 - 0x1e9f  :  255 - 0xff
    "01000000", -- 7840 - 0x1ea0  :   64 - 0x40 -- Background 0xea
    "10100010", -- 7841 - 0x1ea1  :  162 - 0xa2
    "00000101", -- 7842 - 0x1ea2  :    5 - 0x5
    "00000000", -- 7843 - 0x1ea3  :    0 - 0x0
    "00000000", -- 7844 - 0x1ea4  :    0 - 0x0
    "00010000", -- 7845 - 0x1ea5  :   16 - 0x10
    "00101000", -- 7846 - 0x1ea6  :   40 - 0x28
    "00000000", -- 7847 - 0x1ea7  :    0 - 0x0
    "11111111", -- 7848 - 0x1ea8  :  255 - 0xff
    "11111111", -- 7849 - 0x1ea9  :  255 - 0xff
    "11111111", -- 7850 - 0x1eaa  :  255 - 0xff
    "11111111", -- 7851 - 0x1eab  :  255 - 0xff
    "11111111", -- 7852 - 0x1eac  :  255 - 0xff
    "11111111", -- 7853 - 0x1ead  :  255 - 0xff
    "11111111", -- 7854 - 0x1eae  :  255 - 0xff
    "11111111", -- 7855 - 0x1eaf  :  255 - 0xff
    "11111111", -- 7856 - 0x1eb0  :  255 - 0xff -- Background 0xeb
    "11111111", -- 7857 - 0x1eb1  :  255 - 0xff
    "11111111", -- 7858 - 0x1eb2  :  255 - 0xff
    "00000000", -- 7859 - 0x1eb3  :    0 - 0x0
    "00000000", -- 7860 - 0x1eb4  :    0 - 0x0
    "00000000", -- 7861 - 0x1eb5  :    0 - 0x0
    "00000000", -- 7862 - 0x1eb6  :    0 - 0x0
    "11111111", -- 7863 - 0x1eb7  :  255 - 0xff
    "00000000", -- 7864 - 0x1eb8  :    0 - 0x0
    "00000000", -- 7865 - 0x1eb9  :    0 - 0x0
    "00000000", -- 7866 - 0x1eba  :    0 - 0x0
    "00000000", -- 7867 - 0x1ebb  :    0 - 0x0
    "00000000", -- 7868 - 0x1ebc  :    0 - 0x0
    "00000000", -- 7869 - 0x1ebd  :    0 - 0x0
    "00000000", -- 7870 - 0x1ebe  :    0 - 0x0
    "00000000", -- 7871 - 0x1ebf  :    0 - 0x0
    "11100001", -- 7872 - 0x1ec0  :  225 - 0xe1 -- Background 0xec
    "11100001", -- 7873 - 0x1ec1  :  225 - 0xe1
    "11100001", -- 7874 - 0x1ec2  :  225 - 0xe1
    "11100001", -- 7875 - 0x1ec3  :  225 - 0xe1
    "11100001", -- 7876 - 0x1ec4  :  225 - 0xe1
    "11100001", -- 7877 - 0x1ec5  :  225 - 0xe1
    "11100001", -- 7878 - 0x1ec6  :  225 - 0xe1
    "11100001", -- 7879 - 0x1ec7  :  225 - 0xe1
    "00000000", -- 7880 - 0x1ec8  :    0 - 0x0
    "00000000", -- 7881 - 0x1ec9  :    0 - 0x0
    "00000000", -- 7882 - 0x1eca  :    0 - 0x0
    "00000000", -- 7883 - 0x1ecb  :    0 - 0x0
    "00000000", -- 7884 - 0x1ecc  :    0 - 0x0
    "00000000", -- 7885 - 0x1ecd  :    0 - 0x0
    "00000000", -- 7886 - 0x1ece  :    0 - 0x0
    "00000000", -- 7887 - 0x1ecf  :    0 - 0x0
    "11111111", -- 7888 - 0x1ed0  :  255 - 0xff -- Background 0xed
    "11111111", -- 7889 - 0x1ed1  :  255 - 0xff
    "11111111", -- 7890 - 0x1ed2  :  255 - 0xff
    "00000000", -- 7891 - 0x1ed3  :    0 - 0x0
    "00000000", -- 7892 - 0x1ed4  :    0 - 0x0
    "11111111", -- 7893 - 0x1ed5  :  255 - 0xff
    "11111111", -- 7894 - 0x1ed6  :  255 - 0xff
    "11111111", -- 7895 - 0x1ed7  :  255 - 0xff
    "00000000", -- 7896 - 0x1ed8  :    0 - 0x0
    "00000000", -- 7897 - 0x1ed9  :    0 - 0x0
    "00000000", -- 7898 - 0x1eda  :    0 - 0x0
    "11111111", -- 7899 - 0x1edb  :  255 - 0xff
    "11111111", -- 7900 - 0x1edc  :  255 - 0xff
    "00000000", -- 7901 - 0x1edd  :    0 - 0x0
    "00000000", -- 7902 - 0x1ede  :    0 - 0x0
    "00000000", -- 7903 - 0x1edf  :    0 - 0x0
    "11100111", -- 7904 - 0x1ee0  :  231 - 0xe7 -- Background 0xee
    "11100111", -- 7905 - 0x1ee1  :  231 - 0xe7
    "11100111", -- 7906 - 0x1ee2  :  231 - 0xe7
    "11100111", -- 7907 - 0x1ee3  :  231 - 0xe7
    "11100111", -- 7908 - 0x1ee4  :  231 - 0xe7
    "11100111", -- 7909 - 0x1ee5  :  231 - 0xe7
    "11100111", -- 7910 - 0x1ee6  :  231 - 0xe7
    "11100111", -- 7911 - 0x1ee7  :  231 - 0xe7
    "00011000", -- 7912 - 0x1ee8  :   24 - 0x18
    "00011000", -- 7913 - 0x1ee9  :   24 - 0x18
    "00011000", -- 7914 - 0x1eea  :   24 - 0x18
    "00011000", -- 7915 - 0x1eeb  :   24 - 0x18
    "00011000", -- 7916 - 0x1eec  :   24 - 0x18
    "00011000", -- 7917 - 0x1eed  :   24 - 0x18
    "00011000", -- 7918 - 0x1eee  :   24 - 0x18
    "00011000", -- 7919 - 0x1eef  :   24 - 0x18
    "11111111", -- 7920 - 0x1ef0  :  255 - 0xff -- Background 0xef
    "11111111", -- 7921 - 0x1ef1  :  255 - 0xff
    "11111111", -- 7922 - 0x1ef2  :  255 - 0xff
    "11111111", -- 7923 - 0x1ef3  :  255 - 0xff
    "11111111", -- 7924 - 0x1ef4  :  255 - 0xff
    "11111111", -- 7925 - 0x1ef5  :  255 - 0xff
    "11111111", -- 7926 - 0x1ef6  :  255 - 0xff
    "11111111", -- 7927 - 0x1ef7  :  255 - 0xff
    "00110011", -- 7928 - 0x1ef8  :   51 - 0x33
    "00110011", -- 7929 - 0x1ef9  :   51 - 0x33
    "11001100", -- 7930 - 0x1efa  :  204 - 0xcc
    "11001100", -- 7931 - 0x1efb  :  204 - 0xcc
    "00110011", -- 7932 - 0x1efc  :   51 - 0x33
    "00110011", -- 7933 - 0x1efd  :   51 - 0x33
    "11001100", -- 7934 - 0x1efe  :  204 - 0xcc
    "11001100", -- 7935 - 0x1eff  :  204 - 0xcc
    "00000000", -- 7936 - 0x1f00  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 7937 - 0x1f01  :    0 - 0x0
    "00000000", -- 7938 - 0x1f02  :    0 - 0x0
    "00000000", -- 7939 - 0x1f03  :    0 - 0x0
    "00000000", -- 7940 - 0x1f04  :    0 - 0x0
    "00000000", -- 7941 - 0x1f05  :    0 - 0x0
    "00000000", -- 7942 - 0x1f06  :    0 - 0x0
    "00000000", -- 7943 - 0x1f07  :    0 - 0x0
    "00000000", -- 7944 - 0x1f08  :    0 - 0x0
    "00000000", -- 7945 - 0x1f09  :    0 - 0x0
    "00000000", -- 7946 - 0x1f0a  :    0 - 0x0
    "00000000", -- 7947 - 0x1f0b  :    0 - 0x0
    "00000000", -- 7948 - 0x1f0c  :    0 - 0x0
    "00000000", -- 7949 - 0x1f0d  :    0 - 0x0
    "00000000", -- 7950 - 0x1f0e  :    0 - 0x0
    "00000000", -- 7951 - 0x1f0f  :    0 - 0x0
    "00000000", -- 7952 - 0x1f10  :    0 - 0x0 -- Background 0xf1
    "00000000", -- 7953 - 0x1f11  :    0 - 0x0
    "00000000", -- 7954 - 0x1f12  :    0 - 0x0
    "00000000", -- 7955 - 0x1f13  :    0 - 0x0
    "00000000", -- 7956 - 0x1f14  :    0 - 0x0
    "00000000", -- 7957 - 0x1f15  :    0 - 0x0
    "00000000", -- 7958 - 0x1f16  :    0 - 0x0
    "00000000", -- 7959 - 0x1f17  :    0 - 0x0
    "00000000", -- 7960 - 0x1f18  :    0 - 0x0
    "00000000", -- 7961 - 0x1f19  :    0 - 0x0
    "00000000", -- 7962 - 0x1f1a  :    0 - 0x0
    "00000000", -- 7963 - 0x1f1b  :    0 - 0x0
    "00000000", -- 7964 - 0x1f1c  :    0 - 0x0
    "00000000", -- 7965 - 0x1f1d  :    0 - 0x0
    "00000000", -- 7966 - 0x1f1e  :    0 - 0x0
    "00000000", -- 7967 - 0x1f1f  :    0 - 0x0
    "00000000", -- 7968 - 0x1f20  :    0 - 0x0 -- Background 0xf2
    "00000000", -- 7969 - 0x1f21  :    0 - 0x0
    "00000000", -- 7970 - 0x1f22  :    0 - 0x0
    "00000000", -- 7971 - 0x1f23  :    0 - 0x0
    "00000000", -- 7972 - 0x1f24  :    0 - 0x0
    "00000000", -- 7973 - 0x1f25  :    0 - 0x0
    "00000000", -- 7974 - 0x1f26  :    0 - 0x0
    "00000000", -- 7975 - 0x1f27  :    0 - 0x0
    "00000000", -- 7976 - 0x1f28  :    0 - 0x0
    "00000000", -- 7977 - 0x1f29  :    0 - 0x0
    "00000000", -- 7978 - 0x1f2a  :    0 - 0x0
    "00000000", -- 7979 - 0x1f2b  :    0 - 0x0
    "00000000", -- 7980 - 0x1f2c  :    0 - 0x0
    "00000000", -- 7981 - 0x1f2d  :    0 - 0x0
    "00000000", -- 7982 - 0x1f2e  :    0 - 0x0
    "00000000", -- 7983 - 0x1f2f  :    0 - 0x0
    "00000000", -- 7984 - 0x1f30  :    0 - 0x0 -- Background 0xf3
    "00000000", -- 7985 - 0x1f31  :    0 - 0x0
    "00000000", -- 7986 - 0x1f32  :    0 - 0x0
    "00000000", -- 7987 - 0x1f33  :    0 - 0x0
    "00000000", -- 7988 - 0x1f34  :    0 - 0x0
    "00000000", -- 7989 - 0x1f35  :    0 - 0x0
    "00000000", -- 7990 - 0x1f36  :    0 - 0x0
    "00000000", -- 7991 - 0x1f37  :    0 - 0x0
    "00000000", -- 7992 - 0x1f38  :    0 - 0x0
    "00000000", -- 7993 - 0x1f39  :    0 - 0x0
    "00000000", -- 7994 - 0x1f3a  :    0 - 0x0
    "00000000", -- 7995 - 0x1f3b  :    0 - 0x0
    "00000000", -- 7996 - 0x1f3c  :    0 - 0x0
    "00000000", -- 7997 - 0x1f3d  :    0 - 0x0
    "00000000", -- 7998 - 0x1f3e  :    0 - 0x0
    "00000000", -- 7999 - 0x1f3f  :    0 - 0x0
    "11100111", -- 8000 - 0x1f40  :  231 - 0xe7 -- Background 0xf4
    "10011001", -- 8001 - 0x1f41  :  153 - 0x99
    "10000001", -- 8002 - 0x1f42  :  129 - 0x81
    "11000011", -- 8003 - 0x1f43  :  195 - 0xc3
    "11111111", -- 8004 - 0x1f44  :  255 - 0xff
    "10111101", -- 8005 - 0x1f45  :  189 - 0xbd
    "10000001", -- 8006 - 0x1f46  :  129 - 0x81
    "11000011", -- 8007 - 0x1f47  :  195 - 0xc3
    "00100100", -- 8008 - 0x1f48  :   36 - 0x24
    "00011000", -- 8009 - 0x1f49  :   24 - 0x18
    "00000000", -- 8010 - 0x1f4a  :    0 - 0x0
    "01000010", -- 8011 - 0x1f4b  :   66 - 0x42
    "01111110", -- 8012 - 0x1f4c  :  126 - 0x7e
    "00111100", -- 8013 - 0x1f4d  :   60 - 0x3c
    "00000000", -- 8014 - 0x1f4e  :    0 - 0x0
    "00000000", -- 8015 - 0x1f4f  :    0 - 0x0
    "11100001", -- 8016 - 0x1f50  :  225 - 0xe1 -- Background 0xf5
    "11100000", -- 8017 - 0x1f51  :  224 - 0xe0
    "11100000", -- 8018 - 0x1f52  :  224 - 0xe0
    "11100000", -- 8019 - 0x1f53  :  224 - 0xe0
    "11100000", -- 8020 - 0x1f54  :  224 - 0xe0
    "11111111", -- 8021 - 0x1f55  :  255 - 0xff
    "11111111", -- 8022 - 0x1f56  :  255 - 0xff
    "01111111", -- 8023 - 0x1f57  :  127 - 0x7f
    "00000000", -- 8024 - 0x1f58  :    0 - 0x0
    "00000000", -- 8025 - 0x1f59  :    0 - 0x0
    "00000000", -- 8026 - 0x1f5a  :    0 - 0x0
    "00000000", -- 8027 - 0x1f5b  :    0 - 0x0
    "00000000", -- 8028 - 0x1f5c  :    0 - 0x0
    "00000000", -- 8029 - 0x1f5d  :    0 - 0x0
    "00000000", -- 8030 - 0x1f5e  :    0 - 0x0
    "00000000", -- 8031 - 0x1f5f  :    0 - 0x0
    "10000111", -- 8032 - 0x1f60  :  135 - 0x87 -- Background 0xf6
    "00000111", -- 8033 - 0x1f61  :    7 - 0x7
    "00000111", -- 8034 - 0x1f62  :    7 - 0x7
    "00000111", -- 8035 - 0x1f63  :    7 - 0x7
    "00000111", -- 8036 - 0x1f64  :    7 - 0x7
    "11111111", -- 8037 - 0x1f65  :  255 - 0xff
    "11111111", -- 8038 - 0x1f66  :  255 - 0xff
    "11111110", -- 8039 - 0x1f67  :  254 - 0xfe
    "00000000", -- 8040 - 0x1f68  :    0 - 0x0
    "00000000", -- 8041 - 0x1f69  :    0 - 0x0
    "00000000", -- 8042 - 0x1f6a  :    0 - 0x0
    "00000000", -- 8043 - 0x1f6b  :    0 - 0x0
    "00000000", -- 8044 - 0x1f6c  :    0 - 0x0
    "00000000", -- 8045 - 0x1f6d  :    0 - 0x0
    "00000000", -- 8046 - 0x1f6e  :    0 - 0x0
    "00000000", -- 8047 - 0x1f6f  :    0 - 0x0
    "10000111", -- 8048 - 0x1f70  :  135 - 0x87 -- Background 0xf7
    "10000111", -- 8049 - 0x1f71  :  135 - 0x87
    "10000011", -- 8050 - 0x1f72  :  131 - 0x83
    "10000000", -- 8051 - 0x1f73  :  128 - 0x80
    "10000000", -- 8052 - 0x1f74  :  128 - 0x80
    "01000000", -- 8053 - 0x1f75  :   64 - 0x40
    "00100000", -- 8054 - 0x1f76  :   32 - 0x20
    "00011111", -- 8055 - 0x1f77  :   31 - 0x1f
    "00000000", -- 8056 - 0x1f78  :    0 - 0x0
    "00000000", -- 8057 - 0x1f79  :    0 - 0x0
    "00000000", -- 8058 - 0x1f7a  :    0 - 0x0
    "00000000", -- 8059 - 0x1f7b  :    0 - 0x0
    "00000000", -- 8060 - 0x1f7c  :    0 - 0x0
    "10000000", -- 8061 - 0x1f7d  :  128 - 0x80
    "11000000", -- 8062 - 0x1f7e  :  192 - 0xc0
    "11100000", -- 8063 - 0x1f7f  :  224 - 0xe0
    "11100001", -- 8064 - 0x1f80  :  225 - 0xe1 -- Background 0xf8
    "11100001", -- 8065 - 0x1f81  :  225 - 0xe1
    "11000001", -- 8066 - 0x1f82  :  193 - 0xc1
    "00000001", -- 8067 - 0x1f83  :    1 - 0x1
    "00000001", -- 8068 - 0x1f84  :    1 - 0x1
    "00000010", -- 8069 - 0x1f85  :    2 - 0x2
    "00000100", -- 8070 - 0x1f86  :    4 - 0x4
    "11111000", -- 8071 - 0x1f87  :  248 - 0xf8
    "00000000", -- 8072 - 0x1f88  :    0 - 0x0
    "00000000", -- 8073 - 0x1f89  :    0 - 0x0
    "00000000", -- 8074 - 0x1f8a  :    0 - 0x0
    "00000000", -- 8075 - 0x1f8b  :    0 - 0x0
    "00000000", -- 8076 - 0x1f8c  :    0 - 0x0
    "00000001", -- 8077 - 0x1f8d  :    1 - 0x1
    "00000011", -- 8078 - 0x1f8e  :    3 - 0x3
    "00000111", -- 8079 - 0x1f8f  :    7 - 0x7
    "00000000", -- 8080 - 0x1f90  :    0 - 0x0 -- Background 0xf9
    "00000010", -- 8081 - 0x1f91  :    2 - 0x2
    "00000101", -- 8082 - 0x1f92  :    5 - 0x5
    "00000000", -- 8083 - 0x1f93  :    0 - 0x0
    "00100000", -- 8084 - 0x1f94  :   32 - 0x20
    "01010000", -- 8085 - 0x1f95  :   80 - 0x50
    "00000000", -- 8086 - 0x1f96  :    0 - 0x0
    "00000000", -- 8087 - 0x1f97  :    0 - 0x0
    "11111111", -- 8088 - 0x1f98  :  255 - 0xff
    "11111111", -- 8089 - 0x1f99  :  255 - 0xff
    "11111111", -- 8090 - 0x1f9a  :  255 - 0xff
    "11111111", -- 8091 - 0x1f9b  :  255 - 0xff
    "11111111", -- 8092 - 0x1f9c  :  255 - 0xff
    "11111111", -- 8093 - 0x1f9d  :  255 - 0xff
    "11111111", -- 8094 - 0x1f9e  :  255 - 0xff
    "11111111", -- 8095 - 0x1f9f  :  255 - 0xff
    "00000000", -- 8096 - 0x1fa0  :    0 - 0x0 -- Background 0xfa
    "00000000", -- 8097 - 0x1fa1  :    0 - 0x0
    "00000000", -- 8098 - 0x1fa2  :    0 - 0x0
    "00000000", -- 8099 - 0x1fa3  :    0 - 0x0
    "00000000", -- 8100 - 0x1fa4  :    0 - 0x0
    "00000000", -- 8101 - 0x1fa5  :    0 - 0x0
    "00000000", -- 8102 - 0x1fa6  :    0 - 0x0
    "00000000", -- 8103 - 0x1fa7  :    0 - 0x0
    "11111111", -- 8104 - 0x1fa8  :  255 - 0xff
    "11111111", -- 8105 - 0x1fa9  :  255 - 0xff
    "11111111", -- 8106 - 0x1faa  :  255 - 0xff
    "11111111", -- 8107 - 0x1fab  :  255 - 0xff
    "11111111", -- 8108 - 0x1fac  :  255 - 0xff
    "11111111", -- 8109 - 0x1fad  :  255 - 0xff
    "11111111", -- 8110 - 0x1fae  :  255 - 0xff
    "11111111", -- 8111 - 0x1faf  :  255 - 0xff
    "11111111", -- 8112 - 0x1fb0  :  255 - 0xff -- Background 0xfb
    "00000000", -- 8113 - 0x1fb1  :    0 - 0x0
    "00000000", -- 8114 - 0x1fb2  :    0 - 0x0
    "00000000", -- 8115 - 0x1fb3  :    0 - 0x0
    "00000000", -- 8116 - 0x1fb4  :    0 - 0x0
    "11111111", -- 8117 - 0x1fb5  :  255 - 0xff
    "11111111", -- 8118 - 0x1fb6  :  255 - 0xff
    "11111111", -- 8119 - 0x1fb7  :  255 - 0xff
    "00000000", -- 8120 - 0x1fb8  :    0 - 0x0
    "00000000", -- 8121 - 0x1fb9  :    0 - 0x0
    "00000000", -- 8122 - 0x1fba  :    0 - 0x0
    "00000000", -- 8123 - 0x1fbb  :    0 - 0x0
    "00000000", -- 8124 - 0x1fbc  :    0 - 0x0
    "00000000", -- 8125 - 0x1fbd  :    0 - 0x0
    "00000000", -- 8126 - 0x1fbe  :    0 - 0x0
    "00000000", -- 8127 - 0x1fbf  :    0 - 0x0
    "10000111", -- 8128 - 0x1fc0  :  135 - 0x87 -- Background 0xfc
    "10000111", -- 8129 - 0x1fc1  :  135 - 0x87
    "10000111", -- 8130 - 0x1fc2  :  135 - 0x87
    "10000111", -- 8131 - 0x1fc3  :  135 - 0x87
    "10000111", -- 8132 - 0x1fc4  :  135 - 0x87
    "10000111", -- 8133 - 0x1fc5  :  135 - 0x87
    "10000111", -- 8134 - 0x1fc6  :  135 - 0x87
    "10000111", -- 8135 - 0x1fc7  :  135 - 0x87
    "00000000", -- 8136 - 0x1fc8  :    0 - 0x0
    "00000000", -- 8137 - 0x1fc9  :    0 - 0x0
    "00000000", -- 8138 - 0x1fca  :    0 - 0x0
    "00000000", -- 8139 - 0x1fcb  :    0 - 0x0
    "00000000", -- 8140 - 0x1fcc  :    0 - 0x0
    "00000000", -- 8141 - 0x1fcd  :    0 - 0x0
    "00000000", -- 8142 - 0x1fce  :    0 - 0x0
    "00000000", -- 8143 - 0x1fcf  :    0 - 0x0
    "11111111", -- 8144 - 0x1fd0  :  255 - 0xff -- Background 0xfd
    "11111111", -- 8145 - 0x1fd1  :  255 - 0xff
    "11111111", -- 8146 - 0x1fd2  :  255 - 0xff
    "11000011", -- 8147 - 0x1fd3  :  195 - 0xc3
    "11000011", -- 8148 - 0x1fd4  :  195 - 0xc3
    "11111111", -- 8149 - 0x1fd5  :  255 - 0xff
    "11111111", -- 8150 - 0x1fd6  :  255 - 0xff
    "11111111", -- 8151 - 0x1fd7  :  255 - 0xff
    "00000000", -- 8152 - 0x1fd8  :    0 - 0x0
    "00000000", -- 8153 - 0x1fd9  :    0 - 0x0
    "00000000", -- 8154 - 0x1fda  :    0 - 0x0
    "00111100", -- 8155 - 0x1fdb  :   60 - 0x3c
    "00111100", -- 8156 - 0x1fdc  :   60 - 0x3c
    "00000000", -- 8157 - 0x1fdd  :    0 - 0x0
    "00000000", -- 8158 - 0x1fde  :    0 - 0x0
    "00000000", -- 8159 - 0x1fdf  :    0 - 0x0
    "11111111", -- 8160 - 0x1fe0  :  255 - 0xff -- Background 0xfe
    "11111111", -- 8161 - 0x1fe1  :  255 - 0xff
    "11100111", -- 8162 - 0x1fe2  :  231 - 0xe7
    "11100111", -- 8163 - 0x1fe3  :  231 - 0xe7
    "11100111", -- 8164 - 0x1fe4  :  231 - 0xe7
    "11100111", -- 8165 - 0x1fe5  :  231 - 0xe7
    "11111111", -- 8166 - 0x1fe6  :  255 - 0xff
    "11111111", -- 8167 - 0x1fe7  :  255 - 0xff
    "00000000", -- 8168 - 0x1fe8  :    0 - 0x0
    "00000000", -- 8169 - 0x1fe9  :    0 - 0x0
    "00011000", -- 8170 - 0x1fea  :   24 - 0x18
    "00011000", -- 8171 - 0x1feb  :   24 - 0x18
    "00011000", -- 8172 - 0x1fec  :   24 - 0x18
    "00011000", -- 8173 - 0x1fed  :   24 - 0x18
    "00000000", -- 8174 - 0x1fee  :    0 - 0x0
    "00000000", -- 8175 - 0x1fef  :    0 - 0x0
    "11111111", -- 8176 - 0x1ff0  :  255 - 0xff -- Background 0xff
    "11111111", -- 8177 - 0x1ff1  :  255 - 0xff
    "11111111", -- 8178 - 0x1ff2  :  255 - 0xff
    "11111111", -- 8179 - 0x1ff3  :  255 - 0xff
    "11111111", -- 8180 - 0x1ff4  :  255 - 0xff
    "11111111", -- 8181 - 0x1ff5  :  255 - 0xff
    "11111111", -- 8182 - 0x1ff6  :  255 - 0xff
    "11111111", -- 8183 - 0x1ff7  :  255 - 0xff
    "00000000", -- 8184 - 0x1ff8  :    0 - 0x0
    "00000000", -- 8185 - 0x1ff9  :    0 - 0x0
    "00000000", -- 8186 - 0x1ffa  :    0 - 0x0
    "00000000", -- 8187 - 0x1ffb  :    0 - 0x0
    "00000000", -- 8188 - 0x1ffc  :    0 - 0x0
    "00000000", -- 8189 - 0x1ffd  :    0 - 0x0
    "00000000", -- 8190 - 0x1ffe  :    0 - 0x0
    "00000000"  -- 8191 - 0x1fff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
