---   Sprites Pattern table COLOR PLANE 0
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: smario_traspas_patron.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_MARIO_TRASPAS_SPR_PLN0 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_MARIO_TRASPAS_SPR_PLN0;

architecture BEHAVIORAL of ROM_PTABLE_MARIO_TRASPAS_SPR_PLN0 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table COLOR PLANE 0
    "00000011", --    0 -  0x0  :    3 - 0x3 -- Sprite 0x0
    "00001111", --    1 -  0x1  :   15 - 0xf
    "00011111", --    2 -  0x2  :   31 - 0x1f
    "00011111", --    3 -  0x3  :   31 - 0x1f
    "00011100", --    4 -  0x4  :   28 - 0x1c
    "00100100", --    5 -  0x5  :   36 - 0x24
    "00100110", --    6 -  0x6  :   38 - 0x26
    "01100110", --    7 -  0x7  :  102 - 0x66
    "11100000", --    8 -  0x8  :  224 - 0xe0 -- Sprite 0x1
    "11000000", --    9 -  0x9  :  192 - 0xc0
    "10000000", --   10 -  0xa  :  128 - 0x80
    "11111100", --   11 -  0xb  :  252 - 0xfc
    "10000000", --   12 -  0xc  :  128 - 0x80
    "11000000", --   13 -  0xd  :  192 - 0xc0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00100000", --   15 -  0xf  :   32 - 0x20
    "01100000", --   16 - 0x10  :   96 - 0x60 -- Sprite 0x2
    "01110000", --   17 - 0x11  :  112 - 0x70
    "00011000", --   18 - 0x12  :   24 - 0x18
    "00000111", --   19 - 0x13  :    7 - 0x7
    "00001111", --   20 - 0x14  :   15 - 0xf
    "00011111", --   21 - 0x15  :   31 - 0x1f
    "00111111", --   22 - 0x16  :   63 - 0x3f
    "01111111", --   23 - 0x17  :  127 - 0x7f
    "11111100", --   24 - 0x18  :  252 - 0xfc -- Sprite 0x3
    "01111100", --   25 - 0x19  :  124 - 0x7c
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "11100000", --   28 - 0x1c  :  224 - 0xe0
    "11110000", --   29 - 0x1d  :  240 - 0xf0
    "11111000", --   30 - 0x1e  :  248 - 0xf8
    "11111000", --   31 - 0x1f  :  248 - 0xf8
    "01111111", --   32 - 0x20  :  127 - 0x7f -- Sprite 0x4
    "01111111", --   33 - 0x21  :  127 - 0x7f
    "11111111", --   34 - 0x22  :  255 - 0xff
    "11111111", --   35 - 0x23  :  255 - 0xff
    "00000111", --   36 - 0x24  :    7 - 0x7
    "00000111", --   37 - 0x25  :    7 - 0x7
    "00001111", --   38 - 0x26  :   15 - 0xf
    "00001111", --   39 - 0x27  :   15 - 0xf
    "11111101", --   40 - 0x28  :  253 - 0xfd -- Sprite 0x5
    "11111110", --   41 - 0x29  :  254 - 0xfe
    "10110100", --   42 - 0x2a  :  180 - 0xb4
    "11111000", --   43 - 0x2b  :  248 - 0xf8
    "11111000", --   44 - 0x2c  :  248 - 0xf8
    "11111001", --   45 - 0x2d  :  249 - 0xf9
    "11111011", --   46 - 0x2e  :  251 - 0xfb
    "11111111", --   47 - 0x2f  :  255 - 0xff
    "00011111", --   48 - 0x30  :   31 - 0x1f -- Sprite 0x6
    "00111111", --   49 - 0x31  :   63 - 0x3f
    "11111111", --   50 - 0x32  :  255 - 0xff
    "11111111", --   51 - 0x33  :  255 - 0xff
    "11111100", --   52 - 0x34  :  252 - 0xfc
    "01110000", --   53 - 0x35  :  112 - 0x70
    "01110000", --   54 - 0x36  :  112 - 0x70
    "00111000", --   55 - 0x37  :   56 - 0x38
    "11111111", --   56 - 0x38  :  255 - 0xff -- Sprite 0x7
    "11111111", --   57 - 0x39  :  255 - 0xff
    "11111111", --   58 - 0x3a  :  255 - 0xff
    "00011111", --   59 - 0x3b  :   31 - 0x1f
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Sprite 0x8
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000001", --   66 - 0x42  :    1 - 0x1
    "00000111", --   67 - 0x43  :    7 - 0x7
    "00001111", --   68 - 0x44  :   15 - 0xf
    "00001111", --   69 - 0x45  :   15 - 0xf
    "00001110", --   70 - 0x46  :   14 - 0xe
    "00010010", --   71 - 0x47  :   18 - 0x12
    "00000000", --   72 - 0x48  :    0 - 0x0 -- Sprite 0x9
    "00000000", --   73 - 0x49  :    0 - 0x0
    "11110000", --   74 - 0x4a  :  240 - 0xf0
    "11100000", --   75 - 0x4b  :  224 - 0xe0
    "11000000", --   76 - 0x4c  :  192 - 0xc0
    "11111110", --   77 - 0x4d  :  254 - 0xfe
    "01000000", --   78 - 0x4e  :   64 - 0x40
    "01100000", --   79 - 0x4f  :   96 - 0x60
    "00010011", --   80 - 0x50  :   19 - 0x13 -- Sprite 0xa
    "00110011", --   81 - 0x51  :   51 - 0x33
    "00110000", --   82 - 0x52  :   48 - 0x30
    "00011000", --   83 - 0x53  :   24 - 0x18
    "00000100", --   84 - 0x54  :    4 - 0x4
    "00001111", --   85 - 0x55  :   15 - 0xf
    "00011111", --   86 - 0x56  :   31 - 0x1f
    "00011111", --   87 - 0x57  :   31 - 0x1f
    "00000000", --   88 - 0x58  :    0 - 0x0 -- Sprite 0xb
    "00010000", --   89 - 0x59  :   16 - 0x10
    "01111110", --   90 - 0x5a  :  126 - 0x7e
    "00111110", --   91 - 0x5b  :   62 - 0x3e
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "11000000", --   94 - 0x5e  :  192 - 0xc0
    "11100000", --   95 - 0x5f  :  224 - 0xe0
    "00111111", --   96 - 0x60  :   63 - 0x3f -- Sprite 0xc
    "00111111", --   97 - 0x61  :   63 - 0x3f
    "00111111", --   98 - 0x62  :   63 - 0x3f
    "00011111", --   99 - 0x63  :   31 - 0x1f
    "00011111", --  100 - 0x64  :   31 - 0x1f
    "00011111", --  101 - 0x65  :   31 - 0x1f
    "00011111", --  102 - 0x66  :   31 - 0x1f
    "00011111", --  103 - 0x67  :   31 - 0x1f
    "11110000", --  104 - 0x68  :  240 - 0xf0 -- Sprite 0xd
    "11110000", --  105 - 0x69  :  240 - 0xf0
    "11110000", --  106 - 0x6a  :  240 - 0xf0
    "11111000", --  107 - 0x6b  :  248 - 0xf8
    "11111000", --  108 - 0x6c  :  248 - 0xf8
    "11111000", --  109 - 0x6d  :  248 - 0xf8
    "11111000", --  110 - 0x6e  :  248 - 0xf8
    "11111000", --  111 - 0x6f  :  248 - 0xf8
    "11111111", --  112 - 0x70  :  255 - 0xff -- Sprite 0xe
    "11111111", --  113 - 0x71  :  255 - 0xff
    "11111111", --  114 - 0x72  :  255 - 0xff
    "11111110", --  115 - 0x73  :  254 - 0xfe
    "11110000", --  116 - 0x74  :  240 - 0xf0
    "11000000", --  117 - 0x75  :  192 - 0xc0
    "10000000", --  118 - 0x76  :  128 - 0x80
    "00000000", --  119 - 0x77  :    0 - 0x0
    "11111100", --  120 - 0x78  :  252 - 0xfc -- Sprite 0xf
    "11111100", --  121 - 0x79  :  252 - 0xfc
    "11111000", --  122 - 0x7a  :  248 - 0xf8
    "01111000", --  123 - 0x7b  :  120 - 0x78
    "01111000", --  124 - 0x7c  :  120 - 0x78
    "01111000", --  125 - 0x7d  :  120 - 0x78
    "01111110", --  126 - 0x7e  :  126 - 0x7e
    "01111110", --  127 - 0x7f  :  126 - 0x7e
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x10
    "00000011", --  129 - 0x81  :    3 - 0x3
    "00001111", --  130 - 0x82  :   15 - 0xf
    "00011111", --  131 - 0x83  :   31 - 0x1f
    "00011111", --  132 - 0x84  :   31 - 0x1f
    "00011100", --  133 - 0x85  :   28 - 0x1c
    "00100100", --  134 - 0x86  :   36 - 0x24
    "00100110", --  135 - 0x87  :   38 - 0x26
    "00000000", --  136 - 0x88  :    0 - 0x0 -- Sprite 0x11
    "11100000", --  137 - 0x89  :  224 - 0xe0
    "11000000", --  138 - 0x8a  :  192 - 0xc0
    "10000000", --  139 - 0x8b  :  128 - 0x80
    "11111100", --  140 - 0x8c  :  252 - 0xfc
    "10000000", --  141 - 0x8d  :  128 - 0x80
    "11000000", --  142 - 0x8e  :  192 - 0xc0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "01100110", --  144 - 0x90  :  102 - 0x66 -- Sprite 0x12
    "01100000", --  145 - 0x91  :   96 - 0x60
    "00110000", --  146 - 0x92  :   48 - 0x30
    "00011000", --  147 - 0x93  :   24 - 0x18
    "00001111", --  148 - 0x94  :   15 - 0xf
    "00011111", --  149 - 0x95  :   31 - 0x1f
    "00111111", --  150 - 0x96  :   63 - 0x3f
    "00111111", --  151 - 0x97  :   63 - 0x3f
    "00100000", --  152 - 0x98  :   32 - 0x20 -- Sprite 0x13
    "11111100", --  153 - 0x99  :  252 - 0xfc
    "01111100", --  154 - 0x9a  :  124 - 0x7c
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "11100000", --  157 - 0x9d  :  224 - 0xe0
    "11100000", --  158 - 0x9e  :  224 - 0xe0
    "11110000", --  159 - 0x9f  :  240 - 0xf0
    "00111111", --  160 - 0xa0  :   63 - 0x3f -- Sprite 0x14
    "00111111", --  161 - 0xa1  :   63 - 0x3f
    "00111111", --  162 - 0xa2  :   63 - 0x3f
    "00111111", --  163 - 0xa3  :   63 - 0x3f
    "00111111", --  164 - 0xa4  :   63 - 0x3f
    "00111111", --  165 - 0xa5  :   63 - 0x3f
    "00111111", --  166 - 0xa6  :   63 - 0x3f
    "00011111", --  167 - 0xa7  :   31 - 0x1f
    "11110000", --  168 - 0xa8  :  240 - 0xf0 -- Sprite 0x15
    "10010000", --  169 - 0xa9  :  144 - 0x90
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00001000", --  171 - 0xab  :    8 - 0x8
    "00001100", --  172 - 0xac  :   12 - 0xc
    "00011100", --  173 - 0xad  :   28 - 0x1c
    "11111100", --  174 - 0xae  :  252 - 0xfc
    "11111000", --  175 - 0xaf  :  248 - 0xf8
    "00001111", --  176 - 0xb0  :   15 - 0xf -- Sprite 0x16
    "00001111", --  177 - 0xb1  :   15 - 0xf
    "00000111", --  178 - 0xb2  :    7 - 0x7
    "00000111", --  179 - 0xb3  :    7 - 0x7
    "00000111", --  180 - 0xb4  :    7 - 0x7
    "00001111", --  181 - 0xb5  :   15 - 0xf
    "00001111", --  182 - 0xb6  :   15 - 0xf
    "00000011", --  183 - 0xb7  :    3 - 0x3
    "11111000", --  184 - 0xb8  :  248 - 0xf8 -- Sprite 0x17
    "11110000", --  185 - 0xb9  :  240 - 0xf0
    "11100000", --  186 - 0xba  :  224 - 0xe0
    "11110000", --  187 - 0xbb  :  240 - 0xf0
    "10110000", --  188 - 0xbc  :  176 - 0xb0
    "10000000", --  189 - 0xbd  :  128 - 0x80
    "11100000", --  190 - 0xbe  :  224 - 0xe0
    "11100000", --  191 - 0xbf  :  224 - 0xe0
    "00000011", --  192 - 0xc0  :    3 - 0x3 -- Sprite 0x18
    "00111111", --  193 - 0xc1  :   63 - 0x3f
    "01111111", --  194 - 0xc2  :  127 - 0x7f
    "00011001", --  195 - 0xc3  :   25 - 0x19
    "00001001", --  196 - 0xc4  :    9 - 0x9
    "00001001", --  197 - 0xc5  :    9 - 0x9
    "00101000", --  198 - 0xc6  :   40 - 0x28
    "01011100", --  199 - 0xc7  :   92 - 0x5c
    "11111000", --  200 - 0xc8  :  248 - 0xf8 -- Sprite 0x19
    "11100000", --  201 - 0xc9  :  224 - 0xe0
    "11100000", --  202 - 0xca  :  224 - 0xe0
    "11111100", --  203 - 0xcb  :  252 - 0xfc
    "00100110", --  204 - 0xcc  :   38 - 0x26
    "00110000", --  205 - 0xcd  :   48 - 0x30
    "10000000", --  206 - 0xce  :  128 - 0x80
    "00010000", --  207 - 0xcf  :   16 - 0x10
    "00111110", --  208 - 0xd0  :   62 - 0x3e -- Sprite 0x1a
    "00011110", --  209 - 0xd1  :   30 - 0x1e
    "00111111", --  210 - 0xd2  :   63 - 0x3f
    "00111000", --  211 - 0xd3  :   56 - 0x38
    "00110000", --  212 - 0xd4  :   48 - 0x30
    "00110000", --  213 - 0xd5  :   48 - 0x30
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00111010", --  215 - 0xd7  :   58 - 0x3a
    "01111000", --  216 - 0xd8  :  120 - 0x78 -- Sprite 0x1b
    "00011110", --  217 - 0xd9  :   30 - 0x1e
    "10000000", --  218 - 0xda  :  128 - 0x80
    "11111110", --  219 - 0xdb  :  254 - 0xfe
    "01111110", --  220 - 0xdc  :  126 - 0x7e
    "01111110", --  221 - 0xdd  :  126 - 0x7e
    "01111111", --  222 - 0xde  :  127 - 0x7f
    "01111111", --  223 - 0xdf  :  127 - 0x7f
    "00111100", --  224 - 0xe0  :   60 - 0x3c -- Sprite 0x1c
    "00111111", --  225 - 0xe1  :   63 - 0x3f
    "00011111", --  226 - 0xe2  :   31 - 0x1f
    "00001111", --  227 - 0xe3  :   15 - 0xf
    "00000111", --  228 - 0xe4  :    7 - 0x7
    "00111111", --  229 - 0xe5  :   63 - 0x3f
    "00100001", --  230 - 0xe6  :   33 - 0x21
    "00100000", --  231 - 0xe7  :   32 - 0x20
    "11111111", --  232 - 0xe8  :  255 - 0xff -- Sprite 0x1d
    "11111111", --  233 - 0xe9  :  255 - 0xff
    "11111111", --  234 - 0xea  :  255 - 0xff
    "11111110", --  235 - 0xeb  :  254 - 0xfe
    "11111110", --  236 - 0xec  :  254 - 0xfe
    "11111110", --  237 - 0xed  :  254 - 0xfe
    "11111100", --  238 - 0xee  :  252 - 0xfc
    "01110000", --  239 - 0xef  :  112 - 0x70
    "00001111", --  240 - 0xf0  :   15 - 0xf -- Sprite 0x1e
    "10011111", --  241 - 0xf1  :  159 - 0x9f
    "11001111", --  242 - 0xf2  :  207 - 0xcf
    "11111111", --  243 - 0xf3  :  255 - 0xff
    "01111111", --  244 - 0xf4  :  127 - 0x7f
    "00111111", --  245 - 0xf5  :   63 - 0x3f
    "00011110", --  246 - 0xf6  :   30 - 0x1e
    "00001110", --  247 - 0xf7  :   14 - 0xe
    "00100000", --  248 - 0xf8  :   32 - 0x20 -- Sprite 0x1f
    "11000000", --  249 - 0xf9  :  192 - 0xc0
    "10000000", --  250 - 0xfa  :  128 - 0x80
    "10000000", --  251 - 0xfb  :  128 - 0x80
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000011", --  258 - 0x102  :    3 - 0x3
    "00001111", --  259 - 0x103  :   15 - 0xf
    "00011111", --  260 - 0x104  :   31 - 0x1f
    "00011111", --  261 - 0x105  :   31 - 0x1f
    "00011100", --  262 - 0x106  :   28 - 0x1c
    "00100100", --  263 - 0x107  :   36 - 0x24
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Sprite 0x21
    "00000100", --  265 - 0x109  :    4 - 0x4
    "11100110", --  266 - 0x10a  :  230 - 0xe6
    "11100000", --  267 - 0x10b  :  224 - 0xe0
    "11111111", --  268 - 0x10c  :  255 - 0xff
    "11111111", --  269 - 0x10d  :  255 - 0xff
    "10001111", --  270 - 0x10e  :  143 - 0x8f
    "10000011", --  271 - 0x10f  :  131 - 0x83
    "00100110", --  272 - 0x110  :   38 - 0x26 -- Sprite 0x22
    "00100110", --  273 - 0x111  :   38 - 0x26
    "01100000", --  274 - 0x112  :   96 - 0x60
    "01111000", --  275 - 0x113  :  120 - 0x78
    "00011000", --  276 - 0x114  :   24 - 0x18
    "00001111", --  277 - 0x115  :   15 - 0xf
    "01111111", --  278 - 0x116  :  127 - 0x7f
    "11111111", --  279 - 0x117  :  255 - 0xff
    "00000001", --  280 - 0x118  :    1 - 0x1 -- Sprite 0x23
    "00100001", --  281 - 0x119  :   33 - 0x21
    "11111110", --  282 - 0x11a  :  254 - 0xfe
    "01111010", --  283 - 0x11b  :  122 - 0x7a
    "00000110", --  284 - 0x11c  :    6 - 0x6
    "11111110", --  285 - 0x11d  :  254 - 0xfe
    "11111100", --  286 - 0x11e  :  252 - 0xfc
    "11111100", --  287 - 0x11f  :  252 - 0xfc
    "11111111", --  288 - 0x120  :  255 - 0xff -- Sprite 0x24
    "11001111", --  289 - 0x121  :  207 - 0xcf
    "10000111", --  290 - 0x122  :  135 - 0x87
    "00000111", --  291 - 0x123  :    7 - 0x7
    "00000111", --  292 - 0x124  :    7 - 0x7
    "00001111", --  293 - 0x125  :   15 - 0xf
    "00011111", --  294 - 0x126  :   31 - 0x1f
    "00011111", --  295 - 0x127  :   31 - 0x1f
    "11111000", --  296 - 0x128  :  248 - 0xf8 -- Sprite 0x25
    "11111000", --  297 - 0x129  :  248 - 0xf8
    "11110000", --  298 - 0x12a  :  240 - 0xf0
    "10111000", --  299 - 0x12b  :  184 - 0xb8
    "11111000", --  300 - 0x12c  :  248 - 0xf8
    "11111001", --  301 - 0x12d  :  249 - 0xf9
    "11111011", --  302 - 0x12e  :  251 - 0xfb
    "11111111", --  303 - 0x12f  :  255 - 0xff
    "00011111", --  304 - 0x130  :   31 - 0x1f -- Sprite 0x26
    "11111111", --  305 - 0x131  :  255 - 0xff
    "11111111", --  306 - 0x132  :  255 - 0xff
    "11111111", --  307 - 0x133  :  255 - 0xff
    "11111111", --  308 - 0x134  :  255 - 0xff
    "11111110", --  309 - 0x135  :  254 - 0xfe
    "11000000", --  310 - 0x136  :  192 - 0xc0
    "10000000", --  311 - 0x137  :  128 - 0x80
    "11111111", --  312 - 0x138  :  255 - 0xff -- Sprite 0x27
    "11111111", --  313 - 0x139  :  255 - 0xff
    "11111111", --  314 - 0x13a  :  255 - 0xff
    "00111111", --  315 - 0x13b  :   63 - 0x3f
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00010011", --  320 - 0x140  :   19 - 0x13 -- Sprite 0x28
    "00110011", --  321 - 0x141  :   51 - 0x33
    "00110000", --  322 - 0x142  :   48 - 0x30
    "00011000", --  323 - 0x143  :   24 - 0x18
    "00000100", --  324 - 0x144  :    4 - 0x4
    "00001111", --  325 - 0x145  :   15 - 0xf
    "00011111", --  326 - 0x146  :   31 - 0x1f
    "00011111", --  327 - 0x147  :   31 - 0x1f
    "00000000", --  328 - 0x148  :    0 - 0x0 -- Sprite 0x29
    "00010000", --  329 - 0x149  :   16 - 0x10
    "01111110", --  330 - 0x14a  :  126 - 0x7e
    "00110000", --  331 - 0x14b  :   48 - 0x30
    "11100000", --  332 - 0x14c  :  224 - 0xe0
    "11110000", --  333 - 0x14d  :  240 - 0xf0
    "11110000", --  334 - 0x14e  :  240 - 0xf0
    "11100000", --  335 - 0x14f  :  224 - 0xe0
    "00011111", --  336 - 0x150  :   31 - 0x1f -- Sprite 0x2a
    "00011111", --  337 - 0x151  :   31 - 0x1f
    "00001111", --  338 - 0x152  :   15 - 0xf
    "00001111", --  339 - 0x153  :   15 - 0xf
    "00001111", --  340 - 0x154  :   15 - 0xf
    "00011111", --  341 - 0x155  :   31 - 0x1f
    "00011111", --  342 - 0x156  :   31 - 0x1f
    "00011111", --  343 - 0x157  :   31 - 0x1f
    "11110000", --  344 - 0x158  :  240 - 0xf0 -- Sprite 0x2b
    "11110000", --  345 - 0x159  :  240 - 0xf0
    "11111000", --  346 - 0x15a  :  248 - 0xf8
    "11111000", --  347 - 0x15b  :  248 - 0xf8
    "10111000", --  348 - 0x15c  :  184 - 0xb8
    "11111000", --  349 - 0x15d  :  248 - 0xf8
    "11111000", --  350 - 0x15e  :  248 - 0xf8
    "11111000", --  351 - 0x15f  :  248 - 0xf8
    "00111111", --  352 - 0x160  :   63 - 0x3f -- Sprite 0x2c
    "11111111", --  353 - 0x161  :  255 - 0xff
    "11111111", --  354 - 0x162  :  255 - 0xff
    "11111111", --  355 - 0x163  :  255 - 0xff
    "11110110", --  356 - 0x164  :  246 - 0xf6
    "11000110", --  357 - 0x165  :  198 - 0xc6
    "10000100", --  358 - 0x166  :  132 - 0x84
    "00000000", --  359 - 0x167  :    0 - 0x0
    "11110000", --  360 - 0x168  :  240 - 0xf0 -- Sprite 0x2d
    "11100000", --  361 - 0x169  :  224 - 0xe0
    "10000000", --  362 - 0x16a  :  128 - 0x80
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00011111", --  368 - 0x170  :   31 - 0x1f -- Sprite 0x2e
    "00011111", --  369 - 0x171  :   31 - 0x1f
    "00111111", --  370 - 0x172  :   63 - 0x3f
    "00111111", --  371 - 0x173  :   63 - 0x3f
    "00011111", --  372 - 0x174  :   31 - 0x1f
    "00001111", --  373 - 0x175  :   15 - 0xf
    "00001111", --  374 - 0x176  :   15 - 0xf
    "00011111", --  375 - 0x177  :   31 - 0x1f
    "11110000", --  376 - 0x178  :  240 - 0xf0 -- Sprite 0x2f
    "11110000", --  377 - 0x179  :  240 - 0xf0
    "11111000", --  378 - 0x17a  :  248 - 0xf8
    "11111000", --  379 - 0x17b  :  248 - 0xf8
    "10111000", --  380 - 0x17c  :  184 - 0xb8
    "11111000", --  381 - 0x17d  :  248 - 0xf8
    "11111000", --  382 - 0x17e  :  248 - 0xf8
    "11110000", --  383 - 0x17f  :  240 - 0xf0
    "11100000", --  384 - 0x180  :  224 - 0xe0 -- Sprite 0x30
    "11110000", --  385 - 0x181  :  240 - 0xf0
    "11110000", --  386 - 0x182  :  240 - 0xf0
    "11110000", --  387 - 0x183  :  240 - 0xf0
    "11110000", --  388 - 0x184  :  240 - 0xf0
    "11110000", --  389 - 0x185  :  240 - 0xf0
    "11111000", --  390 - 0x186  :  248 - 0xf8
    "11110000", --  391 - 0x187  :  240 - 0xf0
    "00011111", --  392 - 0x188  :   31 - 0x1f -- Sprite 0x31
    "00011111", --  393 - 0x189  :   31 - 0x1f
    "00011111", --  394 - 0x18a  :   31 - 0x1f
    "00111111", --  395 - 0x18b  :   63 - 0x3f
    "00111110", --  396 - 0x18c  :   62 - 0x3e
    "00111100", --  397 - 0x18d  :   60 - 0x3c
    "00111000", --  398 - 0x18e  :   56 - 0x38
    "00011000", --  399 - 0x18f  :   24 - 0x18
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Sprite 0x32
    "00000011", --  401 - 0x191  :    3 - 0x3
    "00000111", --  402 - 0x192  :    7 - 0x7
    "00000111", --  403 - 0x193  :    7 - 0x7
    "00001010", --  404 - 0x194  :   10 - 0xa
    "00001011", --  405 - 0x195  :   11 - 0xb
    "00001100", --  406 - 0x196  :   12 - 0xc
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00000000", --  408 - 0x198  :    0 - 0x0 -- Sprite 0x33
    "11100000", --  409 - 0x199  :  224 - 0xe0
    "11111100", --  410 - 0x19a  :  252 - 0xfc
    "00100000", --  411 - 0x19b  :   32 - 0x20
    "00100000", --  412 - 0x19c  :   32 - 0x20
    "00010000", --  413 - 0x19d  :   16 - 0x10
    "00111100", --  414 - 0x19e  :   60 - 0x3c
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00000111", --  416 - 0x1a0  :    7 - 0x7 -- Sprite 0x34
    "00000111", --  417 - 0x1a1  :    7 - 0x7
    "00000111", --  418 - 0x1a2  :    7 - 0x7
    "00011111", --  419 - 0x1a3  :   31 - 0x1f
    "00011111", --  420 - 0x1a4  :   31 - 0x1f
    "00111110", --  421 - 0x1a5  :   62 - 0x3e
    "00100001", --  422 - 0x1a6  :   33 - 0x21
    "00000001", --  423 - 0x1a7  :    1 - 0x1
    "11100000", --  424 - 0x1a8  :  224 - 0xe0 -- Sprite 0x35
    "11100000", --  425 - 0x1a9  :  224 - 0xe0
    "11100000", --  426 - 0x1aa  :  224 - 0xe0
    "11110000", --  427 - 0x1ab  :  240 - 0xf0
    "11110000", --  428 - 0x1ac  :  240 - 0xf0
    "11100000", --  429 - 0x1ad  :  224 - 0xe0
    "11000000", --  430 - 0x1ae  :  192 - 0xc0
    "11100000", --  431 - 0x1af  :  224 - 0xe0
    "00000111", --  432 - 0x1b0  :    7 - 0x7 -- Sprite 0x36
    "00001111", --  433 - 0x1b1  :   15 - 0xf
    "00001110", --  434 - 0x1b2  :   14 - 0xe
    "00010100", --  435 - 0x1b3  :   20 - 0x14
    "00010110", --  436 - 0x1b4  :   22 - 0x16
    "00011000", --  437 - 0x1b5  :   24 - 0x18
    "00000000", --  438 - 0x1b6  :    0 - 0x0
    "00111111", --  439 - 0x1b7  :   63 - 0x3f
    "11000000", --  440 - 0x1b8  :  192 - 0xc0 -- Sprite 0x37
    "11111000", --  441 - 0x1b9  :  248 - 0xf8
    "01000000", --  442 - 0x1ba  :   64 - 0x40
    "01000000", --  443 - 0x1bb  :   64 - 0x40
    "00100000", --  444 - 0x1bc  :   32 - 0x20
    "01111000", --  445 - 0x1bd  :  120 - 0x78
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "11000000", --  447 - 0x1bf  :  192 - 0xc0
    "00111111", --  448 - 0x1c0  :   63 - 0x3f -- Sprite 0x38
    "00001110", --  449 - 0x1c1  :   14 - 0xe
    "00001111", --  450 - 0x1c2  :   15 - 0xf
    "00011111", --  451 - 0x1c3  :   31 - 0x1f
    "00111111", --  452 - 0x1c4  :   63 - 0x3f
    "01111100", --  453 - 0x1c5  :  124 - 0x7c
    "01110000", --  454 - 0x1c6  :  112 - 0x70
    "00111000", --  455 - 0x1c7  :   56 - 0x38
    "11110000", --  456 - 0x1c8  :  240 - 0xf0 -- Sprite 0x39
    "11111000", --  457 - 0x1c9  :  248 - 0xf8
    "11100100", --  458 - 0x1ca  :  228 - 0xe4
    "11111100", --  459 - 0x1cb  :  252 - 0xfc
    "11111100", --  460 - 0x1cc  :  252 - 0xfc
    "01111100", --  461 - 0x1cd  :  124 - 0x7c
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000111", --  464 - 0x1d0  :    7 - 0x7 -- Sprite 0x3a
    "00001111", --  465 - 0x1d1  :   15 - 0xf
    "00001110", --  466 - 0x1d2  :   14 - 0xe
    "00010100", --  467 - 0x1d3  :   20 - 0x14
    "00010110", --  468 - 0x1d4  :   22 - 0x16
    "00011000", --  469 - 0x1d5  :   24 - 0x18
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00001111", --  471 - 0x1d7  :   15 - 0xf
    "00011111", --  472 - 0x1d8  :   31 - 0x1f -- Sprite 0x3b
    "00011111", --  473 - 0x1d9  :   31 - 0x1f
    "00011111", --  474 - 0x1da  :   31 - 0x1f
    "00011100", --  475 - 0x1db  :   28 - 0x1c
    "00001100", --  476 - 0x1dc  :   12 - 0xc
    "00000111", --  477 - 0x1dd  :    7 - 0x7
    "00000111", --  478 - 0x1de  :    7 - 0x7
    "00000111", --  479 - 0x1df  :    7 - 0x7
    "11100000", --  480 - 0x1e0  :  224 - 0xe0 -- Sprite 0x3c
    "01100000", --  481 - 0x1e1  :   96 - 0x60
    "11110000", --  482 - 0x1e2  :  240 - 0xf0
    "01110000", --  483 - 0x1e3  :  112 - 0x70
    "11100000", --  484 - 0x1e4  :  224 - 0xe0
    "11100000", --  485 - 0x1e5  :  224 - 0xe0
    "11110000", --  486 - 0x1e6  :  240 - 0xf0
    "10000000", --  487 - 0x1e7  :  128 - 0x80
    "00000111", --  488 - 0x1e8  :    7 - 0x7 -- Sprite 0x3d
    "00011111", --  489 - 0x1e9  :   31 - 0x1f
    "00111111", --  490 - 0x1ea  :   63 - 0x3f
    "00010010", --  491 - 0x1eb  :   18 - 0x12
    "00010011", --  492 - 0x1ec  :   19 - 0x13
    "00001000", --  493 - 0x1ed  :    8 - 0x8
    "00011111", --  494 - 0x1ee  :   31 - 0x1f
    "00110001", --  495 - 0x1ef  :   49 - 0x31
    "11000000", --  496 - 0x1f0  :  192 - 0xc0 -- Sprite 0x3e
    "11110000", --  497 - 0x1f1  :  240 - 0xf0
    "01000000", --  498 - 0x1f2  :   64 - 0x40
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00110000", --  500 - 0x1f4  :   48 - 0x30
    "00011000", --  501 - 0x1f5  :   24 - 0x18
    "11000000", --  502 - 0x1f6  :  192 - 0xc0
    "11111000", --  503 - 0x1f7  :  248 - 0xf8
    "00110001", --  504 - 0x1f8  :   49 - 0x31 -- Sprite 0x3f
    "00111001", --  505 - 0x1f9  :   57 - 0x39
    "00011111", --  506 - 0x1fa  :   31 - 0x1f
    "00011111", --  507 - 0x1fb  :   31 - 0x1f
    "00001111", --  508 - 0x1fc  :   15 - 0xf
    "01011111", --  509 - 0x1fd  :   95 - 0x5f
    "01111110", --  510 - 0x1fe  :  126 - 0x7e
    "00111100", --  511 - 0x1ff  :   60 - 0x3c
    "11111000", --  512 - 0x200  :  248 - 0xf8 -- Sprite 0x40
    "11111000", --  513 - 0x201  :  248 - 0xf8
    "11110000", --  514 - 0x202  :  240 - 0xf0
    "11100000", --  515 - 0x203  :  224 - 0xe0
    "11100000", --  516 - 0x204  :  224 - 0xe0
    "11000000", --  517 - 0x205  :  192 - 0xc0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0 -- Sprite 0x41
    "11100000", --  521 - 0x209  :  224 - 0xe0
    "11111100", --  522 - 0x20a  :  252 - 0xfc
    "00100111", --  523 - 0x20b  :   39 - 0x27
    "00100111", --  524 - 0x20c  :   39 - 0x27
    "00010001", --  525 - 0x20d  :   17 - 0x11
    "00111110", --  526 - 0x20e  :   62 - 0x3e
    "00000100", --  527 - 0x20f  :    4 - 0x4
    "00111111", --  528 - 0x210  :   63 - 0x3f -- Sprite 0x42
    "01111111", --  529 - 0x211  :  127 - 0x7f
    "00111111", --  530 - 0x212  :   63 - 0x3f
    "00001111", --  531 - 0x213  :   15 - 0xf
    "00011111", --  532 - 0x214  :   31 - 0x1f
    "00111111", --  533 - 0x215  :   63 - 0x3f
    "01111111", --  534 - 0x216  :  127 - 0x7f
    "01001111", --  535 - 0x217  :   79 - 0x4f
    "11111000", --  536 - 0x218  :  248 - 0xf8 -- Sprite 0x43
    "11111001", --  537 - 0x219  :  249 - 0xf9
    "11111001", --  538 - 0x21a  :  249 - 0xf9
    "10110111", --  539 - 0x21b  :  183 - 0xb7
    "11111111", --  540 - 0x21c  :  255 - 0xff
    "11111111", --  541 - 0x21d  :  255 - 0xff
    "11100000", --  542 - 0x21e  :  224 - 0xe0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000111", --  544 - 0x220  :    7 - 0x7 -- Sprite 0x44
    "00000111", --  545 - 0x221  :    7 - 0x7
    "00001111", --  546 - 0x222  :   15 - 0xf
    "00111111", --  547 - 0x223  :   63 - 0x3f
    "00111111", --  548 - 0x224  :   63 - 0x3f
    "00111111", --  549 - 0x225  :   63 - 0x3f
    "00100110", --  550 - 0x226  :   38 - 0x26
    "00000100", --  551 - 0x227  :    4 - 0x4
    "11110000", --  552 - 0x228  :  240 - 0xf0 -- Sprite 0x45
    "11110000", --  553 - 0x229  :  240 - 0xf0
    "11110000", --  554 - 0x22a  :  240 - 0xf0
    "11100000", --  555 - 0x22b  :  224 - 0xe0
    "11000000", --  556 - 0x22c  :  192 - 0xc0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000111", --  560 - 0x230  :    7 - 0x7 -- Sprite 0x46
    "00000111", --  561 - 0x231  :    7 - 0x7
    "00001111", --  562 - 0x232  :   15 - 0xf
    "00011111", --  563 - 0x233  :   31 - 0x1f
    "00111111", --  564 - 0x234  :   63 - 0x3f
    "00001111", --  565 - 0x235  :   15 - 0xf
    "00011100", --  566 - 0x236  :   28 - 0x1c
    "00011000", --  567 - 0x237  :   24 - 0x18
    "11100000", --  568 - 0x238  :  224 - 0xe0 -- Sprite 0x47
    "11100000", --  569 - 0x239  :  224 - 0xe0
    "11100000", --  570 - 0x23a  :  224 - 0xe0
    "11100000", --  571 - 0x23b  :  224 - 0xe0
    "11000000", --  572 - 0x23c  :  192 - 0xc0
    "10000000", --  573 - 0x23d  :  128 - 0x80
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000111", --  576 - 0x240  :    7 - 0x7 -- Sprite 0x48
    "00001111", --  577 - 0x241  :   15 - 0xf
    "00011111", --  578 - 0x242  :   31 - 0x1f
    "00001111", --  579 - 0x243  :   15 - 0xf
    "00111111", --  580 - 0x244  :   63 - 0x3f
    "00001111", --  581 - 0x245  :   15 - 0xf
    "00011100", --  582 - 0x246  :   28 - 0x1c
    "00011000", --  583 - 0x247  :   24 - 0x18
    "11100000", --  584 - 0x248  :  224 - 0xe0 -- Sprite 0x49
    "11100000", --  585 - 0x249  :  224 - 0xe0
    "11100000", --  586 - 0x24a  :  224 - 0xe0
    "01000000", --  587 - 0x24b  :   64 - 0x40
    "11000000", --  588 - 0x24c  :  192 - 0xc0
    "10000000", --  589 - 0x24d  :  128 - 0x80
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "01111111", --  592 - 0x250  :  127 - 0x7f -- Sprite 0x4a
    "11111111", --  593 - 0x251  :  255 - 0xff
    "11111111", --  594 - 0x252  :  255 - 0xff
    "11111011", --  595 - 0x253  :  251 - 0xfb
    "00001111", --  596 - 0x254  :   15 - 0xf
    "00001111", --  597 - 0x255  :   15 - 0xf
    "00001111", --  598 - 0x256  :   15 - 0xf
    "00011111", --  599 - 0x257  :   31 - 0x1f
    "00111111", --  600 - 0x258  :   63 - 0x3f -- Sprite 0x4b
    "01111110", --  601 - 0x259  :  126 - 0x7e
    "01111100", --  602 - 0x25a  :  124 - 0x7c
    "01111100", --  603 - 0x25b  :  124 - 0x7c
    "00111100", --  604 - 0x25c  :   60 - 0x3c
    "00111100", --  605 - 0x25d  :   60 - 0x3c
    "11111100", --  606 - 0x25e  :  252 - 0xfc
    "11111100", --  607 - 0x25f  :  252 - 0xfc
    "01100000", --  608 - 0x260  :   96 - 0x60 -- Sprite 0x4c
    "01110000", --  609 - 0x261  :  112 - 0x70
    "00011000", --  610 - 0x262  :   24 - 0x18
    "00001000", --  611 - 0x263  :    8 - 0x8
    "00001111", --  612 - 0x264  :   15 - 0xf
    "00011111", --  613 - 0x265  :   31 - 0x1f
    "00111111", --  614 - 0x266  :   63 - 0x3f
    "01111111", --  615 - 0x267  :  127 - 0x7f
    "11111100", --  616 - 0x268  :  252 - 0xfc -- Sprite 0x4d
    "01111100", --  617 - 0x269  :  124 - 0x7c
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00100000", --  619 - 0x26b  :   32 - 0x20
    "11110000", --  620 - 0x26c  :  240 - 0xf0
    "11111000", --  621 - 0x26d  :  248 - 0xf8
    "11111100", --  622 - 0x26e  :  252 - 0xfc
    "11111110", --  623 - 0x26f  :  254 - 0xfe
    "00001011", --  624 - 0x270  :   11 - 0xb -- Sprite 0x4e
    "00001111", --  625 - 0x271  :   15 - 0xf
    "00011111", --  626 - 0x272  :   31 - 0x1f
    "00011110", --  627 - 0x273  :   30 - 0x1e
    "00111100", --  628 - 0x274  :   60 - 0x3c
    "00111100", --  629 - 0x275  :   60 - 0x3c
    "00111100", --  630 - 0x276  :   60 - 0x3c
    "01111100", --  631 - 0x277  :  124 - 0x7c
    "00011111", --  632 - 0x278  :   31 - 0x1f -- Sprite 0x4f
    "00111111", --  633 - 0x279  :   63 - 0x3f
    "00001101", --  634 - 0x27a  :   13 - 0xd
    "00000111", --  635 - 0x27b  :    7 - 0x7
    "00001111", --  636 - 0x27c  :   15 - 0xf
    "00001110", --  637 - 0x27d  :   14 - 0xe
    "00011100", --  638 - 0x27e  :   28 - 0x1c
    "00111100", --  639 - 0x27f  :   60 - 0x3c
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x50
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Sprite 0x51
    "00000111", --  649 - 0x289  :    7 - 0x7
    "00011111", --  650 - 0x28a  :   31 - 0x1f
    "11111111", --  651 - 0x28b  :  255 - 0xff
    "00000111", --  652 - 0x28c  :    7 - 0x7
    "00011111", --  653 - 0x28d  :   31 - 0x1f
    "00001111", --  654 - 0x28e  :   15 - 0xf
    "00000110", --  655 - 0x28f  :    6 - 0x6
    "00111111", --  656 - 0x290  :   63 - 0x3f -- Sprite 0x52
    "11111111", --  657 - 0x291  :  255 - 0xff
    "11111111", --  658 - 0x292  :  255 - 0xff
    "11111111", --  659 - 0x293  :  255 - 0xff
    "11111111", --  660 - 0x294  :  255 - 0xff
    "11111111", --  661 - 0x295  :  255 - 0xff
    "11111011", --  662 - 0x296  :  251 - 0xfb
    "01110110", --  663 - 0x297  :  118 - 0x76
    "00100000", --  664 - 0x298  :   32 - 0x20 -- Sprite 0x53
    "11111000", --  665 - 0x299  :  248 - 0xf8
    "11111111", --  666 - 0x29a  :  255 - 0xff
    "11000011", --  667 - 0x29b  :  195 - 0xc3
    "11111101", --  668 - 0x29c  :  253 - 0xfd
    "11111110", --  669 - 0x29d  :  254 - 0xfe
    "11110000", --  670 - 0x29e  :  240 - 0xf0
    "01000000", --  671 - 0x29f  :   64 - 0x40
    "01000000", --  672 - 0x2a0  :   64 - 0x40 -- Sprite 0x54
    "11100000", --  673 - 0x2a1  :  224 - 0xe0
    "01000000", --  674 - 0x2a2  :   64 - 0x40
    "01000000", --  675 - 0x2a3  :   64 - 0x40
    "01000001", --  676 - 0x2a4  :   65 - 0x41
    "01000001", --  677 - 0x2a5  :   65 - 0x41
    "01001111", --  678 - 0x2a6  :   79 - 0x4f
    "01000111", --  679 - 0x2a7  :   71 - 0x47
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- Sprite 0x55
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "11100000", --  686 - 0x2ae  :  224 - 0xe0
    "11000000", --  687 - 0x2af  :  192 - 0xc0
    "01000011", --  688 - 0x2b0  :   67 - 0x43 -- Sprite 0x56
    "01000110", --  689 - 0x2b1  :   70 - 0x46
    "01000100", --  690 - 0x2b2  :   68 - 0x44
    "01000000", --  691 - 0x2b3  :   64 - 0x40
    "01000000", --  692 - 0x2b4  :   64 - 0x40
    "01000000", --  693 - 0x2b5  :   64 - 0x40
    "01000000", --  694 - 0x2b6  :   64 - 0x40
    "01000000", --  695 - 0x2b7  :   64 - 0x40
    "10000000", --  696 - 0x2b8  :  128 - 0x80 -- Sprite 0x57
    "11000000", --  697 - 0x2b9  :  192 - 0xc0
    "01000000", --  698 - 0x2ba  :   64 - 0x40
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00110001", --  704 - 0x2c0  :   49 - 0x31 -- Sprite 0x58
    "00110000", --  705 - 0x2c1  :   48 - 0x30
    "00111000", --  706 - 0x2c2  :   56 - 0x38
    "01111100", --  707 - 0x2c3  :  124 - 0x7c
    "01111111", --  708 - 0x2c4  :  127 - 0x7f
    "11111111", --  709 - 0x2c5  :  255 - 0xff
    "11111111", --  710 - 0x2c6  :  255 - 0xff
    "11111011", --  711 - 0x2c7  :  251 - 0xfb
    "00010000", --  712 - 0x2c8  :   16 - 0x10 -- Sprite 0x59
    "01111110", --  713 - 0x2c9  :  126 - 0x7e
    "00111110", --  714 - 0x2ca  :   62 - 0x3e
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00011110", --  716 - 0x2cc  :   30 - 0x1e
    "11111110", --  717 - 0x2cd  :  254 - 0xfe
    "11111111", --  718 - 0x2ce  :  255 - 0xff
    "11111111", --  719 - 0x2cf  :  255 - 0xff
    "11111111", --  720 - 0x2d0  :  255 - 0xff -- Sprite 0x5a
    "11111111", --  721 - 0x2d1  :  255 - 0xff
    "11100011", --  722 - 0x2d2  :  227 - 0xe3
    "11000011", --  723 - 0x2d3  :  195 - 0xc3
    "10000111", --  724 - 0x2d4  :  135 - 0x87
    "01001000", --  725 - 0x2d5  :   72 - 0x48
    "00111100", --  726 - 0x2d6  :   60 - 0x3c
    "11111100", --  727 - 0x2d7  :  252 - 0xfc
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Sprite 0x5b
    "11111111", --  729 - 0x2d9  :  255 - 0xff
    "11000011", --  730 - 0x2da  :  195 - 0xc3
    "10000011", --  731 - 0x2db  :  131 - 0x83
    "10000011", --  732 - 0x2dc  :  131 - 0x83
    "11111111", --  733 - 0x2dd  :  255 - 0xff
    "11111111", --  734 - 0x2de  :  255 - 0xff
    "11111111", --  735 - 0x2df  :  255 - 0xff
    "00011111", --  736 - 0x2e0  :   31 - 0x1f -- Sprite 0x5c
    "00011111", --  737 - 0x2e1  :   31 - 0x1f
    "00001111", --  738 - 0x2e2  :   15 - 0xf
    "00000111", --  739 - 0x2e3  :    7 - 0x7
    "00000001", --  740 - 0x2e4  :    1 - 0x1
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "11110000", --  744 - 0x2e8  :  240 - 0xf0 -- Sprite 0x5d
    "11111011", --  745 - 0x2e9  :  251 - 0xfb
    "11111111", --  746 - 0x2ea  :  255 - 0xff
    "11111111", --  747 - 0x2eb  :  255 - 0xff
    "11111110", --  748 - 0x2ec  :  254 - 0xfe
    "00111110", --  749 - 0x2ed  :   62 - 0x3e
    "00001100", --  750 - 0x2ee  :   12 - 0xc
    "00000100", --  751 - 0x2ef  :    4 - 0x4
    "00011111", --  752 - 0x2f0  :   31 - 0x1f -- Sprite 0x5e
    "00011111", --  753 - 0x2f1  :   31 - 0x1f
    "00001111", --  754 - 0x2f2  :   15 - 0xf
    "00001111", --  755 - 0x2f3  :   15 - 0xf
    "00000111", --  756 - 0x2f4  :    7 - 0x7
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "11111011", --  760 - 0x2f8  :  251 - 0xfb -- Sprite 0x5f
    "11111111", --  761 - 0x2f9  :  255 - 0xff
    "11111111", --  762 - 0x2fa  :  255 - 0xff
    "11111111", --  763 - 0x2fb  :  255 - 0xff
    "11111111", --  764 - 0x2fc  :  255 - 0xff
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x60
    "00011000", --  769 - 0x301  :   24 - 0x18
    "00111100", --  770 - 0x302  :   60 - 0x3c
    "01111110", --  771 - 0x303  :  126 - 0x7e
    "01101110", --  772 - 0x304  :  110 - 0x6e
    "11011111", --  773 - 0x305  :  223 - 0xdf
    "11011111", --  774 - 0x306  :  223 - 0xdf
    "11011111", --  775 - 0x307  :  223 - 0xdf
    "00000000", --  776 - 0x308  :    0 - 0x0 -- Sprite 0x61
    "00011000", --  777 - 0x309  :   24 - 0x18
    "00011000", --  778 - 0x30a  :   24 - 0x18
    "00111100", --  779 - 0x30b  :   60 - 0x3c
    "00111100", --  780 - 0x30c  :   60 - 0x3c
    "00111100", --  781 - 0x30d  :   60 - 0x3c
    "00111100", --  782 - 0x30e  :   60 - 0x3c
    "00011100", --  783 - 0x30f  :   28 - 0x1c
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Sprite 0x62
    "00001000", --  785 - 0x311  :    8 - 0x8
    "00001000", --  786 - 0x312  :    8 - 0x8
    "00001000", --  787 - 0x313  :    8 - 0x8
    "00001000", --  788 - 0x314  :    8 - 0x8
    "00001000", --  789 - 0x315  :    8 - 0x8
    "00001000", --  790 - 0x316  :    8 - 0x8
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0 -- Sprite 0x63
    "00001000", --  793 - 0x319  :    8 - 0x8
    "00001000", --  794 - 0x31a  :    8 - 0x8
    "00000100", --  795 - 0x31b  :    4 - 0x4
    "00000100", --  796 - 0x31c  :    4 - 0x4
    "00000100", --  797 - 0x31d  :    4 - 0x4
    "00000100", --  798 - 0x31e  :    4 - 0x4
    "00000100", --  799 - 0x31f  :    4 - 0x4
    "00111100", --  800 - 0x320  :   60 - 0x3c -- Sprite 0x64
    "01111110", --  801 - 0x321  :  126 - 0x7e
    "01110111", --  802 - 0x322  :  119 - 0x77
    "11111011", --  803 - 0x323  :  251 - 0xfb
    "10011111", --  804 - 0x324  :  159 - 0x9f
    "01011111", --  805 - 0x325  :   95 - 0x5f
    "10001110", --  806 - 0x326  :  142 - 0x8e
    "00100000", --  807 - 0x327  :   32 - 0x20
    "01011100", --  808 - 0x328  :   92 - 0x5c -- Sprite 0x65
    "00101110", --  809 - 0x329  :   46 - 0x2e
    "10001111", --  810 - 0x32a  :  143 - 0x8f
    "00111111", --  811 - 0x32b  :   63 - 0x3f
    "01111011", --  812 - 0x32c  :  123 - 0x7b
    "01110111", --  813 - 0x32d  :  119 - 0x77
    "01111110", --  814 - 0x32e  :  126 - 0x7e
    "00111100", --  815 - 0x32f  :   60 - 0x3c
    "00010011", --  816 - 0x330  :   19 - 0x13 -- Sprite 0x66
    "01001111", --  817 - 0x331  :   79 - 0x4f
    "00111111", --  818 - 0x332  :   63 - 0x3f
    "10111111", --  819 - 0x333  :  191 - 0xbf
    "00111111", --  820 - 0x334  :   63 - 0x3f
    "01111010", --  821 - 0x335  :  122 - 0x7a
    "11111000", --  822 - 0x336  :  248 - 0xf8
    "11111000", --  823 - 0x337  :  248 - 0xf8
    "00000000", --  824 - 0x338  :    0 - 0x0 -- Sprite 0x67
    "00001000", --  825 - 0x339  :    8 - 0x8
    "00000101", --  826 - 0x33a  :    5 - 0x5
    "00001111", --  827 - 0x33b  :   15 - 0xf
    "00101111", --  828 - 0x33c  :   47 - 0x2f
    "00011101", --  829 - 0x33d  :   29 - 0x1d
    "00011100", --  830 - 0x33e  :   28 - 0x1c
    "00111100", --  831 - 0x33f  :   60 - 0x3c
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000010", --  836 - 0x344  :    2 - 0x2
    "00001011", --  837 - 0x345  :   11 - 0xb
    "00000111", --  838 - 0x346  :    7 - 0x7
    "00001111", --  839 - 0x347  :   15 - 0xf
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Sprite 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00001000", --  845 - 0x34d  :    8 - 0x8
    "00000100", --  846 - 0x34e  :    4 - 0x4
    "00000100", --  847 - 0x34f  :    4 - 0x4
    "00000010", --  848 - 0x350  :    2 - 0x2 -- Sprite 0x6a
    "00000010", --  849 - 0x351  :    2 - 0x2
    "00000010", --  850 - 0x352  :    2 - 0x2
    "00000101", --  851 - 0x353  :    5 - 0x5
    "01110001", --  852 - 0x354  :  113 - 0x71
    "01111111", --  853 - 0x355  :  127 - 0x7f
    "01111111", --  854 - 0x356  :  127 - 0x7f
    "01111111", --  855 - 0x357  :  127 - 0x7f
    "00000000", --  856 - 0x358  :    0 - 0x0 -- Sprite 0x6b
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000100", --  863 - 0x35f  :    4 - 0x4
    "00000010", --  864 - 0x360  :    2 - 0x2 -- Sprite 0x6c
    "00000010", --  865 - 0x361  :    2 - 0x2
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000001", --  867 - 0x363  :    1 - 0x1
    "00010011", --  868 - 0x364  :   19 - 0x13
    "00111111", --  869 - 0x365  :   63 - 0x3f
    "01111111", --  870 - 0x366  :  127 - 0x7f
    "01111111", --  871 - 0x367  :  127 - 0x7f
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Sprite 0x6d
    "01000000", --  873 - 0x369  :   64 - 0x40
    "01100000", --  874 - 0x36a  :   96 - 0x60
    "01110000", --  875 - 0x36b  :  112 - 0x70
    "01110011", --  876 - 0x36c  :  115 - 0x73
    "00100111", --  877 - 0x36d  :   39 - 0x27
    "00001111", --  878 - 0x36e  :   15 - 0xf
    "00011111", --  879 - 0x36f  :   31 - 0x1f
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000011", --  884 - 0x374  :    3 - 0x3
    "00000111", --  885 - 0x375  :    7 - 0x7
    "00001111", --  886 - 0x376  :   15 - 0xf
    "00011111", --  887 - 0x377  :   31 - 0x1f
    "01111111", --  888 - 0x378  :  127 - 0x7f -- Sprite 0x6f
    "01111111", --  889 - 0x379  :  127 - 0x7f
    "00111111", --  890 - 0x37a  :   63 - 0x3f
    "00111111", --  891 - 0x37b  :   63 - 0x3f
    "00011111", --  892 - 0x37c  :   31 - 0x1f
    "00011111", --  893 - 0x37d  :   31 - 0x1f
    "00001111", --  894 - 0x37e  :   15 - 0xf
    "00000111", --  895 - 0x37f  :    7 - 0x7
    "00000011", --  896 - 0x380  :    3 - 0x3 -- Sprite 0x70
    "00000111", --  897 - 0x381  :    7 - 0x7
    "00001111", --  898 - 0x382  :   15 - 0xf
    "00011111", --  899 - 0x383  :   31 - 0x1f
    "00111111", --  900 - 0x384  :   63 - 0x3f
    "01110111", --  901 - 0x385  :  119 - 0x77
    "01110111", --  902 - 0x386  :  119 - 0x77
    "11110101", --  903 - 0x387  :  245 - 0xf5
    "11000000", --  904 - 0x388  :  192 - 0xc0 -- Sprite 0x71
    "11100000", --  905 - 0x389  :  224 - 0xe0
    "11110000", --  906 - 0x38a  :  240 - 0xf0
    "11111000", --  907 - 0x38b  :  248 - 0xf8
    "11111100", --  908 - 0x38c  :  252 - 0xfc
    "11101110", --  909 - 0x38d  :  238 - 0xee
    "11101110", --  910 - 0x38e  :  238 - 0xee
    "10101111", --  911 - 0x38f  :  175 - 0xaf
    "11110001", --  912 - 0x390  :  241 - 0xf1 -- Sprite 0x72
    "11111111", --  913 - 0x391  :  255 - 0xff
    "01111000", --  914 - 0x392  :  120 - 0x78
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00011000", --  917 - 0x395  :   24 - 0x18
    "00011100", --  918 - 0x396  :   28 - 0x1c
    "00001110", --  919 - 0x397  :   14 - 0xe
    "10001111", --  920 - 0x398  :  143 - 0x8f -- Sprite 0x73
    "11111111", --  921 - 0x399  :  255 - 0xff
    "00011110", --  922 - 0x39a  :   30 - 0x1e
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00001100", --  924 - 0x39c  :   12 - 0xc
    "00111110", --  925 - 0x39d  :   62 - 0x3e
    "01111110", --  926 - 0x39e  :  126 - 0x7e
    "01111100", --  927 - 0x39f  :  124 - 0x7c
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x74
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- Sprite 0x75
    "00000010", --  937 - 0x3a9  :    2 - 0x2
    "01000001", --  938 - 0x3aa  :   65 - 0x41
    "01000001", --  939 - 0x3ab  :   65 - 0x41
    "01100001", --  940 - 0x3ac  :   97 - 0x61
    "00110011", --  941 - 0x3ad  :   51 - 0x33
    "00000110", --  942 - 0x3ae  :    6 - 0x6
    "00111100", --  943 - 0x3af  :   60 - 0x3c
    "00000011", --  944 - 0x3b0  :    3 - 0x3 -- Sprite 0x76
    "00000111", --  945 - 0x3b1  :    7 - 0x7
    "00001111", --  946 - 0x3b2  :   15 - 0xf
    "00011111", --  947 - 0x3b3  :   31 - 0x1f
    "00111111", --  948 - 0x3b4  :   63 - 0x3f
    "01111111", --  949 - 0x3b5  :  127 - 0x7f
    "01111111", --  950 - 0x3b6  :  127 - 0x7f
    "11111111", --  951 - 0x3b7  :  255 - 0xff
    "11000000", --  952 - 0x3b8  :  192 - 0xc0 -- Sprite 0x77
    "11100000", --  953 - 0x3b9  :  224 - 0xe0
    "11110000", --  954 - 0x3ba  :  240 - 0xf0
    "11111000", --  955 - 0x3bb  :  248 - 0xf8
    "11111100", --  956 - 0x3bc  :  252 - 0xfc
    "11111110", --  957 - 0x3bd  :  254 - 0xfe
    "11111110", --  958 - 0x3be  :  254 - 0xfe
    "11111111", --  959 - 0x3bf  :  255 - 0xff
    "11111111", --  960 - 0x3c0  :  255 - 0xff -- Sprite 0x78
    "11111111", --  961 - 0x3c1  :  255 - 0xff
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "01111000", --  963 - 0x3c3  :  120 - 0x78
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "11111111", --  968 - 0x3c8  :  255 - 0xff -- Sprite 0x79
    "11111111", --  969 - 0x3c9  :  255 - 0xff
    "11111111", --  970 - 0x3ca  :  255 - 0xff
    "00011110", --  971 - 0x3cb  :   30 - 0x1e
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00100000", --  973 - 0x3cd  :   32 - 0x20
    "00100000", --  974 - 0x3ce  :   32 - 0x20
    "01000000", --  975 - 0x3cf  :   64 - 0x40
    "00010110", --  976 - 0x3d0  :   22 - 0x16 -- Sprite 0x7a
    "00011111", --  977 - 0x3d1  :   31 - 0x1f
    "00111111", --  978 - 0x3d2  :   63 - 0x3f
    "01111111", --  979 - 0x3d3  :  127 - 0x7f
    "00111101", --  980 - 0x3d4  :   61 - 0x3d
    "00011101", --  981 - 0x3d5  :   29 - 0x1d
    "00111111", --  982 - 0x3d6  :   63 - 0x3f
    "00011111", --  983 - 0x3d7  :   31 - 0x1f
    "10000000", --  984 - 0x3d8  :  128 - 0x80 -- Sprite 0x7b
    "10000000", --  985 - 0x3d9  :  128 - 0x80
    "11000000", --  986 - 0x3da  :  192 - 0xc0
    "11100000", --  987 - 0x3db  :  224 - 0xe0
    "11110000", --  988 - 0x3dc  :  240 - 0xf0
    "11110000", --  989 - 0x3dd  :  240 - 0xf0
    "11110000", --  990 - 0x3de  :  240 - 0xf0
    "11111000", --  991 - 0x3df  :  248 - 0xf8
    "00111100", --  992 - 0x3e0  :   60 - 0x3c -- Sprite 0x7c
    "11111010", --  993 - 0x3e1  :  250 - 0xfa
    "10110001", --  994 - 0x3e2  :  177 - 0xb1
    "01110010", --  995 - 0x3e3  :  114 - 0x72
    "11110010", --  996 - 0x3e4  :  242 - 0xf2
    "11011011", --  997 - 0x3e5  :  219 - 0xdb
    "11011111", --  998 - 0x3e6  :  223 - 0xdf
    "01011111", --  999 - 0x3e7  :   95 - 0x5f
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Sprite 0x7d
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000001", -- 1003 - 0x3eb  :    1 - 0x1
    "00000001", -- 1004 - 0x3ec  :    1 - 0x1
    "00000001", -- 1005 - 0x3ed  :    1 - 0x1
    "00000110", -- 1006 - 0x3ee  :    6 - 0x6
    "00011110", -- 1007 - 0x3ef  :   30 - 0x1e
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Sprite 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- Sprite 0x7f
    "01111100", -- 1017 - 0x3f9  :  124 - 0x7c
    "11010110", -- 1018 - 0x3fa  :  214 - 0xd6
    "10010010", -- 1019 - 0x3fb  :  146 - 0x92
    "10111010", -- 1020 - 0x3fc  :  186 - 0xba
    "11101110", -- 1021 - 0x3fd  :  238 - 0xee
    "11111110", -- 1022 - 0x3fe  :  254 - 0xfe
    "00111000", -- 1023 - 0x3ff  :   56 - 0x38
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Sprite 0x80
    "00010101", -- 1025 - 0x401  :   21 - 0x15
    "00111111", -- 1026 - 0x402  :   63 - 0x3f
    "01100010", -- 1027 - 0x403  :   98 - 0x62
    "01011111", -- 1028 - 0x404  :   95 - 0x5f
    "11111111", -- 1029 - 0x405  :  255 - 0xff
    "10011111", -- 1030 - 0x406  :  159 - 0x9f
    "01111101", -- 1031 - 0x407  :  125 - 0x7d
    "00000000", -- 1032 - 0x408  :    0 - 0x0 -- Sprite 0x81
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00101111", -- 1040 - 0x410  :   47 - 0x2f -- Sprite 0x82
    "00011110", -- 1041 - 0x411  :   30 - 0x1e
    "00101111", -- 1042 - 0x412  :   47 - 0x2f
    "00101111", -- 1043 - 0x413  :   47 - 0x2f
    "00101111", -- 1044 - 0x414  :   47 - 0x2f
    "00010101", -- 1045 - 0x415  :   21 - 0x15
    "00001101", -- 1046 - 0x416  :   13 - 0xd
    "00001110", -- 1047 - 0x417  :   14 - 0xe
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- Sprite 0x83
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00011100", -- 1056 - 0x420  :   28 - 0x1c -- Sprite 0x84
    "00111110", -- 1057 - 0x421  :   62 - 0x3e
    "01111111", -- 1058 - 0x422  :  127 - 0x7f
    "11111111", -- 1059 - 0x423  :  255 - 0xff
    "11111111", -- 1060 - 0x424  :  255 - 0xff
    "11111110", -- 1061 - 0x425  :  254 - 0xfe
    "01111100", -- 1062 - 0x426  :  124 - 0x7c
    "00111000", -- 1063 - 0x427  :   56 - 0x38
    "00000000", -- 1064 - 0x428  :    0 - 0x0 -- Sprite 0x85
    "11111111", -- 1065 - 0x429  :  255 - 0xff
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "11111111", -- 1067 - 0x42b  :  255 - 0xff
    "11111111", -- 1068 - 0x42c  :  255 - 0xff
    "11111111", -- 1069 - 0x42d  :  255 - 0xff
    "11111111", -- 1070 - 0x42e  :  255 - 0xff
    "11111111", -- 1071 - 0x42f  :  255 - 0xff
    "11111111", -- 1072 - 0x430  :  255 - 0xff -- Sprite 0x86
    "11111111", -- 1073 - 0x431  :  255 - 0xff
    "11111111", -- 1074 - 0x432  :  255 - 0xff
    "11111111", -- 1075 - 0x433  :  255 - 0xff
    "11111111", -- 1076 - 0x434  :  255 - 0xff
    "11111111", -- 1077 - 0x435  :  255 - 0xff
    "11111111", -- 1078 - 0x436  :  255 - 0xff
    "11111111", -- 1079 - 0x437  :  255 - 0xff
    "01111111", -- 1080 - 0x438  :  127 - 0x7f -- Sprite 0x87
    "11111111", -- 1081 - 0x439  :  255 - 0xff
    "11111111", -- 1082 - 0x43a  :  255 - 0xff
    "11111111", -- 1083 - 0x43b  :  255 - 0xff
    "11111111", -- 1084 - 0x43c  :  255 - 0xff
    "11111111", -- 1085 - 0x43d  :  255 - 0xff
    "11111111", -- 1086 - 0x43e  :  255 - 0xff
    "11111111", -- 1087 - 0x43f  :  255 - 0xff
    "01101000", -- 1088 - 0x440  :  104 - 0x68 -- Sprite 0x88
    "01001110", -- 1089 - 0x441  :   78 - 0x4e
    "11100000", -- 1090 - 0x442  :  224 - 0xe0
    "11100000", -- 1091 - 0x443  :  224 - 0xe0
    "11100000", -- 1092 - 0x444  :  224 - 0xe0
    "11110000", -- 1093 - 0x445  :  240 - 0xf0
    "11111000", -- 1094 - 0x446  :  248 - 0xf8
    "11111100", -- 1095 - 0x447  :  252 - 0xfc
    "00111111", -- 1096 - 0x448  :   63 - 0x3f -- Sprite 0x89
    "01011100", -- 1097 - 0x449  :   92 - 0x5c
    "00111001", -- 1098 - 0x44a  :   57 - 0x39
    "00111011", -- 1099 - 0x44b  :   59 - 0x3b
    "10111011", -- 1100 - 0x44c  :  187 - 0xbb
    "11111001", -- 1101 - 0x44d  :  249 - 0xf9
    "11111100", -- 1102 - 0x44e  :  252 - 0xfc
    "11111110", -- 1103 - 0x44f  :  254 - 0xfe
    "11000000", -- 1104 - 0x450  :  192 - 0xc0 -- Sprite 0x8a
    "11110000", -- 1105 - 0x451  :  240 - 0xf0
    "11110000", -- 1106 - 0x452  :  240 - 0xf0
    "11110000", -- 1107 - 0x453  :  240 - 0xf0
    "11110000", -- 1108 - 0x454  :  240 - 0xf0
    "11100000", -- 1109 - 0x455  :  224 - 0xe0
    "11000000", -- 1110 - 0x456  :  192 - 0xc0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "11111110", -- 1112 - 0x458  :  254 - 0xfe -- Sprite 0x8b
    "11111100", -- 1113 - 0x459  :  252 - 0xfc
    "01100001", -- 1114 - 0x45a  :   97 - 0x61
    "00001111", -- 1115 - 0x45b  :   15 - 0xf
    "11111111", -- 1116 - 0x45c  :  255 - 0xff
    "11111110", -- 1117 - 0x45d  :  254 - 0xfe
    "11110000", -- 1118 - 0x45e  :  240 - 0xf0
    "11100000", -- 1119 - 0x45f  :  224 - 0xe0
    "01101110", -- 1120 - 0x460  :  110 - 0x6e -- Sprite 0x8c
    "01000000", -- 1121 - 0x461  :   64 - 0x40
    "11100000", -- 1122 - 0x462  :  224 - 0xe0
    "11100000", -- 1123 - 0x463  :  224 - 0xe0
    "11100000", -- 1124 - 0x464  :  224 - 0xe0
    "11100000", -- 1125 - 0x465  :  224 - 0xe0
    "11100000", -- 1126 - 0x466  :  224 - 0xe0
    "11000000", -- 1127 - 0x467  :  192 - 0xc0
    "00000001", -- 1128 - 0x468  :    1 - 0x1 -- Sprite 0x8d
    "00000001", -- 1129 - 0x469  :    1 - 0x1
    "00000011", -- 1130 - 0x46a  :    3 - 0x3
    "00000011", -- 1131 - 0x46b  :    3 - 0x3
    "00000111", -- 1132 - 0x46c  :    7 - 0x7
    "01111111", -- 1133 - 0x46d  :  127 - 0x7f
    "01111111", -- 1134 - 0x46e  :  127 - 0x7f
    "00111111", -- 1135 - 0x46f  :   63 - 0x3f
    "00000110", -- 1136 - 0x470  :    6 - 0x6 -- Sprite 0x8e
    "00000111", -- 1137 - 0x471  :    7 - 0x7
    "00111111", -- 1138 - 0x472  :   63 - 0x3f
    "00111100", -- 1139 - 0x473  :   60 - 0x3c
    "00011001", -- 1140 - 0x474  :   25 - 0x19
    "01111011", -- 1141 - 0x475  :  123 - 0x7b
    "01111111", -- 1142 - 0x476  :  127 - 0x7f
    "00111111", -- 1143 - 0x477  :   63 - 0x3f
    "00111111", -- 1144 - 0x478  :   63 - 0x3f -- Sprite 0x8f
    "01111111", -- 1145 - 0x479  :  127 - 0x7f
    "01111111", -- 1146 - 0x47a  :  127 - 0x7f
    "00011111", -- 1147 - 0x47b  :   31 - 0x1f
    "00111111", -- 1148 - 0x47c  :   63 - 0x3f
    "00111111", -- 1149 - 0x47d  :   63 - 0x3f
    "00000111", -- 1150 - 0x47e  :    7 - 0x7
    "00000110", -- 1151 - 0x47f  :    6 - 0x6
    "00000011", -- 1152 - 0x480  :    3 - 0x3 -- Sprite 0x90
    "00000111", -- 1153 - 0x481  :    7 - 0x7
    "00001111", -- 1154 - 0x482  :   15 - 0xf
    "00001111", -- 1155 - 0x483  :   15 - 0xf
    "00001111", -- 1156 - 0x484  :   15 - 0xf
    "00001111", -- 1157 - 0x485  :   15 - 0xf
    "00000111", -- 1158 - 0x486  :    7 - 0x7
    "00000011", -- 1159 - 0x487  :    3 - 0x3
    "11111000", -- 1160 - 0x488  :  248 - 0xf8 -- Sprite 0x91
    "11111000", -- 1161 - 0x489  :  248 - 0xf8
    "11111000", -- 1162 - 0x48a  :  248 - 0xf8
    "10100000", -- 1163 - 0x48b  :  160 - 0xa0
    "11100001", -- 1164 - 0x48c  :  225 - 0xe1
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "11111111", -- 1166 - 0x48e  :  255 - 0xff
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "00001111", -- 1168 - 0x490  :   15 - 0xf -- Sprite 0x92
    "00001111", -- 1169 - 0x491  :   15 - 0xf
    "00001111", -- 1170 - 0x492  :   15 - 0xf
    "00011111", -- 1171 - 0x493  :   31 - 0x1f
    "00011111", -- 1172 - 0x494  :   31 - 0x1f
    "00011111", -- 1173 - 0x495  :   31 - 0x1f
    "00001111", -- 1174 - 0x496  :   15 - 0xf
    "00000111", -- 1175 - 0x497  :    7 - 0x7
    "11100000", -- 1176 - 0x498  :  224 - 0xe0 -- Sprite 0x93
    "11111000", -- 1177 - 0x499  :  248 - 0xf8
    "11111000", -- 1178 - 0x49a  :  248 - 0xf8
    "11111000", -- 1179 - 0x49b  :  248 - 0xf8
    "11111111", -- 1180 - 0x49c  :  255 - 0xff
    "11111110", -- 1181 - 0x49d  :  254 - 0xfe
    "11110000", -- 1182 - 0x49e  :  240 - 0xf0
    "11000000", -- 1183 - 0x49f  :  192 - 0xc0
    "00000001", -- 1184 - 0x4a0  :    1 - 0x1 -- Sprite 0x94
    "00001111", -- 1185 - 0x4a1  :   15 - 0xf
    "00001111", -- 1186 - 0x4a2  :   15 - 0xf
    "00011111", -- 1187 - 0x4a3  :   31 - 0x1f
    "00111001", -- 1188 - 0x4a4  :   57 - 0x39
    "00110011", -- 1189 - 0x4a5  :   51 - 0x33
    "00110111", -- 1190 - 0x4a6  :   55 - 0x37
    "01111111", -- 1191 - 0x4a7  :  127 - 0x7f
    "01111111", -- 1192 - 0x4a8  :  127 - 0x7f -- Sprite 0x95
    "00111111", -- 1193 - 0x4a9  :   63 - 0x3f
    "00111111", -- 1194 - 0x4aa  :   63 - 0x3f
    "00111111", -- 1195 - 0x4ab  :   63 - 0x3f
    "00011111", -- 1196 - 0x4ac  :   31 - 0x1f
    "00001111", -- 1197 - 0x4ad  :   15 - 0xf
    "00001111", -- 1198 - 0x4ae  :   15 - 0xf
    "00000001", -- 1199 - 0x4af  :    1 - 0x1
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0 -- Sprite 0x96
    "00000000", -- 1201 - 0x4b1  :    0 - 0x0
    "00000011", -- 1202 - 0x4b2  :    3 - 0x3
    "00000011", -- 1203 - 0x4b3  :    3 - 0x3
    "01000111", -- 1204 - 0x4b4  :   71 - 0x47
    "01100111", -- 1205 - 0x4b5  :  103 - 0x67
    "01110111", -- 1206 - 0x4b6  :  119 - 0x77
    "01110111", -- 1207 - 0x4b7  :  119 - 0x77
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0 -- Sprite 0x97
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "10001000", -- 1212 - 0x4bc  :  136 - 0x88
    "10011000", -- 1213 - 0x4bd  :  152 - 0x98
    "11111000", -- 1214 - 0x4be  :  248 - 0xf8
    "11110000", -- 1215 - 0x4bf  :  240 - 0xf0
    "01111110", -- 1216 - 0x4c0  :  126 - 0x7e -- Sprite 0x98
    "01111111", -- 1217 - 0x4c1  :  127 - 0x7f
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "00011111", -- 1219 - 0x4c3  :   31 - 0x1f
    "00000111", -- 1220 - 0x4c4  :    7 - 0x7
    "00110000", -- 1221 - 0x4c5  :   48 - 0x30
    "00011100", -- 1222 - 0x4c6  :   28 - 0x1c
    "00001100", -- 1223 - 0x4c7  :   12 - 0xc
    "01111110", -- 1224 - 0x4c8  :  126 - 0x7e -- Sprite 0x99
    "00111000", -- 1225 - 0x4c9  :   56 - 0x38
    "11110110", -- 1226 - 0x4ca  :  246 - 0xf6
    "11101101", -- 1227 - 0x4cb  :  237 - 0xed
    "11011111", -- 1228 - 0x4cc  :  223 - 0xdf
    "00111000", -- 1229 - 0x4cd  :   56 - 0x38
    "01110000", -- 1230 - 0x4ce  :  112 - 0x70
    "01100000", -- 1231 - 0x4cf  :   96 - 0x60
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Sprite 0x9a
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00000011", -- 1235 - 0x4d3  :    3 - 0x3
    "00000011", -- 1236 - 0x4d4  :    3 - 0x3
    "01000111", -- 1237 - 0x4d5  :   71 - 0x47
    "01100111", -- 1238 - 0x4d6  :  103 - 0x67
    "01110111", -- 1239 - 0x4d7  :  119 - 0x77
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0 -- Sprite 0x9b
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "10001000", -- 1245 - 0x4dd  :  136 - 0x88
    "10011000", -- 1246 - 0x4de  :  152 - 0x98
    "11111000", -- 1247 - 0x4df  :  248 - 0xf8
    "01110111", -- 1248 - 0x4e0  :  119 - 0x77 -- Sprite 0x9c
    "01111110", -- 1249 - 0x4e1  :  126 - 0x7e
    "01111111", -- 1250 - 0x4e2  :  127 - 0x7f
    "11111111", -- 1251 - 0x4e3  :  255 - 0xff
    "00011111", -- 1252 - 0x4e4  :   31 - 0x1f
    "00000111", -- 1253 - 0x4e5  :    7 - 0x7
    "01110000", -- 1254 - 0x4e6  :  112 - 0x70
    "11110000", -- 1255 - 0x4e7  :  240 - 0xf0
    "11110000", -- 1256 - 0x4e8  :  240 - 0xf0 -- Sprite 0x9d
    "01111110", -- 1257 - 0x4e9  :  126 - 0x7e
    "00111000", -- 1258 - 0x4ea  :   56 - 0x38
    "11110110", -- 1259 - 0x4eb  :  246 - 0xf6
    "11101101", -- 1260 - 0x4ec  :  237 - 0xed
    "11011111", -- 1261 - 0x4ed  :  223 - 0xdf
    "00111000", -- 1262 - 0x4ee  :   56 - 0x38
    "00111100", -- 1263 - 0x4ef  :   60 - 0x3c
    "00000011", -- 1264 - 0x4f0  :    3 - 0x3 -- Sprite 0x9e
    "00000111", -- 1265 - 0x4f1  :    7 - 0x7
    "00001010", -- 1266 - 0x4f2  :   10 - 0xa
    "00011010", -- 1267 - 0x4f3  :   26 - 0x1a
    "00011100", -- 1268 - 0x4f4  :   28 - 0x1c
    "00011110", -- 1269 - 0x4f5  :   30 - 0x1e
    "00001011", -- 1270 - 0x4f6  :   11 - 0xb
    "00001000", -- 1271 - 0x4f7  :    8 - 0x8
    "00011100", -- 1272 - 0x4f8  :   28 - 0x1c -- Sprite 0x9f
    "00111111", -- 1273 - 0x4f9  :   63 - 0x3f
    "00111111", -- 1274 - 0x4fa  :   63 - 0x3f
    "00111101", -- 1275 - 0x4fb  :   61 - 0x3d
    "00111111", -- 1276 - 0x4fc  :   63 - 0x3f
    "00011111", -- 1277 - 0x4fd  :   31 - 0x1f
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- Sprite 0xa0
    "00000000", -- 1281 - 0x501  :    0 - 0x0
    "00000100", -- 1282 - 0x502  :    4 - 0x4
    "01001100", -- 1283 - 0x503  :   76 - 0x4c
    "01001110", -- 1284 - 0x504  :   78 - 0x4e
    "01001110", -- 1285 - 0x505  :   78 - 0x4e
    "01000110", -- 1286 - 0x506  :   70 - 0x46
    "01101111", -- 1287 - 0x507  :  111 - 0x6f
    "00000000", -- 1288 - 0x508  :    0 - 0x0 -- Sprite 0xa1
    "00011111", -- 1289 - 0x509  :   31 - 0x1f
    "00111111", -- 1290 - 0x50a  :   63 - 0x3f
    "00111111", -- 1291 - 0x50b  :   63 - 0x3f
    "01001111", -- 1292 - 0x50c  :   79 - 0x4f
    "01011111", -- 1293 - 0x50d  :   95 - 0x5f
    "01111111", -- 1294 - 0x50e  :  127 - 0x7f
    "01111111", -- 1295 - 0x50f  :  127 - 0x7f
    "01111111", -- 1296 - 0x510  :  127 - 0x7f -- Sprite 0xa2
    "01100111", -- 1297 - 0x511  :  103 - 0x67
    "10100011", -- 1298 - 0x512  :  163 - 0xa3
    "10110000", -- 1299 - 0x513  :  176 - 0xb0
    "11011000", -- 1300 - 0x514  :  216 - 0xd8
    "11011110", -- 1301 - 0x515  :  222 - 0xde
    "11011100", -- 1302 - 0x516  :  220 - 0xdc
    "11001000", -- 1303 - 0x517  :  200 - 0xc8
    "01111111", -- 1304 - 0x518  :  127 - 0x7f -- Sprite 0xa3
    "01111111", -- 1305 - 0x519  :  127 - 0x7f
    "01111111", -- 1306 - 0x51a  :  127 - 0x7f
    "00011111", -- 1307 - 0x51b  :   31 - 0x1f
    "01000111", -- 1308 - 0x51c  :   71 - 0x47
    "01110000", -- 1309 - 0x51d  :  112 - 0x70
    "01110000", -- 1310 - 0x51e  :  112 - 0x70
    "00111001", -- 1311 - 0x51f  :   57 - 0x39
    "11101000", -- 1312 - 0x520  :  232 - 0xe8 -- Sprite 0xa4
    "11101000", -- 1313 - 0x521  :  232 - 0xe8
    "11100000", -- 1314 - 0x522  :  224 - 0xe0
    "11000000", -- 1315 - 0x523  :  192 - 0xc0
    "00010000", -- 1316 - 0x524  :   16 - 0x10
    "01110000", -- 1317 - 0x525  :  112 - 0x70
    "11100000", -- 1318 - 0x526  :  224 - 0xe0
    "11000000", -- 1319 - 0x527  :  192 - 0xc0
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- Sprite 0xa5
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00100000", -- 1323 - 0x52b  :   32 - 0x20
    "01100110", -- 1324 - 0x52c  :  102 - 0x66
    "01100110", -- 1325 - 0x52d  :  102 - 0x66
    "01100110", -- 1326 - 0x52e  :  102 - 0x66
    "01100010", -- 1327 - 0x52f  :   98 - 0x62
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Sprite 0xa6
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00011111", -- 1330 - 0x532  :   31 - 0x1f
    "00111111", -- 1331 - 0x533  :   63 - 0x3f
    "01111111", -- 1332 - 0x534  :  127 - 0x7f
    "01001111", -- 1333 - 0x535  :   79 - 0x4f
    "01011111", -- 1334 - 0x536  :   95 - 0x5f
    "01111111", -- 1335 - 0x537  :  127 - 0x7f
    "01110111", -- 1336 - 0x538  :  119 - 0x77 -- Sprite 0xa7
    "01111111", -- 1337 - 0x539  :  127 - 0x7f
    "00111111", -- 1338 - 0x53a  :   63 - 0x3f
    "10110111", -- 1339 - 0x53b  :  183 - 0xb7
    "10110011", -- 1340 - 0x53c  :  179 - 0xb3
    "11011011", -- 1341 - 0x53d  :  219 - 0xdb
    "11011010", -- 1342 - 0x53e  :  218 - 0xda
    "11011000", -- 1343 - 0x53f  :  216 - 0xd8
    "01111111", -- 1344 - 0x540  :  127 - 0x7f -- Sprite 0xa8
    "01111111", -- 1345 - 0x541  :  127 - 0x7f
    "01111111", -- 1346 - 0x542  :  127 - 0x7f
    "01111111", -- 1347 - 0x543  :  127 - 0x7f
    "00011111", -- 1348 - 0x544  :   31 - 0x1f
    "00000111", -- 1349 - 0x545  :    7 - 0x7
    "01110000", -- 1350 - 0x546  :  112 - 0x70
    "11110000", -- 1351 - 0x547  :  240 - 0xf0
    "11001100", -- 1352 - 0x548  :  204 - 0xcc -- Sprite 0xa9
    "11101000", -- 1353 - 0x549  :  232 - 0xe8
    "11101000", -- 1354 - 0x54a  :  232 - 0xe8
    "11100000", -- 1355 - 0x54b  :  224 - 0xe0
    "11000000", -- 1356 - 0x54c  :  192 - 0xc0
    "00011000", -- 1357 - 0x54d  :   24 - 0x18
    "01111100", -- 1358 - 0x54e  :  124 - 0x7c
    "00111110", -- 1359 - 0x54f  :   62 - 0x3e
    "00000011", -- 1360 - 0x550  :    3 - 0x3 -- Sprite 0xaa
    "00001111", -- 1361 - 0x551  :   15 - 0xf
    "00011111", -- 1362 - 0x552  :   31 - 0x1f
    "00111111", -- 1363 - 0x553  :   63 - 0x3f
    "00111011", -- 1364 - 0x554  :   59 - 0x3b
    "00111111", -- 1365 - 0x555  :   63 - 0x3f
    "01111111", -- 1366 - 0x556  :  127 - 0x7f
    "01111111", -- 1367 - 0x557  :  127 - 0x7f
    "10000000", -- 1368 - 0x558  :  128 - 0x80 -- Sprite 0xab
    "11110000", -- 1369 - 0x559  :  240 - 0xf0
    "11111000", -- 1370 - 0x55a  :  248 - 0xf8
    "11111100", -- 1371 - 0x55b  :  252 - 0xfc
    "11111110", -- 1372 - 0x55c  :  254 - 0xfe
    "11111110", -- 1373 - 0x55d  :  254 - 0xfe
    "11111111", -- 1374 - 0x55e  :  255 - 0xff
    "11111110", -- 1375 - 0x55f  :  254 - 0xfe
    "01111111", -- 1376 - 0x560  :  127 - 0x7f -- Sprite 0xac
    "01111111", -- 1377 - 0x561  :  127 - 0x7f
    "01111111", -- 1378 - 0x562  :  127 - 0x7f
    "01111111", -- 1379 - 0x563  :  127 - 0x7f
    "11111111", -- 1380 - 0x564  :  255 - 0xff
    "00001111", -- 1381 - 0x565  :   15 - 0xf
    "00000011", -- 1382 - 0x566  :    3 - 0x3
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "11111110", -- 1384 - 0x568  :  254 - 0xfe -- Sprite 0xad
    "11111011", -- 1385 - 0x569  :  251 - 0xfb
    "11111111", -- 1386 - 0x56a  :  255 - 0xff
    "11111111", -- 1387 - 0x56b  :  255 - 0xff
    "11110110", -- 1388 - 0x56c  :  246 - 0xf6
    "11100000", -- 1389 - 0x56d  :  224 - 0xe0
    "11000000", -- 1390 - 0x56e  :  192 - 0xc0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0xae
    "00000011", -- 1393 - 0x571  :    3 - 0x3
    "00001111", -- 1394 - 0x572  :   15 - 0xf
    "00011111", -- 1395 - 0x573  :   31 - 0x1f
    "00111111", -- 1396 - 0x574  :   63 - 0x3f
    "00111011", -- 1397 - 0x575  :   59 - 0x3b
    "00111111", -- 1398 - 0x576  :   63 - 0x3f
    "01111111", -- 1399 - 0x577  :  127 - 0x7f
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Sprite 0xaf
    "11000000", -- 1401 - 0x579  :  192 - 0xc0
    "11110000", -- 1402 - 0x57a  :  240 - 0xf0
    "11111000", -- 1403 - 0x57b  :  248 - 0xf8
    "11111100", -- 1404 - 0x57c  :  252 - 0xfc
    "11111110", -- 1405 - 0x57d  :  254 - 0xfe
    "11111110", -- 1406 - 0x57e  :  254 - 0xfe
    "11111111", -- 1407 - 0x57f  :  255 - 0xff
    "01111111", -- 1408 - 0x580  :  127 - 0x7f -- Sprite 0xb0
    "01111111", -- 1409 - 0x581  :  127 - 0x7f
    "01111111", -- 1410 - 0x582  :  127 - 0x7f
    "01111111", -- 1411 - 0x583  :  127 - 0x7f
    "01111111", -- 1412 - 0x584  :  127 - 0x7f
    "11111111", -- 1413 - 0x585  :  255 - 0xff
    "00001111", -- 1414 - 0x586  :   15 - 0xf
    "00000011", -- 1415 - 0x587  :    3 - 0x3
    "11111110", -- 1416 - 0x588  :  254 - 0xfe -- Sprite 0xb1
    "11111110", -- 1417 - 0x589  :  254 - 0xfe
    "11111011", -- 1418 - 0x58a  :  251 - 0xfb
    "11111111", -- 1419 - 0x58b  :  255 - 0xff
    "11111111", -- 1420 - 0x58c  :  255 - 0xff
    "11110110", -- 1421 - 0x58d  :  246 - 0xf6
    "11100000", -- 1422 - 0x58e  :  224 - 0xe0
    "11000000", -- 1423 - 0x58f  :  192 - 0xc0
    "00000000", -- 1424 - 0x590  :    0 - 0x0 -- Sprite 0xb2
    "00000001", -- 1425 - 0x591  :    1 - 0x1
    "00000001", -- 1426 - 0x592  :    1 - 0x1
    "00000001", -- 1427 - 0x593  :    1 - 0x1
    "00000001", -- 1428 - 0x594  :    1 - 0x1
    "00000000", -- 1429 - 0x595  :    0 - 0x0
    "00000000", -- 1430 - 0x596  :    0 - 0x0
    "00001000", -- 1431 - 0x597  :    8 - 0x8
    "01111000", -- 1432 - 0x598  :  120 - 0x78 -- Sprite 0xb3
    "11110000", -- 1433 - 0x599  :  240 - 0xf0
    "11111000", -- 1434 - 0x59a  :  248 - 0xf8
    "11100100", -- 1435 - 0x59b  :  228 - 0xe4
    "11000000", -- 1436 - 0x59c  :  192 - 0xc0
    "11001010", -- 1437 - 0x59d  :  202 - 0xca
    "11001010", -- 1438 - 0x59e  :  202 - 0xca
    "11000000", -- 1439 - 0x59f  :  192 - 0xc0
    "00001111", -- 1440 - 0x5a0  :   15 - 0xf -- Sprite 0xb4
    "00011111", -- 1441 - 0x5a1  :   31 - 0x1f
    "10011111", -- 1442 - 0x5a2  :  159 - 0x9f
    "11111111", -- 1443 - 0x5a3  :  255 - 0xff
    "11111111", -- 1444 - 0x5a4  :  255 - 0xff
    "01111111", -- 1445 - 0x5a5  :  127 - 0x7f
    "01110100", -- 1446 - 0x5a6  :  116 - 0x74
    "00100000", -- 1447 - 0x5a7  :   32 - 0x20
    "11100100", -- 1448 - 0x5a8  :  228 - 0xe4 -- Sprite 0xb5
    "11111111", -- 1449 - 0x5a9  :  255 - 0xff
    "11111110", -- 1450 - 0x5aa  :  254 - 0xfe
    "11111100", -- 1451 - 0x5ab  :  252 - 0xfc
    "10011100", -- 1452 - 0x5ac  :  156 - 0x9c
    "00011110", -- 1453 - 0x5ad  :   30 - 0x1e
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0xb6
    "00000001", -- 1457 - 0x5b1  :    1 - 0x1
    "00000011", -- 1458 - 0x5b2  :    3 - 0x3
    "00000011", -- 1459 - 0x5b3  :    3 - 0x3
    "00000111", -- 1460 - 0x5b4  :    7 - 0x7
    "00000011", -- 1461 - 0x5b5  :    3 - 0x3
    "00000001", -- 1462 - 0x5b6  :    1 - 0x1
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0 -- Sprite 0xb7
    "01011111", -- 1465 - 0x5b9  :   95 - 0x5f
    "01111111", -- 1466 - 0x5ba  :  127 - 0x7f
    "01111111", -- 1467 - 0x5bb  :  127 - 0x7f
    "00111111", -- 1468 - 0x5bc  :   63 - 0x3f
    "00111111", -- 1469 - 0x5bd  :   63 - 0x3f
    "00010100", -- 1470 - 0x5be  :   20 - 0x14
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "11000000", -- 1472 - 0x5c0  :  192 - 0xc0 -- Sprite 0xb8
    "11100000", -- 1473 - 0x5c1  :  224 - 0xe0
    "11110000", -- 1474 - 0x5c2  :  240 - 0xf0
    "00110000", -- 1475 - 0x5c3  :   48 - 0x30
    "00111000", -- 1476 - 0x5c4  :   56 - 0x38
    "00111100", -- 1477 - 0x5c5  :   60 - 0x3c
    "00111100", -- 1478 - 0x5c6  :   60 - 0x3c
    "11111100", -- 1479 - 0x5c7  :  252 - 0xfc
    "00000111", -- 1480 - 0x5c8  :    7 - 0x7 -- Sprite 0xb9
    "00001111", -- 1481 - 0x5c9  :   15 - 0xf
    "00011111", -- 1482 - 0x5ca  :   31 - 0x1f
    "00100010", -- 1483 - 0x5cb  :   34 - 0x22
    "00100000", -- 1484 - 0x5cc  :   32 - 0x20
    "00100101", -- 1485 - 0x5cd  :   37 - 0x25
    "00100101", -- 1486 - 0x5ce  :   37 - 0x25
    "00011111", -- 1487 - 0x5cf  :   31 - 0x1f
    "11111110", -- 1488 - 0x5d0  :  254 - 0xfe -- Sprite 0xba
    "11111110", -- 1489 - 0x5d1  :  254 - 0xfe
    "01111110", -- 1490 - 0x5d2  :  126 - 0x7e
    "00111010", -- 1491 - 0x5d3  :   58 - 0x3a
    "00000010", -- 1492 - 0x5d4  :    2 - 0x2
    "00000001", -- 1493 - 0x5d5  :    1 - 0x1
    "01000001", -- 1494 - 0x5d6  :   65 - 0x41
    "01000001", -- 1495 - 0x5d7  :   65 - 0x41
    "00011111", -- 1496 - 0x5d8  :   31 - 0x1f -- Sprite 0xbb
    "00111111", -- 1497 - 0x5d9  :   63 - 0x3f
    "01111110", -- 1498 - 0x5da  :  126 - 0x7e
    "01011100", -- 1499 - 0x5db  :   92 - 0x5c
    "01000000", -- 1500 - 0x5dc  :   64 - 0x40
    "10000000", -- 1501 - 0x5dd  :  128 - 0x80
    "10000010", -- 1502 - 0x5de  :  130 - 0x82
    "10000010", -- 1503 - 0x5df  :  130 - 0x82
    "10000010", -- 1504 - 0x5e0  :  130 - 0x82 -- Sprite 0xbc
    "10000000", -- 1505 - 0x5e1  :  128 - 0x80
    "10100000", -- 1506 - 0x5e2  :  160 - 0xa0
    "01000100", -- 1507 - 0x5e3  :   68 - 0x44
    "01000011", -- 1508 - 0x5e4  :   67 - 0x43
    "01000000", -- 1509 - 0x5e5  :   64 - 0x40
    "00100001", -- 1510 - 0x5e6  :   33 - 0x21
    "00011110", -- 1511 - 0x5e7  :   30 - 0x1e
    "00011100", -- 1512 - 0x5e8  :   28 - 0x1c -- Sprite 0xbd
    "00111111", -- 1513 - 0x5e9  :   63 - 0x3f
    "00111110", -- 1514 - 0x5ea  :   62 - 0x3e
    "00111100", -- 1515 - 0x5eb  :   60 - 0x3c
    "01000000", -- 1516 - 0x5ec  :   64 - 0x40
    "10000000", -- 1517 - 0x5ed  :  128 - 0x80
    "10000010", -- 1518 - 0x5ee  :  130 - 0x82
    "10000010", -- 1519 - 0x5ef  :  130 - 0x82
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Sprite 0xbe
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "10000000", -- 1522 - 0x5f2  :  128 - 0x80
    "10000000", -- 1523 - 0x5f3  :  128 - 0x80
    "10010010", -- 1524 - 0x5f4  :  146 - 0x92
    "10011101", -- 1525 - 0x5f5  :  157 - 0x9d
    "11000111", -- 1526 - 0x5f6  :  199 - 0xc7
    "11101111", -- 1527 - 0x5f7  :  239 - 0xef
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Sprite 0xbf
    "00100011", -- 1529 - 0x5f9  :   35 - 0x23
    "00110011", -- 1530 - 0x5fa  :   51 - 0x33
    "00111111", -- 1531 - 0x5fb  :   63 - 0x3f
    "00111111", -- 1532 - 0x5fc  :   63 - 0x3f
    "01111111", -- 1533 - 0x5fd  :  127 - 0x7f
    "01111111", -- 1534 - 0x5fe  :  127 - 0x7f
    "01111111", -- 1535 - 0x5ff  :  127 - 0x7f
    "11111110", -- 1536 - 0x600  :  254 - 0xfe -- Sprite 0xc0
    "11111000", -- 1537 - 0x601  :  248 - 0xf8
    "10100000", -- 1538 - 0x602  :  160 - 0xa0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "10000000", -- 1542 - 0x606  :  128 - 0x80
    "10000000", -- 1543 - 0x607  :  128 - 0x80
    "01111110", -- 1544 - 0x608  :  126 - 0x7e -- Sprite 0xc1
    "01111111", -- 1545 - 0x609  :  127 - 0x7f
    "01111101", -- 1546 - 0x60a  :  125 - 0x7d
    "00111111", -- 1547 - 0x60b  :   63 - 0x3f
    "00011110", -- 1548 - 0x60c  :   30 - 0x1e
    "10001111", -- 1549 - 0x60d  :  143 - 0x8f
    "10001111", -- 1550 - 0x60e  :  143 - 0x8f
    "00011001", -- 1551 - 0x60f  :   25 - 0x19
    "11100000", -- 1552 - 0x610  :  224 - 0xe0 -- Sprite 0xc2
    "00001110", -- 1553 - 0x611  :   14 - 0xe
    "01110011", -- 1554 - 0x612  :  115 - 0x73
    "11110011", -- 1555 - 0x613  :  243 - 0xf3
    "11111001", -- 1556 - 0x614  :  249 - 0xf9
    "11111001", -- 1557 - 0x615  :  249 - 0xf9
    "11111000", -- 1558 - 0x616  :  248 - 0xf8
    "01110000", -- 1559 - 0x617  :  112 - 0x70
    "00001110", -- 1560 - 0x618  :   14 - 0xe -- Sprite 0xc3
    "01100110", -- 1561 - 0x619  :  102 - 0x66
    "11100010", -- 1562 - 0x61a  :  226 - 0xe2
    "11110110", -- 1563 - 0x61b  :  246 - 0xf6
    "11111111", -- 1564 - 0x61c  :  255 - 0xff
    "11111111", -- 1565 - 0x61d  :  255 - 0xff
    "00011111", -- 1566 - 0x61e  :   31 - 0x1f
    "10011000", -- 1567 - 0x61f  :  152 - 0x98
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000100", -- 1571 - 0x623  :    4 - 0x4
    "00001111", -- 1572 - 0x624  :   15 - 0xf
    "00001111", -- 1573 - 0x625  :   15 - 0xf
    "00011111", -- 1574 - 0x626  :   31 - 0x1f
    "00000111", -- 1575 - 0x627  :    7 - 0x7
    "11110011", -- 1576 - 0x628  :  243 - 0xf3 -- Sprite 0xc5
    "11100111", -- 1577 - 0x629  :  231 - 0xe7
    "11101110", -- 1578 - 0x62a  :  238 - 0xee
    "11101100", -- 1579 - 0x62b  :  236 - 0xec
    "11001101", -- 1580 - 0x62c  :  205 - 0xcd
    "11001111", -- 1581 - 0x62d  :  207 - 0xcf
    "11001111", -- 1582 - 0x62e  :  207 - 0xcf
    "11011111", -- 1583 - 0x62f  :  223 - 0xdf
    "00100111", -- 1584 - 0x630  :   39 - 0x27 -- Sprite 0xc6
    "00111111", -- 1585 - 0x631  :   63 - 0x3f
    "00111111", -- 1586 - 0x632  :   63 - 0x3f
    "01111000", -- 1587 - 0x633  :  120 - 0x78
    "00111100", -- 1588 - 0x634  :   60 - 0x3c
    "00011111", -- 1589 - 0x635  :   31 - 0x1f
    "00011111", -- 1590 - 0x636  :   31 - 0x1f
    "01110011", -- 1591 - 0x637  :  115 - 0x73
    "10011111", -- 1592 - 0x638  :  159 - 0x9f -- Sprite 0xc7
    "00111110", -- 1593 - 0x639  :   62 - 0x3e
    "01111100", -- 1594 - 0x63a  :  124 - 0x7c
    "11111100", -- 1595 - 0x63b  :  252 - 0xfc
    "11111000", -- 1596 - 0x63c  :  248 - 0xf8
    "11111000", -- 1597 - 0x63d  :  248 - 0xf8
    "11000000", -- 1598 - 0x63e  :  192 - 0xc0
    "01000000", -- 1599 - 0x63f  :   64 - 0x40
    "01111111", -- 1600 - 0x640  :  127 - 0x7f -- Sprite 0xc8
    "01111110", -- 1601 - 0x641  :  126 - 0x7e
    "01111000", -- 1602 - 0x642  :  120 - 0x78
    "00000001", -- 1603 - 0x643  :    1 - 0x1
    "00000111", -- 1604 - 0x644  :    7 - 0x7
    "00011111", -- 1605 - 0x645  :   31 - 0x1f
    "00111100", -- 1606 - 0x646  :   60 - 0x3c
    "01111100", -- 1607 - 0x647  :  124 - 0x7c
    "11111100", -- 1608 - 0x648  :  252 - 0xfc -- Sprite 0xc9
    "11111000", -- 1609 - 0x649  :  248 - 0xf8
    "10100000", -- 1610 - 0x64a  :  160 - 0xa0
    "11111110", -- 1611 - 0x64b  :  254 - 0xfe
    "11111100", -- 1612 - 0x64c  :  252 - 0xfc
    "11110000", -- 1613 - 0x64d  :  240 - 0xf0
    "10000000", -- 1614 - 0x64e  :  128 - 0x80
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "01111110", -- 1616 - 0x650  :  126 - 0x7e -- Sprite 0xca
    "01111111", -- 1617 - 0x651  :  127 - 0x7f
    "01111111", -- 1618 - 0x652  :  127 - 0x7f
    "00111111", -- 1619 - 0x653  :   63 - 0x3f
    "00011111", -- 1620 - 0x654  :   31 - 0x1f
    "10001111", -- 1621 - 0x655  :  143 - 0x8f
    "10001111", -- 1622 - 0x656  :  143 - 0x8f
    "00011000", -- 1623 - 0x657  :   24 - 0x18
    "10011111", -- 1624 - 0x658  :  159 - 0x9f -- Sprite 0xcb
    "00111110", -- 1625 - 0x659  :   62 - 0x3e
    "01111100", -- 1626 - 0x65a  :  124 - 0x7c
    "11111000", -- 1627 - 0x65b  :  248 - 0xf8
    "11111000", -- 1628 - 0x65c  :  248 - 0xf8
    "00111100", -- 1629 - 0x65d  :   60 - 0x3c
    "00011000", -- 1630 - 0x65e  :   24 - 0x18
    "11111000", -- 1631 - 0x65f  :  248 - 0xf8
    "01111111", -- 1632 - 0x660  :  127 - 0x7f -- Sprite 0xcc
    "01111111", -- 1633 - 0x661  :  127 - 0x7f
    "01111000", -- 1634 - 0x662  :  120 - 0x78
    "00000001", -- 1635 - 0x663  :    1 - 0x1
    "00000111", -- 1636 - 0x664  :    7 - 0x7
    "00010011", -- 1637 - 0x665  :   19 - 0x13
    "11110001", -- 1638 - 0x666  :  241 - 0xf1
    "00000011", -- 1639 - 0x667  :    3 - 0x3
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00011100", -- 1642 - 0x66a  :   28 - 0x1c
    "00011101", -- 1643 - 0x66b  :   29 - 0x1d
    "00011011", -- 1644 - 0x66c  :   27 - 0x1b
    "11000011", -- 1645 - 0x66d  :  195 - 0xc3
    "11100011", -- 1646 - 0x66e  :  227 - 0xe3
    "11100001", -- 1647 - 0x66f  :  225 - 0xe1
    "11100000", -- 1648 - 0x670  :  224 - 0xe0 -- Sprite 0xce
    "11001101", -- 1649 - 0x671  :  205 - 0xcd
    "00011101", -- 1650 - 0x672  :   29 - 0x1d
    "01001111", -- 1651 - 0x673  :   79 - 0x4f
    "11101110", -- 1652 - 0x674  :  238 - 0xee
    "11111111", -- 1653 - 0x675  :  255 - 0xff
    "00111111", -- 1654 - 0x676  :   63 - 0x3f
    "00111111", -- 1655 - 0x677  :   63 - 0x3f
    "00111111", -- 1656 - 0x678  :   63 - 0x3f -- Sprite 0xcf
    "00111111", -- 1657 - 0x679  :   63 - 0x3f
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "01110000", -- 1660 - 0x67c  :  112 - 0x70
    "10111000", -- 1661 - 0x67d  :  184 - 0xb8
    "11111100", -- 1662 - 0x67e  :  252 - 0xfc
    "11111100", -- 1663 - 0x67f  :  252 - 0xfc
    "00000111", -- 1664 - 0x680  :    7 - 0x7 -- Sprite 0xd0
    "00001111", -- 1665 - 0x681  :   15 - 0xf
    "00011111", -- 1666 - 0x682  :   31 - 0x1f
    "00111111", -- 1667 - 0x683  :   63 - 0x3f
    "00111110", -- 1668 - 0x684  :   62 - 0x3e
    "01111100", -- 1669 - 0x685  :  124 - 0x7c
    "01111000", -- 1670 - 0x686  :  120 - 0x78
    "01111000", -- 1671 - 0x687  :  120 - 0x78
    "00111111", -- 1672 - 0x688  :   63 - 0x3f -- Sprite 0xd1
    "01011100", -- 1673 - 0x689  :   92 - 0x5c
    "00111001", -- 1674 - 0x68a  :   57 - 0x39
    "00111011", -- 1675 - 0x68b  :   59 - 0x3b
    "10111111", -- 1676 - 0x68c  :  191 - 0xbf
    "11111111", -- 1677 - 0x68d  :  255 - 0xff
    "11111110", -- 1678 - 0x68e  :  254 - 0xfe
    "11111110", -- 1679 - 0x68f  :  254 - 0xfe
    "11000000", -- 1680 - 0x690  :  192 - 0xc0 -- Sprite 0xd2
    "11000000", -- 1681 - 0x691  :  192 - 0xc0
    "10000000", -- 1682 - 0x692  :  128 - 0x80
    "10000000", -- 1683 - 0x693  :  128 - 0x80
    "10000000", -- 1684 - 0x694  :  128 - 0x80
    "10000000", -- 1685 - 0x695  :  128 - 0x80
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "11111110", -- 1688 - 0x698  :  254 - 0xfe -- Sprite 0xd3
    "11111100", -- 1689 - 0x699  :  252 - 0xfc
    "01100001", -- 1690 - 0x69a  :   97 - 0x61
    "00001111", -- 1691 - 0x69b  :   15 - 0xf
    "01111111", -- 1692 - 0x69c  :  127 - 0x7f
    "00111111", -- 1693 - 0x69d  :   63 - 0x3f
    "00011111", -- 1694 - 0x69e  :   31 - 0x1f
    "00011110", -- 1695 - 0x69f  :   30 - 0x1e
    "11110000", -- 1696 - 0x6a0  :  240 - 0xf0 -- Sprite 0xd4
    "01111000", -- 1697 - 0x6a1  :  120 - 0x78
    "11100100", -- 1698 - 0x6a2  :  228 - 0xe4
    "11001000", -- 1699 - 0x6a3  :  200 - 0xc8
    "11001100", -- 1700 - 0x6a4  :  204 - 0xcc
    "10111110", -- 1701 - 0x6a5  :  190 - 0xbe
    "10111110", -- 1702 - 0x6a6  :  190 - 0xbe
    "00111110", -- 1703 - 0x6a7  :   62 - 0x3e
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0 -- Sprite 0xd5
    "00000001", -- 1705 - 0x6a9  :    1 - 0x1
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000111", -- 1707 - 0x6ab  :    7 - 0x7
    "00000111", -- 1708 - 0x6ac  :    7 - 0x7
    "00000111", -- 1709 - 0x6ad  :    7 - 0x7
    "00000111", -- 1710 - 0x6ae  :    7 - 0x7
    "00011111", -- 1711 - 0x6af  :   31 - 0x1f
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00001111", -- 1714 - 0x6b2  :   15 - 0xf
    "00111111", -- 1715 - 0x6b3  :   63 - 0x3f
    "00111111", -- 1716 - 0x6b4  :   63 - 0x3f
    "00001111", -- 1717 - 0x6b5  :   15 - 0xf
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "01111000", -- 1720 - 0x6b8  :  120 - 0x78 -- Sprite 0xd7
    "01111100", -- 1721 - 0x6b9  :  124 - 0x7c
    "01111110", -- 1722 - 0x6ba  :  126 - 0x7e
    "01111111", -- 1723 - 0x6bb  :  127 - 0x7f
    "00111111", -- 1724 - 0x6bc  :   63 - 0x3f
    "00111111", -- 1725 - 0x6bd  :   63 - 0x3f
    "00011011", -- 1726 - 0x6be  :   27 - 0x1b
    "00001001", -- 1727 - 0x6bf  :    9 - 0x9
    "00001100", -- 1728 - 0x6c0  :   12 - 0xc -- Sprite 0xd8
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000111", -- 1732 - 0x6c4  :    7 - 0x7
    "01111111", -- 1733 - 0x6c5  :  127 - 0x7f
    "01111100", -- 1734 - 0x6c6  :  124 - 0x7c
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "00000001", -- 1736 - 0x6c8  :    1 - 0x1 -- Sprite 0xd9
    "11100001", -- 1737 - 0x6c9  :  225 - 0xe1
    "01110001", -- 1738 - 0x6ca  :  113 - 0x71
    "01111001", -- 1739 - 0x6cb  :  121 - 0x79
    "00111101", -- 1740 - 0x6cc  :   61 - 0x3d
    "00111101", -- 1741 - 0x6cd  :   61 - 0x3d
    "00011111", -- 1742 - 0x6ce  :   31 - 0x1f
    "00000011", -- 1743 - 0x6cf  :    3 - 0x3
    "00111111", -- 1744 - 0x6d0  :   63 - 0x3f -- Sprite 0xda
    "00111111", -- 1745 - 0x6d1  :   63 - 0x3f
    "00011111", -- 1746 - 0x6d2  :   31 - 0x1f
    "00011011", -- 1747 - 0x6d3  :   27 - 0x1b
    "00110110", -- 1748 - 0x6d4  :   54 - 0x36
    "00110000", -- 1749 - 0x6d5  :   48 - 0x30
    "01111111", -- 1750 - 0x6d6  :  127 - 0x7f
    "00111111", -- 1751 - 0x6d7  :   63 - 0x3f
    "11111000", -- 1752 - 0x6d8  :  248 - 0xf8 -- Sprite 0xdb
    "11111000", -- 1753 - 0x6d9  :  248 - 0xf8
    "11111000", -- 1754 - 0x6da  :  248 - 0xf8
    "10111000", -- 1755 - 0x6db  :  184 - 0xb8
    "00011000", -- 1756 - 0x6dc  :   24 - 0x18
    "11011000", -- 1757 - 0x6dd  :  216 - 0xd8
    "11011000", -- 1758 - 0x6de  :  216 - 0xd8
    "10111000", -- 1759 - 0x6df  :  184 - 0xb8
    "00000001", -- 1760 - 0x6e0  :    1 - 0x1 -- Sprite 0xdc
    "00000010", -- 1761 - 0x6e1  :    2 - 0x2
    "00000100", -- 1762 - 0x6e2  :    4 - 0x4
    "00000100", -- 1763 - 0x6e3  :    4 - 0x4
    "00001000", -- 1764 - 0x6e4  :    8 - 0x8
    "00001000", -- 1765 - 0x6e5  :    8 - 0x8
    "00010000", -- 1766 - 0x6e6  :   16 - 0x10
    "00010000", -- 1767 - 0x6e7  :   16 - 0x10
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- Sprite 0xdd
    "00001111", -- 1769 - 0x6e9  :   15 - 0xf
    "00010011", -- 1770 - 0x6ea  :   19 - 0x13
    "00001101", -- 1771 - 0x6eb  :   13 - 0xd
    "00001101", -- 1772 - 0x6ec  :   13 - 0xd
    "00010011", -- 1773 - 0x6ed  :   19 - 0x13
    "00001100", -- 1774 - 0x6ee  :   12 - 0xc
    "00100000", -- 1775 - 0x6ef  :   32 - 0x20
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0 -- Sprite 0xde
    "00100100", -- 1777 - 0x6f1  :   36 - 0x24
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00100100", -- 1779 - 0x6f3  :   36 - 0x24
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "00000100", -- 1781 - 0x6f5  :    4 - 0x4
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "00001111", -- 1784 - 0x6f8  :   15 - 0xf -- Sprite 0xdf
    "01000001", -- 1785 - 0x6f9  :   65 - 0x41
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "10001000", -- 1787 - 0x6fb  :  136 - 0x88
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "01000100", -- 1789 - 0x6fd  :   68 - 0x44
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00111000", -- 1792 - 0x700  :   56 - 0x38 -- Sprite 0xe0
    "01111100", -- 1793 - 0x701  :  124 - 0x7c
    "11111110", -- 1794 - 0x702  :  254 - 0xfe
    "11111110", -- 1795 - 0x703  :  254 - 0xfe
    "00111011", -- 1796 - 0x704  :   59 - 0x3b
    "00000011", -- 1797 - 0x705  :    3 - 0x3
    "00000011", -- 1798 - 0x706  :    3 - 0x3
    "00000011", -- 1799 - 0x707  :    3 - 0x3
    "00000011", -- 1800 - 0x708  :    3 - 0x3 -- Sprite 0xe1
    "00110011", -- 1801 - 0x709  :   51 - 0x33
    "01111011", -- 1802 - 0x70a  :  123 - 0x7b
    "01111111", -- 1803 - 0x70b  :  127 - 0x7f
    "11111111", -- 1804 - 0x70c  :  255 - 0xff
    "11111011", -- 1805 - 0x70d  :  251 - 0xfb
    "00000011", -- 1806 - 0x70e  :    3 - 0x3
    "00000011", -- 1807 - 0x70f  :    3 - 0x3
    "11011100", -- 1808 - 0x710  :  220 - 0xdc -- Sprite 0xe2
    "11000000", -- 1809 - 0x711  :  192 - 0xc0
    "11100000", -- 1810 - 0x712  :  224 - 0xe0
    "11100000", -- 1811 - 0x713  :  224 - 0xe0
    "11100000", -- 1812 - 0x714  :  224 - 0xe0
    "11100000", -- 1813 - 0x715  :  224 - 0xe0
    "11100000", -- 1814 - 0x716  :  224 - 0xe0
    "11000000", -- 1815 - 0x717  :  192 - 0xc0
    "00111111", -- 1816 - 0x718  :   63 - 0x3f -- Sprite 0xe3
    "01011111", -- 1817 - 0x719  :   95 - 0x5f
    "00111111", -- 1818 - 0x71a  :   63 - 0x3f
    "00111111", -- 1819 - 0x71b  :   63 - 0x3f
    "10111011", -- 1820 - 0x71c  :  187 - 0xbb
    "11111000", -- 1821 - 0x71d  :  248 - 0xf8
    "11111110", -- 1822 - 0x71e  :  254 - 0xfe
    "11111110", -- 1823 - 0x71f  :  254 - 0xfe
    "00011111", -- 1824 - 0x720  :   31 - 0x1f -- Sprite 0xe4
    "00001111", -- 1825 - 0x721  :   15 - 0xf
    "00001111", -- 1826 - 0x722  :   15 - 0xf
    "00011111", -- 1827 - 0x723  :   31 - 0x1f
    "00011111", -- 1828 - 0x724  :   31 - 0x1f
    "00011110", -- 1829 - 0x725  :   30 - 0x1e
    "00111000", -- 1830 - 0x726  :   56 - 0x38
    "00110000", -- 1831 - 0x727  :   48 - 0x30
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- Sprite 0xe5
    "00100000", -- 1833 - 0x729  :   32 - 0x20
    "01100000", -- 1834 - 0x72a  :   96 - 0x60
    "01100000", -- 1835 - 0x72b  :   96 - 0x60
    "01110000", -- 1836 - 0x72c  :  112 - 0x70
    "11110000", -- 1837 - 0x72d  :  240 - 0xf0
    "11111000", -- 1838 - 0x72e  :  248 - 0xf8
    "11111000", -- 1839 - 0x72f  :  248 - 0xf8
    "11111000", -- 1840 - 0x730  :  248 - 0xf8 -- Sprite 0xe6
    "11111100", -- 1841 - 0x731  :  252 - 0xfc
    "11111100", -- 1842 - 0x732  :  252 - 0xfc
    "01111110", -- 1843 - 0x733  :  126 - 0x7e
    "01111110", -- 1844 - 0x734  :  126 - 0x7e
    "00111110", -- 1845 - 0x735  :   62 - 0x3e
    "00011111", -- 1846 - 0x736  :   31 - 0x1f
    "00000111", -- 1847 - 0x737  :    7 - 0x7
    "00000000", -- 1848 - 0x738  :    0 - 0x0 -- Sprite 0xe7
    "11000000", -- 1849 - 0x739  :  192 - 0xc0
    "01110000", -- 1850 - 0x73a  :  112 - 0x70
    "10111000", -- 1851 - 0x73b  :  184 - 0xb8
    "11110100", -- 1852 - 0x73c  :  244 - 0xf4
    "11110010", -- 1853 - 0x73d  :  242 - 0xf2
    "11110101", -- 1854 - 0x73e  :  245 - 0xf5
    "01111011", -- 1855 - 0x73f  :  123 - 0x7b
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0xe8
    "11011111", -- 1857 - 0x741  :  223 - 0xdf
    "00010000", -- 1858 - 0x742  :   16 - 0x10
    "11111111", -- 1859 - 0x743  :  255 - 0xff
    "11011111", -- 1860 - 0x744  :  223 - 0xdf
    "11111111", -- 1861 - 0x745  :  255 - 0xff
    "11111111", -- 1862 - 0x746  :  255 - 0xff
    "11111001", -- 1863 - 0x747  :  249 - 0xf9
    "00011111", -- 1864 - 0x748  :   31 - 0x1f -- Sprite 0xe9
    "00011111", -- 1865 - 0x749  :   31 - 0x1f
    "00111110", -- 1866 - 0x74a  :   62 - 0x3e
    "11111100", -- 1867 - 0x74b  :  252 - 0xfc
    "11111000", -- 1868 - 0x74c  :  248 - 0xf8
    "11110000", -- 1869 - 0x74d  :  240 - 0xf0
    "11000000", -- 1870 - 0x74e  :  192 - 0xc0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "11111000", -- 1872 - 0x750  :  248 - 0xf8 -- Sprite 0xea
    "11111100", -- 1873 - 0x751  :  252 - 0xfc
    "11111110", -- 1874 - 0x752  :  254 - 0xfe
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "11111111", -- 1876 - 0x754  :  255 - 0xff
    "11011111", -- 1877 - 0x755  :  223 - 0xdf
    "11011111", -- 1878 - 0x756  :  223 - 0xdf
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "11000001", -- 1880 - 0x758  :  193 - 0xc1 -- Sprite 0xeb
    "11110001", -- 1881 - 0x759  :  241 - 0xf1
    "01111001", -- 1882 - 0x75a  :  121 - 0x79
    "01111101", -- 1883 - 0x75b  :  125 - 0x7d
    "00111101", -- 1884 - 0x75c  :   61 - 0x3d
    "00111111", -- 1885 - 0x75d  :   63 - 0x3f
    "00011111", -- 1886 - 0x75e  :   31 - 0x1f
    "00000011", -- 1887 - 0x75f  :    3 - 0x3
    "00000010", -- 1888 - 0x760  :    2 - 0x2 -- Sprite 0xec
    "00000110", -- 1889 - 0x761  :    6 - 0x6
    "00001110", -- 1890 - 0x762  :   14 - 0xe
    "00001110", -- 1891 - 0x763  :   14 - 0xe
    "00011110", -- 1892 - 0x764  :   30 - 0x1e
    "00011110", -- 1893 - 0x765  :   30 - 0x1e
    "00111110", -- 1894 - 0x766  :   62 - 0x3e
    "00111110", -- 1895 - 0x767  :   62 - 0x3e
    "00111110", -- 1896 - 0x768  :   62 - 0x3e -- Sprite 0xed
    "00111110", -- 1897 - 0x769  :   62 - 0x3e
    "00111110", -- 1898 - 0x76a  :   62 - 0x3e
    "00111110", -- 1899 - 0x76b  :   62 - 0x3e
    "00011110", -- 1900 - 0x76c  :   30 - 0x1e
    "00011110", -- 1901 - 0x76d  :   30 - 0x1e
    "00001110", -- 1902 - 0x76e  :   14 - 0xe
    "00000010", -- 1903 - 0x76f  :    2 - 0x2
    "11000001", -- 1904 - 0x770  :  193 - 0xc1 -- Sprite 0xee
    "11110001", -- 1905 - 0x771  :  241 - 0xf1
    "01111001", -- 1906 - 0x772  :  121 - 0x79
    "01111101", -- 1907 - 0x773  :  125 - 0x7d
    "00111101", -- 1908 - 0x774  :   61 - 0x3d
    "00111111", -- 1909 - 0x775  :   63 - 0x3f
    "00011111", -- 1910 - 0x776  :   31 - 0x1f
    "00000011", -- 1911 - 0x777  :    3 - 0x3
    "01111100", -- 1912 - 0x778  :  124 - 0x7c -- Sprite 0xef
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "11000011", -- 1916 - 0x77c  :  195 - 0xc3
    "01111111", -- 1917 - 0x77d  :  127 - 0x7f
    "00011111", -- 1918 - 0x77e  :   31 - 0x1f
    "00000011", -- 1919 - 0x77f  :    3 - 0x3
    "11111111", -- 1920 - 0x780  :  255 - 0xff -- Sprite 0xf0
    "11111111", -- 1921 - 0x781  :  255 - 0xff
    "01111100", -- 1922 - 0x782  :  124 - 0x7c
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "01111100", -- 1925 - 0x785  :  124 - 0x7c
    "11111111", -- 1926 - 0x786  :  255 - 0xff
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11111111", -- 1928 - 0x788  :  255 - 0xff -- Sprite 0xf1
    "11111111", -- 1929 - 0x789  :  255 - 0xff
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000100", -- 1931 - 0x78b  :    4 - 0x4
    "00001100", -- 1932 - 0x78c  :   12 - 0xc
    "00011000", -- 1933 - 0x78d  :   24 - 0x18
    "00110000", -- 1934 - 0x78e  :   48 - 0x30
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "11111111", -- 1936 - 0x790  :  255 - 0xff -- Sprite 0xf2
    "11111111", -- 1937 - 0x791  :  255 - 0xff
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000100", -- 1939 - 0x793  :    4 - 0x4
    "00000100", -- 1940 - 0x794  :    4 - 0x4
    "00000100", -- 1941 - 0x795  :    4 - 0x4
    "00001000", -- 1942 - 0x796  :    8 - 0x8
    "00001000", -- 1943 - 0x797  :    8 - 0x8
    "00001000", -- 1944 - 0x798  :    8 - 0x8 -- Sprite 0xf3
    "00010000", -- 1945 - 0x799  :   16 - 0x10
    "00010000", -- 1946 - 0x79a  :   16 - 0x10
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00010000", -- 1949 - 0x79d  :   16 - 0x10
    "00010000", -- 1950 - 0x79e  :   16 - 0x10
    "00001000", -- 1951 - 0x79f  :    8 - 0x8
    "01111111", -- 1952 - 0x7a0  :  127 - 0x7f -- Sprite 0xf4
    "00111111", -- 1953 - 0x7a1  :   63 - 0x3f
    "00111111", -- 1954 - 0x7a2  :   63 - 0x3f
    "00111110", -- 1955 - 0x7a3  :   62 - 0x3e
    "00011111", -- 1956 - 0x7a4  :   31 - 0x1f
    "00001111", -- 1957 - 0x7a5  :   15 - 0xf
    "00000011", -- 1958 - 0x7a6  :    3 - 0x3
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000011", -- 1960 - 0x7a8  :    3 - 0x3 -- Sprite 0xf5
    "00001111", -- 1961 - 0x7a9  :   15 - 0xf
    "11111111", -- 1962 - 0x7aa  :  255 - 0xff
    "01111111", -- 1963 - 0x7ab  :  127 - 0x7f
    "01111111", -- 1964 - 0x7ac  :  127 - 0x7f
    "01111111", -- 1965 - 0x7ad  :  127 - 0x7f
    "01111111", -- 1966 - 0x7ae  :  127 - 0x7f
    "01111111", -- 1967 - 0x7af  :  127 - 0x7f
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0xf6
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- Sprite 0xf7
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0xf8
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- Sprite 0xf9
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Sprite 0xfa
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- Sprite 0xfb
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0xfc
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- Sprite 0xfd
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Sprite 0xfe
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Sprite 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "01111100", -- 2045 - 0x7fd  :  124 - 0x7c
    "00111000", -- 2046 - 0x7fe  :   56 - 0x38
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
