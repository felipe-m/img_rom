---   Background Pattern table COLOR PLANE 1
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: nova_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_NOVA_BG_PLN1 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_NOVA_BG_PLN1;

architecture BEHAVIORAL of ROM_PTABLE_NOVA_BG_PLN1 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table COLOR PLANE 1
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Background 0x0
    "01111111", --    1 -  0x1  :  127 - 0x7f
    "01111111", --    2 -  0x2  :  127 - 0x7f
    "01111111", --    3 -  0x3  :  127 - 0x7f
    "01111111", --    4 -  0x4  :  127 - 0x7f
    "01111111", --    5 -  0x5  :  127 - 0x7f
    "01101010", --    6 -  0x6  :  106 - 0x6a
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Background 0x1
    "01111011", --    9 -  0x9  :  123 - 0x7b
    "01110011", --   10 -  0xa  :  115 - 0x73
    "01111011", --   11 -  0xb  :  123 - 0x7b
    "01110011", --   12 -  0xc  :  115 - 0x73
    "01111011", --   13 -  0xd  :  123 - 0x7b
    "01010011", --   14 -  0xe  :   83 - 0x53
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Background 0x2
    "11011110", --   17 - 0x11  :  222 - 0xde
    "10011110", --   18 - 0x12  :  158 - 0x9e
    "11011100", --   19 - 0x13  :  220 - 0xdc
    "10011110", --   20 - 0x14  :  158 - 0x9e
    "11011100", --   21 - 0x15  :  220 - 0xdc
    "10011010", --   22 - 0x16  :  154 - 0x9a
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- Background 0x3
    "11111110", --   25 - 0x19  :  254 - 0xfe
    "11111100", --   26 - 0x1a  :  252 - 0xfc
    "11111110", --   27 - 0x1b  :  254 - 0xfe
    "11111100", --   28 - 0x1c  :  252 - 0xfc
    "11111110", --   29 - 0x1d  :  254 - 0xfe
    "01010100", --   30 - 0x1e  :   84 - 0x54
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Background 0x4
    "01111111", --   33 - 0x21  :  127 - 0x7f
    "01011111", --   34 - 0x22  :   95 - 0x5f
    "01111001", --   35 - 0x23  :  121 - 0x79
    "01111001", --   36 - 0x24  :  121 - 0x79
    "01001001", --   37 - 0x25  :   73 - 0x49
    "01001111", --   38 - 0x26  :   79 - 0x4f
    "01001110", --   39 - 0x27  :   78 - 0x4e
    "01111000", --   40 - 0x28  :  120 - 0x78 -- Background 0x5
    "01110000", --   41 - 0x29  :  112 - 0x70
    "01100000", --   42 - 0x2a  :   96 - 0x60
    "01100000", --   43 - 0x2b  :   96 - 0x60
    "01110001", --   44 - 0x2c  :  113 - 0x71
    "01011111", --   45 - 0x2d  :   95 - 0x5f
    "01111111", --   46 - 0x2e  :  127 - 0x7f
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Background 0x6
    "11111110", --   49 - 0x31  :  254 - 0xfe
    "11111010", --   50 - 0x32  :  250 - 0xfa
    "10011110", --   51 - 0x33  :  158 - 0x9e
    "10011110", --   52 - 0x34  :  158 - 0x9e
    "10010010", --   53 - 0x35  :  146 - 0x92
    "11110010", --   54 - 0x36  :  242 - 0xf2
    "01110010", --   55 - 0x37  :  114 - 0x72
    "00011110", --   56 - 0x38  :   30 - 0x1e -- Background 0x7
    "00001110", --   57 - 0x39  :   14 - 0xe
    "00000110", --   58 - 0x3a  :    6 - 0x6
    "00000110", --   59 - 0x3b  :    6 - 0x6
    "10001110", --   60 - 0x3c  :  142 - 0x8e
    "11111010", --   61 - 0x3d  :  250 - 0xfa
    "11111110", --   62 - 0x3e  :  254 - 0xfe
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Background 0x8
    "01111111", --   65 - 0x41  :  127 - 0x7f
    "01011111", --   66 - 0x42  :   95 - 0x5f
    "01111111", --   67 - 0x43  :  127 - 0x7f
    "01111111", --   68 - 0x44  :  127 - 0x7f
    "01111111", --   69 - 0x45  :  127 - 0x7f
    "01111111", --   70 - 0x46  :  127 - 0x7f
    "01111111", --   71 - 0x47  :  127 - 0x7f
    "01111111", --   72 - 0x48  :  127 - 0x7f -- Background 0x9
    "01111111", --   73 - 0x49  :  127 - 0x7f
    "01111111", --   74 - 0x4a  :  127 - 0x7f
    "01111111", --   75 - 0x4b  :  127 - 0x7f
    "01111111", --   76 - 0x4c  :  127 - 0x7f
    "01011111", --   77 - 0x4d  :   95 - 0x5f
    "01111111", --   78 - 0x4e  :  127 - 0x7f
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Background 0xa
    "11111110", --   81 - 0x51  :  254 - 0xfe
    "11111010", --   82 - 0x52  :  250 - 0xfa
    "11111110", --   83 - 0x53  :  254 - 0xfe
    "11111110", --   84 - 0x54  :  254 - 0xfe
    "11111110", --   85 - 0x55  :  254 - 0xfe
    "11111110", --   86 - 0x56  :  254 - 0xfe
    "11111110", --   87 - 0x57  :  254 - 0xfe
    "11111110", --   88 - 0x58  :  254 - 0xfe -- Background 0xb
    "11111110", --   89 - 0x59  :  254 - 0xfe
    "11111110", --   90 - 0x5a  :  254 - 0xfe
    "11111110", --   91 - 0x5b  :  254 - 0xfe
    "11111110", --   92 - 0x5c  :  254 - 0xfe
    "11111010", --   93 - 0x5d  :  250 - 0xfa
    "11111110", --   94 - 0x5e  :  254 - 0xfe
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Background 0xc
    "00111111", --   97 - 0x61  :   63 - 0x3f
    "01011111", --   98 - 0x62  :   95 - 0x5f
    "01101111", --   99 - 0x63  :  111 - 0x6f
    "01110000", --  100 - 0x64  :  112 - 0x70
    "01110111", --  101 - 0x65  :  119 - 0x77
    "01110111", --  102 - 0x66  :  119 - 0x77
    "01110111", --  103 - 0x67  :  119 - 0x77
    "01110111", --  104 - 0x68  :  119 - 0x77 -- Background 0xd
    "01110111", --  105 - 0x69  :  119 - 0x77
    "01110111", --  106 - 0x6a  :  119 - 0x77
    "01110000", --  107 - 0x6b  :  112 - 0x70
    "01101111", --  108 - 0x6c  :  111 - 0x6f
    "01011111", --  109 - 0x6d  :   95 - 0x5f
    "00010101", --  110 - 0x6e  :   21 - 0x15
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Background 0xe
    "11111100", --  113 - 0x71  :  252 - 0xfc
    "11111000", --  114 - 0x72  :  248 - 0xf8
    "11110110", --  115 - 0x73  :  246 - 0xf6
    "00001100", --  116 - 0x74  :   12 - 0xc
    "11101110", --  117 - 0x75  :  238 - 0xee
    "11101100", --  118 - 0x76  :  236 - 0xec
    "11101110", --  119 - 0x77  :  238 - 0xee
    "11101100", --  120 - 0x78  :  236 - 0xec -- Background 0xf
    "11101110", --  121 - 0x79  :  238 - 0xee
    "11101100", --  122 - 0x7a  :  236 - 0xec
    "00001110", --  123 - 0x7b  :   14 - 0xe
    "11110100", --  124 - 0x7c  :  244 - 0xf4
    "11111010", --  125 - 0x7d  :  250 - 0xfa
    "01010100", --  126 - 0x7e  :   84 - 0x54
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "01100000", --  128 - 0x80  :   96 - 0x60 -- Background 0x10
    "01100000", --  129 - 0x81  :   96 - 0x60
    "01100000", --  130 - 0x82  :   96 - 0x60
    "01101111", --  131 - 0x83  :  111 - 0x6f
    "01101010", --  132 - 0x84  :  106 - 0x6a
    "01100000", --  133 - 0x85  :   96 - 0x60
    "01100000", --  134 - 0x86  :   96 - 0x60
    "01100000", --  135 - 0x87  :   96 - 0x60
    "00000110", --  136 - 0x88  :    6 - 0x6 -- Background 0x11
    "00000100", --  137 - 0x89  :    4 - 0x4
    "00000110", --  138 - 0x8a  :    6 - 0x6
    "11110100", --  139 - 0x8b  :  244 - 0xf4
    "10100110", --  140 - 0x8c  :  166 - 0xa6
    "00000100", --  141 - 0x8d  :    4 - 0x4
    "00000110", --  142 - 0x8e  :    6 - 0x6
    "00000100", --  143 - 0x8f  :    4 - 0x4
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Background 0x12
    "00001000", --  145 - 0x91  :    8 - 0x8
    "00001000", --  146 - 0x92  :    8 - 0x8
    "00011100", --  147 - 0x93  :   28 - 0x1c
    "00011100", --  148 - 0x94  :   28 - 0x1c
    "00111100", --  149 - 0x95  :   60 - 0x3c
    "00111100", --  150 - 0x96  :   60 - 0x3c
    "00111100", --  151 - 0x97  :   60 - 0x3c
    "00111100", --  152 - 0x98  :   60 - 0x3c -- Background 0x13
    "01111110", --  153 - 0x99  :  126 - 0x7e
    "01111110", --  154 - 0x9a  :  126 - 0x7e
    "01111110", --  155 - 0x9b  :  126 - 0x7e
    "01111110", --  156 - 0x9c  :  126 - 0x7e
    "01111110", --  157 - 0x9d  :  126 - 0x7e
    "01111110", --  158 - 0x9e  :  126 - 0x7e
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Background 0x14
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000101", --  162 - 0xa2  :    5 - 0x5
    "00000011", --  163 - 0xa3  :    3 - 0x3
    "00000000", --  164 - 0xa4  :    0 - 0x0
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000010", --  166 - 0xa6  :    2 - 0x2
    "00001111", --  167 - 0xa7  :   15 - 0xf
    "00011100", --  168 - 0xa8  :   28 - 0x1c -- Background 0x15
    "00111010", --  169 - 0xa9  :   58 - 0x3a
    "00111100", --  170 - 0xaa  :   60 - 0x3c
    "00111111", --  171 - 0xab  :   63 - 0x3f
    "00111000", --  172 - 0xac  :   56 - 0x38
    "00011110", --  173 - 0xad  :   30 - 0x1e
    "00001111", --  174 - 0xae  :   15 - 0xf
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Background 0x16
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "01000000", --  178 - 0xb2  :   64 - 0x40
    "11000000", --  179 - 0xb3  :  192 - 0xc0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "10000000", --  181 - 0xb5  :  128 - 0x80
    "11000000", --  182 - 0xb6  :  192 - 0xc0
    "01110000", --  183 - 0xb7  :  112 - 0x70
    "00011000", --  184 - 0xb8  :   24 - 0x18 -- Background 0x17
    "11111100", --  185 - 0xb9  :  252 - 0xfc
    "00111100", --  186 - 0xba  :   60 - 0x3c
    "01011100", --  187 - 0xbb  :   92 - 0x5c
    "00111100", --  188 - 0xbc  :   60 - 0x3c
    "11111000", --  189 - 0xbd  :  248 - 0xf8
    "11110000", --  190 - 0xbe  :  240 - 0xf0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Background 0x18
    "00111111", --  193 - 0xc1  :   63 - 0x3f
    "00111111", --  194 - 0xc2  :   63 - 0x3f
    "01111111", --  195 - 0xc3  :  127 - 0x7f
    "01111111", --  196 - 0xc4  :  127 - 0x7f
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- Background 0x19
    "11111100", --  201 - 0xc9  :  252 - 0xfc
    "11111100", --  202 - 0xca  :  252 - 0xfc
    "11111110", --  203 - 0xcb  :  254 - 0xfe
    "11111110", --  204 - 0xcc  :  254 - 0xfe
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Background 0x1a
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00111111", --  211 - 0xd3  :   63 - 0x3f
    "00111111", --  212 - 0xd4  :   63 - 0x3f
    "01111111", --  213 - 0xd5  :  127 - 0x7f
    "01111111", --  214 - 0xd6  :  127 - 0x7f
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Background 0x1b
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "11111100", --  219 - 0xdb  :  252 - 0xfc
    "11111100", --  220 - 0xdc  :  252 - 0xfc
    "11111110", --  221 - 0xdd  :  254 - 0xfe
    "11111110", --  222 - 0xde  :  254 - 0xfe
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Background 0x1c
    "01111111", --  225 - 0xe1  :  127 - 0x7f
    "01111111", --  226 - 0xe2  :  127 - 0x7f
    "01111111", --  227 - 0xe3  :  127 - 0x7f
    "01100100", --  228 - 0xe4  :  100 - 0x64
    "01011011", --  229 - 0xe5  :   91 - 0x5b
    "01011001", --  230 - 0xe6  :   89 - 0x59
    "01111111", --  231 - 0xe7  :  127 - 0x7f
    "01111111", --  232 - 0xe8  :  127 - 0x7f -- Background 0x1d
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000001", --  234 - 0xea  :    1 - 0x1
    "00000001", --  235 - 0xeb  :    1 - 0x1
    "00000001", --  236 - 0xec  :    1 - 0x1
    "00000001", --  237 - 0xed  :    1 - 0x1
    "00000001", --  238 - 0xee  :    1 - 0x1
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Background 0x1e
    "11111110", --  241 - 0xf1  :  254 - 0xfe
    "11111110", --  242 - 0xf2  :  254 - 0xfe
    "11111110", --  243 - 0xf3  :  254 - 0xfe
    "10111110", --  244 - 0xf4  :  190 - 0xbe
    "00001010", --  245 - 0xf5  :   10 - 0xa
    "11100010", --  246 - 0xf6  :  226 - 0xe2
    "11111110", --  247 - 0xf7  :  254 - 0xfe
    "11111110", --  248 - 0xf8  :  254 - 0xfe -- Background 0x1f
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "10000000", --  250 - 0xfa  :  128 - 0x80
    "10000000", --  251 - 0xfb  :  128 - 0x80
    "10000000", --  252 - 0xfc  :  128 - 0x80
    "10000000", --  253 - 0xfd  :  128 - 0x80
    "10000000", --  254 - 0xfe  :  128 - 0x80
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Background 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Background 0x21
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00000000", --  272 - 0x110  :    0 - 0x0 -- Background 0x22
    "00000000", --  273 - 0x111  :    0 - 0x0
    "00011000", --  274 - 0x112  :   24 - 0x18
    "00010000", --  275 - 0x113  :   16 - 0x10
    "00011010", --  276 - 0x114  :   26 - 0x1a
    "00010001", --  277 - 0x115  :   17 - 0x11
    "00011010", --  278 - 0x116  :   26 - 0x1a
    "00000000", --  279 - 0x117  :    0 - 0x0
    "00000000", --  280 - 0x118  :    0 - 0x0 -- Background 0x23
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00101000", --  283 - 0x11b  :   40 - 0x28
    "10001100", --  284 - 0x11c  :  140 - 0x8c
    "00101000", --  285 - 0x11d  :   40 - 0x28
    "10101100", --  286 - 0x11e  :  172 - 0xac
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Background 0x24
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00011100", --  296 - 0x128  :   28 - 0x1c -- Background 0x25
    "00111001", --  297 - 0x129  :   57 - 0x39
    "00111111", --  298 - 0x12a  :   63 - 0x3f
    "00111110", --  299 - 0x12b  :   62 - 0x3e
    "00111111", --  300 - 0x12c  :   63 - 0x3f
    "00011110", --  301 - 0x12d  :   30 - 0x1e
    "00001111", --  302 - 0x12e  :   15 - 0xf
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Background 0x26
    "00000000", --  305 - 0x131  :    0 - 0x0
    "01000000", --  306 - 0x132  :   64 - 0x40
    "11000000", --  307 - 0x133  :  192 - 0xc0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "10000000", --  309 - 0x135  :  128 - 0x80
    "11000000", --  310 - 0x136  :  192 - 0xc0
    "11110000", --  311 - 0x137  :  240 - 0xf0
    "00111000", --  312 - 0x138  :   56 - 0x38 -- Background 0x27
    "10011100", --  313 - 0x139  :  156 - 0x9c
    "10011100", --  314 - 0x13a  :  156 - 0x9c
    "00111100", --  315 - 0x13b  :   60 - 0x3c
    "11111100", --  316 - 0x13c  :  252 - 0xfc
    "01111000", --  317 - 0x13d  :  120 - 0x78
    "11110000", --  318 - 0x13e  :  240 - 0xf0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Background 0x28
    "00111110", --  321 - 0x141  :   62 - 0x3e
    "01011101", --  322 - 0x142  :   93 - 0x5d
    "01101011", --  323 - 0x143  :  107 - 0x6b
    "01110101", --  324 - 0x144  :  117 - 0x75
    "01110001", --  325 - 0x145  :  113 - 0x71
    "01110101", --  326 - 0x146  :  117 - 0x75
    "01110100", --  327 - 0x147  :  116 - 0x74
    "01110000", --  328 - 0x148  :  112 - 0x70 -- Background 0x29
    "01110111", --  329 - 0x149  :  119 - 0x77
    "01110111", --  330 - 0x14a  :  119 - 0x77
    "01110000", --  331 - 0x14b  :  112 - 0x70
    "01101111", --  332 - 0x14c  :  111 - 0x6f
    "01011111", --  333 - 0x14d  :   95 - 0x5f
    "00010101", --  334 - 0x14e  :   21 - 0x15
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00000000", --  336 - 0x150  :    0 - 0x0 -- Background 0x2a
    "01111100", --  337 - 0x151  :  124 - 0x7c
    "10111000", --  338 - 0x152  :  184 - 0xb8
    "11010110", --  339 - 0x153  :  214 - 0xd6
    "10101100", --  340 - 0x154  :  172 - 0xac
    "10001110", --  341 - 0x155  :  142 - 0x8e
    "10101100", --  342 - 0x156  :  172 - 0xac
    "00101110", --  343 - 0x157  :   46 - 0x2e
    "00001100", --  344 - 0x158  :   12 - 0xc -- Background 0x2b
    "11101110", --  345 - 0x159  :  238 - 0xee
    "11101100", --  346 - 0x15a  :  236 - 0xec
    "00001110", --  347 - 0x15b  :   14 - 0xe
    "11110100", --  348 - 0x15c  :  244 - 0xf4
    "11111010", --  349 - 0x15d  :  250 - 0xfa
    "01010100", --  350 - 0x15e  :   84 - 0x54
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Background 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00011110", --  360 - 0x168  :   30 - 0x1e -- Background 0x2d
    "00111110", --  361 - 0x169  :   62 - 0x3e
    "00111110", --  362 - 0x16a  :   62 - 0x3e
    "00111110", --  363 - 0x16b  :   62 - 0x3e
    "00111111", --  364 - 0x16c  :   63 - 0x3f
    "00011110", --  365 - 0x16d  :   30 - 0x1e
    "00001111", --  366 - 0x16e  :   15 - 0xf
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Background 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "01111000", --  376 - 0x178  :  120 - 0x78 -- Background 0x2f
    "01111100", --  377 - 0x179  :  124 - 0x7c
    "01111100", --  378 - 0x17a  :  124 - 0x7c
    "01111100", --  379 - 0x17b  :  124 - 0x7c
    "11111100", --  380 - 0x17c  :  252 - 0xfc
    "01111000", --  381 - 0x17d  :  120 - 0x78
    "11110000", --  382 - 0x17e  :  240 - 0xf0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000000", --  384 - 0x180  :    0 - 0x0 -- Background 0x30
    "00011000", --  385 - 0x181  :   24 - 0x18
    "00111100", --  386 - 0x182  :   60 - 0x3c
    "01011010", --  387 - 0x183  :   90 - 0x5a
    "00011000", --  388 - 0x184  :   24 - 0x18
    "00011000", --  389 - 0x185  :   24 - 0x18
    "00011000", --  390 - 0x186  :   24 - 0x18
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0 -- Background 0x31
    "00011000", --  393 - 0x189  :   24 - 0x18
    "00011000", --  394 - 0x18a  :   24 - 0x18
    "00011000", --  395 - 0x18b  :   24 - 0x18
    "01011010", --  396 - 0x18c  :   90 - 0x5a
    "00111100", --  397 - 0x18d  :   60 - 0x3c
    "00011000", --  398 - 0x18e  :   24 - 0x18
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00000001", --  400 - 0x190  :    1 - 0x1 -- Background 0x32
    "00000001", --  401 - 0x191  :    1 - 0x1
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000001", --  403 - 0x193  :    1 - 0x1
    "00000001", --  404 - 0x194  :    1 - 0x1
    "00000001", --  405 - 0x195  :    1 - 0x1
    "00000000", --  406 - 0x196  :    0 - 0x0
    "00000001", --  407 - 0x197  :    1 - 0x1
    "10000000", --  408 - 0x198  :  128 - 0x80 -- Background 0x33
    "00000000", --  409 - 0x199  :    0 - 0x0
    "10000000", --  410 - 0x19a  :  128 - 0x80
    "10000000", --  411 - 0x19b  :  128 - 0x80
    "10000000", --  412 - 0x19c  :  128 - 0x80
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "10000000", --  414 - 0x19e  :  128 - 0x80
    "10000000", --  415 - 0x19f  :  128 - 0x80
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- Background 0x34
    "00000000", --  417 - 0x1a1  :    0 - 0x0
    "00011000", --  418 - 0x1a2  :   24 - 0x18
    "00111100", --  419 - 0x1a3  :   60 - 0x3c
    "00111110", --  420 - 0x1a4  :   62 - 0x3e
    "01111111", --  421 - 0x1a5  :  127 - 0x7f
    "01111111", --  422 - 0x1a6  :  127 - 0x7f
    "01111111", --  423 - 0x1a7  :  127 - 0x7f
    "00111111", --  424 - 0x1a8  :   63 - 0x3f -- Background 0x35
    "00111111", --  425 - 0x1a9  :   63 - 0x3f
    "00011111", --  426 - 0x1aa  :   31 - 0x1f
    "00001111", --  427 - 0x1ab  :   15 - 0xf
    "00000111", --  428 - 0x1ac  :    7 - 0x7
    "00000011", --  429 - 0x1ad  :    3 - 0x3
    "00000001", --  430 - 0x1ae  :    1 - 0x1
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Background 0x36
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00011000", --  434 - 0x1b2  :   24 - 0x18
    "00111100", --  435 - 0x1b3  :   60 - 0x3c
    "01111100", --  436 - 0x1b4  :  124 - 0x7c
    "11111110", --  437 - 0x1b5  :  254 - 0xfe
    "11111110", --  438 - 0x1b6  :  254 - 0xfe
    "11111110", --  439 - 0x1b7  :  254 - 0xfe
    "11111100", --  440 - 0x1b8  :  252 - 0xfc -- Background 0x37
    "11111100", --  441 - 0x1b9  :  252 - 0xfc
    "11111000", --  442 - 0x1ba  :  248 - 0xf8
    "11110000", --  443 - 0x1bb  :  240 - 0xf0
    "11100000", --  444 - 0x1bc  :  224 - 0xe0
    "11000000", --  445 - 0x1bd  :  192 - 0xc0
    "10000000", --  446 - 0x1be  :  128 - 0x80
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Background 0x38
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000110", --  450 - 0x1c2  :    6 - 0x6
    "00000111", --  451 - 0x1c3  :    7 - 0x7
    "00000111", --  452 - 0x1c4  :    7 - 0x7
    "00000011", --  453 - 0x1c5  :    3 - 0x3
    "00000001", --  454 - 0x1c6  :    1 - 0x1
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- Background 0x39
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Background 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "01100000", --  466 - 0x1d2  :   96 - 0x60
    "11100000", --  467 - 0x1d3  :  224 - 0xe0
    "11100000", --  468 - 0x1d4  :  224 - 0xe0
    "11000000", --  469 - 0x1d5  :  192 - 0xc0
    "10000000", --  470 - 0x1d6  :  128 - 0x80
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Background 0x3b
    "00101010", --  473 - 0x1d9  :   42 - 0x2a
    "01000000", --  474 - 0x1da  :   64 - 0x40
    "00000010", --  475 - 0x1db  :    2 - 0x2
    "01000000", --  476 - 0x1dc  :   64 - 0x40
    "00000010", --  477 - 0x1dd  :    2 - 0x2
    "01010100", --  478 - 0x1de  :   84 - 0x54
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Background 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "00000000", --  485 - 0x1e5  :    0 - 0x0
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "11111111", --  488 - 0x1e8  :  255 - 0xff -- Background 0x3d
    "11111111", --  489 - 0x1e9  :  255 - 0xff
    "11111111", --  490 - 0x1ea  :  255 - 0xff
    "11111111", --  491 - 0x1eb  :  255 - 0xff
    "11111111", --  492 - 0x1ec  :  255 - 0xff
    "11111111", --  493 - 0x1ed  :  255 - 0xff
    "11111111", --  494 - 0x1ee  :  255 - 0xff
    "11111111", --  495 - 0x1ef  :  255 - 0xff
    "11111111", --  496 - 0x1f0  :  255 - 0xff -- Background 0x3e
    "11111111", --  497 - 0x1f1  :  255 - 0xff
    "11111111", --  498 - 0x1f2  :  255 - 0xff
    "11111111", --  499 - 0x1f3  :  255 - 0xff
    "11111111", --  500 - 0x1f4  :  255 - 0xff
    "11111111", --  501 - 0x1f5  :  255 - 0xff
    "11111111", --  502 - 0x1f6  :  255 - 0xff
    "11111111", --  503 - 0x1f7  :  255 - 0xff
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- Background 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Background 0x40
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0 -- Background 0x41
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Background 0x42
    "00000000", --  529 - 0x211  :    0 - 0x0
    "00000000", --  530 - 0x212  :    0 - 0x0
    "00000000", --  531 - 0x213  :    0 - 0x0
    "00000000", --  532 - 0x214  :    0 - 0x0
    "00000000", --  533 - 0x215  :    0 - 0x0
    "00000000", --  534 - 0x216  :    0 - 0x0
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00000000", --  536 - 0x218  :    0 - 0x0 -- Background 0x43
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Background 0x44
    "00000000", --  545 - 0x221  :    0 - 0x0
    "00000000", --  546 - 0x222  :    0 - 0x0
    "00000000", --  547 - 0x223  :    0 - 0x0
    "00000000", --  548 - 0x224  :    0 - 0x0
    "00000000", --  549 - 0x225  :    0 - 0x0
    "00000000", --  550 - 0x226  :    0 - 0x0
    "00000000", --  551 - 0x227  :    0 - 0x0
    "00000000", --  552 - 0x228  :    0 - 0x0 -- Background 0x45
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000000", --  560 - 0x230  :    0 - 0x0 -- Background 0x46
    "00000000", --  561 - 0x231  :    0 - 0x0
    "00000000", --  562 - 0x232  :    0 - 0x0
    "00000000", --  563 - 0x233  :    0 - 0x0
    "00000000", --  564 - 0x234  :    0 - 0x0
    "00000000", --  565 - 0x235  :    0 - 0x0
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00000000", --  568 - 0x238  :    0 - 0x0 -- Background 0x47
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Background 0x48
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00000000", --  584 - 0x248  :    0 - 0x0 -- Background 0x49
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000000", --  592 - 0x250  :    0 - 0x0 -- Background 0x4a
    "00000000", --  593 - 0x251  :    0 - 0x0
    "00000000", --  594 - 0x252  :    0 - 0x0
    "00000000", --  595 - 0x253  :    0 - 0x0
    "00000000", --  596 - 0x254  :    0 - 0x0
    "00000000", --  597 - 0x255  :    0 - 0x0
    "00000000", --  598 - 0x256  :    0 - 0x0
    "00000000", --  599 - 0x257  :    0 - 0x0
    "00000000", --  600 - 0x258  :    0 - 0x0 -- Background 0x4b
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Background 0x4c
    "00000000", --  609 - 0x261  :    0 - 0x0
    "00000000", --  610 - 0x262  :    0 - 0x0
    "00000000", --  611 - 0x263  :    0 - 0x0
    "00000000", --  612 - 0x264  :    0 - 0x0
    "00000000", --  613 - 0x265  :    0 - 0x0
    "00000000", --  614 - 0x266  :    0 - 0x0
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0 -- Background 0x4d
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Background 0x4e
    "00000000", --  625 - 0x271  :    0 - 0x0
    "00000000", --  626 - 0x272  :    0 - 0x0
    "00000000", --  627 - 0x273  :    0 - 0x0
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000000", --  629 - 0x275  :    0 - 0x0
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0 -- Background 0x4f
    "00000000", --  633 - 0x279  :    0 - 0x0
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "00000000", --  635 - 0x27b  :    0 - 0x0
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Background 0x50
    "00111111", --  641 - 0x281  :   63 - 0x3f
    "01111111", --  642 - 0x282  :  127 - 0x7f
    "01111111", --  643 - 0x283  :  127 - 0x7f
    "01111111", --  644 - 0x284  :  127 - 0x7f
    "00111100", --  645 - 0x285  :   60 - 0x3c
    "00000000", --  646 - 0x286  :    0 - 0x0
    "01000000", --  647 - 0x287  :   64 - 0x40
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Background 0x51
    "11111100", --  649 - 0x289  :  252 - 0xfc
    "11111110", --  650 - 0x28a  :  254 - 0xfe
    "11111110", --  651 - 0x28b  :  254 - 0xfe
    "11111110", --  652 - 0x28c  :  254 - 0xfe
    "00111100", --  653 - 0x28d  :   60 - 0x3c
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000010", --  655 - 0x28f  :    2 - 0x2
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Background 0x52
    "00000000", --  657 - 0x291  :    0 - 0x0
    "00000011", --  658 - 0x292  :    3 - 0x3
    "00000111", --  659 - 0x293  :    7 - 0x7
    "00001111", --  660 - 0x294  :   15 - 0xf
    "00011111", --  661 - 0x295  :   31 - 0x1f
    "00111111", --  662 - 0x296  :   63 - 0x3f
    "00110000", --  663 - 0x297  :   48 - 0x30
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Background 0x53
    "00000000", --  665 - 0x299  :    0 - 0x0
    "10100000", --  666 - 0x29a  :  160 - 0xa0
    "10110000", --  667 - 0x29b  :  176 - 0xb0
    "10110000", --  668 - 0x29c  :  176 - 0xb0
    "10111000", --  669 - 0x29d  :  184 - 0xb8
    "01111100", --  670 - 0x29e  :  124 - 0x7c
    "01111100", --  671 - 0x29f  :  124 - 0x7c
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Background 0x54
    "00100001", --  673 - 0x2a1  :   33 - 0x21
    "01110001", --  674 - 0x2a2  :  113 - 0x71
    "00111010", --  675 - 0x2a3  :   58 - 0x3a
    "01101101", --  676 - 0x2a4  :  109 - 0x6d
    "00111000", --  677 - 0x2a5  :   56 - 0x38
    "00011101", --  678 - 0x2a6  :   29 - 0x1d
    "00101111", --  679 - 0x2a7  :   47 - 0x2f
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- Background 0x55
    "00100001", --  681 - 0x2a9  :   33 - 0x21
    "01110001", --  682 - 0x2aa  :  113 - 0x71
    "00111010", --  683 - 0x2ab  :   58 - 0x3a
    "01101101", --  684 - 0x2ac  :  109 - 0x6d
    "10111000", --  685 - 0x2ad  :  184 - 0xb8
    "00011101", --  686 - 0x2ae  :   29 - 0x1d
    "10101111", --  687 - 0x2af  :  175 - 0xaf
    "00000000", --  688 - 0x2b0  :    0 - 0x0 -- Background 0x56
    "00100000", --  689 - 0x2b1  :   32 - 0x20
    "01110000", --  690 - 0x2b2  :  112 - 0x70
    "00111010", --  691 - 0x2b3  :   58 - 0x3a
    "01101100", --  692 - 0x2b4  :  108 - 0x6c
    "10111000", --  693 - 0x2b5  :  184 - 0xb8
    "00011100", --  694 - 0x2b6  :   28 - 0x1c
    "10101110", --  695 - 0x2b7  :  174 - 0xae
    "00000000", --  696 - 0x2b8  :    0 - 0x0 -- Background 0x57
    "01111111", --  697 - 0x2b9  :  127 - 0x7f
    "01001100", --  698 - 0x2ba  :   76 - 0x4c
    "00110011", --  699 - 0x2bb  :   51 - 0x33
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Background 0x58
    "11111111", --  705 - 0x2c1  :  255 - 0xff
    "11001100", --  706 - 0x2c2  :  204 - 0xcc
    "00110011", --  707 - 0x2c3  :   51 - 0x33
    "11001100", --  708 - 0x2c4  :  204 - 0xcc
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0 -- Background 0x59
    "11111110", --  713 - 0x2c9  :  254 - 0xfe
    "11001100", --  714 - 0x2ca  :  204 - 0xcc
    "00110000", --  715 - 0x2cb  :   48 - 0x30
    "11000000", --  716 - 0x2cc  :  192 - 0xc0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Background 0x5a
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Background 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000001", --  732 - 0x2dc  :    1 - 0x1
    "00000001", --  733 - 0x2dd  :    1 - 0x1
    "00000011", --  734 - 0x2de  :    3 - 0x3
    "00000011", --  735 - 0x2df  :    3 - 0x3
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Background 0x5c
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000001", --  738 - 0x2e2  :    1 - 0x1
    "01111110", --  739 - 0x2e3  :  126 - 0x7e
    "11111111", --  740 - 0x2e4  :  255 - 0xff
    "11111111", --  741 - 0x2e5  :  255 - 0xff
    "11111111", --  742 - 0x2e6  :  255 - 0xff
    "11111111", --  743 - 0x2e7  :  255 - 0xff
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- Background 0x5d
    "11111111", --  745 - 0x2e9  :  255 - 0xff
    "11111111", --  746 - 0x2ea  :  255 - 0xff
    "11111111", --  747 - 0x2eb  :  255 - 0xff
    "01111111", --  748 - 0x2ec  :  127 - 0x7f
    "11111111", --  749 - 0x2ed  :  255 - 0xff
    "11111111", --  750 - 0x2ee  :  255 - 0xff
    "11111111", --  751 - 0x2ef  :  255 - 0xff
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Background 0x5e
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "10000000", --  754 - 0x2f2  :  128 - 0x80
    "01111110", --  755 - 0x2f3  :  126 - 0x7e
    "10111111", --  756 - 0x2f4  :  191 - 0xbf
    "11111111", --  757 - 0x2f5  :  255 - 0xff
    "11111111", --  758 - 0x2f6  :  255 - 0xff
    "11111111", --  759 - 0x2f7  :  255 - 0xff
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- Background 0x5f
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "10000000", --  764 - 0x2fc  :  128 - 0x80
    "10000000", --  765 - 0x2fd  :  128 - 0x80
    "11000000", --  766 - 0x2fe  :  192 - 0xc0
    "11000000", --  767 - 0x2ff  :  192 - 0xc0
    "01111111", --  768 - 0x300  :  127 - 0x7f -- Background 0x60
    "01111111", --  769 - 0x301  :  127 - 0x7f
    "01111101", --  770 - 0x302  :  125 - 0x7d
    "01111111", --  771 - 0x303  :  127 - 0x7f
    "00111111", --  772 - 0x304  :   63 - 0x3f
    "01111111", --  773 - 0x305  :  127 - 0x7f
    "01111111", --  774 - 0x306  :  127 - 0x7f
    "01110111", --  775 - 0x307  :  119 - 0x77
    "11111110", --  776 - 0x308  :  254 - 0xfe -- Background 0x61
    "11111110", --  777 - 0x309  :  254 - 0xfe
    "11111100", --  778 - 0x30a  :  252 - 0xfc
    "11111110", --  779 - 0x30b  :  254 - 0xfe
    "10111110", --  780 - 0x30c  :  190 - 0xbe
    "11111110", --  781 - 0x30d  :  254 - 0xfe
    "11111110", --  782 - 0x30e  :  254 - 0xfe
    "11110110", --  783 - 0x30f  :  246 - 0xf6
    "00000111", --  784 - 0x310  :    7 - 0x7 -- Background 0x62
    "00011111", --  785 - 0x311  :   31 - 0x1f
    "00111111", --  786 - 0x312  :   63 - 0x3f
    "00111111", --  787 - 0x313  :   63 - 0x3f
    "00111111", --  788 - 0x314  :   63 - 0x3f
    "00011111", --  789 - 0x315  :   31 - 0x1f
    "00001111", --  790 - 0x316  :   15 - 0xf
    "00000000", --  791 - 0x317  :    0 - 0x0
    "01111110", --  792 - 0x318  :  126 - 0x7e -- Background 0x63
    "01111100", --  793 - 0x319  :  124 - 0x7c
    "00111110", --  794 - 0x31a  :   62 - 0x3e
    "10111100", --  795 - 0x31b  :  188 - 0xbc
    "10111110", --  796 - 0x31c  :  190 - 0xbe
    "10011100", --  797 - 0x31d  :  156 - 0x9c
    "11011000", --  798 - 0x31e  :  216 - 0xd8
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "01000110", --  800 - 0x320  :   70 - 0x46 -- Background 0x64
    "01101011", --  801 - 0x321  :  107 - 0x6b
    "01110001", --  802 - 0x322  :  113 - 0x71
    "00111010", --  803 - 0x323  :   58 - 0x3a
    "01101101", --  804 - 0x324  :  109 - 0x6d
    "00111000", --  805 - 0x325  :   56 - 0x38
    "00011101", --  806 - 0x326  :   29 - 0x1d
    "00101111", --  807 - 0x327  :   47 - 0x2f
    "01000110", --  808 - 0x328  :   70 - 0x46 -- Background 0x65
    "11101011", --  809 - 0x329  :  235 - 0xeb
    "01110001", --  810 - 0x32a  :  113 - 0x71
    "00111010", --  811 - 0x32b  :   58 - 0x3a
    "01101101", --  812 - 0x32c  :  109 - 0x6d
    "10111000", --  813 - 0x32d  :  184 - 0xb8
    "00011101", --  814 - 0x32e  :   29 - 0x1d
    "10101111", --  815 - 0x32f  :  175 - 0xaf
    "01000110", --  816 - 0x330  :   70 - 0x46 -- Background 0x66
    "11101010", --  817 - 0x331  :  234 - 0xea
    "01110000", --  818 - 0x332  :  112 - 0x70
    "00111010", --  819 - 0x333  :   58 - 0x3a
    "01101100", --  820 - 0x334  :  108 - 0x6c
    "10111000", --  821 - 0x335  :  184 - 0xb8
    "00011100", --  822 - 0x336  :   28 - 0x1c
    "10101110", --  823 - 0x337  :  174 - 0xae
    "00000000", --  824 - 0x338  :    0 - 0x0 -- Background 0x67
    "01111111", --  825 - 0x339  :  127 - 0x7f
    "01111111", --  826 - 0x33a  :  127 - 0x7f
    "00110011", --  827 - 0x33b  :   51 - 0x33
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Background 0x68
    "11111111", --  833 - 0x341  :  255 - 0xff
    "11111111", --  834 - 0x342  :  255 - 0xff
    "11111111", --  835 - 0x343  :  255 - 0xff
    "11001100", --  836 - 0x344  :  204 - 0xcc
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Background 0x69
    "11111110", --  841 - 0x349  :  254 - 0xfe
    "11111110", --  842 - 0x34a  :  254 - 0xfe
    "11110000", --  843 - 0x34b  :  240 - 0xf0
    "11000000", --  844 - 0x34c  :  192 - 0xc0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Background 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00111101", --  856 - 0x358  :   61 - 0x3d -- Background 0x6b
    "01111111", --  857 - 0x359  :  127 - 0x7f
    "01111111", --  858 - 0x35a  :  127 - 0x7f
    "01111111", --  859 - 0x35b  :  127 - 0x7f
    "00111111", --  860 - 0x35c  :   63 - 0x3f
    "00001111", --  861 - 0x35d  :   15 - 0xf
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "11111111", --  864 - 0x360  :  255 - 0xff -- Background 0x6c
    "11111111", --  865 - 0x361  :  255 - 0xff
    "11111111", --  866 - 0x362  :  255 - 0xff
    "11111111", --  867 - 0x363  :  255 - 0xff
    "11111111", --  868 - 0x364  :  255 - 0xff
    "11111111", --  869 - 0x365  :  255 - 0xff
    "11111110", --  870 - 0x366  :  254 - 0xfe
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Background 0x6d
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Background 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "10111000", --  888 - 0x378  :  184 - 0xb8 -- Background 0x6f
    "11111100", --  889 - 0x379  :  252 - 0xfc
    "11111110", --  890 - 0x37a  :  254 - 0xfe
    "11111110", --  891 - 0x37b  :  254 - 0xfe
    "11111100", --  892 - 0x37c  :  252 - 0xfc
    "11110000", --  893 - 0x37d  :  240 - 0xf0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Background 0x70
    "00111111", --  897 - 0x381  :   63 - 0x3f
    "01111111", --  898 - 0x382  :  127 - 0x7f
    "01111111", --  899 - 0x383  :  127 - 0x7f
    "00011100", --  900 - 0x384  :   28 - 0x1c
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0 -- Background 0x71
    "11111111", --  905 - 0x389  :  255 - 0xff
    "11111111", --  906 - 0x38a  :  255 - 0xff
    "11111111", --  907 - 0x38b  :  255 - 0xff
    "11111111", --  908 - 0x38c  :  255 - 0xff
    "00111100", --  909 - 0x38d  :   60 - 0x3c
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Background 0x72
    "11111100", --  913 - 0x391  :  252 - 0xfc
    "11111110", --  914 - 0x392  :  254 - 0xfe
    "11111110", --  915 - 0x393  :  254 - 0xfe
    "00111000", --  916 - 0x394  :   56 - 0x38
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "11111111", --  920 - 0x398  :  255 - 0xff -- Background 0x73
    "11111111", --  921 - 0x399  :  255 - 0xff
    "11111101", --  922 - 0x39a  :  253 - 0xfd
    "11111111", --  923 - 0x39b  :  255 - 0xff
    "10111111", --  924 - 0x39c  :  191 - 0xbf
    "11111111", --  925 - 0x39d  :  255 - 0xff
    "11111111", --  926 - 0x39e  :  255 - 0xff
    "11110111", --  927 - 0x39f  :  247 - 0xf7
    "01000110", --  928 - 0x3a0  :   70 - 0x46 -- Background 0x74
    "01101011", --  929 - 0x3a1  :  107 - 0x6b
    "01110001", --  930 - 0x3a2  :  113 - 0x71
    "00111010", --  931 - 0x3a3  :   58 - 0x3a
    "01101101", --  932 - 0x3a4  :  109 - 0x6d
    "00111000", --  933 - 0x3a5  :   56 - 0x38
    "00011101", --  934 - 0x3a6  :   29 - 0x1d
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "01000110", --  936 - 0x3a8  :   70 - 0x46 -- Background 0x75
    "11101011", --  937 - 0x3a9  :  235 - 0xeb
    "01110001", --  938 - 0x3aa  :  113 - 0x71
    "00111010", --  939 - 0x3ab  :   58 - 0x3a
    "01101101", --  940 - 0x3ac  :  109 - 0x6d
    "10111000", --  941 - 0x3ad  :  184 - 0xb8
    "00011101", --  942 - 0x3ae  :   29 - 0x1d
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "01000110", --  944 - 0x3b0  :   70 - 0x46 -- Background 0x76
    "11101010", --  945 - 0x3b1  :  234 - 0xea
    "01110000", --  946 - 0x3b2  :  112 - 0x70
    "00111010", --  947 - 0x3b3  :   58 - 0x3a
    "01101100", --  948 - 0x3b4  :  108 - 0x6c
    "10111000", --  949 - 0x3b5  :  184 - 0xb8
    "00011100", --  950 - 0x3b6  :   28 - 0x1c
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "10000001", --  952 - 0x3b8  :  129 - 0x81 -- Background 0x77
    "11111111", --  953 - 0x3b9  :  255 - 0xff
    "11111101", --  954 - 0x3ba  :  253 - 0xfd
    "11111111", --  955 - 0x3bb  :  255 - 0xff
    "10111111", --  956 - 0x3bc  :  191 - 0xbf
    "11111111", --  957 - 0x3bd  :  255 - 0xff
    "11111111", --  958 - 0x3be  :  255 - 0xff
    "11110111", --  959 - 0x3bf  :  247 - 0xf7
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Background 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Background 0x79
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Background 0x7a
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Background 0x7b
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Background 0x7c
    "00100010", --  993 - 0x3e1  :   34 - 0x22
    "01110111", --  994 - 0x3e2  :  119 - 0x77
    "11111111", --  995 - 0x3e3  :  255 - 0xff
    "11111011", --  996 - 0x3e4  :  251 - 0xfb
    "11110101", --  997 - 0x3e5  :  245 - 0xf5
    "11101111", --  998 - 0x3e6  :  239 - 0xef
    "11111111", --  999 - 0x3e7  :  255 - 0xff
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Background 0x7d
    "01110011", -- 1001 - 0x3e9  :  115 - 0x73
    "11111111", -- 1002 - 0x3ea  :  255 - 0xff
    "11111111", -- 1003 - 0x3eb  :  255 - 0xff
    "11111011", -- 1004 - 0x3ec  :  251 - 0xfb
    "11111101", -- 1005 - 0x3ed  :  253 - 0xfd
    "11101111", -- 1006 - 0x3ee  :  239 - 0xef
    "11111111", -- 1007 - 0x3ef  :  255 - 0xff
    "11011111", -- 1008 - 0x3f0  :  223 - 0xdf -- Background 0x7e
    "10101111", -- 1009 - 0x3f1  :  175 - 0xaf
    "01111111", -- 1010 - 0x3f2  :  127 - 0x7f
    "11111111", -- 1011 - 0x3f3  :  255 - 0xff
    "11111011", -- 1012 - 0x3f4  :  251 - 0xfb
    "11110101", -- 1013 - 0x3f5  :  245 - 0xf5
    "11101111", -- 1014 - 0x3f6  :  239 - 0xef
    "11111111", -- 1015 - 0x3f7  :  255 - 0xff
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- Background 0x7f
    "10101111", -- 1017 - 0x3f9  :  175 - 0xaf
    "01111111", -- 1018 - 0x3fa  :  127 - 0x7f
    "11111111", -- 1019 - 0x3fb  :  255 - 0xff
    "11111011", -- 1020 - 0x3fc  :  251 - 0xfb
    "11110101", -- 1021 - 0x3fd  :  245 - 0xf5
    "11101111", -- 1022 - 0x3fe  :  239 - 0xef
    "11111111", -- 1023 - 0x3ff  :  255 - 0xff
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Background 0x80
    "01111111", -- 1025 - 0x401  :  127 - 0x7f
    "00110000", -- 1026 - 0x402  :   48 - 0x30
    "00110000", -- 1027 - 0x403  :   48 - 0x30
    "00110000", -- 1028 - 0x404  :   48 - 0x30
    "01111111", -- 1029 - 0x405  :  127 - 0x7f
    "00110000", -- 1030 - 0x406  :   48 - 0x30
    "00110000", -- 1031 - 0x407  :   48 - 0x30
    "00000000", -- 1032 - 0x408  :    0 - 0x0 -- Background 0x81
    "01111111", -- 1033 - 0x409  :  127 - 0x7f
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "01111111", -- 1035 - 0x40b  :  127 - 0x7f
    "01111111", -- 1036 - 0x40c  :  127 - 0x7f
    "00100000", -- 1037 - 0x40d  :   32 - 0x20
    "01000000", -- 1038 - 0x40e  :   64 - 0x40
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Background 0x82
    "11111110", -- 1041 - 0x411  :  254 - 0xfe
    "00001100", -- 1042 - 0x412  :   12 - 0xc
    "00001100", -- 1043 - 0x413  :   12 - 0xc
    "00001100", -- 1044 - 0x414  :   12 - 0xc
    "11111110", -- 1045 - 0x415  :  254 - 0xfe
    "00001100", -- 1046 - 0x416  :   12 - 0xc
    "00001100", -- 1047 - 0x417  :   12 - 0xc
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- Background 0x83
    "11111111", -- 1049 - 0x419  :  255 - 0xff
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "11111111", -- 1051 - 0x41b  :  255 - 0xff
    "11111111", -- 1052 - 0x41c  :  255 - 0xff
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- Background 0x84
    "11111111", -- 1057 - 0x421  :  255 - 0xff
    "11111111", -- 1058 - 0x422  :  255 - 0xff
    "11111111", -- 1059 - 0x423  :  255 - 0xff
    "11111111", -- 1060 - 0x424  :  255 - 0xff
    "11101111", -- 1061 - 0x425  :  239 - 0xef
    "10111011", -- 1062 - 0x426  :  187 - 0xbb
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0 -- Background 0x85
    "11111110", -- 1065 - 0x429  :  254 - 0xfe
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "11111110", -- 1067 - 0x42b  :  254 - 0xfe
    "11111110", -- 1068 - 0x42c  :  254 - 0xfe
    "00001100", -- 1069 - 0x42d  :   12 - 0xc
    "00000010", -- 1070 - 0x42e  :    2 - 0x2
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Background 0x86
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- Background 0x87
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Background 0x88
    "00000111", -- 1089 - 0x441  :    7 - 0x7
    "00011111", -- 1090 - 0x442  :   31 - 0x1f
    "00111100", -- 1091 - 0x443  :   60 - 0x3c
    "00110001", -- 1092 - 0x444  :   49 - 0x31
    "01110100", -- 1093 - 0x445  :  116 - 0x74
    "01100101", -- 1094 - 0x446  :  101 - 0x65
    "01101010", -- 1095 - 0x447  :  106 - 0x6a
    "01100100", -- 1096 - 0x448  :  100 - 0x64 -- Background 0x89
    "01101101", -- 1097 - 0x449  :  109 - 0x6d
    "01110010", -- 1098 - 0x44a  :  114 - 0x72
    "00110000", -- 1099 - 0x44b  :   48 - 0x30
    "00111100", -- 1100 - 0x44c  :   60 - 0x3c
    "00011111", -- 1101 - 0x44d  :   31 - 0x1f
    "00000111", -- 1102 - 0x44e  :    7 - 0x7
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Background 0x8a
    "11100000", -- 1105 - 0x451  :  224 - 0xe0
    "11111000", -- 1106 - 0x452  :  248 - 0xf8
    "00111100", -- 1107 - 0x453  :   60 - 0x3c
    "01001100", -- 1108 - 0x454  :   76 - 0x4c
    "01101110", -- 1109 - 0x455  :  110 - 0x6e
    "00100110", -- 1110 - 0x456  :   38 - 0x26
    "01000110", -- 1111 - 0x457  :   70 - 0x46
    "10010110", -- 1112 - 0x458  :  150 - 0x96 -- Background 0x8b
    "01100110", -- 1113 - 0x459  :  102 - 0x66
    "10101110", -- 1114 - 0x45a  :  174 - 0xae
    "01001100", -- 1115 - 0x45b  :   76 - 0x4c
    "00111100", -- 1116 - 0x45c  :   60 - 0x3c
    "11111000", -- 1117 - 0x45d  :  248 - 0xf8
    "11100000", -- 1118 - 0x45e  :  224 - 0xe0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Background 0x8c
    "00000111", -- 1121 - 0x461  :    7 - 0x7
    "00011111", -- 1122 - 0x462  :   31 - 0x1f
    "00111111", -- 1123 - 0x463  :   63 - 0x3f
    "00111111", -- 1124 - 0x464  :   63 - 0x3f
    "01111111", -- 1125 - 0x465  :  127 - 0x7f
    "01111111", -- 1126 - 0x466  :  127 - 0x7f
    "01111111", -- 1127 - 0x467  :  127 - 0x7f
    "01111111", -- 1128 - 0x468  :  127 - 0x7f -- Background 0x8d
    "01111111", -- 1129 - 0x469  :  127 - 0x7f
    "01111111", -- 1130 - 0x46a  :  127 - 0x7f
    "00111111", -- 1131 - 0x46b  :   63 - 0x3f
    "00111111", -- 1132 - 0x46c  :   63 - 0x3f
    "00011111", -- 1133 - 0x46d  :   31 - 0x1f
    "00000111", -- 1134 - 0x46e  :    7 - 0x7
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0 -- Background 0x8e
    "11100000", -- 1137 - 0x471  :  224 - 0xe0
    "11111000", -- 1138 - 0x472  :  248 - 0xf8
    "11111100", -- 1139 - 0x473  :  252 - 0xfc
    "11111100", -- 1140 - 0x474  :  252 - 0xfc
    "11111110", -- 1141 - 0x475  :  254 - 0xfe
    "11111110", -- 1142 - 0x476  :  254 - 0xfe
    "11111110", -- 1143 - 0x477  :  254 - 0xfe
    "11111110", -- 1144 - 0x478  :  254 - 0xfe -- Background 0x8f
    "11111110", -- 1145 - 0x479  :  254 - 0xfe
    "11111110", -- 1146 - 0x47a  :  254 - 0xfe
    "11111100", -- 1147 - 0x47b  :  252 - 0xfc
    "11111100", -- 1148 - 0x47c  :  252 - 0xfc
    "11111000", -- 1149 - 0x47d  :  248 - 0xf8
    "11100000", -- 1150 - 0x47e  :  224 - 0xe0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Background 0x90
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00010000", -- 1156 - 0x484  :   16 - 0x10
    "00011100", -- 1157 - 0x485  :   28 - 0x1c
    "00001110", -- 1158 - 0x486  :   14 - 0xe
    "00000111", -- 1159 - 0x487  :    7 - 0x7
    "00000011", -- 1160 - 0x488  :    3 - 0x3 -- Background 0x91
    "00000001", -- 1161 - 0x489  :    1 - 0x1
    "00110000", -- 1162 - 0x48a  :   48 - 0x30
    "00001111", -- 1163 - 0x48b  :   15 - 0xf
    "00000011", -- 1164 - 0x48c  :    3 - 0x3
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "01111111", -- 1166 - 0x48e  :  127 - 0x7f
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0 -- Background 0x92
    "01000010", -- 1169 - 0x491  :   66 - 0x42
    "01000010", -- 1170 - 0x492  :   66 - 0x42
    "01100110", -- 1171 - 0x493  :  102 - 0x66
    "01100110", -- 1172 - 0x494  :  102 - 0x66
    "01100110", -- 1173 - 0x495  :  102 - 0x66
    "11111110", -- 1174 - 0x496  :  254 - 0xfe
    "11111111", -- 1175 - 0x497  :  255 - 0xff
    "01111110", -- 1176 - 0x498  :  126 - 0x7e -- Background 0x93
    "01111110", -- 1177 - 0x499  :  126 - 0x7e
    "01111110", -- 1178 - 0x49a  :  126 - 0x7e
    "01111110", -- 1179 - 0x49b  :  126 - 0x7e
    "01111110", -- 1180 - 0x49c  :  126 - 0x7e
    "01111110", -- 1181 - 0x49d  :  126 - 0x7e
    "01111110", -- 1182 - 0x49e  :  126 - 0x7e
    "01111110", -- 1183 - 0x49f  :  126 - 0x7e
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- Background 0x94
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000000", -- 1186 - 0x4a2  :    0 - 0x0
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00001000", -- 1188 - 0x4a4  :    8 - 0x8
    "00111000", -- 1189 - 0x4a5  :   56 - 0x38
    "01110000", -- 1190 - 0x4a6  :  112 - 0x70
    "11100000", -- 1191 - 0x4a7  :  224 - 0xe0
    "11000000", -- 1192 - 0x4a8  :  192 - 0xc0 -- Background 0x95
    "10000000", -- 1193 - 0x4a9  :  128 - 0x80
    "00001100", -- 1194 - 0x4aa  :   12 - 0xc
    "11110000", -- 1195 - 0x4ab  :  240 - 0xf0
    "11000000", -- 1196 - 0x4ac  :  192 - 0xc0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "11111110", -- 1198 - 0x4ae  :  254 - 0xfe
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0 -- Background 0x96
    "00111111", -- 1201 - 0x4b1  :   63 - 0x3f
    "01111111", -- 1202 - 0x4b2  :  127 - 0x7f
    "01111111", -- 1203 - 0x4b3  :  127 - 0x7f
    "01111111", -- 1204 - 0x4b4  :  127 - 0x7f
    "01111111", -- 1205 - 0x4b5  :  127 - 0x7f
    "01111111", -- 1206 - 0x4b6  :  127 - 0x7f
    "01111111", -- 1207 - 0x4b7  :  127 - 0x7f
    "01111111", -- 1208 - 0x4b8  :  127 - 0x7f -- Background 0x97
    "01111111", -- 1209 - 0x4b9  :  127 - 0x7f
    "00111111", -- 1210 - 0x4ba  :   63 - 0x3f
    "01111111", -- 1211 - 0x4bb  :  127 - 0x7f
    "01111111", -- 1212 - 0x4bc  :  127 - 0x7f
    "01111111", -- 1213 - 0x4bd  :  127 - 0x7f
    "01111111", -- 1214 - 0x4be  :  127 - 0x7f
    "01111111", -- 1215 - 0x4bf  :  127 - 0x7f
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- Background 0x98
    "11011111", -- 1217 - 0x4c1  :  223 - 0xdf
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111111", -- 1219 - 0x4c3  :  255 - 0xff
    "11111111", -- 1220 - 0x4c4  :  255 - 0xff
    "11111111", -- 1221 - 0x4c5  :  255 - 0xff
    "11111111", -- 1222 - 0x4c6  :  255 - 0xff
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "11111111", -- 1224 - 0x4c8  :  255 - 0xff -- Background 0x99
    "11111111", -- 1225 - 0x4c9  :  255 - 0xff
    "10111111", -- 1226 - 0x4ca  :  191 - 0xbf
    "11111111", -- 1227 - 0x4cb  :  255 - 0xff
    "11111111", -- 1228 - 0x4cc  :  255 - 0xff
    "11111111", -- 1229 - 0x4cd  :  255 - 0xff
    "11111111", -- 1230 - 0x4ce  :  255 - 0xff
    "11111111", -- 1231 - 0x4cf  :  255 - 0xff
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Background 0x9a
    "10111100", -- 1233 - 0x4d1  :  188 - 0xbc
    "11111110", -- 1234 - 0x4d2  :  254 - 0xfe
    "11111110", -- 1235 - 0x4d3  :  254 - 0xfe
    "11111110", -- 1236 - 0x4d4  :  254 - 0xfe
    "11111110", -- 1237 - 0x4d5  :  254 - 0xfe
    "11111110", -- 1238 - 0x4d6  :  254 - 0xfe
    "11111110", -- 1239 - 0x4d7  :  254 - 0xfe
    "11111110", -- 1240 - 0x4d8  :  254 - 0xfe -- Background 0x9b
    "11111110", -- 1241 - 0x4d9  :  254 - 0xfe
    "10111110", -- 1242 - 0x4da  :  190 - 0xbe
    "11111110", -- 1243 - 0x4db  :  254 - 0xfe
    "11111110", -- 1244 - 0x4dc  :  254 - 0xfe
    "11111110", -- 1245 - 0x4dd  :  254 - 0xfe
    "11111110", -- 1246 - 0x4de  :  254 - 0xfe
    "11111110", -- 1247 - 0x4df  :  254 - 0xfe
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0 -- Background 0x9c
    "00111111", -- 1249 - 0x4e1  :   63 - 0x3f
    "01011111", -- 1250 - 0x4e2  :   95 - 0x5f
    "01101111", -- 1251 - 0x4e3  :  111 - 0x6f
    "01110111", -- 1252 - 0x4e4  :  119 - 0x77
    "01111011", -- 1253 - 0x4e5  :  123 - 0x7b
    "00010101", -- 1254 - 0x4e6  :   21 - 0x15
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0 -- Background 0x9d
    "10111110", -- 1257 - 0x4e9  :  190 - 0xbe
    "11011110", -- 1258 - 0x4ea  :  222 - 0xde
    "11101110", -- 1259 - 0x4eb  :  238 - 0xee
    "11110110", -- 1260 - 0x4ec  :  246 - 0xf6
    "11111010", -- 1261 - 0x4ed  :  250 - 0xfa
    "01010100", -- 1262 - 0x4ee  :   84 - 0x54
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0 -- Background 0x9e
    "10111111", -- 1265 - 0x4f1  :  191 - 0xbf
    "11011111", -- 1266 - 0x4f2  :  223 - 0xdf
    "11101111", -- 1267 - 0x4f3  :  239 - 0xef
    "11110111", -- 1268 - 0x4f4  :  247 - 0xf7
    "11111011", -- 1269 - 0x4f5  :  251 - 0xfb
    "01010101", -- 1270 - 0x4f6  :   85 - 0x55
    "00000000", -- 1271 - 0x4f7  :    0 - 0x0
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- Background 0x9f
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- Background 0xa0
    "01111111", -- 1281 - 0x501  :  127 - 0x7f
    "00000000", -- 1282 - 0x502  :    0 - 0x0
    "00000001", -- 1283 - 0x503  :    1 - 0x1
    "00000001", -- 1284 - 0x504  :    1 - 0x1
    "00000001", -- 1285 - 0x505  :    1 - 0x1
    "00000001", -- 1286 - 0x506  :    1 - 0x1
    "00000001", -- 1287 - 0x507  :    1 - 0x1
    "00000001", -- 1288 - 0x508  :    1 - 0x1 -- Background 0xa1
    "00000001", -- 1289 - 0x509  :    1 - 0x1
    "00000001", -- 1290 - 0x50a  :    1 - 0x1
    "00000001", -- 1291 - 0x50b  :    1 - 0x1
    "00000001", -- 1292 - 0x50c  :    1 - 0x1
    "00000001", -- 1293 - 0x50d  :    1 - 0x1
    "00000001", -- 1294 - 0x50e  :    1 - 0x1
    "00000001", -- 1295 - 0x50f  :    1 - 0x1
    "00000000", -- 1296 - 0x510  :    0 - 0x0 -- Background 0xa2
    "11111110", -- 1297 - 0x511  :  254 - 0xfe
    "00000000", -- 1298 - 0x512  :    0 - 0x0
    "10000000", -- 1299 - 0x513  :  128 - 0x80
    "10000000", -- 1300 - 0x514  :  128 - 0x80
    "10000000", -- 1301 - 0x515  :  128 - 0x80
    "10000000", -- 1302 - 0x516  :  128 - 0x80
    "10000000", -- 1303 - 0x517  :  128 - 0x80
    "10000000", -- 1304 - 0x518  :  128 - 0x80 -- Background 0xa3
    "10000000", -- 1305 - 0x519  :  128 - 0x80
    "10000000", -- 1306 - 0x51a  :  128 - 0x80
    "10000000", -- 1307 - 0x51b  :  128 - 0x80
    "10000000", -- 1308 - 0x51c  :  128 - 0x80
    "10000000", -- 1309 - 0x51d  :  128 - 0x80
    "10000000", -- 1310 - 0x51e  :  128 - 0x80
    "10000000", -- 1311 - 0x51f  :  128 - 0x80
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Background 0xa4
    "00110000", -- 1313 - 0x521  :   48 - 0x30
    "00111000", -- 1314 - 0x522  :   56 - 0x38
    "01111000", -- 1315 - 0x523  :  120 - 0x78
    "01111100", -- 1316 - 0x524  :  124 - 0x7c
    "01111101", -- 1317 - 0x525  :  125 - 0x7d
    "00011101", -- 1318 - 0x526  :   29 - 0x1d
    "00001101", -- 1319 - 0x527  :   13 - 0xd
    "00001101", -- 1320 - 0x528  :   13 - 0xd -- Background 0xa5
    "00011101", -- 1321 - 0x529  :   29 - 0x1d
    "00111101", -- 1322 - 0x52a  :   61 - 0x3d
    "00111111", -- 1323 - 0x52b  :   63 - 0x3f
    "00111111", -- 1324 - 0x52c  :   63 - 0x3f
    "00011111", -- 1325 - 0x52d  :   31 - 0x1f
    "00000001", -- 1326 - 0x52e  :    1 - 0x1
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Background 0xa6
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "11100000", -- 1330 - 0x532  :  224 - 0xe0
    "11111000", -- 1331 - 0x533  :  248 - 0xf8
    "11111000", -- 1332 - 0x534  :  248 - 0xf8
    "11110000", -- 1333 - 0x535  :  240 - 0xf0
    "11000000", -- 1334 - 0x536  :  192 - 0xc0
    "11000000", -- 1335 - 0x537  :  192 - 0xc0
    "11000000", -- 1336 - 0x538  :  192 - 0xc0 -- Background 0xa7
    "11110000", -- 1337 - 0x539  :  240 - 0xf0
    "11110000", -- 1338 - 0x53a  :  240 - 0xf0
    "11000000", -- 1339 - 0x53b  :  192 - 0xc0
    "11000000", -- 1340 - 0x53c  :  192 - 0xc0
    "11000000", -- 1341 - 0x53d  :  192 - 0xc0
    "11000000", -- 1342 - 0x53e  :  192 - 0xc0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Background 0xa8
    "01100000", -- 1345 - 0x541  :   96 - 0x60
    "01100000", -- 1346 - 0x542  :   96 - 0x60
    "01100000", -- 1347 - 0x543  :   96 - 0x60
    "01100000", -- 1348 - 0x544  :   96 - 0x60
    "01100000", -- 1349 - 0x545  :   96 - 0x60
    "01100000", -- 1350 - 0x546  :   96 - 0x60
    "01100000", -- 1351 - 0x547  :   96 - 0x60
    "01100000", -- 1352 - 0x548  :   96 - 0x60 -- Background 0xa9
    "01100000", -- 1353 - 0x549  :   96 - 0x60
    "01100000", -- 1354 - 0x54a  :   96 - 0x60
    "01100000", -- 1355 - 0x54b  :   96 - 0x60
    "01100000", -- 1356 - 0x54c  :   96 - 0x60
    "01100000", -- 1357 - 0x54d  :   96 - 0x60
    "01100000", -- 1358 - 0x54e  :   96 - 0x60
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Background 0xaa
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- Background 0xab
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Background 0xac
    "00000110", -- 1377 - 0x561  :    6 - 0x6
    "00000110", -- 1378 - 0x562  :    6 - 0x6
    "00000110", -- 1379 - 0x563  :    6 - 0x6
    "00000110", -- 1380 - 0x564  :    6 - 0x6
    "00000110", -- 1381 - 0x565  :    6 - 0x6
    "00000110", -- 1382 - 0x566  :    6 - 0x6
    "00000110", -- 1383 - 0x567  :    6 - 0x6
    "00000110", -- 1384 - 0x568  :    6 - 0x6 -- Background 0xad
    "00000110", -- 1385 - 0x569  :    6 - 0x6
    "00000110", -- 1386 - 0x56a  :    6 - 0x6
    "00000110", -- 1387 - 0x56b  :    6 - 0x6
    "00000110", -- 1388 - 0x56c  :    6 - 0x6
    "00000110", -- 1389 - 0x56d  :    6 - 0x6
    "00000110", -- 1390 - 0x56e  :    6 - 0x6
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Background 0xae
    "00000001", -- 1393 - 0x571  :    1 - 0x1
    "00000011", -- 1394 - 0x572  :    3 - 0x3
    "00000010", -- 1395 - 0x573  :    2 - 0x2
    "00000010", -- 1396 - 0x574  :    2 - 0x2
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000011", -- 1398 - 0x576  :    3 - 0x3
    "00000010", -- 1399 - 0x577  :    2 - 0x2
    "00000001", -- 1400 - 0x578  :    1 - 0x1 -- Background 0xaf
    "00000011", -- 1401 - 0x579  :    3 - 0x3
    "00000101", -- 1402 - 0x57a  :    5 - 0x5
    "00000100", -- 1403 - 0x57b  :    4 - 0x4
    "00000101", -- 1404 - 0x57c  :    5 - 0x5
    "00001101", -- 1405 - 0x57d  :   13 - 0xd
    "00001100", -- 1406 - 0x57e  :   12 - 0xc
    "00000001", -- 1407 - 0x57f  :    1 - 0x1
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Background 0xb0
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "01000000", -- 1410 - 0x582  :   64 - 0x40
    "11110000", -- 1411 - 0x583  :  240 - 0xf0
    "11101000", -- 1412 - 0x584  :  232 - 0xe8
    "10010000", -- 1413 - 0x585  :  144 - 0x90
    "01010000", -- 1414 - 0x586  :   80 - 0x50
    "11010000", -- 1415 - 0x587  :  208 - 0xd0
    "11111000", -- 1416 - 0x588  :  248 - 0xf8 -- Background 0xb1
    "11000000", -- 1417 - 0x589  :  192 - 0xc0
    "11100000", -- 1418 - 0x58a  :  224 - 0xe0
    "01000000", -- 1419 - 0x58b  :   64 - 0x40
    "10000000", -- 1420 - 0x58c  :  128 - 0x80
    "11000000", -- 1421 - 0x58d  :  192 - 0xc0
    "11100000", -- 1422 - 0x58e  :  224 - 0xe0
    "01110000", -- 1423 - 0x58f  :  112 - 0x70
    "00000001", -- 1424 - 0x590  :    1 - 0x1 -- Background 0xb2
    "00001101", -- 1425 - 0x591  :   13 - 0xd
    "00001101", -- 1426 - 0x592  :   13 - 0xd
    "00000011", -- 1427 - 0x593  :    3 - 0x3
    "00000011", -- 1428 - 0x594  :    3 - 0x3
    "00000111", -- 1429 - 0x595  :    7 - 0x7
    "00000111", -- 1430 - 0x596  :    7 - 0x7
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00111111", -- 1432 - 0x598  :   63 - 0x3f -- Background 0xb3
    "00111111", -- 1433 - 0x599  :   63 - 0x3f
    "00111111", -- 1434 - 0x59a  :   63 - 0x3f
    "00111111", -- 1435 - 0x59b  :   63 - 0x3f
    "00111111", -- 1436 - 0x59c  :   63 - 0x3f
    "00111111", -- 1437 - 0x59d  :   63 - 0x3f
    "00110101", -- 1438 - 0x59e  :   53 - 0x35
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "10110000", -- 1440 - 0x5a0  :  176 - 0xb0 -- Background 0xb4
    "11000000", -- 1441 - 0x5a1  :  192 - 0xc0
    "11100000", -- 1442 - 0x5a2  :  224 - 0xe0
    "11100000", -- 1443 - 0x5a3  :  224 - 0xe0
    "11110000", -- 1444 - 0x5a4  :  240 - 0xf0
    "11110000", -- 1445 - 0x5a5  :  240 - 0xf0
    "11110000", -- 1446 - 0x5a6  :  240 - 0xf0
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "11111100", -- 1448 - 0x5a8  :  252 - 0xfc -- Background 0xb5
    "11111000", -- 1449 - 0x5a9  :  248 - 0xf8
    "11111100", -- 1450 - 0x5aa  :  252 - 0xfc
    "11111000", -- 1451 - 0x5ab  :  248 - 0xf8
    "11111100", -- 1452 - 0x5ac  :  252 - 0xfc
    "11111000", -- 1453 - 0x5ad  :  248 - 0xf8
    "01010100", -- 1454 - 0x5ae  :   84 - 0x54
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Background 0xb6
    "01111111", -- 1457 - 0x5b1  :  127 - 0x7f
    "01111111", -- 1458 - 0x5b2  :  127 - 0x7f
    "01111111", -- 1459 - 0x5b3  :  127 - 0x7f
    "01111111", -- 1460 - 0x5b4  :  127 - 0x7f
    "01111111", -- 1461 - 0x5b5  :  127 - 0x7f
    "01101010", -- 1462 - 0x5b6  :  106 - 0x6a
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0 -- Background 0xb7
    "01111011", -- 1465 - 0x5b9  :  123 - 0x7b
    "01110011", -- 1466 - 0x5ba  :  115 - 0x73
    "01111011", -- 1467 - 0x5bb  :  123 - 0x7b
    "01110011", -- 1468 - 0x5bc  :  115 - 0x73
    "01111011", -- 1469 - 0x5bd  :  123 - 0x7b
    "01010011", -- 1470 - 0x5be  :   83 - 0x53
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Background 0xb8
    "11011110", -- 1473 - 0x5c1  :  222 - 0xde
    "10011110", -- 1474 - 0x5c2  :  158 - 0x9e
    "11011100", -- 1475 - 0x5c3  :  220 - 0xdc
    "10011110", -- 1476 - 0x5c4  :  158 - 0x9e
    "11011100", -- 1477 - 0x5c5  :  220 - 0xdc
    "10011010", -- 1478 - 0x5c6  :  154 - 0x9a
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0 -- Background 0xb9
    "11111110", -- 1481 - 0x5c9  :  254 - 0xfe
    "11111100", -- 1482 - 0x5ca  :  252 - 0xfc
    "11111110", -- 1483 - 0x5cb  :  254 - 0xfe
    "11111100", -- 1484 - 0x5cc  :  252 - 0xfc
    "11111110", -- 1485 - 0x5cd  :  254 - 0xfe
    "01010100", -- 1486 - 0x5ce  :   84 - 0x54
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Background 0xba
    "01111111", -- 1489 - 0x5d1  :  127 - 0x7f
    "01111111", -- 1490 - 0x5d2  :  127 - 0x7f
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "01111111", -- 1492 - 0x5d4  :  127 - 0x7f
    "01111111", -- 1493 - 0x5d5  :  127 - 0x7f
    "01101010", -- 1494 - 0x5d6  :  106 - 0x6a
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0 -- Background 0xbb
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Background 0xbc
    "11111110", -- 1505 - 0x5e1  :  254 - 0xfe
    "11111110", -- 1506 - 0x5e2  :  254 - 0xfe
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "10011110", -- 1508 - 0x5e4  :  158 - 0x9e
    "11011100", -- 1509 - 0x5e5  :  220 - 0xdc
    "10011010", -- 1510 - 0x5e6  :  154 - 0x9a
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- Background 0xbd
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00000000", -- 1514 - 0x5ea  :    0 - 0x0
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "00000000", -- 1516 - 0x5ec  :    0 - 0x0
    "00000000", -- 1517 - 0x5ed  :    0 - 0x0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Background 0xbe
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Background 0xbf
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000000", -- 1542 - 0x606  :    0 - 0x0
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00000000", -- 1544 - 0x608  :    0 - 0x0 -- Background 0xc1
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- Background 0xc3
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Background 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0 -- Background 0xc5
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000000", -- 1578 - 0x62a  :    0 - 0x0
    "00000001", -- 1579 - 0x62b  :    1 - 0x1
    "00000111", -- 1580 - 0x62c  :    7 - 0x7
    "00001111", -- 1581 - 0x62d  :   15 - 0xf
    "00001111", -- 1582 - 0x62e  :   15 - 0xf
    "00011111", -- 1583 - 0x62f  :   31 - 0x1f
    "00000000", -- 1584 - 0x630  :    0 - 0x0 -- Background 0xc6
    "00011111", -- 1585 - 0x631  :   31 - 0x1f
    "01111111", -- 1586 - 0x632  :  127 - 0x7f
    "11111111", -- 1587 - 0x633  :  255 - 0xff
    "11111111", -- 1588 - 0x634  :  255 - 0xff
    "11111111", -- 1589 - 0x635  :  255 - 0xff
    "11111111", -- 1590 - 0x636  :  255 - 0xff
    "11111111", -- 1591 - 0x637  :  255 - 0xff
    "00011111", -- 1592 - 0x638  :   31 - 0x1f -- Background 0xc7
    "00111111", -- 1593 - 0x639  :   63 - 0x3f
    "00111111", -- 1594 - 0x63a  :   63 - 0x3f
    "01111111", -- 1595 - 0x63b  :  127 - 0x7f
    "01111111", -- 1596 - 0x63c  :  127 - 0x7f
    "01111111", -- 1597 - 0x63d  :  127 - 0x7f
    "01111111", -- 1598 - 0x63e  :  127 - 0x7f
    "01111111", -- 1599 - 0x63f  :  127 - 0x7f
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Background 0xc8
    "11111111", -- 1601 - 0x641  :  255 - 0xff
    "11111111", -- 1602 - 0x642  :  255 - 0xff
    "11111111", -- 1603 - 0x643  :  255 - 0xff
    "11111111", -- 1604 - 0x644  :  255 - 0xff
    "11111111", -- 1605 - 0x645  :  255 - 0xff
    "11111111", -- 1606 - 0x646  :  255 - 0xff
    "11111111", -- 1607 - 0x647  :  255 - 0xff
    "11101000", -- 1608 - 0x648  :  232 - 0xe8 -- Background 0xc9
    "11010100", -- 1609 - 0x649  :  212 - 0xd4
    "11101000", -- 1610 - 0x64a  :  232 - 0xe8
    "11010100", -- 1611 - 0x64b  :  212 - 0xd4
    "11101010", -- 1612 - 0x64c  :  234 - 0xea
    "11010100", -- 1613 - 0x64d  :  212 - 0xd4
    "11101010", -- 1614 - 0x64e  :  234 - 0xea
    "11010100", -- 1615 - 0x64f  :  212 - 0xd4
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Background 0xca
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "00000000", -- 1622 - 0x656  :    0 - 0x0
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- Background 0xcb
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000101", -- 1636 - 0x664  :    5 - 0x5
    "00000010", -- 1637 - 0x665  :    2 - 0x2
    "00000001", -- 1638 - 0x666  :    1 - 0x1
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "10000000", -- 1643 - 0x66b  :  128 - 0x80
    "01010000", -- 1644 - 0x66c  :   80 - 0x50
    "10100000", -- 1645 - 0x66d  :  160 - 0xa0
    "01000000", -- 1646 - 0x66e  :   64 - 0x40
    "10000000", -- 1647 - 0x66f  :  128 - 0x80
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Background 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00110000", -- 1652 - 0x674  :   48 - 0x30
    "01111111", -- 1653 - 0x675  :  127 - 0x7f
    "00110000", -- 1654 - 0x676  :   48 - 0x30
    "00110000", -- 1655 - 0x677  :   48 - 0x30
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00001100", -- 1660 - 0x67c  :   12 - 0xc
    "11111110", -- 1661 - 0x67d  :  254 - 0xfe
    "00001100", -- 1662 - 0x67e  :   12 - 0xc
    "00001100", -- 1663 - 0x67f  :   12 - 0xc
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Background 0xd0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- Background 0xd1
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00000111", -- 1680 - 0x690  :    7 - 0x7 -- Background 0xd2
    "00000111", -- 1681 - 0x691  :    7 - 0x7
    "00000111", -- 1682 - 0x692  :    7 - 0x7
    "00000111", -- 1683 - 0x693  :    7 - 0x7
    "00000111", -- 1684 - 0x694  :    7 - 0x7
    "00000111", -- 1685 - 0x695  :    7 - 0x7
    "00000111", -- 1686 - 0x696  :    7 - 0x7
    "00000111", -- 1687 - 0x697  :    7 - 0x7
    "11100000", -- 1688 - 0x698  :  224 - 0xe0 -- Background 0xd3
    "11100000", -- 1689 - 0x699  :  224 - 0xe0
    "11000000", -- 1690 - 0x69a  :  192 - 0xc0
    "11100000", -- 1691 - 0x69b  :  224 - 0xe0
    "10100000", -- 1692 - 0x69c  :  160 - 0xa0
    "11100000", -- 1693 - 0x69d  :  224 - 0xe0
    "11000000", -- 1694 - 0x69e  :  192 - 0xc0
    "11100000", -- 1695 - 0x69f  :  224 - 0xe0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0 -- Background 0xd5
    "11111000", -- 1705 - 0x6a9  :  248 - 0xf8
    "11111110", -- 1706 - 0x6aa  :  254 - 0xfe
    "11111111", -- 1707 - 0x6ab  :  255 - 0xff
    "11111111", -- 1708 - 0x6ac  :  255 - 0xff
    "11111111", -- 1709 - 0x6ad  :  255 - 0xff
    "11111111", -- 1710 - 0x6ae  :  255 - 0xff
    "11111111", -- 1711 - 0x6af  :  255 - 0xff
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "10000000", -- 1715 - 0x6b3  :  128 - 0x80
    "10100000", -- 1716 - 0x6b4  :  160 - 0xa0
    "01010000", -- 1717 - 0x6b5  :   80 - 0x50
    "10100000", -- 1718 - 0x6b6  :  160 - 0xa0
    "11010000", -- 1719 - 0x6b7  :  208 - 0xd0
    "01111111", -- 1720 - 0x6b8  :  127 - 0x7f -- Background 0xd7
    "01111111", -- 1721 - 0x6b9  :  127 - 0x7f
    "01111111", -- 1722 - 0x6ba  :  127 - 0x7f
    "00111111", -- 1723 - 0x6bb  :   63 - 0x3f
    "00111111", -- 1724 - 0x6bc  :   63 - 0x3f
    "00001111", -- 1725 - 0x6bd  :   15 - 0xf
    "00000111", -- 1726 - 0x6be  :    7 - 0x7
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "11111111", -- 1728 - 0x6c0  :  255 - 0xff -- Background 0xd8
    "11111111", -- 1729 - 0x6c1  :  255 - 0xff
    "11111111", -- 1730 - 0x6c2  :  255 - 0xff
    "11111111", -- 1731 - 0x6c3  :  255 - 0xff
    "11111111", -- 1732 - 0x6c4  :  255 - 0xff
    "11111111", -- 1733 - 0x6c5  :  255 - 0xff
    "11111111", -- 1734 - 0x6c6  :  255 - 0xff
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "11101010", -- 1736 - 0x6c8  :  234 - 0xea -- Background 0xd9
    "11010100", -- 1737 - 0x6c9  :  212 - 0xd4
    "11101010", -- 1738 - 0x6ca  :  234 - 0xea
    "11010100", -- 1739 - 0x6cb  :  212 - 0xd4
    "10101000", -- 1740 - 0x6cc  :  168 - 0xa8
    "01010000", -- 1741 - 0x6cd  :   80 - 0x50
    "10100000", -- 1742 - 0x6ce  :  160 - 0xa0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Background 0xda
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00001100", -- 1746 - 0x6d2  :   12 - 0xc
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0 -- Background 0xdb
    "10000000", -- 1753 - 0x6d9  :  128 - 0x80
    "10000000", -- 1754 - 0x6da  :  128 - 0x80
    "10000000", -- 1755 - 0x6db  :  128 - 0x80
    "10011000", -- 1756 - 0x6dc  :  152 - 0x98
    "10000000", -- 1757 - 0x6dd  :  128 - 0x80
    "10000000", -- 1758 - 0x6de  :  128 - 0x80
    "10000000", -- 1759 - 0x6df  :  128 - 0x80
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000010", -- 1764 - 0x6e4  :    2 - 0x2
    "00000011", -- 1765 - 0x6e5  :    3 - 0x3
    "00000011", -- 1766 - 0x6e6  :    3 - 0x3
    "00000001", -- 1767 - 0x6e7  :    1 - 0x1
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- Background 0xdd
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "10100000", -- 1772 - 0x6ec  :  160 - 0xa0
    "11100000", -- 1773 - 0x6ed  :  224 - 0xe0
    "11100000", -- 1774 - 0x6ee  :  224 - 0xe0
    "11000000", -- 1775 - 0x6ef  :  192 - 0xc0
    "00110000", -- 1776 - 0x6f0  :   48 - 0x30 -- Background 0xde
    "01111111", -- 1777 - 0x6f1  :  127 - 0x7f
    "00110000", -- 1778 - 0x6f2  :   48 - 0x30
    "00110000", -- 1779 - 0x6f3  :   48 - 0x30
    "00110000", -- 1780 - 0x6f4  :   48 - 0x30
    "00110000", -- 1781 - 0x6f5  :   48 - 0x30
    "00110000", -- 1782 - 0x6f6  :   48 - 0x30
    "00110000", -- 1783 - 0x6f7  :   48 - 0x30
    "00001100", -- 1784 - 0x6f8  :   12 - 0xc -- Background 0xdf
    "11111110", -- 1785 - 0x6f9  :  254 - 0xfe
    "00001100", -- 1786 - 0x6fa  :   12 - 0xc
    "00001100", -- 1787 - 0x6fb  :   12 - 0xc
    "00001100", -- 1788 - 0x6fc  :   12 - 0xc
    "00001100", -- 1789 - 0x6fd  :   12 - 0xc
    "00001100", -- 1790 - 0x6fe  :   12 - 0xc
    "00001100", -- 1791 - 0x6ff  :   12 - 0xc
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Background 0xe0
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0 -- Background 0xe1
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0 -- Background 0xe2
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000000", -- 1816 - 0x718  :    0 - 0x0 -- Background 0xe3
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Background 0xe4
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000000", -- 1828 - 0x724  :    0 - 0x0
    "00000000", -- 1829 - 0x725  :    0 - 0x0
    "00000000", -- 1830 - 0x726  :    0 - 0x0
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- Background 0xe5
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "00000000", -- 1840 - 0x730  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "00000000", -- 1845 - 0x735  :    0 - 0x0
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0 -- Background 0xe7
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0 -- Background 0xe9
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Background 0xea
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- Background 0xeb
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Background 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0 -- Background 0xed
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Background 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- Background 0xef
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- Background 0xf1
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Background 0xf2
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- Background 0xf3
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Background 0xf4
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0 -- Background 0xf5
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Background 0xf6
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- Background 0xf7
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Background 0xf8
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- Background 0xf9
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Background 0xfa
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- Background 0xfb
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Background 0xfc
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- Background 0xfd
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Background 0xfe
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Background 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
