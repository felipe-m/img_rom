//-   Sprites Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: smario_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_SMARIO_SPR
  (
     //input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table both color planes
      12'h0: dout  = 8'b00000011; //    0 :   3 - 0x3 -- Sprite 0x0
      12'h1: dout  = 8'b00001111; //    1 :  15 - 0xf
      12'h2: dout  = 8'b00011111; //    2 :  31 - 0x1f
      12'h3: dout  = 8'b00011111; //    3 :  31 - 0x1f
      12'h4: dout  = 8'b00011100; //    4 :  28 - 0x1c
      12'h5: dout  = 8'b00100100; //    5 :  36 - 0x24
      12'h6: dout  = 8'b00100110; //    6 :  38 - 0x26
      12'h7: dout  = 8'b01100110; //    7 : 102 - 0x66
      12'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- plane 1
      12'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      12'hA: dout  = 8'b00000000; //   10 :   0 - 0x0
      12'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      12'hC: dout  = 8'b00011111; //   12 :  31 - 0x1f
      12'hD: dout  = 8'b00111111; //   13 :  63 - 0x3f
      12'hE: dout  = 8'b00111111; //   14 :  63 - 0x3f
      12'hF: dout  = 8'b01111111; //   15 : 127 - 0x7f
      12'h10: dout  = 8'b11100000; //   16 : 224 - 0xe0 -- Sprite 0x1
      12'h11: dout  = 8'b11000000; //   17 : 192 - 0xc0
      12'h12: dout  = 8'b10000000; //   18 : 128 - 0x80
      12'h13: dout  = 8'b11111100; //   19 : 252 - 0xfc
      12'h14: dout  = 8'b10000000; //   20 : 128 - 0x80
      12'h15: dout  = 8'b11000000; //   21 : 192 - 0xc0
      12'h16: dout  = 8'b00000000; //   22 :   0 - 0x0
      12'h17: dout  = 8'b00100000; //   23 :  32 - 0x20
      12'h18: dout  = 8'b00000000; //   24 :   0 - 0x0 -- plane 1
      12'h19: dout  = 8'b00100000; //   25 :  32 - 0x20
      12'h1A: dout  = 8'b01100000; //   26 :  96 - 0x60
      12'h1B: dout  = 8'b00000000; //   27 :   0 - 0x0
      12'h1C: dout  = 8'b11110000; //   28 : 240 - 0xf0
      12'h1D: dout  = 8'b11111100; //   29 : 252 - 0xfc
      12'h1E: dout  = 8'b11111110; //   30 : 254 - 0xfe
      12'h1F: dout  = 8'b11111110; //   31 : 254 - 0xfe
      12'h20: dout  = 8'b01100000; //   32 :  96 - 0x60 -- Sprite 0x2
      12'h21: dout  = 8'b01110000; //   33 : 112 - 0x70
      12'h22: dout  = 8'b00011000; //   34 :  24 - 0x18
      12'h23: dout  = 8'b00000111; //   35 :   7 - 0x7
      12'h24: dout  = 8'b00001111; //   36 :  15 - 0xf
      12'h25: dout  = 8'b00011111; //   37 :  31 - 0x1f
      12'h26: dout  = 8'b00111111; //   38 :  63 - 0x3f
      12'h27: dout  = 8'b01111111; //   39 : 127 - 0x7f
      12'h28: dout  = 8'b01111111; //   40 : 127 - 0x7f -- plane 1
      12'h29: dout  = 8'b01111111; //   41 : 127 - 0x7f
      12'h2A: dout  = 8'b00011111; //   42 :  31 - 0x1f
      12'h2B: dout  = 8'b00000111; //   43 :   7 - 0x7
      12'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout  = 8'b00011110; //   45 :  30 - 0x1e
      12'h2E: dout  = 8'b00111111; //   46 :  63 - 0x3f
      12'h2F: dout  = 8'b01111111; //   47 : 127 - 0x7f
      12'h30: dout  = 8'b11111100; //   48 : 252 - 0xfc -- Sprite 0x3
      12'h31: dout  = 8'b01111100; //   49 : 124 - 0x7c
      12'h32: dout  = 8'b00000000; //   50 :   0 - 0x0
      12'h33: dout  = 8'b00000000; //   51 :   0 - 0x0
      12'h34: dout  = 8'b11100000; //   52 : 224 - 0xe0
      12'h35: dout  = 8'b11110000; //   53 : 240 - 0xf0
      12'h36: dout  = 8'b11111000; //   54 : 248 - 0xf8
      12'h37: dout  = 8'b11111000; //   55 : 248 - 0xf8
      12'h38: dout  = 8'b11111100; //   56 : 252 - 0xfc -- plane 1
      12'h39: dout  = 8'b11111100; //   57 : 252 - 0xfc
      12'h3A: dout  = 8'b11111000; //   58 : 248 - 0xf8
      12'h3B: dout  = 8'b11000000; //   59 : 192 - 0xc0
      12'h3C: dout  = 8'b11000010; //   60 : 194 - 0xc2
      12'h3D: dout  = 8'b01100111; //   61 : 103 - 0x67
      12'h3E: dout  = 8'b00101111; //   62 :  47 - 0x2f
      12'h3F: dout  = 8'b00110111; //   63 :  55 - 0x37
      12'h40: dout  = 8'b01111111; //   64 : 127 - 0x7f -- Sprite 0x4
      12'h41: dout  = 8'b01111111; //   65 : 127 - 0x7f
      12'h42: dout  = 8'b11111111; //   66 : 255 - 0xff
      12'h43: dout  = 8'b11111111; //   67 : 255 - 0xff
      12'h44: dout  = 8'b00000111; //   68 :   7 - 0x7
      12'h45: dout  = 8'b00000111; //   69 :   7 - 0x7
      12'h46: dout  = 8'b00001111; //   70 :  15 - 0xf
      12'h47: dout  = 8'b00001111; //   71 :  15 - 0xf
      12'h48: dout  = 8'b01111111; //   72 : 127 - 0x7f -- plane 1
      12'h49: dout  = 8'b01111110; //   73 : 126 - 0x7e
      12'h4A: dout  = 8'b11111100; //   74 : 252 - 0xfc
      12'h4B: dout  = 8'b11110000; //   75 : 240 - 0xf0
      12'h4C: dout  = 8'b11111000; //   76 : 248 - 0xf8
      12'h4D: dout  = 8'b11111000; //   77 : 248 - 0xf8
      12'h4E: dout  = 8'b11110000; //   78 : 240 - 0xf0
      12'h4F: dout  = 8'b01110000; //   79 : 112 - 0x70
      12'h50: dout  = 8'b11111101; //   80 : 253 - 0xfd -- Sprite 0x5
      12'h51: dout  = 8'b11111110; //   81 : 254 - 0xfe
      12'h52: dout  = 8'b10110100; //   82 : 180 - 0xb4
      12'h53: dout  = 8'b11111000; //   83 : 248 - 0xf8
      12'h54: dout  = 8'b11111000; //   84 : 248 - 0xf8
      12'h55: dout  = 8'b11111001; //   85 : 249 - 0xf9
      12'h56: dout  = 8'b11111011; //   86 : 251 - 0xfb
      12'h57: dout  = 8'b11111111; //   87 : 255 - 0xff
      12'h58: dout  = 8'b00110111; //   88 :  55 - 0x37 -- plane 1
      12'h59: dout  = 8'b00110110; //   89 :  54 - 0x36
      12'h5A: dout  = 8'b01011100; //   90 :  92 - 0x5c
      12'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      12'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      12'h5D: dout  = 8'b00000001; //   93 :   1 - 0x1
      12'h5E: dout  = 8'b00000011; //   94 :   3 - 0x3
      12'h5F: dout  = 8'b00011111; //   95 :  31 - 0x1f
      12'h60: dout  = 8'b00011111; //   96 :  31 - 0x1f -- Sprite 0x6
      12'h61: dout  = 8'b00111111; //   97 :  63 - 0x3f
      12'h62: dout  = 8'b11111111; //   98 : 255 - 0xff
      12'h63: dout  = 8'b11111111; //   99 : 255 - 0xff
      12'h64: dout  = 8'b11111100; //  100 : 252 - 0xfc
      12'h65: dout  = 8'b01110000; //  101 : 112 - 0x70
      12'h66: dout  = 8'b01110000; //  102 : 112 - 0x70
      12'h67: dout  = 8'b00111000; //  103 :  56 - 0x38
      12'h68: dout  = 8'b00001000; //  104 :   8 - 0x8 -- plane 1
      12'h69: dout  = 8'b00100100; //  105 :  36 - 0x24
      12'h6A: dout  = 8'b11100011; //  106 : 227 - 0xe3
      12'h6B: dout  = 8'b11110000; //  107 : 240 - 0xf0
      12'h6C: dout  = 8'b11111000; //  108 : 248 - 0xf8
      12'h6D: dout  = 8'b01110000; //  109 : 112 - 0x70
      12'h6E: dout  = 8'b01110000; //  110 : 112 - 0x70
      12'h6F: dout  = 8'b00111000; //  111 :  56 - 0x38
      12'h70: dout  = 8'b11111111; //  112 : 255 - 0xff -- Sprite 0x7
      12'h71: dout  = 8'b11111111; //  113 : 255 - 0xff
      12'h72: dout  = 8'b11111111; //  114 : 255 - 0xff
      12'h73: dout  = 8'b00011111; //  115 :  31 - 0x1f
      12'h74: dout  = 8'b00000000; //  116 :   0 - 0x0
      12'h75: dout  = 8'b00000000; //  117 :   0 - 0x0
      12'h76: dout  = 8'b00000000; //  118 :   0 - 0x0
      12'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      12'h78: dout  = 8'b00011111; //  120 :  31 - 0x1f -- plane 1
      12'h79: dout  = 8'b00011111; //  121 :  31 - 0x1f
      12'h7A: dout  = 8'b00011111; //  122 :  31 - 0x1f
      12'h7B: dout  = 8'b00011111; //  123 :  31 - 0x1f
      12'h7C: dout  = 8'b00000000; //  124 :   0 - 0x0
      12'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      12'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      12'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x8
      12'h81: dout  = 8'b00000000; //  129 :   0 - 0x0
      12'h82: dout  = 8'b00000001; //  130 :   1 - 0x1
      12'h83: dout  = 8'b00000111; //  131 :   7 - 0x7
      12'h84: dout  = 8'b00001111; //  132 :  15 - 0xf
      12'h85: dout  = 8'b00001111; //  133 :  15 - 0xf
      12'h86: dout  = 8'b00001110; //  134 :  14 - 0xe
      12'h87: dout  = 8'b00010010; //  135 :  18 - 0x12
      12'h88: dout  = 8'b00000000; //  136 :   0 - 0x0 -- plane 1
      12'h89: dout  = 8'b00000000; //  137 :   0 - 0x0
      12'h8A: dout  = 8'b00000000; //  138 :   0 - 0x0
      12'h8B: dout  = 8'b00000000; //  139 :   0 - 0x0
      12'h8C: dout  = 8'b00000000; //  140 :   0 - 0x0
      12'h8D: dout  = 8'b00000000; //  141 :   0 - 0x0
      12'h8E: dout  = 8'b00001111; //  142 :  15 - 0xf
      12'h8F: dout  = 8'b00011111; //  143 :  31 - 0x1f
      12'h90: dout  = 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x9
      12'h91: dout  = 8'b00000000; //  145 :   0 - 0x0
      12'h92: dout  = 8'b11110000; //  146 : 240 - 0xf0
      12'h93: dout  = 8'b11100000; //  147 : 224 - 0xe0
      12'h94: dout  = 8'b11000000; //  148 : 192 - 0xc0
      12'h95: dout  = 8'b11111110; //  149 : 254 - 0xfe
      12'h96: dout  = 8'b01000000; //  150 :  64 - 0x40
      12'h97: dout  = 8'b01100000; //  151 :  96 - 0x60
      12'h98: dout  = 8'b00000000; //  152 :   0 - 0x0 -- plane 1
      12'h99: dout  = 8'b00000000; //  153 :   0 - 0x0
      12'h9A: dout  = 8'b00000000; //  154 :   0 - 0x0
      12'h9B: dout  = 8'b00010000; //  155 :  16 - 0x10
      12'h9C: dout  = 8'b00110000; //  156 :  48 - 0x30
      12'h9D: dout  = 8'b00000000; //  157 :   0 - 0x0
      12'h9E: dout  = 8'b11111000; //  158 : 248 - 0xf8
      12'h9F: dout  = 8'b11111110; //  159 : 254 - 0xfe
      12'hA0: dout  = 8'b00010011; //  160 :  19 - 0x13 -- Sprite 0xa
      12'hA1: dout  = 8'b00110011; //  161 :  51 - 0x33
      12'hA2: dout  = 8'b00110000; //  162 :  48 - 0x30
      12'hA3: dout  = 8'b00011000; //  163 :  24 - 0x18
      12'hA4: dout  = 8'b00000100; //  164 :   4 - 0x4
      12'hA5: dout  = 8'b00001111; //  165 :  15 - 0xf
      12'hA6: dout  = 8'b00011111; //  166 :  31 - 0x1f
      12'hA7: dout  = 8'b00011111; //  167 :  31 - 0x1f
      12'hA8: dout  = 8'b00011111; //  168 :  31 - 0x1f -- plane 1
      12'hA9: dout  = 8'b00111111; //  169 :  63 - 0x3f
      12'hAA: dout  = 8'b00111111; //  170 :  63 - 0x3f
      12'hAB: dout  = 8'b00011111; //  171 :  31 - 0x1f
      12'hAC: dout  = 8'b00000111; //  172 :   7 - 0x7
      12'hAD: dout  = 8'b00001000; //  173 :   8 - 0x8
      12'hAE: dout  = 8'b00010111; //  174 :  23 - 0x17
      12'hAF: dout  = 8'b00010111; //  175 :  23 - 0x17
      12'hB0: dout  = 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0xb
      12'hB1: dout  = 8'b00010000; //  177 :  16 - 0x10
      12'hB2: dout  = 8'b01111110; //  178 : 126 - 0x7e
      12'hB3: dout  = 8'b00111110; //  179 :  62 - 0x3e
      12'hB4: dout  = 8'b00000000; //  180 :   0 - 0x0
      12'hB5: dout  = 8'b00000000; //  181 :   0 - 0x0
      12'hB6: dout  = 8'b11000000; //  182 : 192 - 0xc0
      12'hB7: dout  = 8'b11100000; //  183 : 224 - 0xe0
      12'hB8: dout  = 8'b11111111; //  184 : 255 - 0xff -- plane 1
      12'hB9: dout  = 8'b11111111; //  185 : 255 - 0xff
      12'hBA: dout  = 8'b11111110; //  186 : 254 - 0xfe
      12'hBB: dout  = 8'b11111110; //  187 : 254 - 0xfe
      12'hBC: dout  = 8'b11111100; //  188 : 252 - 0xfc
      12'hBD: dout  = 8'b11100000; //  189 : 224 - 0xe0
      12'hBE: dout  = 8'b01000000; //  190 :  64 - 0x40
      12'hBF: dout  = 8'b10100000; //  191 : 160 - 0xa0
      12'hC0: dout  = 8'b00111111; //  192 :  63 - 0x3f -- Sprite 0xc
      12'hC1: dout  = 8'b00111111; //  193 :  63 - 0x3f
      12'hC2: dout  = 8'b00111111; //  194 :  63 - 0x3f
      12'hC3: dout  = 8'b00011111; //  195 :  31 - 0x1f
      12'hC4: dout  = 8'b00011111; //  196 :  31 - 0x1f
      12'hC5: dout  = 8'b00011111; //  197 :  31 - 0x1f
      12'hC6: dout  = 8'b00011111; //  198 :  31 - 0x1f
      12'hC7: dout  = 8'b00011111; //  199 :  31 - 0x1f
      12'hC8: dout  = 8'b00110111; //  200 :  55 - 0x37 -- plane 1
      12'hC9: dout  = 8'b00100111; //  201 :  39 - 0x27
      12'hCA: dout  = 8'b00100011; //  202 :  35 - 0x23
      12'hCB: dout  = 8'b00000011; //  203 :   3 - 0x3
      12'hCC: dout  = 8'b00000001; //  204 :   1 - 0x1
      12'hCD: dout  = 8'b00000000; //  205 :   0 - 0x0
      12'hCE: dout  = 8'b00000000; //  206 :   0 - 0x0
      12'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      12'hD0: dout  = 8'b11110000; //  208 : 240 - 0xf0 -- Sprite 0xd
      12'hD1: dout  = 8'b11110000; //  209 : 240 - 0xf0
      12'hD2: dout  = 8'b11110000; //  210 : 240 - 0xf0
      12'hD3: dout  = 8'b11111000; //  211 : 248 - 0xf8
      12'hD4: dout  = 8'b11111000; //  212 : 248 - 0xf8
      12'hD5: dout  = 8'b11111000; //  213 : 248 - 0xf8
      12'hD6: dout  = 8'b11111000; //  214 : 248 - 0xf8
      12'hD7: dout  = 8'b11111000; //  215 : 248 - 0xf8
      12'hD8: dout  = 8'b11001100; //  216 : 204 - 0xcc -- plane 1
      12'hD9: dout  = 8'b11111111; //  217 : 255 - 0xff
      12'hDA: dout  = 8'b11111111; //  218 : 255 - 0xff
      12'hDB: dout  = 8'b11111111; //  219 : 255 - 0xff
      12'hDC: dout  = 8'b11111111; //  220 : 255 - 0xff
      12'hDD: dout  = 8'b01110000; //  221 : 112 - 0x70
      12'hDE: dout  = 8'b00000000; //  222 :   0 - 0x0
      12'hDF: dout  = 8'b00001000; //  223 :   8 - 0x8
      12'hE0: dout  = 8'b11111111; //  224 : 255 - 0xff -- Sprite 0xe
      12'hE1: dout  = 8'b11111111; //  225 : 255 - 0xff
      12'hE2: dout  = 8'b11111111; //  226 : 255 - 0xff
      12'hE3: dout  = 8'b11111110; //  227 : 254 - 0xfe
      12'hE4: dout  = 8'b11110000; //  228 : 240 - 0xf0
      12'hE5: dout  = 8'b11000000; //  229 : 192 - 0xc0
      12'hE6: dout  = 8'b10000000; //  230 : 128 - 0x80
      12'hE7: dout  = 8'b00000000; //  231 :   0 - 0x0
      12'hE8: dout  = 8'b11110000; //  232 : 240 - 0xf0 -- plane 1
      12'hE9: dout  = 8'b11110000; //  233 : 240 - 0xf0
      12'hEA: dout  = 8'b11110000; //  234 : 240 - 0xf0
      12'hEB: dout  = 8'b11110000; //  235 : 240 - 0xf0
      12'hEC: dout  = 8'b11110000; //  236 : 240 - 0xf0
      12'hED: dout  = 8'b11000000; //  237 : 192 - 0xc0
      12'hEE: dout  = 8'b10000000; //  238 : 128 - 0x80
      12'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      12'hF0: dout  = 8'b11111100; //  240 : 252 - 0xfc -- Sprite 0xf
      12'hF1: dout  = 8'b11111100; //  241 : 252 - 0xfc
      12'hF2: dout  = 8'b11111000; //  242 : 248 - 0xf8
      12'hF3: dout  = 8'b01111000; //  243 : 120 - 0x78
      12'hF4: dout  = 8'b01111000; //  244 : 120 - 0x78
      12'hF5: dout  = 8'b01111000; //  245 : 120 - 0x78
      12'hF6: dout  = 8'b01111110; //  246 : 126 - 0x7e
      12'hF7: dout  = 8'b01111110; //  247 : 126 - 0x7e
      12'hF8: dout  = 8'b00010000; //  248 :  16 - 0x10 -- plane 1
      12'hF9: dout  = 8'b01100000; //  249 :  96 - 0x60
      12'hFA: dout  = 8'b10000000; //  250 : 128 - 0x80
      12'hFB: dout  = 8'b00000000; //  251 :   0 - 0x0
      12'hFC: dout  = 8'b01111000; //  252 : 120 - 0x78
      12'hFD: dout  = 8'b01111000; //  253 : 120 - 0x78
      12'hFE: dout  = 8'b01111110; //  254 : 126 - 0x7e
      12'hFF: dout  = 8'b01111110; //  255 : 126 - 0x7e
      12'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x10
      12'h101: dout  = 8'b00000011; //  257 :   3 - 0x3
      12'h102: dout  = 8'b00001111; //  258 :  15 - 0xf
      12'h103: dout  = 8'b00011111; //  259 :  31 - 0x1f
      12'h104: dout  = 8'b00011111; //  260 :  31 - 0x1f
      12'h105: dout  = 8'b00011100; //  261 :  28 - 0x1c
      12'h106: dout  = 8'b00100100; //  262 :  36 - 0x24
      12'h107: dout  = 8'b00100110; //  263 :  38 - 0x26
      12'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- plane 1
      12'h109: dout  = 8'b00000000; //  265 :   0 - 0x0
      12'h10A: dout  = 8'b00000000; //  266 :   0 - 0x0
      12'h10B: dout  = 8'b00000000; //  267 :   0 - 0x0
      12'h10C: dout  = 8'b00000000; //  268 :   0 - 0x0
      12'h10D: dout  = 8'b00011111; //  269 :  31 - 0x1f
      12'h10E: dout  = 8'b00111111; //  270 :  63 - 0x3f
      12'h10F: dout  = 8'b00111111; //  271 :  63 - 0x3f
      12'h110: dout  = 8'b00000000; //  272 :   0 - 0x0 -- Sprite 0x11
      12'h111: dout  = 8'b11100000; //  273 : 224 - 0xe0
      12'h112: dout  = 8'b11000000; //  274 : 192 - 0xc0
      12'h113: dout  = 8'b10000000; //  275 : 128 - 0x80
      12'h114: dout  = 8'b11111100; //  276 : 252 - 0xfc
      12'h115: dout  = 8'b10000000; //  277 : 128 - 0x80
      12'h116: dout  = 8'b11000000; //  278 : 192 - 0xc0
      12'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      12'h118: dout  = 8'b00000000; //  280 :   0 - 0x0 -- plane 1
      12'h119: dout  = 8'b00000000; //  281 :   0 - 0x0
      12'h11A: dout  = 8'b00100000; //  282 :  32 - 0x20
      12'h11B: dout  = 8'b01100000; //  283 :  96 - 0x60
      12'h11C: dout  = 8'b00000000; //  284 :   0 - 0x0
      12'h11D: dout  = 8'b11110000; //  285 : 240 - 0xf0
      12'h11E: dout  = 8'b11111100; //  286 : 252 - 0xfc
      12'h11F: dout  = 8'b11111110; //  287 : 254 - 0xfe
      12'h120: dout  = 8'b01100110; //  288 : 102 - 0x66 -- Sprite 0x12
      12'h121: dout  = 8'b01100000; //  289 :  96 - 0x60
      12'h122: dout  = 8'b00110000; //  290 :  48 - 0x30
      12'h123: dout  = 8'b00011000; //  291 :  24 - 0x18
      12'h124: dout  = 8'b00001111; //  292 :  15 - 0xf
      12'h125: dout  = 8'b00011111; //  293 :  31 - 0x1f
      12'h126: dout  = 8'b00111111; //  294 :  63 - 0x3f
      12'h127: dout  = 8'b00111111; //  295 :  63 - 0x3f
      12'h128: dout  = 8'b01111111; //  296 : 127 - 0x7f -- plane 1
      12'h129: dout  = 8'b01111111; //  297 : 127 - 0x7f
      12'h12A: dout  = 8'b00111111; //  298 :  63 - 0x3f
      12'h12B: dout  = 8'b00011111; //  299 :  31 - 0x1f
      12'h12C: dout  = 8'b00000000; //  300 :   0 - 0x0
      12'h12D: dout  = 8'b00010110; //  301 :  22 - 0x16
      12'h12E: dout  = 8'b00101111; //  302 :  47 - 0x2f
      12'h12F: dout  = 8'b00101111; //  303 :  47 - 0x2f
      12'h130: dout  = 8'b00100000; //  304 :  32 - 0x20 -- Sprite 0x13
      12'h131: dout  = 8'b11111100; //  305 : 252 - 0xfc
      12'h132: dout  = 8'b01111100; //  306 : 124 - 0x7c
      12'h133: dout  = 8'b00000000; //  307 :   0 - 0x0
      12'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      12'h135: dout  = 8'b11100000; //  309 : 224 - 0xe0
      12'h136: dout  = 8'b11100000; //  310 : 224 - 0xe0
      12'h137: dout  = 8'b11110000; //  311 : 240 - 0xf0
      12'h138: dout  = 8'b11111110; //  312 : 254 - 0xfe -- plane 1
      12'h139: dout  = 8'b11111100; //  313 : 252 - 0xfc
      12'h13A: dout  = 8'b11111100; //  314 : 252 - 0xfc
      12'h13B: dout  = 8'b11111000; //  315 : 248 - 0xf8
      12'h13C: dout  = 8'b11000000; //  316 : 192 - 0xc0
      12'h13D: dout  = 8'b01100000; //  317 :  96 - 0x60
      12'h13E: dout  = 8'b00100000; //  318 :  32 - 0x20
      12'h13F: dout  = 8'b00110000; //  319 :  48 - 0x30
      12'h140: dout  = 8'b00111111; //  320 :  63 - 0x3f -- Sprite 0x14
      12'h141: dout  = 8'b00111111; //  321 :  63 - 0x3f
      12'h142: dout  = 8'b00111111; //  322 :  63 - 0x3f
      12'h143: dout  = 8'b00111111; //  323 :  63 - 0x3f
      12'h144: dout  = 8'b00111111; //  324 :  63 - 0x3f
      12'h145: dout  = 8'b00111111; //  325 :  63 - 0x3f
      12'h146: dout  = 8'b00111111; //  326 :  63 - 0x3f
      12'h147: dout  = 8'b00011111; //  327 :  31 - 0x1f
      12'h148: dout  = 8'b00101111; //  328 :  47 - 0x2f -- plane 1
      12'h149: dout  = 8'b00101111; //  329 :  47 - 0x2f
      12'h14A: dout  = 8'b00101111; //  330 :  47 - 0x2f
      12'h14B: dout  = 8'b00001111; //  331 :  15 - 0xf
      12'h14C: dout  = 8'b00000111; //  332 :   7 - 0x7
      12'h14D: dout  = 8'b00000011; //  333 :   3 - 0x3
      12'h14E: dout  = 8'b00000000; //  334 :   0 - 0x0
      12'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      12'h150: dout  = 8'b11110000; //  336 : 240 - 0xf0 -- Sprite 0x15
      12'h151: dout  = 8'b10010000; //  337 : 144 - 0x90
      12'h152: dout  = 8'b00000000; //  338 :   0 - 0x0
      12'h153: dout  = 8'b00001000; //  339 :   8 - 0x8
      12'h154: dout  = 8'b00001100; //  340 :  12 - 0xc
      12'h155: dout  = 8'b00011100; //  341 :  28 - 0x1c
      12'h156: dout  = 8'b11111100; //  342 : 252 - 0xfc
      12'h157: dout  = 8'b11111000; //  343 : 248 - 0xf8
      12'h158: dout  = 8'b00010000; //  344 :  16 - 0x10 -- plane 1
      12'h159: dout  = 8'b11110000; //  345 : 240 - 0xf0
      12'h15A: dout  = 8'b11110000; //  346 : 240 - 0xf0
      12'h15B: dout  = 8'b11110000; //  347 : 240 - 0xf0
      12'h15C: dout  = 8'b11110000; //  348 : 240 - 0xf0
      12'h15D: dout  = 8'b11100000; //  349 : 224 - 0xe0
      12'h15E: dout  = 8'b11000000; //  350 : 192 - 0xc0
      12'h15F: dout  = 8'b11100000; //  351 : 224 - 0xe0
      12'h160: dout  = 8'b00001111; //  352 :  15 - 0xf -- Sprite 0x16
      12'h161: dout  = 8'b00001111; //  353 :  15 - 0xf
      12'h162: dout  = 8'b00000111; //  354 :   7 - 0x7
      12'h163: dout  = 8'b00000111; //  355 :   7 - 0x7
      12'h164: dout  = 8'b00000111; //  356 :   7 - 0x7
      12'h165: dout  = 8'b00001111; //  357 :  15 - 0xf
      12'h166: dout  = 8'b00001111; //  358 :  15 - 0xf
      12'h167: dout  = 8'b00000011; //  359 :   3 - 0x3
      12'h168: dout  = 8'b00000001; //  360 :   1 - 0x1 -- plane 1
      12'h169: dout  = 8'b00000011; //  361 :   3 - 0x3
      12'h16A: dout  = 8'b00000001; //  362 :   1 - 0x1
      12'h16B: dout  = 8'b00000100; //  363 :   4 - 0x4
      12'h16C: dout  = 8'b00000111; //  364 :   7 - 0x7
      12'h16D: dout  = 8'b00001111; //  365 :  15 - 0xf
      12'h16E: dout  = 8'b00001111; //  366 :  15 - 0xf
      12'h16F: dout  = 8'b00000011; //  367 :   3 - 0x3
      12'h170: dout  = 8'b11111000; //  368 : 248 - 0xf8 -- Sprite 0x17
      12'h171: dout  = 8'b11110000; //  369 : 240 - 0xf0
      12'h172: dout  = 8'b11100000; //  370 : 224 - 0xe0
      12'h173: dout  = 8'b11110000; //  371 : 240 - 0xf0
      12'h174: dout  = 8'b10110000; //  372 : 176 - 0xb0
      12'h175: dout  = 8'b10000000; //  373 : 128 - 0x80
      12'h176: dout  = 8'b11100000; //  374 : 224 - 0xe0
      12'h177: dout  = 8'b11100000; //  375 : 224 - 0xe0
      12'h178: dout  = 8'b11111000; //  376 : 248 - 0xf8 -- plane 1
      12'h179: dout  = 8'b11110000; //  377 : 240 - 0xf0
      12'h17A: dout  = 8'b11100000; //  378 : 224 - 0xe0
      12'h17B: dout  = 8'b01110000; //  379 : 112 - 0x70
      12'h17C: dout  = 8'b10110000; //  380 : 176 - 0xb0
      12'h17D: dout  = 8'b10000000; //  381 : 128 - 0x80
      12'h17E: dout  = 8'b11100000; //  382 : 224 - 0xe0
      12'h17F: dout  = 8'b11100000; //  383 : 224 - 0xe0
      12'h180: dout  = 8'b00000011; //  384 :   3 - 0x3 -- Sprite 0x18
      12'h181: dout  = 8'b00111111; //  385 :  63 - 0x3f
      12'h182: dout  = 8'b01111111; //  386 : 127 - 0x7f
      12'h183: dout  = 8'b00011001; //  387 :  25 - 0x19
      12'h184: dout  = 8'b00001001; //  388 :   9 - 0x9
      12'h185: dout  = 8'b00001001; //  389 :   9 - 0x9
      12'h186: dout  = 8'b00101000; //  390 :  40 - 0x28
      12'h187: dout  = 8'b01011100; //  391 :  92 - 0x5c
      12'h188: dout  = 8'b00000000; //  392 :   0 - 0x0 -- plane 1
      12'h189: dout  = 8'b00110000; //  393 :  48 - 0x30
      12'h18A: dout  = 8'b01110000; //  394 : 112 - 0x70
      12'h18B: dout  = 8'b01111111; //  395 : 127 - 0x7f
      12'h18C: dout  = 8'b11111111; //  396 : 255 - 0xff
      12'h18D: dout  = 8'b11111111; //  397 : 255 - 0xff
      12'h18E: dout  = 8'b11110111; //  398 : 247 - 0xf7
      12'h18F: dout  = 8'b11110011; //  399 : 243 - 0xf3
      12'h190: dout  = 8'b11111000; //  400 : 248 - 0xf8 -- Sprite 0x19
      12'h191: dout  = 8'b11100000; //  401 : 224 - 0xe0
      12'h192: dout  = 8'b11100000; //  402 : 224 - 0xe0
      12'h193: dout  = 8'b11111100; //  403 : 252 - 0xfc
      12'h194: dout  = 8'b00100110; //  404 :  38 - 0x26
      12'h195: dout  = 8'b00110000; //  405 :  48 - 0x30
      12'h196: dout  = 8'b10000000; //  406 : 128 - 0x80
      12'h197: dout  = 8'b00010000; //  407 :  16 - 0x10
      12'h198: dout  = 8'b00000000; //  408 :   0 - 0x0 -- plane 1
      12'h199: dout  = 8'b00011000; //  409 :  24 - 0x18
      12'h19A: dout  = 8'b00010000; //  410 :  16 - 0x10
      12'h19B: dout  = 8'b00000000; //  411 :   0 - 0x0
      12'h19C: dout  = 8'b11111000; //  412 : 248 - 0xf8
      12'h19D: dout  = 8'b11111000; //  413 : 248 - 0xf8
      12'h19E: dout  = 8'b11111110; //  414 : 254 - 0xfe
      12'h19F: dout  = 8'b11111111; //  415 : 255 - 0xff
      12'h1A0: dout  = 8'b00111110; //  416 :  62 - 0x3e -- Sprite 0x1a
      12'h1A1: dout  = 8'b00011110; //  417 :  30 - 0x1e
      12'h1A2: dout  = 8'b00111111; //  418 :  63 - 0x3f
      12'h1A3: dout  = 8'b00111000; //  419 :  56 - 0x38
      12'h1A4: dout  = 8'b00110000; //  420 :  48 - 0x30
      12'h1A5: dout  = 8'b00110000; //  421 :  48 - 0x30
      12'h1A6: dout  = 8'b00000000; //  422 :   0 - 0x0
      12'h1A7: dout  = 8'b00111010; //  423 :  58 - 0x3a
      12'h1A8: dout  = 8'b11100111; //  424 : 231 - 0xe7 -- plane 1
      12'h1A9: dout  = 8'b00001111; //  425 :  15 - 0xf
      12'h1AA: dout  = 8'b00001111; //  426 :  15 - 0xf
      12'h1AB: dout  = 8'b00011111; //  427 :  31 - 0x1f
      12'h1AC: dout  = 8'b00011111; //  428 :  31 - 0x1f
      12'h1AD: dout  = 8'b00011111; //  429 :  31 - 0x1f
      12'h1AE: dout  = 8'b00001111; //  430 :  15 - 0xf
      12'h1AF: dout  = 8'b00000111; //  431 :   7 - 0x7
      12'h1B0: dout  = 8'b01111000; //  432 : 120 - 0x78 -- Sprite 0x1b
      12'h1B1: dout  = 8'b00011110; //  433 :  30 - 0x1e
      12'h1B2: dout  = 8'b10000000; //  434 : 128 - 0x80
      12'h1B3: dout  = 8'b11111110; //  435 : 254 - 0xfe
      12'h1B4: dout  = 8'b01111110; //  436 : 126 - 0x7e
      12'h1B5: dout  = 8'b01111110; //  437 : 126 - 0x7e
      12'h1B6: dout  = 8'b01111111; //  438 : 127 - 0x7f
      12'h1B7: dout  = 8'b01111111; //  439 : 127 - 0x7f
      12'h1B8: dout  = 8'b11111111; //  440 : 255 - 0xff -- plane 1
      12'h1B9: dout  = 8'b11111110; //  441 : 254 - 0xfe
      12'h1BA: dout  = 8'b11111100; //  442 : 252 - 0xfc
      12'h1BB: dout  = 8'b11000110; //  443 : 198 - 0xc6
      12'h1BC: dout  = 8'b10001110; //  444 : 142 - 0x8e
      12'h1BD: dout  = 8'b11101110; //  445 : 238 - 0xee
      12'h1BE: dout  = 8'b11111111; //  446 : 255 - 0xff
      12'h1BF: dout  = 8'b11111111; //  447 : 255 - 0xff
      12'h1C0: dout  = 8'b00111100; //  448 :  60 - 0x3c -- Sprite 0x1c
      12'h1C1: dout  = 8'b00111111; //  449 :  63 - 0x3f
      12'h1C2: dout  = 8'b00011111; //  450 :  31 - 0x1f
      12'h1C3: dout  = 8'b00001111; //  451 :  15 - 0xf
      12'h1C4: dout  = 8'b00000111; //  452 :   7 - 0x7
      12'h1C5: dout  = 8'b00111111; //  453 :  63 - 0x3f
      12'h1C6: dout  = 8'b00100001; //  454 :  33 - 0x21
      12'h1C7: dout  = 8'b00100000; //  455 :  32 - 0x20
      12'h1C8: dout  = 8'b00000011; //  456 :   3 - 0x3 -- plane 1
      12'h1C9: dout  = 8'b00000000; //  457 :   0 - 0x0
      12'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout  = 8'b00001110; //  459 :  14 - 0xe
      12'h1CC: dout  = 8'b00000111; //  460 :   7 - 0x7
      12'h1CD: dout  = 8'b00111111; //  461 :  63 - 0x3f
      12'h1CE: dout  = 8'b00111111; //  462 :  63 - 0x3f
      12'h1CF: dout  = 8'b00111111; //  463 :  63 - 0x3f
      12'h1D0: dout  = 8'b11111111; //  464 : 255 - 0xff -- Sprite 0x1d
      12'h1D1: dout  = 8'b11111111; //  465 : 255 - 0xff
      12'h1D2: dout  = 8'b11111111; //  466 : 255 - 0xff
      12'h1D3: dout  = 8'b11111110; //  467 : 254 - 0xfe
      12'h1D4: dout  = 8'b11111110; //  468 : 254 - 0xfe
      12'h1D5: dout  = 8'b11111110; //  469 : 254 - 0xfe
      12'h1D6: dout  = 8'b11111100; //  470 : 252 - 0xfc
      12'h1D7: dout  = 8'b01110000; //  471 : 112 - 0x70
      12'h1D8: dout  = 8'b11111111; //  472 : 255 - 0xff -- plane 1
      12'h1D9: dout  = 8'b01111111; //  473 : 127 - 0x7f
      12'h1DA: dout  = 8'b00111111; //  474 :  63 - 0x3f
      12'h1DB: dout  = 8'b00001110; //  475 :  14 - 0xe
      12'h1DC: dout  = 8'b11000000; //  476 : 192 - 0xc0
      12'h1DD: dout  = 8'b11000000; //  477 : 192 - 0xc0
      12'h1DE: dout  = 8'b11100000; //  478 : 224 - 0xe0
      12'h1DF: dout  = 8'b11100000; //  479 : 224 - 0xe0
      12'h1E0: dout  = 8'b00001111; //  480 :  15 - 0xf -- Sprite 0x1e
      12'h1E1: dout  = 8'b10011111; //  481 : 159 - 0x9f
      12'h1E2: dout  = 8'b11001111; //  482 : 207 - 0xcf
      12'h1E3: dout  = 8'b11111111; //  483 : 255 - 0xff
      12'h1E4: dout  = 8'b01111111; //  484 : 127 - 0x7f
      12'h1E5: dout  = 8'b00111111; //  485 :  63 - 0x3f
      12'h1E6: dout  = 8'b00011110; //  486 :  30 - 0x1e
      12'h1E7: dout  = 8'b00001110; //  487 :  14 - 0xe
      12'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0 -- plane 1
      12'h1E9: dout  = 8'b10000000; //  489 : 128 - 0x80
      12'h1EA: dout  = 8'b11001000; //  490 : 200 - 0xc8
      12'h1EB: dout  = 8'b11111110; //  491 : 254 - 0xfe
      12'h1EC: dout  = 8'b01111111; //  492 : 127 - 0x7f
      12'h1ED: dout  = 8'b00111111; //  493 :  63 - 0x3f
      12'h1EE: dout  = 8'b00011110; //  494 :  30 - 0x1e
      12'h1EF: dout  = 8'b00001110; //  495 :  14 - 0xe
      12'h1F0: dout  = 8'b00100000; //  496 :  32 - 0x20 -- Sprite 0x1f
      12'h1F1: dout  = 8'b11000000; //  497 : 192 - 0xc0
      12'h1F2: dout  = 8'b10000000; //  498 : 128 - 0x80
      12'h1F3: dout  = 8'b10000000; //  499 : 128 - 0x80
      12'h1F4: dout  = 8'b00000000; //  500 :   0 - 0x0
      12'h1F5: dout  = 8'b00000000; //  501 :   0 - 0x0
      12'h1F6: dout  = 8'b00000000; //  502 :   0 - 0x0
      12'h1F7: dout  = 8'b00000000; //  503 :   0 - 0x0
      12'h1F8: dout  = 8'b11100000; //  504 : 224 - 0xe0 -- plane 1
      12'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout  = 8'b00000000; //  507 :   0 - 0x0
      12'h1FC: dout  = 8'b00000000; //  508 :   0 - 0x0
      12'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      12'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout  = 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x20
      12'h201: dout  = 8'b00000000; //  513 :   0 - 0x0
      12'h202: dout  = 8'b00000011; //  514 :   3 - 0x3
      12'h203: dout  = 8'b00001111; //  515 :  15 - 0xf
      12'h204: dout  = 8'b00011111; //  516 :  31 - 0x1f
      12'h205: dout  = 8'b00011111; //  517 :  31 - 0x1f
      12'h206: dout  = 8'b00011100; //  518 :  28 - 0x1c
      12'h207: dout  = 8'b00100100; //  519 :  36 - 0x24
      12'h208: dout  = 8'b00000000; //  520 :   0 - 0x0 -- plane 1
      12'h209: dout  = 8'b00000000; //  521 :   0 - 0x0
      12'h20A: dout  = 8'b00000000; //  522 :   0 - 0x0
      12'h20B: dout  = 8'b00000000; //  523 :   0 - 0x0
      12'h20C: dout  = 8'b00000000; //  524 :   0 - 0x0
      12'h20D: dout  = 8'b00000000; //  525 :   0 - 0x0
      12'h20E: dout  = 8'b00011111; //  526 :  31 - 0x1f
      12'h20F: dout  = 8'b00111111; //  527 :  63 - 0x3f
      12'h210: dout  = 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x21
      12'h211: dout  = 8'b00000100; //  529 :   4 - 0x4
      12'h212: dout  = 8'b11100110; //  530 : 230 - 0xe6
      12'h213: dout  = 8'b11100000; //  531 : 224 - 0xe0
      12'h214: dout  = 8'b11111111; //  532 : 255 - 0xff
      12'h215: dout  = 8'b11111111; //  533 : 255 - 0xff
      12'h216: dout  = 8'b10001111; //  534 : 143 - 0x8f
      12'h217: dout  = 8'b10000011; //  535 : 131 - 0x83
      12'h218: dout  = 8'b00001110; //  536 :  14 - 0xe -- plane 1
      12'h219: dout  = 8'b00011111; //  537 :  31 - 0x1f
      12'h21A: dout  = 8'b00011111; //  538 :  31 - 0x1f
      12'h21B: dout  = 8'b00011111; //  539 :  31 - 0x1f
      12'h21C: dout  = 8'b00011111; //  540 :  31 - 0x1f
      12'h21D: dout  = 8'b00000011; //  541 :   3 - 0x3
      12'h21E: dout  = 8'b11111111; //  542 : 255 - 0xff
      12'h21F: dout  = 8'b11111111; //  543 : 255 - 0xff
      12'h220: dout  = 8'b00100110; //  544 :  38 - 0x26 -- Sprite 0x22
      12'h221: dout  = 8'b00100110; //  545 :  38 - 0x26
      12'h222: dout  = 8'b01100000; //  546 :  96 - 0x60
      12'h223: dout  = 8'b01111000; //  547 : 120 - 0x78
      12'h224: dout  = 8'b00011000; //  548 :  24 - 0x18
      12'h225: dout  = 8'b00001111; //  549 :  15 - 0xf
      12'h226: dout  = 8'b01111111; //  550 : 127 - 0x7f
      12'h227: dout  = 8'b11111111; //  551 : 255 - 0xff
      12'h228: dout  = 8'b00111111; //  552 :  63 - 0x3f -- plane 1
      12'h229: dout  = 8'b00111111; //  553 :  63 - 0x3f
      12'h22A: dout  = 8'b01111111; //  554 : 127 - 0x7f
      12'h22B: dout  = 8'b01111111; //  555 : 127 - 0x7f
      12'h22C: dout  = 8'b00011111; //  556 :  31 - 0x1f
      12'h22D: dout  = 8'b00000000; //  557 :   0 - 0x0
      12'h22E: dout  = 8'b01111110; //  558 : 126 - 0x7e
      12'h22F: dout  = 8'b11111111; //  559 : 255 - 0xff
      12'h230: dout  = 8'b00000001; //  560 :   1 - 0x1 -- Sprite 0x23
      12'h231: dout  = 8'b00100001; //  561 :  33 - 0x21
      12'h232: dout  = 8'b11111110; //  562 : 254 - 0xfe
      12'h233: dout  = 8'b01111010; //  563 : 122 - 0x7a
      12'h234: dout  = 8'b00000110; //  564 :   6 - 0x6
      12'h235: dout  = 8'b11111110; //  565 : 254 - 0xfe
      12'h236: dout  = 8'b11111100; //  566 : 252 - 0xfc
      12'h237: dout  = 8'b11111100; //  567 : 252 - 0xfc
      12'h238: dout  = 8'b11111111; //  568 : 255 - 0xff -- plane 1
      12'h239: dout  = 8'b11111111; //  569 : 255 - 0xff
      12'h23A: dout  = 8'b11111110; //  570 : 254 - 0xfe
      12'h23B: dout  = 8'b11111110; //  571 : 254 - 0xfe
      12'h23C: dout  = 8'b11111110; //  572 : 254 - 0xfe
      12'h23D: dout  = 8'b11011110; //  573 : 222 - 0xde
      12'h23E: dout  = 8'b01011100; //  574 :  92 - 0x5c
      12'h23F: dout  = 8'b01101100; //  575 : 108 - 0x6c
      12'h240: dout  = 8'b11111111; //  576 : 255 - 0xff -- Sprite 0x24
      12'h241: dout  = 8'b11001111; //  577 : 207 - 0xcf
      12'h242: dout  = 8'b10000111; //  578 : 135 - 0x87
      12'h243: dout  = 8'b00000111; //  579 :   7 - 0x7
      12'h244: dout  = 8'b00000111; //  580 :   7 - 0x7
      12'h245: dout  = 8'b00001111; //  581 :  15 - 0xf
      12'h246: dout  = 8'b00011111; //  582 :  31 - 0x1f
      12'h247: dout  = 8'b00011111; //  583 :  31 - 0x1f
      12'h248: dout  = 8'b11111111; //  584 : 255 - 0xff -- plane 1
      12'h249: dout  = 8'b11111111; //  585 : 255 - 0xff
      12'h24A: dout  = 8'b11111110; //  586 : 254 - 0xfe
      12'h24B: dout  = 8'b11111100; //  587 : 252 - 0xfc
      12'h24C: dout  = 8'b11111000; //  588 : 248 - 0xf8
      12'h24D: dout  = 8'b10110000; //  589 : 176 - 0xb0
      12'h24E: dout  = 8'b01100000; //  590 :  96 - 0x60
      12'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout  = 8'b11111000; //  592 : 248 - 0xf8 -- Sprite 0x25
      12'h251: dout  = 8'b11111000; //  593 : 248 - 0xf8
      12'h252: dout  = 8'b11110000; //  594 : 240 - 0xf0
      12'h253: dout  = 8'b10111000; //  595 : 184 - 0xb8
      12'h254: dout  = 8'b11111000; //  596 : 248 - 0xf8
      12'h255: dout  = 8'b11111001; //  597 : 249 - 0xf9
      12'h256: dout  = 8'b11111011; //  598 : 251 - 0xfb
      12'h257: dout  = 8'b11111111; //  599 : 255 - 0xff
      12'h258: dout  = 8'b00101000; //  600 :  40 - 0x28 -- plane 1
      12'h259: dout  = 8'b00110000; //  601 :  48 - 0x30
      12'h25A: dout  = 8'b00011000; //  602 :  24 - 0x18
      12'h25B: dout  = 8'b01000000; //  603 :  64 - 0x40
      12'h25C: dout  = 8'b00000000; //  604 :   0 - 0x0
      12'h25D: dout  = 8'b00000001; //  605 :   1 - 0x1
      12'h25E: dout  = 8'b00000011; //  606 :   3 - 0x3
      12'h25F: dout  = 8'b00001111; //  607 :  15 - 0xf
      12'h260: dout  = 8'b00011111; //  608 :  31 - 0x1f -- Sprite 0x26
      12'h261: dout  = 8'b11111111; //  609 : 255 - 0xff
      12'h262: dout  = 8'b11111111; //  610 : 255 - 0xff
      12'h263: dout  = 8'b11111111; //  611 : 255 - 0xff
      12'h264: dout  = 8'b11111111; //  612 : 255 - 0xff
      12'h265: dout  = 8'b11111110; //  613 : 254 - 0xfe
      12'h266: dout  = 8'b11000000; //  614 : 192 - 0xc0
      12'h267: dout  = 8'b10000000; //  615 : 128 - 0x80
      12'h268: dout  = 8'b00010000; //  616 :  16 - 0x10 -- plane 1
      12'h269: dout  = 8'b11101100; //  617 : 236 - 0xec
      12'h26A: dout  = 8'b11100011; //  618 : 227 - 0xe3
      12'h26B: dout  = 8'b11100000; //  619 : 224 - 0xe0
      12'h26C: dout  = 8'b11100000; //  620 : 224 - 0xe0
      12'h26D: dout  = 8'b11100000; //  621 : 224 - 0xe0
      12'h26E: dout  = 8'b11000000; //  622 : 192 - 0xc0
      12'h26F: dout  = 8'b10000000; //  623 : 128 - 0x80
      12'h270: dout  = 8'b11111111; //  624 : 255 - 0xff -- Sprite 0x27
      12'h271: dout  = 8'b11111111; //  625 : 255 - 0xff
      12'h272: dout  = 8'b11111111; //  626 : 255 - 0xff
      12'h273: dout  = 8'b00111111; //  627 :  63 - 0x3f
      12'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      12'h275: dout  = 8'b00000000; //  629 :   0 - 0x0
      12'h276: dout  = 8'b00000000; //  630 :   0 - 0x0
      12'h277: dout  = 8'b00000000; //  631 :   0 - 0x0
      12'h278: dout  = 8'b00001111; //  632 :  15 - 0xf -- plane 1
      12'h279: dout  = 8'b00001111; //  633 :  15 - 0xf
      12'h27A: dout  = 8'b00001111; //  634 :  15 - 0xf
      12'h27B: dout  = 8'b00001111; //  635 :  15 - 0xf
      12'h27C: dout  = 8'b00000000; //  636 :   0 - 0x0
      12'h27D: dout  = 8'b00000000; //  637 :   0 - 0x0
      12'h27E: dout  = 8'b00000000; //  638 :   0 - 0x0
      12'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout  = 8'b00010011; //  640 :  19 - 0x13 -- Sprite 0x28
      12'h281: dout  = 8'b00110011; //  641 :  51 - 0x33
      12'h282: dout  = 8'b00110000; //  642 :  48 - 0x30
      12'h283: dout  = 8'b00011000; //  643 :  24 - 0x18
      12'h284: dout  = 8'b00000100; //  644 :   4 - 0x4
      12'h285: dout  = 8'b00001111; //  645 :  15 - 0xf
      12'h286: dout  = 8'b00011111; //  646 :  31 - 0x1f
      12'h287: dout  = 8'b00011111; //  647 :  31 - 0x1f
      12'h288: dout  = 8'b00011111; //  648 :  31 - 0x1f -- plane 1
      12'h289: dout  = 8'b00111111; //  649 :  63 - 0x3f
      12'h28A: dout  = 8'b00111111; //  650 :  63 - 0x3f
      12'h28B: dout  = 8'b00011111; //  651 :  31 - 0x1f
      12'h28C: dout  = 8'b00000111; //  652 :   7 - 0x7
      12'h28D: dout  = 8'b00001001; //  653 :   9 - 0x9
      12'h28E: dout  = 8'b00010011; //  654 :  19 - 0x13
      12'h28F: dout  = 8'b00010111; //  655 :  23 - 0x17
      12'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x29
      12'h291: dout  = 8'b00010000; //  657 :  16 - 0x10
      12'h292: dout  = 8'b01111110; //  658 : 126 - 0x7e
      12'h293: dout  = 8'b00110000; //  659 :  48 - 0x30
      12'h294: dout  = 8'b11100000; //  660 : 224 - 0xe0
      12'h295: dout  = 8'b11110000; //  661 : 240 - 0xf0
      12'h296: dout  = 8'b11110000; //  662 : 240 - 0xf0
      12'h297: dout  = 8'b11100000; //  663 : 224 - 0xe0
      12'h298: dout  = 8'b11111111; //  664 : 255 - 0xff -- plane 1
      12'h299: dout  = 8'b11111111; //  665 : 255 - 0xff
      12'h29A: dout  = 8'b11111110; //  666 : 254 - 0xfe
      12'h29B: dout  = 8'b11111111; //  667 : 255 - 0xff
      12'h29C: dout  = 8'b11111110; //  668 : 254 - 0xfe
      12'h29D: dout  = 8'b11111100; //  669 : 252 - 0xfc
      12'h29E: dout  = 8'b11111000; //  670 : 248 - 0xf8
      12'h29F: dout  = 8'b11100000; //  671 : 224 - 0xe0
      12'h2A0: dout  = 8'b00011111; //  672 :  31 - 0x1f -- Sprite 0x2a
      12'h2A1: dout  = 8'b00011111; //  673 :  31 - 0x1f
      12'h2A2: dout  = 8'b00001111; //  674 :  15 - 0xf
      12'h2A3: dout  = 8'b00001111; //  675 :  15 - 0xf
      12'h2A4: dout  = 8'b00001111; //  676 :  15 - 0xf
      12'h2A5: dout  = 8'b00011111; //  677 :  31 - 0x1f
      12'h2A6: dout  = 8'b00011111; //  678 :  31 - 0x1f
      12'h2A7: dout  = 8'b00011111; //  679 :  31 - 0x1f
      12'h2A8: dout  = 8'b00010111; //  680 :  23 - 0x17 -- plane 1
      12'h2A9: dout  = 8'b00010111; //  681 :  23 - 0x17
      12'h2AA: dout  = 8'b00000011; //  682 :   3 - 0x3
      12'h2AB: dout  = 8'b00000000; //  683 :   0 - 0x0
      12'h2AC: dout  = 8'b00000000; //  684 :   0 - 0x0
      12'h2AD: dout  = 8'b00000000; //  685 :   0 - 0x0
      12'h2AE: dout  = 8'b00000000; //  686 :   0 - 0x0
      12'h2AF: dout  = 8'b00000000; //  687 :   0 - 0x0
      12'h2B0: dout  = 8'b11110000; //  688 : 240 - 0xf0 -- Sprite 0x2b
      12'h2B1: dout  = 8'b11110000; //  689 : 240 - 0xf0
      12'h2B2: dout  = 8'b11111000; //  690 : 248 - 0xf8
      12'h2B3: dout  = 8'b11111000; //  691 : 248 - 0xf8
      12'h2B4: dout  = 8'b10111000; //  692 : 184 - 0xb8
      12'h2B5: dout  = 8'b11111000; //  693 : 248 - 0xf8
      12'h2B6: dout  = 8'b11111000; //  694 : 248 - 0xf8
      12'h2B7: dout  = 8'b11111000; //  695 : 248 - 0xf8
      12'h2B8: dout  = 8'b11010000; //  696 : 208 - 0xd0 -- plane 1
      12'h2B9: dout  = 8'b10010000; //  697 : 144 - 0x90
      12'h2BA: dout  = 8'b00011000; //  698 :  24 - 0x18
      12'h2BB: dout  = 8'b00001000; //  699 :   8 - 0x8
      12'h2BC: dout  = 8'b01000000; //  700 :  64 - 0x40
      12'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout  = 8'b00111111; //  704 :  63 - 0x3f -- Sprite 0x2c
      12'h2C1: dout  = 8'b11111111; //  705 : 255 - 0xff
      12'h2C2: dout  = 8'b11111111; //  706 : 255 - 0xff
      12'h2C3: dout  = 8'b11111111; //  707 : 255 - 0xff
      12'h2C4: dout  = 8'b11110110; //  708 : 246 - 0xf6
      12'h2C5: dout  = 8'b11000110; //  709 : 198 - 0xc6
      12'h2C6: dout  = 8'b10000100; //  710 : 132 - 0x84
      12'h2C7: dout  = 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout  = 8'b00110000; //  712 :  48 - 0x30 -- plane 1
      12'h2C9: dout  = 8'b11110000; //  713 : 240 - 0xf0
      12'h2CA: dout  = 8'b11110000; //  714 : 240 - 0xf0
      12'h2CB: dout  = 8'b11110001; //  715 : 241 - 0xf1
      12'h2CC: dout  = 8'b11110110; //  716 : 246 - 0xf6
      12'h2CD: dout  = 8'b11000110; //  717 : 198 - 0xc6
      12'h2CE: dout  = 8'b10000100; //  718 : 132 - 0x84
      12'h2CF: dout  = 8'b00000000; //  719 :   0 - 0x0
      12'h2D0: dout  = 8'b11110000; //  720 : 240 - 0xf0 -- Sprite 0x2d
      12'h2D1: dout  = 8'b11100000; //  721 : 224 - 0xe0
      12'h2D2: dout  = 8'b10000000; //  722 : 128 - 0x80
      12'h2D3: dout  = 8'b00000000; //  723 :   0 - 0x0
      12'h2D4: dout  = 8'b00000000; //  724 :   0 - 0x0
      12'h2D5: dout  = 8'b00000000; //  725 :   0 - 0x0
      12'h2D6: dout  = 8'b00000000; //  726 :   0 - 0x0
      12'h2D7: dout  = 8'b00000000; //  727 :   0 - 0x0
      12'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- plane 1
      12'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      12'h2DA: dout  = 8'b00000000; //  730 :   0 - 0x0
      12'h2DB: dout  = 8'b00000000; //  731 :   0 - 0x0
      12'h2DC: dout  = 8'b00000000; //  732 :   0 - 0x0
      12'h2DD: dout  = 8'b00000000; //  733 :   0 - 0x0
      12'h2DE: dout  = 8'b00000000; //  734 :   0 - 0x0
      12'h2DF: dout  = 8'b00000000; //  735 :   0 - 0x0
      12'h2E0: dout  = 8'b00011111; //  736 :  31 - 0x1f -- Sprite 0x2e
      12'h2E1: dout  = 8'b00011111; //  737 :  31 - 0x1f
      12'h2E2: dout  = 8'b00111111; //  738 :  63 - 0x3f
      12'h2E3: dout  = 8'b00111111; //  739 :  63 - 0x3f
      12'h2E4: dout  = 8'b00011111; //  740 :  31 - 0x1f
      12'h2E5: dout  = 8'b00001111; //  741 :  15 - 0xf
      12'h2E6: dout  = 8'b00001111; //  742 :  15 - 0xf
      12'h2E7: dout  = 8'b00011111; //  743 :  31 - 0x1f
      12'h2E8: dout  = 8'b00011111; //  744 :  31 - 0x1f -- plane 1
      12'h2E9: dout  = 8'b00011111; //  745 :  31 - 0x1f
      12'h2EA: dout  = 8'b00111111; //  746 :  63 - 0x3f
      12'h2EB: dout  = 8'b00111110; //  747 :  62 - 0x3e
      12'h2EC: dout  = 8'b01111100; //  748 : 124 - 0x7c
      12'h2ED: dout  = 8'b01111000; //  749 : 120 - 0x78
      12'h2EE: dout  = 8'b11110000; //  750 : 240 - 0xf0
      12'h2EF: dout  = 8'b11100000; //  751 : 224 - 0xe0
      12'h2F0: dout  = 8'b11110000; //  752 : 240 - 0xf0 -- Sprite 0x2f
      12'h2F1: dout  = 8'b11110000; //  753 : 240 - 0xf0
      12'h2F2: dout  = 8'b11111000; //  754 : 248 - 0xf8
      12'h2F3: dout  = 8'b11111000; //  755 : 248 - 0xf8
      12'h2F4: dout  = 8'b10111000; //  756 : 184 - 0xb8
      12'h2F5: dout  = 8'b11111000; //  757 : 248 - 0xf8
      12'h2F6: dout  = 8'b11111000; //  758 : 248 - 0xf8
      12'h2F7: dout  = 8'b11110000; //  759 : 240 - 0xf0
      12'h2F8: dout  = 8'b10110000; //  760 : 176 - 0xb0 -- plane 1
      12'h2F9: dout  = 8'b10010000; //  761 : 144 - 0x90
      12'h2FA: dout  = 8'b00011000; //  762 :  24 - 0x18
      12'h2FB: dout  = 8'b00001000; //  763 :   8 - 0x8
      12'h2FC: dout  = 8'b01000000; //  764 :  64 - 0x40
      12'h2FD: dout  = 8'b00000000; //  765 :   0 - 0x0
      12'h2FE: dout  = 8'b00000000; //  766 :   0 - 0x0
      12'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout  = 8'b11100000; //  768 : 224 - 0xe0 -- Sprite 0x30
      12'h301: dout  = 8'b11110000; //  769 : 240 - 0xf0
      12'h302: dout  = 8'b11110000; //  770 : 240 - 0xf0
      12'h303: dout  = 8'b11110000; //  771 : 240 - 0xf0
      12'h304: dout  = 8'b11110000; //  772 : 240 - 0xf0
      12'h305: dout  = 8'b11110000; //  773 : 240 - 0xf0
      12'h306: dout  = 8'b11111000; //  774 : 248 - 0xf8
      12'h307: dout  = 8'b11110000; //  775 : 240 - 0xf0
      12'h308: dout  = 8'b11000000; //  776 : 192 - 0xc0 -- plane 1
      12'h309: dout  = 8'b11100000; //  777 : 224 - 0xe0
      12'h30A: dout  = 8'b11111100; //  778 : 252 - 0xfc
      12'h30B: dout  = 8'b11111110; //  779 : 254 - 0xfe
      12'h30C: dout  = 8'b11111111; //  780 : 255 - 0xff
      12'h30D: dout  = 8'b01111111; //  781 : 127 - 0x7f
      12'h30E: dout  = 8'b00000011; //  782 :   3 - 0x3
      12'h30F: dout  = 8'b00000000; //  783 :   0 - 0x0
      12'h310: dout  = 8'b00011111; //  784 :  31 - 0x1f -- Sprite 0x31
      12'h311: dout  = 8'b00011111; //  785 :  31 - 0x1f
      12'h312: dout  = 8'b00011111; //  786 :  31 - 0x1f
      12'h313: dout  = 8'b00111111; //  787 :  63 - 0x3f
      12'h314: dout  = 8'b00111110; //  788 :  62 - 0x3e
      12'h315: dout  = 8'b00111100; //  789 :  60 - 0x3c
      12'h316: dout  = 8'b00111000; //  790 :  56 - 0x38
      12'h317: dout  = 8'b00011000; //  791 :  24 - 0x18
      12'h318: dout  = 8'b00000000; //  792 :   0 - 0x0 -- plane 1
      12'h319: dout  = 8'b00000000; //  793 :   0 - 0x0
      12'h31A: dout  = 8'b00010000; //  794 :  16 - 0x10
      12'h31B: dout  = 8'b00111000; //  795 :  56 - 0x38
      12'h31C: dout  = 8'b00111110; //  796 :  62 - 0x3e
      12'h31D: dout  = 8'b00111100; //  797 :  60 - 0x3c
      12'h31E: dout  = 8'b00111000; //  798 :  56 - 0x38
      12'h31F: dout  = 8'b00011000; //  799 :  24 - 0x18
      12'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x32
      12'h321: dout  = 8'b00000011; //  801 :   3 - 0x3
      12'h322: dout  = 8'b00000111; //  802 :   7 - 0x7
      12'h323: dout  = 8'b00000111; //  803 :   7 - 0x7
      12'h324: dout  = 8'b00001010; //  804 :  10 - 0xa
      12'h325: dout  = 8'b00001011; //  805 :  11 - 0xb
      12'h326: dout  = 8'b00001100; //  806 :  12 - 0xc
      12'h327: dout  = 8'b00000000; //  807 :   0 - 0x0
      12'h328: dout  = 8'b00000000; //  808 :   0 - 0x0 -- plane 1
      12'h329: dout  = 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout  = 8'b00000000; //  810 :   0 - 0x0
      12'h32B: dout  = 8'b00000111; //  811 :   7 - 0x7
      12'h32C: dout  = 8'b00001111; //  812 :  15 - 0xf
      12'h32D: dout  = 8'b00001111; //  813 :  15 - 0xf
      12'h32E: dout  = 8'b00001111; //  814 :  15 - 0xf
      12'h32F: dout  = 8'b00000011; //  815 :   3 - 0x3
      12'h330: dout  = 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x33
      12'h331: dout  = 8'b11100000; //  817 : 224 - 0xe0
      12'h332: dout  = 8'b11111100; //  818 : 252 - 0xfc
      12'h333: dout  = 8'b00100000; //  819 :  32 - 0x20
      12'h334: dout  = 8'b00100000; //  820 :  32 - 0x20
      12'h335: dout  = 8'b00010000; //  821 :  16 - 0x10
      12'h336: dout  = 8'b00111100; //  822 :  60 - 0x3c
      12'h337: dout  = 8'b00000000; //  823 :   0 - 0x0
      12'h338: dout  = 8'b00000000; //  824 :   0 - 0x0 -- plane 1
      12'h339: dout  = 8'b00000000; //  825 :   0 - 0x0
      12'h33A: dout  = 8'b00000000; //  826 :   0 - 0x0
      12'h33B: dout  = 8'b11110000; //  827 : 240 - 0xf0
      12'h33C: dout  = 8'b11111100; //  828 : 252 - 0xfc
      12'h33D: dout  = 8'b11111110; //  829 : 254 - 0xfe
      12'h33E: dout  = 8'b11111100; //  830 : 252 - 0xfc
      12'h33F: dout  = 8'b11111000; //  831 : 248 - 0xf8
      12'h340: dout  = 8'b00000111; //  832 :   7 - 0x7 -- Sprite 0x34
      12'h341: dout  = 8'b00000111; //  833 :   7 - 0x7
      12'h342: dout  = 8'b00000111; //  834 :   7 - 0x7
      12'h343: dout  = 8'b00011111; //  835 :  31 - 0x1f
      12'h344: dout  = 8'b00011111; //  836 :  31 - 0x1f
      12'h345: dout  = 8'b00111110; //  837 :  62 - 0x3e
      12'h346: dout  = 8'b00100001; //  838 :  33 - 0x21
      12'h347: dout  = 8'b00000001; //  839 :   1 - 0x1
      12'h348: dout  = 8'b00000111; //  840 :   7 - 0x7 -- plane 1
      12'h349: dout  = 8'b00001111; //  841 :  15 - 0xf
      12'h34A: dout  = 8'b00011011; //  842 :  27 - 0x1b
      12'h34B: dout  = 8'b00011000; //  843 :  24 - 0x18
      12'h34C: dout  = 8'b00010000; //  844 :  16 - 0x10
      12'h34D: dout  = 8'b00110000; //  845 :  48 - 0x30
      12'h34E: dout  = 8'b00100001; //  846 :  33 - 0x21
      12'h34F: dout  = 8'b00000001; //  847 :   1 - 0x1
      12'h350: dout  = 8'b11100000; //  848 : 224 - 0xe0 -- Sprite 0x35
      12'h351: dout  = 8'b11100000; //  849 : 224 - 0xe0
      12'h352: dout  = 8'b11100000; //  850 : 224 - 0xe0
      12'h353: dout  = 8'b11110000; //  851 : 240 - 0xf0
      12'h354: dout  = 8'b11110000; //  852 : 240 - 0xf0
      12'h355: dout  = 8'b11100000; //  853 : 224 - 0xe0
      12'h356: dout  = 8'b11000000; //  854 : 192 - 0xc0
      12'h357: dout  = 8'b11100000; //  855 : 224 - 0xe0
      12'h358: dout  = 8'b10101000; //  856 : 168 - 0xa8 -- plane 1
      12'h359: dout  = 8'b11111100; //  857 : 252 - 0xfc
      12'h35A: dout  = 8'b11111000; //  858 : 248 - 0xf8
      12'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout  = 8'b11000000; //  862 : 192 - 0xc0
      12'h35F: dout  = 8'b11100000; //  863 : 224 - 0xe0
      12'h360: dout  = 8'b00000111; //  864 :   7 - 0x7 -- Sprite 0x36
      12'h361: dout  = 8'b00001111; //  865 :  15 - 0xf
      12'h362: dout  = 8'b00001110; //  866 :  14 - 0xe
      12'h363: dout  = 8'b00010100; //  867 :  20 - 0x14
      12'h364: dout  = 8'b00010110; //  868 :  22 - 0x16
      12'h365: dout  = 8'b00011000; //  869 :  24 - 0x18
      12'h366: dout  = 8'b00000000; //  870 :   0 - 0x0
      12'h367: dout  = 8'b00111111; //  871 :  63 - 0x3f
      12'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- plane 1
      12'h369: dout  = 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout  = 8'b00001111; //  874 :  15 - 0xf
      12'h36B: dout  = 8'b00011111; //  875 :  31 - 0x1f
      12'h36C: dout  = 8'b00011111; //  876 :  31 - 0x1f
      12'h36D: dout  = 8'b00011111; //  877 :  31 - 0x1f
      12'h36E: dout  = 8'b00000111; //  878 :   7 - 0x7
      12'h36F: dout  = 8'b00111100; //  879 :  60 - 0x3c
      12'h370: dout  = 8'b11000000; //  880 : 192 - 0xc0 -- Sprite 0x37
      12'h371: dout  = 8'b11111000; //  881 : 248 - 0xf8
      12'h372: dout  = 8'b01000000; //  882 :  64 - 0x40
      12'h373: dout  = 8'b01000000; //  883 :  64 - 0x40
      12'h374: dout  = 8'b00100000; //  884 :  32 - 0x20
      12'h375: dout  = 8'b01111000; //  885 : 120 - 0x78
      12'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout  = 8'b11000000; //  887 : 192 - 0xc0
      12'h378: dout  = 8'b00000000; //  888 :   0 - 0x0 -- plane 1
      12'h379: dout  = 8'b00000000; //  889 :   0 - 0x0
      12'h37A: dout  = 8'b11100000; //  890 : 224 - 0xe0
      12'h37B: dout  = 8'b11111000; //  891 : 248 - 0xf8
      12'h37C: dout  = 8'b11111100; //  892 : 252 - 0xfc
      12'h37D: dout  = 8'b11111000; //  893 : 248 - 0xf8
      12'h37E: dout  = 8'b11110000; //  894 : 240 - 0xf0
      12'h37F: dout  = 8'b11000000; //  895 : 192 - 0xc0
      12'h380: dout  = 8'b00111111; //  896 :  63 - 0x3f -- Sprite 0x38
      12'h381: dout  = 8'b00001110; //  897 :  14 - 0xe
      12'h382: dout  = 8'b00001111; //  898 :  15 - 0xf
      12'h383: dout  = 8'b00011111; //  899 :  31 - 0x1f
      12'h384: dout  = 8'b00111111; //  900 :  63 - 0x3f
      12'h385: dout  = 8'b01111100; //  901 : 124 - 0x7c
      12'h386: dout  = 8'b01110000; //  902 : 112 - 0x70
      12'h387: dout  = 8'b00111000; //  903 :  56 - 0x38
      12'h388: dout  = 8'b11111100; //  904 : 252 - 0xfc -- plane 1
      12'h389: dout  = 8'b11101101; //  905 : 237 - 0xed
      12'h38A: dout  = 8'b11000000; //  906 : 192 - 0xc0
      12'h38B: dout  = 8'b00000000; //  907 :   0 - 0x0
      12'h38C: dout  = 8'b00000000; //  908 :   0 - 0x0
      12'h38D: dout  = 8'b01100000; //  909 :  96 - 0x60
      12'h38E: dout  = 8'b01110000; //  910 : 112 - 0x70
      12'h38F: dout  = 8'b00111000; //  911 :  56 - 0x38
      12'h390: dout  = 8'b11110000; //  912 : 240 - 0xf0 -- Sprite 0x39
      12'h391: dout  = 8'b11111000; //  913 : 248 - 0xf8
      12'h392: dout  = 8'b11100100; //  914 : 228 - 0xe4
      12'h393: dout  = 8'b11111100; //  915 : 252 - 0xfc
      12'h394: dout  = 8'b11111100; //  916 : 252 - 0xfc
      12'h395: dout  = 8'b01111100; //  917 : 124 - 0x7c
      12'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      12'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout  = 8'b01111110; //  920 : 126 - 0x7e -- plane 1
      12'h399: dout  = 8'b00011110; //  921 :  30 - 0x1e
      12'h39A: dout  = 8'b00000100; //  922 :   4 - 0x4
      12'h39B: dout  = 8'b00001100; //  923 :  12 - 0xc
      12'h39C: dout  = 8'b00001100; //  924 :  12 - 0xc
      12'h39D: dout  = 8'b00001100; //  925 :  12 - 0xc
      12'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout  = 8'b00000111; //  928 :   7 - 0x7 -- Sprite 0x3a
      12'h3A1: dout  = 8'b00001111; //  929 :  15 - 0xf
      12'h3A2: dout  = 8'b00001110; //  930 :  14 - 0xe
      12'h3A3: dout  = 8'b00010100; //  931 :  20 - 0x14
      12'h3A4: dout  = 8'b00010110; //  932 :  22 - 0x16
      12'h3A5: dout  = 8'b00011000; //  933 :  24 - 0x18
      12'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout  = 8'b00001111; //  935 :  15 - 0xf
      12'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0 -- plane 1
      12'h3A9: dout  = 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout  = 8'b00001111; //  938 :  15 - 0xf
      12'h3AB: dout  = 8'b00011111; //  939 :  31 - 0x1f
      12'h3AC: dout  = 8'b00011111; //  940 :  31 - 0x1f
      12'h3AD: dout  = 8'b00011111; //  941 :  31 - 0x1f
      12'h3AE: dout  = 8'b00000111; //  942 :   7 - 0x7
      12'h3AF: dout  = 8'b00001101; //  943 :  13 - 0xd
      12'h3B0: dout  = 8'b00011111; //  944 :  31 - 0x1f -- Sprite 0x3b
      12'h3B1: dout  = 8'b00011111; //  945 :  31 - 0x1f
      12'h3B2: dout  = 8'b00011111; //  946 :  31 - 0x1f
      12'h3B3: dout  = 8'b00011100; //  947 :  28 - 0x1c
      12'h3B4: dout  = 8'b00001100; //  948 :  12 - 0xc
      12'h3B5: dout  = 8'b00000111; //  949 :   7 - 0x7
      12'h3B6: dout  = 8'b00000111; //  950 :   7 - 0x7
      12'h3B7: dout  = 8'b00000111; //  951 :   7 - 0x7
      12'h3B8: dout  = 8'b00011110; //  952 :  30 - 0x1e -- plane 1
      12'h3B9: dout  = 8'b00011100; //  953 :  28 - 0x1c
      12'h3BA: dout  = 8'b00011110; //  954 :  30 - 0x1e
      12'h3BB: dout  = 8'b00001111; //  955 :  15 - 0xf
      12'h3BC: dout  = 8'b00000111; //  956 :   7 - 0x7
      12'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout  = 8'b00000111; //  958 :   7 - 0x7
      12'h3BF: dout  = 8'b00000111; //  959 :   7 - 0x7
      12'h3C0: dout  = 8'b11100000; //  960 : 224 - 0xe0 -- Sprite 0x3c
      12'h3C1: dout  = 8'b01100000; //  961 :  96 - 0x60
      12'h3C2: dout  = 8'b11110000; //  962 : 240 - 0xf0
      12'h3C3: dout  = 8'b01110000; //  963 : 112 - 0x70
      12'h3C4: dout  = 8'b11100000; //  964 : 224 - 0xe0
      12'h3C5: dout  = 8'b11100000; //  965 : 224 - 0xe0
      12'h3C6: dout  = 8'b11110000; //  966 : 240 - 0xf0
      12'h3C7: dout  = 8'b10000000; //  967 : 128 - 0x80
      12'h3C8: dout  = 8'b01100000; //  968 :  96 - 0x60 -- plane 1
      12'h3C9: dout  = 8'b10010000; //  969 : 144 - 0x90
      12'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout  = 8'b10000000; //  971 : 128 - 0x80
      12'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout  = 8'b11100000; //  973 : 224 - 0xe0
      12'h3CE: dout  = 8'b11110000; //  974 : 240 - 0xf0
      12'h3CF: dout  = 8'b10000000; //  975 : 128 - 0x80
      12'h3D0: dout  = 8'b00000111; //  976 :   7 - 0x7 -- Sprite 0x3d
      12'h3D1: dout  = 8'b00011111; //  977 :  31 - 0x1f
      12'h3D2: dout  = 8'b00111111; //  978 :  63 - 0x3f
      12'h3D3: dout  = 8'b00010010; //  979 :  18 - 0x12
      12'h3D4: dout  = 8'b00010011; //  980 :  19 - 0x13
      12'h3D5: dout  = 8'b00001000; //  981 :   8 - 0x8
      12'h3D6: dout  = 8'b00011111; //  982 :  31 - 0x1f
      12'h3D7: dout  = 8'b00110001; //  983 :  49 - 0x31
      12'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0 -- plane 1
      12'h3D9: dout  = 8'b00010000; //  985 :  16 - 0x10
      12'h3DA: dout  = 8'b00111111; //  986 :  63 - 0x3f
      12'h3DB: dout  = 8'b01111111; //  987 : 127 - 0x7f
      12'h3DC: dout  = 8'b01111111; //  988 : 127 - 0x7f
      12'h3DD: dout  = 8'b00111111; //  989 :  63 - 0x3f
      12'h3DE: dout  = 8'b00000011; //  990 :   3 - 0x3
      12'h3DF: dout  = 8'b00001111; //  991 :  15 - 0xf
      12'h3E0: dout  = 8'b11000000; //  992 : 192 - 0xc0 -- Sprite 0x3e
      12'h3E1: dout  = 8'b11110000; //  993 : 240 - 0xf0
      12'h3E2: dout  = 8'b01000000; //  994 :  64 - 0x40
      12'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      12'h3E4: dout  = 8'b00110000; //  996 :  48 - 0x30
      12'h3E5: dout  = 8'b00011000; //  997 :  24 - 0x18
      12'h3E6: dout  = 8'b11000000; //  998 : 192 - 0xc0
      12'h3E7: dout  = 8'b11111000; //  999 : 248 - 0xf8
      12'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- plane 1
      12'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout  = 8'b11100000; // 1002 : 224 - 0xe0
      12'h3EB: dout  = 8'b11111000; // 1003 : 248 - 0xf8
      12'h3EC: dout  = 8'b11111100; // 1004 : 252 - 0xfc
      12'h3ED: dout  = 8'b11111000; // 1005 : 248 - 0xf8
      12'h3EE: dout  = 8'b10110000; // 1006 : 176 - 0xb0
      12'h3EF: dout  = 8'b00111000; // 1007 :  56 - 0x38
      12'h3F0: dout  = 8'b00110001; // 1008 :  49 - 0x31 -- Sprite 0x3f
      12'h3F1: dout  = 8'b00111001; // 1009 :  57 - 0x39
      12'h3F2: dout  = 8'b00011111; // 1010 :  31 - 0x1f
      12'h3F3: dout  = 8'b00011111; // 1011 :  31 - 0x1f
      12'h3F4: dout  = 8'b00001111; // 1012 :  15 - 0xf
      12'h3F5: dout  = 8'b01011111; // 1013 :  95 - 0x5f
      12'h3F6: dout  = 8'b01111110; // 1014 : 126 - 0x7e
      12'h3F7: dout  = 8'b00111100; // 1015 :  60 - 0x3c
      12'h3F8: dout  = 8'b00011111; // 1016 :  31 - 0x1f -- plane 1
      12'h3F9: dout  = 8'b00000111; // 1017 :   7 - 0x7
      12'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      12'h3FB: dout  = 8'b00001110; // 1019 :  14 - 0xe
      12'h3FC: dout  = 8'b00001111; // 1020 :  15 - 0xf
      12'h3FD: dout  = 8'b01010011; // 1021 :  83 - 0x53
      12'h3FE: dout  = 8'b01111100; // 1022 : 124 - 0x7c
      12'h3FF: dout  = 8'b00111100; // 1023 :  60 - 0x3c
      12'h400: dout  = 8'b11111000; // 1024 : 248 - 0xf8 -- Sprite 0x40
      12'h401: dout  = 8'b11111000; // 1025 : 248 - 0xf8
      12'h402: dout  = 8'b11110000; // 1026 : 240 - 0xf0
      12'h403: dout  = 8'b11100000; // 1027 : 224 - 0xe0
      12'h404: dout  = 8'b11100000; // 1028 : 224 - 0xe0
      12'h405: dout  = 8'b11000000; // 1029 : 192 - 0xc0
      12'h406: dout  = 8'b00000000; // 1030 :   0 - 0x0
      12'h407: dout  = 8'b00000000; // 1031 :   0 - 0x0
      12'h408: dout  = 8'b11111000; // 1032 : 248 - 0xf8 -- plane 1
      12'h409: dout  = 8'b11111000; // 1033 : 248 - 0xf8
      12'h40A: dout  = 8'b11110000; // 1034 : 240 - 0xf0
      12'h40B: dout  = 8'b00000000; // 1035 :   0 - 0x0
      12'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout  = 8'b10000000; // 1037 : 128 - 0x80
      12'h40E: dout  = 8'b00000000; // 1038 :   0 - 0x0
      12'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x41
      12'h411: dout  = 8'b11100000; // 1041 : 224 - 0xe0
      12'h412: dout  = 8'b11111100; // 1042 : 252 - 0xfc
      12'h413: dout  = 8'b00100111; // 1043 :  39 - 0x27
      12'h414: dout  = 8'b00100111; // 1044 :  39 - 0x27
      12'h415: dout  = 8'b00010001; // 1045 :  17 - 0x11
      12'h416: dout  = 8'b00111110; // 1046 :  62 - 0x3e
      12'h417: dout  = 8'b00000100; // 1047 :   4 - 0x4
      12'h418: dout  = 8'b00000111; // 1048 :   7 - 0x7 -- plane 1
      12'h419: dout  = 8'b00000111; // 1049 :   7 - 0x7
      12'h41A: dout  = 8'b00000011; // 1050 :   3 - 0x3
      12'h41B: dout  = 8'b11110111; // 1051 : 247 - 0xf7
      12'h41C: dout  = 8'b11111111; // 1052 : 255 - 0xff
      12'h41D: dout  = 8'b11111111; // 1053 : 255 - 0xff
      12'h41E: dout  = 8'b11111110; // 1054 : 254 - 0xfe
      12'h41F: dout  = 8'b11111100; // 1055 : 252 - 0xfc
      12'h420: dout  = 8'b00111111; // 1056 :  63 - 0x3f -- Sprite 0x42
      12'h421: dout  = 8'b01111111; // 1057 : 127 - 0x7f
      12'h422: dout  = 8'b00111111; // 1058 :  63 - 0x3f
      12'h423: dout  = 8'b00001111; // 1059 :  15 - 0xf
      12'h424: dout  = 8'b00011111; // 1060 :  31 - 0x1f
      12'h425: dout  = 8'b00111111; // 1061 :  63 - 0x3f
      12'h426: dout  = 8'b01111111; // 1062 : 127 - 0x7f
      12'h427: dout  = 8'b01001111; // 1063 :  79 - 0x4f
      12'h428: dout  = 8'b00111110; // 1064 :  62 - 0x3e -- plane 1
      12'h429: dout  = 8'b01111111; // 1065 : 127 - 0x7f
      12'h42A: dout  = 8'b11111111; // 1066 : 255 - 0xff
      12'h42B: dout  = 8'b11100010; // 1067 : 226 - 0xe2
      12'h42C: dout  = 8'b01010000; // 1068 :  80 - 0x50
      12'h42D: dout  = 8'b00111000; // 1069 :  56 - 0x38
      12'h42E: dout  = 8'b01110000; // 1070 : 112 - 0x70
      12'h42F: dout  = 8'b01000000; // 1071 :  64 - 0x40
      12'h430: dout  = 8'b11111000; // 1072 : 248 - 0xf8 -- Sprite 0x43
      12'h431: dout  = 8'b11111001; // 1073 : 249 - 0xf9
      12'h432: dout  = 8'b11111001; // 1074 : 249 - 0xf9
      12'h433: dout  = 8'b10110111; // 1075 : 183 - 0xb7
      12'h434: dout  = 8'b11111111; // 1076 : 255 - 0xff
      12'h435: dout  = 8'b11111111; // 1077 : 255 - 0xff
      12'h436: dout  = 8'b11100000; // 1078 : 224 - 0xe0
      12'h437: dout  = 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout  = 8'b11101000; // 1080 : 232 - 0xe8 -- plane 1
      12'h439: dout  = 8'b01110001; // 1081 : 113 - 0x71
      12'h43A: dout  = 8'b00000001; // 1082 :   1 - 0x1
      12'h43B: dout  = 8'b01001011; // 1083 :  75 - 0x4b
      12'h43C: dout  = 8'b00000011; // 1084 :   3 - 0x3
      12'h43D: dout  = 8'b00000011; // 1085 :   3 - 0x3
      12'h43E: dout  = 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout  = 8'b00000111; // 1088 :   7 - 0x7 -- Sprite 0x44
      12'h441: dout  = 8'b00000111; // 1089 :   7 - 0x7
      12'h442: dout  = 8'b00001111; // 1090 :  15 - 0xf
      12'h443: dout  = 8'b00111111; // 1091 :  63 - 0x3f
      12'h444: dout  = 8'b00111111; // 1092 :  63 - 0x3f
      12'h445: dout  = 8'b00111111; // 1093 :  63 - 0x3f
      12'h446: dout  = 8'b00100110; // 1094 :  38 - 0x26
      12'h447: dout  = 8'b00000100; // 1095 :   4 - 0x4
      12'h448: dout  = 8'b00000101; // 1096 :   5 - 0x5 -- plane 1
      12'h449: dout  = 8'b00000011; // 1097 :   3 - 0x3
      12'h44A: dout  = 8'b00000001; // 1098 :   1 - 0x1
      12'h44B: dout  = 8'b00110000; // 1099 :  48 - 0x30
      12'h44C: dout  = 8'b00110000; // 1100 :  48 - 0x30
      12'h44D: dout  = 8'b00110000; // 1101 :  48 - 0x30
      12'h44E: dout  = 8'b00100110; // 1102 :  38 - 0x26
      12'h44F: dout  = 8'b00000100; // 1103 :   4 - 0x4
      12'h450: dout  = 8'b11110000; // 1104 : 240 - 0xf0 -- Sprite 0x45
      12'h451: dout  = 8'b11110000; // 1105 : 240 - 0xf0
      12'h452: dout  = 8'b11110000; // 1106 : 240 - 0xf0
      12'h453: dout  = 8'b11100000; // 1107 : 224 - 0xe0
      12'h454: dout  = 8'b11000000; // 1108 : 192 - 0xc0
      12'h455: dout  = 8'b00000000; // 1109 :   0 - 0x0
      12'h456: dout  = 8'b00000000; // 1110 :   0 - 0x0
      12'h457: dout  = 8'b00000000; // 1111 :   0 - 0x0
      12'h458: dout  = 8'b11111110; // 1112 : 254 - 0xfe -- plane 1
      12'h459: dout  = 8'b11111100; // 1113 : 252 - 0xfc
      12'h45A: dout  = 8'b11100000; // 1114 : 224 - 0xe0
      12'h45B: dout  = 8'b00000000; // 1115 :   0 - 0x0
      12'h45C: dout  = 8'b00000000; // 1116 :   0 - 0x0
      12'h45D: dout  = 8'b00000000; // 1117 :   0 - 0x0
      12'h45E: dout  = 8'b00000000; // 1118 :   0 - 0x0
      12'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout  = 8'b00000111; // 1120 :   7 - 0x7 -- Sprite 0x46
      12'h461: dout  = 8'b00000111; // 1121 :   7 - 0x7
      12'h462: dout  = 8'b00001111; // 1122 :  15 - 0xf
      12'h463: dout  = 8'b00011111; // 1123 :  31 - 0x1f
      12'h464: dout  = 8'b00111111; // 1124 :  63 - 0x3f
      12'h465: dout  = 8'b00001111; // 1125 :  15 - 0xf
      12'h466: dout  = 8'b00011100; // 1126 :  28 - 0x1c
      12'h467: dout  = 8'b00011000; // 1127 :  24 - 0x18
      12'h468: dout  = 8'b00000101; // 1128 :   5 - 0x5 -- plane 1
      12'h469: dout  = 8'b00000011; // 1129 :   3 - 0x3
      12'h46A: dout  = 8'b00000001; // 1130 :   1 - 0x1
      12'h46B: dout  = 8'b00010000; // 1131 :  16 - 0x10
      12'h46C: dout  = 8'b00110000; // 1132 :  48 - 0x30
      12'h46D: dout  = 8'b00001100; // 1133 :  12 - 0xc
      12'h46E: dout  = 8'b00011100; // 1134 :  28 - 0x1c
      12'h46F: dout  = 8'b00011000; // 1135 :  24 - 0x18
      12'h470: dout  = 8'b11100000; // 1136 : 224 - 0xe0 -- Sprite 0x47
      12'h471: dout  = 8'b11100000; // 1137 : 224 - 0xe0
      12'h472: dout  = 8'b11100000; // 1138 : 224 - 0xe0
      12'h473: dout  = 8'b11100000; // 1139 : 224 - 0xe0
      12'h474: dout  = 8'b11000000; // 1140 : 192 - 0xc0
      12'h475: dout  = 8'b10000000; // 1141 : 128 - 0x80
      12'h476: dout  = 8'b00000000; // 1142 :   0 - 0x0
      12'h477: dout  = 8'b00000000; // 1143 :   0 - 0x0
      12'h478: dout  = 8'b11000000; // 1144 : 192 - 0xc0 -- plane 1
      12'h479: dout  = 8'b11100000; // 1145 : 224 - 0xe0
      12'h47A: dout  = 8'b11110000; // 1146 : 240 - 0xf0
      12'h47B: dout  = 8'b01111000; // 1147 : 120 - 0x78
      12'h47C: dout  = 8'b00011000; // 1148 :  24 - 0x18
      12'h47D: dout  = 8'b00001000; // 1149 :   8 - 0x8
      12'h47E: dout  = 8'b00000000; // 1150 :   0 - 0x0
      12'h47F: dout  = 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout  = 8'b00000111; // 1152 :   7 - 0x7 -- Sprite 0x48
      12'h481: dout  = 8'b00001111; // 1153 :  15 - 0xf
      12'h482: dout  = 8'b00011111; // 1154 :  31 - 0x1f
      12'h483: dout  = 8'b00001111; // 1155 :  15 - 0xf
      12'h484: dout  = 8'b00111111; // 1156 :  63 - 0x3f
      12'h485: dout  = 8'b00001111; // 1157 :  15 - 0xf
      12'h486: dout  = 8'b00011100; // 1158 :  28 - 0x1c
      12'h487: dout  = 8'b00011000; // 1159 :  24 - 0x18
      12'h488: dout  = 8'b00000111; // 1160 :   7 - 0x7 -- plane 1
      12'h489: dout  = 8'b00001111; // 1161 :  15 - 0xf
      12'h48A: dout  = 8'b00111110; // 1162 :  62 - 0x3e
      12'h48B: dout  = 8'b01111100; // 1163 : 124 - 0x7c
      12'h48C: dout  = 8'b00110000; // 1164 :  48 - 0x30
      12'h48D: dout  = 8'b00001100; // 1165 :  12 - 0xc
      12'h48E: dout  = 8'b00011100; // 1166 :  28 - 0x1c
      12'h48F: dout  = 8'b00011000; // 1167 :  24 - 0x18
      12'h490: dout  = 8'b11100000; // 1168 : 224 - 0xe0 -- Sprite 0x49
      12'h491: dout  = 8'b11100000; // 1169 : 224 - 0xe0
      12'h492: dout  = 8'b11100000; // 1170 : 224 - 0xe0
      12'h493: dout  = 8'b01000000; // 1171 :  64 - 0x40
      12'h494: dout  = 8'b11000000; // 1172 : 192 - 0xc0
      12'h495: dout  = 8'b10000000; // 1173 : 128 - 0x80
      12'h496: dout  = 8'b00000000; // 1174 :   0 - 0x0
      12'h497: dout  = 8'b00000000; // 1175 :   0 - 0x0
      12'h498: dout  = 8'b01100000; // 1176 :  96 - 0x60 -- plane 1
      12'h499: dout  = 8'b01100000; // 1177 :  96 - 0x60
      12'h49A: dout  = 8'b01100000; // 1178 :  96 - 0x60
      12'h49B: dout  = 8'b10000000; // 1179 : 128 - 0x80
      12'h49C: dout  = 8'b00000000; // 1180 :   0 - 0x0
      12'h49D: dout  = 8'b00000000; // 1181 :   0 - 0x0
      12'h49E: dout  = 8'b00000000; // 1182 :   0 - 0x0
      12'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      12'h4A0: dout  = 8'b01111111; // 1184 : 127 - 0x7f -- Sprite 0x4a
      12'h4A1: dout  = 8'b11111111; // 1185 : 255 - 0xff
      12'h4A2: dout  = 8'b11111111; // 1186 : 255 - 0xff
      12'h4A3: dout  = 8'b11111011; // 1187 : 251 - 0xfb
      12'h4A4: dout  = 8'b00001111; // 1188 :  15 - 0xf
      12'h4A5: dout  = 8'b00001111; // 1189 :  15 - 0xf
      12'h4A6: dout  = 8'b00001111; // 1190 :  15 - 0xf
      12'h4A7: dout  = 8'b00011111; // 1191 :  31 - 0x1f
      12'h4A8: dout  = 8'b01110011; // 1192 : 115 - 0x73 -- plane 1
      12'h4A9: dout  = 8'b11110011; // 1193 : 243 - 0xf3
      12'h4AA: dout  = 8'b11110000; // 1194 : 240 - 0xf0
      12'h4AB: dout  = 8'b11110100; // 1195 : 244 - 0xf4
      12'h4AC: dout  = 8'b11110000; // 1196 : 240 - 0xf0
      12'h4AD: dout  = 8'b11110000; // 1197 : 240 - 0xf0
      12'h4AE: dout  = 8'b01110000; // 1198 : 112 - 0x70
      12'h4AF: dout  = 8'b01100000; // 1199 :  96 - 0x60
      12'h4B0: dout  = 8'b00111111; // 1200 :  63 - 0x3f -- Sprite 0x4b
      12'h4B1: dout  = 8'b01111110; // 1201 : 126 - 0x7e
      12'h4B2: dout  = 8'b01111100; // 1202 : 124 - 0x7c
      12'h4B3: dout  = 8'b01111100; // 1203 : 124 - 0x7c
      12'h4B4: dout  = 8'b00111100; // 1204 :  60 - 0x3c
      12'h4B5: dout  = 8'b00111100; // 1205 :  60 - 0x3c
      12'h4B6: dout  = 8'b11111100; // 1206 : 252 - 0xfc
      12'h4B7: dout  = 8'b11111100; // 1207 : 252 - 0xfc
      12'h4B8: dout  = 8'b00000000; // 1208 :   0 - 0x0 -- plane 1
      12'h4B9: dout  = 8'b00000000; // 1209 :   0 - 0x0
      12'h4BA: dout  = 8'b00000000; // 1210 :   0 - 0x0
      12'h4BB: dout  = 8'b00000000; // 1211 :   0 - 0x0
      12'h4BC: dout  = 8'b00111100; // 1212 :  60 - 0x3c
      12'h4BD: dout  = 8'b00111100; // 1213 :  60 - 0x3c
      12'h4BE: dout  = 8'b11111100; // 1214 : 252 - 0xfc
      12'h4BF: dout  = 8'b11111100; // 1215 : 252 - 0xfc
      12'h4C0: dout  = 8'b01100000; // 1216 :  96 - 0x60 -- Sprite 0x4c
      12'h4C1: dout  = 8'b01110000; // 1217 : 112 - 0x70
      12'h4C2: dout  = 8'b00011000; // 1218 :  24 - 0x18
      12'h4C3: dout  = 8'b00001000; // 1219 :   8 - 0x8
      12'h4C4: dout  = 8'b00001111; // 1220 :  15 - 0xf
      12'h4C5: dout  = 8'b00011111; // 1221 :  31 - 0x1f
      12'h4C6: dout  = 8'b00111111; // 1222 :  63 - 0x3f
      12'h4C7: dout  = 8'b01111111; // 1223 : 127 - 0x7f
      12'h4C8: dout  = 8'b01111111; // 1224 : 127 - 0x7f -- plane 1
      12'h4C9: dout  = 8'b01111111; // 1225 : 127 - 0x7f
      12'h4CA: dout  = 8'b00011111; // 1226 :  31 - 0x1f
      12'h4CB: dout  = 8'b00000111; // 1227 :   7 - 0x7
      12'h4CC: dout  = 8'b00001011; // 1228 :  11 - 0xb
      12'h4CD: dout  = 8'b00011011; // 1229 :  27 - 0x1b
      12'h4CE: dout  = 8'b00111011; // 1230 :  59 - 0x3b
      12'h4CF: dout  = 8'b01111011; // 1231 : 123 - 0x7b
      12'h4D0: dout  = 8'b11111100; // 1232 : 252 - 0xfc -- Sprite 0x4d
      12'h4D1: dout  = 8'b01111100; // 1233 : 124 - 0x7c
      12'h4D2: dout  = 8'b00000000; // 1234 :   0 - 0x0
      12'h4D3: dout  = 8'b00100000; // 1235 :  32 - 0x20
      12'h4D4: dout  = 8'b11110000; // 1236 : 240 - 0xf0
      12'h4D5: dout  = 8'b11111000; // 1237 : 248 - 0xf8
      12'h4D6: dout  = 8'b11111100; // 1238 : 252 - 0xfc
      12'h4D7: dout  = 8'b11111110; // 1239 : 254 - 0xfe
      12'h4D8: dout  = 8'b11111100; // 1240 : 252 - 0xfc -- plane 1
      12'h4D9: dout  = 8'b11111100; // 1241 : 252 - 0xfc
      12'h4DA: dout  = 8'b11111000; // 1242 : 248 - 0xf8
      12'h4DB: dout  = 8'b11100000; // 1243 : 224 - 0xe0
      12'h4DC: dout  = 8'b11010000; // 1244 : 208 - 0xd0
      12'h4DD: dout  = 8'b11011000; // 1245 : 216 - 0xd8
      12'h4DE: dout  = 8'b11011100; // 1246 : 220 - 0xdc
      12'h4DF: dout  = 8'b11011110; // 1247 : 222 - 0xde
      12'h4E0: dout  = 8'b00001011; // 1248 :  11 - 0xb -- Sprite 0x4e
      12'h4E1: dout  = 8'b00001111; // 1249 :  15 - 0xf
      12'h4E2: dout  = 8'b00011111; // 1250 :  31 - 0x1f
      12'h4E3: dout  = 8'b00011110; // 1251 :  30 - 0x1e
      12'h4E4: dout  = 8'b00111100; // 1252 :  60 - 0x3c
      12'h4E5: dout  = 8'b00111100; // 1253 :  60 - 0x3c
      12'h4E6: dout  = 8'b00111100; // 1254 :  60 - 0x3c
      12'h4E7: dout  = 8'b01111100; // 1255 : 124 - 0x7c
      12'h4E8: dout  = 8'b11000100; // 1256 : 196 - 0xc4 -- plane 1
      12'h4E9: dout  = 8'b11100000; // 1257 : 224 - 0xe0
      12'h4EA: dout  = 8'b11100000; // 1258 : 224 - 0xe0
      12'h4EB: dout  = 8'b01000000; // 1259 :  64 - 0x40
      12'h4EC: dout  = 8'b00000000; // 1260 :   0 - 0x0
      12'h4ED: dout  = 8'b00111100; // 1261 :  60 - 0x3c
      12'h4EE: dout  = 8'b00111100; // 1262 :  60 - 0x3c
      12'h4EF: dout  = 8'b01111100; // 1263 : 124 - 0x7c
      12'h4F0: dout  = 8'b00011111; // 1264 :  31 - 0x1f -- Sprite 0x4f
      12'h4F1: dout  = 8'b00111111; // 1265 :  63 - 0x3f
      12'h4F2: dout  = 8'b00001101; // 1266 :  13 - 0xd
      12'h4F3: dout  = 8'b00000111; // 1267 :   7 - 0x7
      12'h4F4: dout  = 8'b00001111; // 1268 :  15 - 0xf
      12'h4F5: dout  = 8'b00001110; // 1269 :  14 - 0xe
      12'h4F6: dout  = 8'b00011100; // 1270 :  28 - 0x1c
      12'h4F7: dout  = 8'b00111100; // 1271 :  60 - 0x3c
      12'h4F8: dout  = 8'b00011101; // 1272 :  29 - 0x1d -- plane 1
      12'h4F9: dout  = 8'b00111100; // 1273 :  60 - 0x3c
      12'h4FA: dout  = 8'b00111010; // 1274 :  58 - 0x3a
      12'h4FB: dout  = 8'b00111000; // 1275 :  56 - 0x38
      12'h4FC: dout  = 8'b00110000; // 1276 :  48 - 0x30
      12'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      12'h4FE: dout  = 8'b00011100; // 1278 :  28 - 0x1c
      12'h4FF: dout  = 8'b00111100; // 1279 :  60 - 0x3c
      12'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0x50
      12'h501: dout  = 8'b00000000; // 1281 :   0 - 0x0
      12'h502: dout  = 8'b00000000; // 1282 :   0 - 0x0
      12'h503: dout  = 8'b00000000; // 1283 :   0 - 0x0
      12'h504: dout  = 8'b00000000; // 1284 :   0 - 0x0
      12'h505: dout  = 8'b00000000; // 1285 :   0 - 0x0
      12'h506: dout  = 8'b00000000; // 1286 :   0 - 0x0
      12'h507: dout  = 8'b00000000; // 1287 :   0 - 0x0
      12'h508: dout  = 8'b00100010; // 1288 :  34 - 0x22 -- plane 1
      12'h509: dout  = 8'b01010101; // 1289 :  85 - 0x55
      12'h50A: dout  = 8'b01010101; // 1290 :  85 - 0x55
      12'h50B: dout  = 8'b01010101; // 1291 :  85 - 0x55
      12'h50C: dout  = 8'b01010101; // 1292 :  85 - 0x55
      12'h50D: dout  = 8'b01010101; // 1293 :  85 - 0x55
      12'h50E: dout  = 8'b01110111; // 1294 : 119 - 0x77
      12'h50F: dout  = 8'b00100010; // 1295 :  34 - 0x22
      12'h510: dout  = 8'b00000000; // 1296 :   0 - 0x0 -- Sprite 0x51
      12'h511: dout  = 8'b00000111; // 1297 :   7 - 0x7
      12'h512: dout  = 8'b00011111; // 1298 :  31 - 0x1f
      12'h513: dout  = 8'b11111111; // 1299 : 255 - 0xff
      12'h514: dout  = 8'b00000111; // 1300 :   7 - 0x7
      12'h515: dout  = 8'b00011111; // 1301 :  31 - 0x1f
      12'h516: dout  = 8'b00001111; // 1302 :  15 - 0xf
      12'h517: dout  = 8'b00000110; // 1303 :   6 - 0x6
      12'h518: dout  = 8'b00000000; // 1304 :   0 - 0x0 -- plane 1
      12'h519: dout  = 8'b00000000; // 1305 :   0 - 0x0
      12'h51A: dout  = 8'b00000000; // 1306 :   0 - 0x0
      12'h51B: dout  = 8'b00000000; // 1307 :   0 - 0x0
      12'h51C: dout  = 8'b00000000; // 1308 :   0 - 0x0
      12'h51D: dout  = 8'b00000000; // 1309 :   0 - 0x0
      12'h51E: dout  = 8'b00000000; // 1310 :   0 - 0x0
      12'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      12'h520: dout  = 8'b00111111; // 1312 :  63 - 0x3f -- Sprite 0x52
      12'h521: dout  = 8'b11111111; // 1313 : 255 - 0xff
      12'h522: dout  = 8'b11111111; // 1314 : 255 - 0xff
      12'h523: dout  = 8'b11111111; // 1315 : 255 - 0xff
      12'h524: dout  = 8'b11111111; // 1316 : 255 - 0xff
      12'h525: dout  = 8'b11111111; // 1317 : 255 - 0xff
      12'h526: dout  = 8'b11111011; // 1318 : 251 - 0xfb
      12'h527: dout  = 8'b01110110; // 1319 : 118 - 0x76
      12'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- plane 1
      12'h529: dout  = 8'b00000000; // 1321 :   0 - 0x0
      12'h52A: dout  = 8'b11001111; // 1322 : 207 - 0xcf
      12'h52B: dout  = 8'b00000111; // 1323 :   7 - 0x7
      12'h52C: dout  = 8'b01111111; // 1324 : 127 - 0x7f
      12'h52D: dout  = 8'b00000000; // 1325 :   0 - 0x0
      12'h52E: dout  = 8'b00000000; // 1326 :   0 - 0x0
      12'h52F: dout  = 8'b00000000; // 1327 :   0 - 0x0
      12'h530: dout  = 8'b00100000; // 1328 :  32 - 0x20 -- Sprite 0x53
      12'h531: dout  = 8'b11111000; // 1329 : 248 - 0xf8
      12'h532: dout  = 8'b11111111; // 1330 : 255 - 0xff
      12'h533: dout  = 8'b11000011; // 1331 : 195 - 0xc3
      12'h534: dout  = 8'b11111101; // 1332 : 253 - 0xfd
      12'h535: dout  = 8'b11111110; // 1333 : 254 - 0xfe
      12'h536: dout  = 8'b11110000; // 1334 : 240 - 0xf0
      12'h537: dout  = 8'b01000000; // 1335 :  64 - 0x40
      12'h538: dout  = 8'b00000000; // 1336 :   0 - 0x0 -- plane 1
      12'h539: dout  = 8'b00000000; // 1337 :   0 - 0x0
      12'h53A: dout  = 8'b00111100; // 1338 :  60 - 0x3c
      12'h53B: dout  = 8'b11111100; // 1339 : 252 - 0xfc
      12'h53C: dout  = 8'b11111110; // 1340 : 254 - 0xfe
      12'h53D: dout  = 8'b11100000; // 1341 : 224 - 0xe0
      12'h53E: dout  = 8'b00000000; // 1342 :   0 - 0x0
      12'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      12'h540: dout  = 8'b01000000; // 1344 :  64 - 0x40 -- Sprite 0x54
      12'h541: dout  = 8'b11100000; // 1345 : 224 - 0xe0
      12'h542: dout  = 8'b01000000; // 1346 :  64 - 0x40
      12'h543: dout  = 8'b01000000; // 1347 :  64 - 0x40
      12'h544: dout  = 8'b01000001; // 1348 :  65 - 0x41
      12'h545: dout  = 8'b01000001; // 1349 :  65 - 0x41
      12'h546: dout  = 8'b01001111; // 1350 :  79 - 0x4f
      12'h547: dout  = 8'b01000111; // 1351 :  71 - 0x47
      12'h548: dout  = 8'b01000000; // 1352 :  64 - 0x40 -- plane 1
      12'h549: dout  = 8'b11100000; // 1353 : 224 - 0xe0
      12'h54A: dout  = 8'b01000000; // 1354 :  64 - 0x40
      12'h54B: dout  = 8'b00111111; // 1355 :  63 - 0x3f
      12'h54C: dout  = 8'b00111110; // 1356 :  62 - 0x3e
      12'h54D: dout  = 8'b00111110; // 1357 :  62 - 0x3e
      12'h54E: dout  = 8'b00110000; // 1358 :  48 - 0x30
      12'h54F: dout  = 8'b00111000; // 1359 :  56 - 0x38
      12'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0x55
      12'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      12'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      12'h553: dout  = 8'b00000000; // 1363 :   0 - 0x0
      12'h554: dout  = 8'b00000000; // 1364 :   0 - 0x0
      12'h555: dout  = 8'b00000000; // 1365 :   0 - 0x0
      12'h556: dout  = 8'b11100000; // 1366 : 224 - 0xe0
      12'h557: dout  = 8'b11000000; // 1367 : 192 - 0xc0
      12'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0 -- plane 1
      12'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout  = 8'b11111000; // 1371 : 248 - 0xf8
      12'h55C: dout  = 8'b11111000; // 1372 : 248 - 0xf8
      12'h55D: dout  = 8'b11111000; // 1373 : 248 - 0xf8
      12'h55E: dout  = 8'b00011000; // 1374 :  24 - 0x18
      12'h55F: dout  = 8'b00111000; // 1375 :  56 - 0x38
      12'h560: dout  = 8'b01000011; // 1376 :  67 - 0x43 -- Sprite 0x56
      12'h561: dout  = 8'b01000110; // 1377 :  70 - 0x46
      12'h562: dout  = 8'b01000100; // 1378 :  68 - 0x44
      12'h563: dout  = 8'b01000000; // 1379 :  64 - 0x40
      12'h564: dout  = 8'b01000000; // 1380 :  64 - 0x40
      12'h565: dout  = 8'b01000000; // 1381 :  64 - 0x40
      12'h566: dout  = 8'b01000000; // 1382 :  64 - 0x40
      12'h567: dout  = 8'b01000000; // 1383 :  64 - 0x40
      12'h568: dout  = 8'b00111100; // 1384 :  60 - 0x3c -- plane 1
      12'h569: dout  = 8'b00111001; // 1385 :  57 - 0x39
      12'h56A: dout  = 8'b00111011; // 1386 :  59 - 0x3b
      12'h56B: dout  = 8'b00111111; // 1387 :  63 - 0x3f
      12'h56C: dout  = 8'b00000000; // 1388 :   0 - 0x0
      12'h56D: dout  = 8'b00000000; // 1389 :   0 - 0x0
      12'h56E: dout  = 8'b00000000; // 1390 :   0 - 0x0
      12'h56F: dout  = 8'b00000000; // 1391 :   0 - 0x0
      12'h570: dout  = 8'b10000000; // 1392 : 128 - 0x80 -- Sprite 0x57
      12'h571: dout  = 8'b11000000; // 1393 : 192 - 0xc0
      12'h572: dout  = 8'b01000000; // 1394 :  64 - 0x40
      12'h573: dout  = 8'b00000000; // 1395 :   0 - 0x0
      12'h574: dout  = 8'b00000000; // 1396 :   0 - 0x0
      12'h575: dout  = 8'b00000000; // 1397 :   0 - 0x0
      12'h576: dout  = 8'b00000000; // 1398 :   0 - 0x0
      12'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout  = 8'b01111000; // 1400 : 120 - 0x78 -- plane 1
      12'h579: dout  = 8'b00111000; // 1401 :  56 - 0x38
      12'h57A: dout  = 8'b10111000; // 1402 : 184 - 0xb8
      12'h57B: dout  = 8'b11111000; // 1403 : 248 - 0xf8
      12'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      12'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      12'h57E: dout  = 8'b00000000; // 1406 :   0 - 0x0
      12'h57F: dout  = 8'b00000000; // 1407 :   0 - 0x0
      12'h580: dout  = 8'b00110001; // 1408 :  49 - 0x31 -- Sprite 0x58
      12'h581: dout  = 8'b00110000; // 1409 :  48 - 0x30
      12'h582: dout  = 8'b00111000; // 1410 :  56 - 0x38
      12'h583: dout  = 8'b01111100; // 1411 : 124 - 0x7c
      12'h584: dout  = 8'b01111111; // 1412 : 127 - 0x7f
      12'h585: dout  = 8'b11111111; // 1413 : 255 - 0xff
      12'h586: dout  = 8'b11111111; // 1414 : 255 - 0xff
      12'h587: dout  = 8'b11111011; // 1415 : 251 - 0xfb
      12'h588: dout  = 8'b00111111; // 1416 :  63 - 0x3f -- plane 1
      12'h589: dout  = 8'b00111111; // 1417 :  63 - 0x3f
      12'h58A: dout  = 8'b00001111; // 1418 :  15 - 0xf
      12'h58B: dout  = 8'b01110111; // 1419 : 119 - 0x77
      12'h58C: dout  = 8'b01110111; // 1420 : 119 - 0x77
      12'h58D: dout  = 8'b11110111; // 1421 : 247 - 0xf7
      12'h58E: dout  = 8'b11110111; // 1422 : 247 - 0xf7
      12'h58F: dout  = 8'b11110111; // 1423 : 247 - 0xf7
      12'h590: dout  = 8'b00010000; // 1424 :  16 - 0x10 -- Sprite 0x59
      12'h591: dout  = 8'b01111110; // 1425 : 126 - 0x7e
      12'h592: dout  = 8'b00111110; // 1426 :  62 - 0x3e
      12'h593: dout  = 8'b00000000; // 1427 :   0 - 0x0
      12'h594: dout  = 8'b00011110; // 1428 :  30 - 0x1e
      12'h595: dout  = 8'b11111110; // 1429 : 254 - 0xfe
      12'h596: dout  = 8'b11111111; // 1430 : 255 - 0xff
      12'h597: dout  = 8'b11111111; // 1431 : 255 - 0xff
      12'h598: dout  = 8'b11111111; // 1432 : 255 - 0xff -- plane 1
      12'h599: dout  = 8'b11111110; // 1433 : 254 - 0xfe
      12'h59A: dout  = 8'b11111110; // 1434 : 254 - 0xfe
      12'h59B: dout  = 8'b11111110; // 1435 : 254 - 0xfe
      12'h59C: dout  = 8'b11111010; // 1436 : 250 - 0xfa
      12'h59D: dout  = 8'b11111010; // 1437 : 250 - 0xfa
      12'h59E: dout  = 8'b11110011; // 1438 : 243 - 0xf3
      12'h59F: dout  = 8'b11100111; // 1439 : 231 - 0xe7
      12'h5A0: dout  = 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0x5a
      12'h5A1: dout  = 8'b11111111; // 1441 : 255 - 0xff
      12'h5A2: dout  = 8'b11100011; // 1442 : 227 - 0xe3
      12'h5A3: dout  = 8'b11000011; // 1443 : 195 - 0xc3
      12'h5A4: dout  = 8'b10000111; // 1444 : 135 - 0x87
      12'h5A5: dout  = 8'b01001000; // 1445 :  72 - 0x48
      12'h5A6: dout  = 8'b00111100; // 1446 :  60 - 0x3c
      12'h5A7: dout  = 8'b11111100; // 1447 : 252 - 0xfc
      12'h5A8: dout  = 8'b11110000; // 1448 : 240 - 0xf0 -- plane 1
      12'h5A9: dout  = 8'b11111000; // 1449 : 248 - 0xf8
      12'h5AA: dout  = 8'b11111100; // 1450 : 252 - 0xfc
      12'h5AB: dout  = 8'b01111100; // 1451 : 124 - 0x7c
      12'h5AC: dout  = 8'b01111000; // 1452 : 120 - 0x78
      12'h5AD: dout  = 8'b00111000; // 1453 :  56 - 0x38
      12'h5AE: dout  = 8'b00111100; // 1454 :  60 - 0x3c
      12'h5AF: dout  = 8'b11111100; // 1455 : 252 - 0xfc
      12'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0x5b
      12'h5B1: dout  = 8'b11111111; // 1457 : 255 - 0xff
      12'h5B2: dout  = 8'b11000011; // 1458 : 195 - 0xc3
      12'h5B3: dout  = 8'b10000011; // 1459 : 131 - 0x83
      12'h5B4: dout  = 8'b10000011; // 1460 : 131 - 0x83
      12'h5B5: dout  = 8'b11111111; // 1461 : 255 - 0xff
      12'h5B6: dout  = 8'b11111111; // 1462 : 255 - 0xff
      12'h5B7: dout  = 8'b11111111; // 1463 : 255 - 0xff
      12'h5B8: dout  = 8'b11111111; // 1464 : 255 - 0xff -- plane 1
      12'h5B9: dout  = 8'b00000000; // 1465 :   0 - 0x0
      12'h5BA: dout  = 8'b11000011; // 1466 : 195 - 0xc3
      12'h5BB: dout  = 8'b10000001; // 1467 : 129 - 0x81
      12'h5BC: dout  = 8'b10000001; // 1468 : 129 - 0x81
      12'h5BD: dout  = 8'b11000011; // 1469 : 195 - 0xc3
      12'h5BE: dout  = 8'b11111111; // 1470 : 255 - 0xff
      12'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout  = 8'b00011111; // 1472 :  31 - 0x1f -- Sprite 0x5c
      12'h5C1: dout  = 8'b00011111; // 1473 :  31 - 0x1f
      12'h5C2: dout  = 8'b00001111; // 1474 :  15 - 0xf
      12'h5C3: dout  = 8'b00000111; // 1475 :   7 - 0x7
      12'h5C4: dout  = 8'b00000001; // 1476 :   1 - 0x1
      12'h5C5: dout  = 8'b00000000; // 1477 :   0 - 0x0
      12'h5C6: dout  = 8'b00000000; // 1478 :   0 - 0x0
      12'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout  = 8'b00000000; // 1480 :   0 - 0x0 -- plane 1
      12'h5C9: dout  = 8'b00000000; // 1481 :   0 - 0x0
      12'h5CA: dout  = 8'b00000000; // 1482 :   0 - 0x0
      12'h5CB: dout  = 8'b00000000; // 1483 :   0 - 0x0
      12'h5CC: dout  = 8'b00000000; // 1484 :   0 - 0x0
      12'h5CD: dout  = 8'b00000000; // 1485 :   0 - 0x0
      12'h5CE: dout  = 8'b00000000; // 1486 :   0 - 0x0
      12'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout  = 8'b11110000; // 1488 : 240 - 0xf0 -- Sprite 0x5d
      12'h5D1: dout  = 8'b11111011; // 1489 : 251 - 0xfb
      12'h5D2: dout  = 8'b11111111; // 1490 : 255 - 0xff
      12'h5D3: dout  = 8'b11111111; // 1491 : 255 - 0xff
      12'h5D4: dout  = 8'b11111110; // 1492 : 254 - 0xfe
      12'h5D5: dout  = 8'b00111110; // 1493 :  62 - 0x3e
      12'h5D6: dout  = 8'b00001100; // 1494 :  12 - 0xc
      12'h5D7: dout  = 8'b00000100; // 1495 :   4 - 0x4
      12'h5D8: dout  = 8'b00000000; // 1496 :   0 - 0x0 -- plane 1
      12'h5D9: dout  = 8'b00001011; // 1497 :  11 - 0xb
      12'h5DA: dout  = 8'b00011111; // 1498 :  31 - 0x1f
      12'h5DB: dout  = 8'b00011111; // 1499 :  31 - 0x1f
      12'h5DC: dout  = 8'b00011110; // 1500 :  30 - 0x1e
      12'h5DD: dout  = 8'b00111110; // 1501 :  62 - 0x3e
      12'h5DE: dout  = 8'b00001100; // 1502 :  12 - 0xc
      12'h5DF: dout  = 8'b00000100; // 1503 :   4 - 0x4
      12'h5E0: dout  = 8'b00011111; // 1504 :  31 - 0x1f -- Sprite 0x5e
      12'h5E1: dout  = 8'b00011111; // 1505 :  31 - 0x1f
      12'h5E2: dout  = 8'b00001111; // 1506 :  15 - 0xf
      12'h5E3: dout  = 8'b00001111; // 1507 :  15 - 0xf
      12'h5E4: dout  = 8'b00000111; // 1508 :   7 - 0x7
      12'h5E5: dout  = 8'b00000000; // 1509 :   0 - 0x0
      12'h5E6: dout  = 8'b00000000; // 1510 :   0 - 0x0
      12'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout  = 8'b00000000; // 1512 :   0 - 0x0 -- plane 1
      12'h5E9: dout  = 8'b00000000; // 1513 :   0 - 0x0
      12'h5EA: dout  = 8'b00000000; // 1514 :   0 - 0x0
      12'h5EB: dout  = 8'b00000000; // 1515 :   0 - 0x0
      12'h5EC: dout  = 8'b00000000; // 1516 :   0 - 0x0
      12'h5ED: dout  = 8'b00000000; // 1517 :   0 - 0x0
      12'h5EE: dout  = 8'b00000000; // 1518 :   0 - 0x0
      12'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout  = 8'b11111011; // 1520 : 251 - 0xfb -- Sprite 0x5f
      12'h5F1: dout  = 8'b11111111; // 1521 : 255 - 0xff
      12'h5F2: dout  = 8'b11111111; // 1522 : 255 - 0xff
      12'h5F3: dout  = 8'b11111111; // 1523 : 255 - 0xff
      12'h5F4: dout  = 8'b11111111; // 1524 : 255 - 0xff
      12'h5F5: dout  = 8'b00000000; // 1525 :   0 - 0x0
      12'h5F6: dout  = 8'b00000000; // 1526 :   0 - 0x0
      12'h5F7: dout  = 8'b00000000; // 1527 :   0 - 0x0
      12'h5F8: dout  = 8'b00000011; // 1528 :   3 - 0x3 -- plane 1
      12'h5F9: dout  = 8'b00001111; // 1529 :  15 - 0xf
      12'h5FA: dout  = 8'b00001111; // 1530 :  15 - 0xf
      12'h5FB: dout  = 8'b00001111; // 1531 :  15 - 0xf
      12'h5FC: dout  = 8'b00001111; // 1532 :  15 - 0xf
      12'h5FD: dout  = 8'b00000000; // 1533 :   0 - 0x0
      12'h5FE: dout  = 8'b00000000; // 1534 :   0 - 0x0
      12'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0x60
      12'h601: dout  = 8'b00011000; // 1537 :  24 - 0x18
      12'h602: dout  = 8'b00111100; // 1538 :  60 - 0x3c
      12'h603: dout  = 8'b01111110; // 1539 : 126 - 0x7e
      12'h604: dout  = 8'b01101110; // 1540 : 110 - 0x6e
      12'h605: dout  = 8'b11011111; // 1541 : 223 - 0xdf
      12'h606: dout  = 8'b11011111; // 1542 : 223 - 0xdf
      12'h607: dout  = 8'b11011111; // 1543 : 223 - 0xdf
      12'h608: dout  = 8'b00000000; // 1544 :   0 - 0x0 -- plane 1
      12'h609: dout  = 8'b00011000; // 1545 :  24 - 0x18
      12'h60A: dout  = 8'b00111100; // 1546 :  60 - 0x3c
      12'h60B: dout  = 8'b01111110; // 1547 : 126 - 0x7e
      12'h60C: dout  = 8'b01110110; // 1548 : 118 - 0x76
      12'h60D: dout  = 8'b11111011; // 1549 : 251 - 0xfb
      12'h60E: dout  = 8'b11111011; // 1550 : 251 - 0xfb
      12'h60F: dout  = 8'b11111011; // 1551 : 251 - 0xfb
      12'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0x61
      12'h611: dout  = 8'b00011000; // 1553 :  24 - 0x18
      12'h612: dout  = 8'b00011000; // 1554 :  24 - 0x18
      12'h613: dout  = 8'b00111100; // 1555 :  60 - 0x3c
      12'h614: dout  = 8'b00111100; // 1556 :  60 - 0x3c
      12'h615: dout  = 8'b00111100; // 1557 :  60 - 0x3c
      12'h616: dout  = 8'b00111100; // 1558 :  60 - 0x3c
      12'h617: dout  = 8'b00011100; // 1559 :  28 - 0x1c
      12'h618: dout  = 8'b00000000; // 1560 :   0 - 0x0 -- plane 1
      12'h619: dout  = 8'b00010000; // 1561 :  16 - 0x10
      12'h61A: dout  = 8'b00010000; // 1562 :  16 - 0x10
      12'h61B: dout  = 8'b00100000; // 1563 :  32 - 0x20
      12'h61C: dout  = 8'b00100000; // 1564 :  32 - 0x20
      12'h61D: dout  = 8'b00100000; // 1565 :  32 - 0x20
      12'h61E: dout  = 8'b00100000; // 1566 :  32 - 0x20
      12'h61F: dout  = 8'b00100000; // 1567 :  32 - 0x20
      12'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0x62
      12'h621: dout  = 8'b00001000; // 1569 :   8 - 0x8
      12'h622: dout  = 8'b00001000; // 1570 :   8 - 0x8
      12'h623: dout  = 8'b00001000; // 1571 :   8 - 0x8
      12'h624: dout  = 8'b00001000; // 1572 :   8 - 0x8
      12'h625: dout  = 8'b00001000; // 1573 :   8 - 0x8
      12'h626: dout  = 8'b00001000; // 1574 :   8 - 0x8
      12'h627: dout  = 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout  = 8'b00000000; // 1576 :   0 - 0x0 -- plane 1
      12'h629: dout  = 8'b00001000; // 1577 :   8 - 0x8
      12'h62A: dout  = 8'b00001000; // 1578 :   8 - 0x8
      12'h62B: dout  = 8'b00001000; // 1579 :   8 - 0x8
      12'h62C: dout  = 8'b00001000; // 1580 :   8 - 0x8
      12'h62D: dout  = 8'b00001000; // 1581 :   8 - 0x8
      12'h62E: dout  = 8'b00001000; // 1582 :   8 - 0x8
      12'h62F: dout  = 8'b00001000; // 1583 :   8 - 0x8
      12'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0x63
      12'h631: dout  = 8'b00001000; // 1585 :   8 - 0x8
      12'h632: dout  = 8'b00001000; // 1586 :   8 - 0x8
      12'h633: dout  = 8'b00000100; // 1587 :   4 - 0x4
      12'h634: dout  = 8'b00000100; // 1588 :   4 - 0x4
      12'h635: dout  = 8'b00000100; // 1589 :   4 - 0x4
      12'h636: dout  = 8'b00000100; // 1590 :   4 - 0x4
      12'h637: dout  = 8'b00000100; // 1591 :   4 - 0x4
      12'h638: dout  = 8'b00000000; // 1592 :   0 - 0x0 -- plane 1
      12'h639: dout  = 8'b00010000; // 1593 :  16 - 0x10
      12'h63A: dout  = 8'b00010000; // 1594 :  16 - 0x10
      12'h63B: dout  = 8'b00111000; // 1595 :  56 - 0x38
      12'h63C: dout  = 8'b00111000; // 1596 :  56 - 0x38
      12'h63D: dout  = 8'b00111000; // 1597 :  56 - 0x38
      12'h63E: dout  = 8'b00111000; // 1598 :  56 - 0x38
      12'h63F: dout  = 8'b00111000; // 1599 :  56 - 0x38
      12'h640: dout  = 8'b00111100; // 1600 :  60 - 0x3c -- Sprite 0x64
      12'h641: dout  = 8'b01111110; // 1601 : 126 - 0x7e
      12'h642: dout  = 8'b01110111; // 1602 : 119 - 0x77
      12'h643: dout  = 8'b11111011; // 1603 : 251 - 0xfb
      12'h644: dout  = 8'b10011111; // 1604 : 159 - 0x9f
      12'h645: dout  = 8'b01011111; // 1605 :  95 - 0x5f
      12'h646: dout  = 8'b10001110; // 1606 : 142 - 0x8e
      12'h647: dout  = 8'b00100000; // 1607 :  32 - 0x20
      12'h648: dout  = 8'b00000000; // 1608 :   0 - 0x0 -- plane 1
      12'h649: dout  = 8'b00011000; // 1609 :  24 - 0x18
      12'h64A: dout  = 8'b00111100; // 1610 :  60 - 0x3c
      12'h64B: dout  = 8'b00001110; // 1611 :  14 - 0xe
      12'h64C: dout  = 8'b00001110; // 1612 :  14 - 0xe
      12'h64D: dout  = 8'b00000100; // 1613 :   4 - 0x4
      12'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout  = 8'b01011100; // 1616 :  92 - 0x5c -- Sprite 0x65
      12'h651: dout  = 8'b00101110; // 1617 :  46 - 0x2e
      12'h652: dout  = 8'b10001111; // 1618 : 143 - 0x8f
      12'h653: dout  = 8'b00111111; // 1619 :  63 - 0x3f
      12'h654: dout  = 8'b01111011; // 1620 : 123 - 0x7b
      12'h655: dout  = 8'b01110111; // 1621 : 119 - 0x77
      12'h656: dout  = 8'b01111110; // 1622 : 126 - 0x7e
      12'h657: dout  = 8'b00111100; // 1623 :  60 - 0x3c
      12'h658: dout  = 8'b00000000; // 1624 :   0 - 0x0 -- plane 1
      12'h659: dout  = 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout  = 8'b00000100; // 1626 :   4 - 0x4
      12'h65B: dout  = 8'b00000110; // 1627 :   6 - 0x6
      12'h65C: dout  = 8'b00011110; // 1628 :  30 - 0x1e
      12'h65D: dout  = 8'b00111100; // 1629 :  60 - 0x3c
      12'h65E: dout  = 8'b00011000; // 1630 :  24 - 0x18
      12'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout  = 8'b00010011; // 1632 :  19 - 0x13 -- Sprite 0x66
      12'h661: dout  = 8'b01001111; // 1633 :  79 - 0x4f
      12'h662: dout  = 8'b00111111; // 1634 :  63 - 0x3f
      12'h663: dout  = 8'b10111111; // 1635 : 191 - 0xbf
      12'h664: dout  = 8'b00111111; // 1636 :  63 - 0x3f
      12'h665: dout  = 8'b01111010; // 1637 : 122 - 0x7a
      12'h666: dout  = 8'b11111000; // 1638 : 248 - 0xf8
      12'h667: dout  = 8'b11111000; // 1639 : 248 - 0xf8
      12'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0 -- plane 1
      12'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout  = 8'b00000001; // 1642 :   1 - 0x1
      12'h66B: dout  = 8'b00001010; // 1643 :  10 - 0xa
      12'h66C: dout  = 8'b00010111; // 1644 :  23 - 0x17
      12'h66D: dout  = 8'b00001111; // 1645 :  15 - 0xf
      12'h66E: dout  = 8'b00101111; // 1646 :  47 - 0x2f
      12'h66F: dout  = 8'b00011111; // 1647 :  31 - 0x1f
      12'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0x67
      12'h671: dout  = 8'b00001000; // 1649 :   8 - 0x8
      12'h672: dout  = 8'b00000101; // 1650 :   5 - 0x5
      12'h673: dout  = 8'b00001111; // 1651 :  15 - 0xf
      12'h674: dout  = 8'b00101111; // 1652 :  47 - 0x2f
      12'h675: dout  = 8'b00011101; // 1653 :  29 - 0x1d
      12'h676: dout  = 8'b00011100; // 1654 :  28 - 0x1c
      12'h677: dout  = 8'b00111100; // 1655 :  60 - 0x3c
      12'h678: dout  = 8'b00000000; // 1656 :   0 - 0x0 -- plane 1
      12'h679: dout  = 8'b00000000; // 1657 :   0 - 0x0
      12'h67A: dout  = 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout  = 8'b00000101; // 1660 :   5 - 0x5
      12'h67D: dout  = 8'b00000111; // 1661 :   7 - 0x7
      12'h67E: dout  = 8'b00001111; // 1662 :  15 - 0xf
      12'h67F: dout  = 8'b00000111; // 1663 :   7 - 0x7
      12'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0x68
      12'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout  = 8'b00000000; // 1666 :   0 - 0x0
      12'h683: dout  = 8'b00000000; // 1667 :   0 - 0x0
      12'h684: dout  = 8'b00000010; // 1668 :   2 - 0x2
      12'h685: dout  = 8'b00001011; // 1669 :  11 - 0xb
      12'h686: dout  = 8'b00000111; // 1670 :   7 - 0x7
      12'h687: dout  = 8'b00001111; // 1671 :  15 - 0xf
      12'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0 -- plane 1
      12'h689: dout  = 8'b00000000; // 1673 :   0 - 0x0
      12'h68A: dout  = 8'b00000000; // 1674 :   0 - 0x0
      12'h68B: dout  = 8'b00000000; // 1675 :   0 - 0x0
      12'h68C: dout  = 8'b00000000; // 1676 :   0 - 0x0
      12'h68D: dout  = 8'b00000000; // 1677 :   0 - 0x0
      12'h68E: dout  = 8'b00000001; // 1678 :   1 - 0x1
      12'h68F: dout  = 8'b00000011; // 1679 :   3 - 0x3
      12'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0x69
      12'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      12'h692: dout  = 8'b00000000; // 1682 :   0 - 0x0
      12'h693: dout  = 8'b00000000; // 1683 :   0 - 0x0
      12'h694: dout  = 8'b00000000; // 1684 :   0 - 0x0
      12'h695: dout  = 8'b00001000; // 1685 :   8 - 0x8
      12'h696: dout  = 8'b00000100; // 1686 :   4 - 0x4
      12'h697: dout  = 8'b00000100; // 1687 :   4 - 0x4
      12'h698: dout  = 8'b00000000; // 1688 :   0 - 0x0 -- plane 1
      12'h699: dout  = 8'b01100000; // 1689 :  96 - 0x60
      12'h69A: dout  = 8'b11110000; // 1690 : 240 - 0xf0
      12'h69B: dout  = 8'b11111000; // 1691 : 248 - 0xf8
      12'h69C: dout  = 8'b01111100; // 1692 : 124 - 0x7c
      12'h69D: dout  = 8'b00111110; // 1693 :  62 - 0x3e
      12'h69E: dout  = 8'b01111110; // 1694 : 126 - 0x7e
      12'h69F: dout  = 8'b01111111; // 1695 : 127 - 0x7f
      12'h6A0: dout  = 8'b00000010; // 1696 :   2 - 0x2 -- Sprite 0x6a
      12'h6A1: dout  = 8'b00000010; // 1697 :   2 - 0x2
      12'h6A2: dout  = 8'b00000010; // 1698 :   2 - 0x2
      12'h6A3: dout  = 8'b00000101; // 1699 :   5 - 0x5
      12'h6A4: dout  = 8'b01110001; // 1700 : 113 - 0x71
      12'h6A5: dout  = 8'b01111111; // 1701 : 127 - 0x7f
      12'h6A6: dout  = 8'b01111111; // 1702 : 127 - 0x7f
      12'h6A7: dout  = 8'b01111111; // 1703 : 127 - 0x7f
      12'h6A8: dout  = 8'b00111111; // 1704 :  63 - 0x3f -- plane 1
      12'h6A9: dout  = 8'b01011111; // 1705 :  95 - 0x5f
      12'h6AA: dout  = 8'b01111111; // 1706 : 127 - 0x7f
      12'h6AB: dout  = 8'b00111110; // 1707 :  62 - 0x3e
      12'h6AC: dout  = 8'b00001110; // 1708 :  14 - 0xe
      12'h6AD: dout  = 8'b00001010; // 1709 :  10 - 0xa
      12'h6AE: dout  = 8'b01010001; // 1710 :  81 - 0x51
      12'h6AF: dout  = 8'b00100000; // 1711 :  32 - 0x20
      12'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0x6b
      12'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      12'h6B3: dout  = 8'b00000000; // 1715 :   0 - 0x0
      12'h6B4: dout  = 8'b00000000; // 1716 :   0 - 0x0
      12'h6B5: dout  = 8'b00000000; // 1717 :   0 - 0x0
      12'h6B6: dout  = 8'b00000000; // 1718 :   0 - 0x0
      12'h6B7: dout  = 8'b00000100; // 1719 :   4 - 0x4
      12'h6B8: dout  = 8'b00000000; // 1720 :   0 - 0x0 -- plane 1
      12'h6B9: dout  = 8'b00000000; // 1721 :   0 - 0x0
      12'h6BA: dout  = 8'b00000000; // 1722 :   0 - 0x0
      12'h6BB: dout  = 8'b00000000; // 1723 :   0 - 0x0
      12'h6BC: dout  = 8'b00000000; // 1724 :   0 - 0x0
      12'h6BD: dout  = 8'b00000000; // 1725 :   0 - 0x0
      12'h6BE: dout  = 8'b00001110; // 1726 :  14 - 0xe
      12'h6BF: dout  = 8'b00011111; // 1727 :  31 - 0x1f
      12'h6C0: dout  = 8'b00000010; // 1728 :   2 - 0x2 -- Sprite 0x6c
      12'h6C1: dout  = 8'b00000010; // 1729 :   2 - 0x2
      12'h6C2: dout  = 8'b00000000; // 1730 :   0 - 0x0
      12'h6C3: dout  = 8'b00000001; // 1731 :   1 - 0x1
      12'h6C4: dout  = 8'b00010011; // 1732 :  19 - 0x13
      12'h6C5: dout  = 8'b00111111; // 1733 :  63 - 0x3f
      12'h6C6: dout  = 8'b01111111; // 1734 : 127 - 0x7f
      12'h6C7: dout  = 8'b01111111; // 1735 : 127 - 0x7f
      12'h6C8: dout  = 8'b00111111; // 1736 :  63 - 0x3f -- plane 1
      12'h6C9: dout  = 8'b01111111; // 1737 : 127 - 0x7f
      12'h6CA: dout  = 8'b01111111; // 1738 : 127 - 0x7f
      12'h6CB: dout  = 8'b11111110; // 1739 : 254 - 0xfe
      12'h6CC: dout  = 8'b11101100; // 1740 : 236 - 0xec
      12'h6CD: dout  = 8'b11001010; // 1741 : 202 - 0xca
      12'h6CE: dout  = 8'b01010001; // 1742 :  81 - 0x51
      12'h6CF: dout  = 8'b00100000; // 1743 :  32 - 0x20
      12'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0x6d
      12'h6D1: dout  = 8'b01000000; // 1745 :  64 - 0x40
      12'h6D2: dout  = 8'b01100000; // 1746 :  96 - 0x60
      12'h6D3: dout  = 8'b01110000; // 1747 : 112 - 0x70
      12'h6D4: dout  = 8'b01110011; // 1748 : 115 - 0x73
      12'h6D5: dout  = 8'b00100111; // 1749 :  39 - 0x27
      12'h6D6: dout  = 8'b00001111; // 1750 :  15 - 0xf
      12'h6D7: dout  = 8'b00011111; // 1751 :  31 - 0x1f
      12'h6D8: dout  = 8'b00000000; // 1752 :   0 - 0x0 -- plane 1
      12'h6D9: dout  = 8'b01000000; // 1753 :  64 - 0x40
      12'h6DA: dout  = 8'b01100011; // 1754 :  99 - 0x63
      12'h6DB: dout  = 8'b01110111; // 1755 : 119 - 0x77
      12'h6DC: dout  = 8'b01111100; // 1756 : 124 - 0x7c
      12'h6DD: dout  = 8'b00111000; // 1757 :  56 - 0x38
      12'h6DE: dout  = 8'b11111000; // 1758 : 248 - 0xf8
      12'h6DF: dout  = 8'b11100100; // 1759 : 228 - 0xe4
      12'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0x6e
      12'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout  = 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout  = 8'b00000011; // 1764 :   3 - 0x3
      12'h6E5: dout  = 8'b00000111; // 1765 :   7 - 0x7
      12'h6E6: dout  = 8'b00001111; // 1766 :  15 - 0xf
      12'h6E7: dout  = 8'b00011111; // 1767 :  31 - 0x1f
      12'h6E8: dout  = 8'b00000000; // 1768 :   0 - 0x0 -- plane 1
      12'h6E9: dout  = 8'b00000000; // 1769 :   0 - 0x0
      12'h6EA: dout  = 8'b00000011; // 1770 :   3 - 0x3
      12'h6EB: dout  = 8'b00000111; // 1771 :   7 - 0x7
      12'h6EC: dout  = 8'b00001100; // 1772 :  12 - 0xc
      12'h6ED: dout  = 8'b00011000; // 1773 :  24 - 0x18
      12'h6EE: dout  = 8'b11111000; // 1774 : 248 - 0xf8
      12'h6EF: dout  = 8'b11100100; // 1775 : 228 - 0xe4
      12'h6F0: dout  = 8'b01111111; // 1776 : 127 - 0x7f -- Sprite 0x6f
      12'h6F1: dout  = 8'b01111111; // 1777 : 127 - 0x7f
      12'h6F2: dout  = 8'b00111111; // 1778 :  63 - 0x3f
      12'h6F3: dout  = 8'b00111111; // 1779 :  63 - 0x3f
      12'h6F4: dout  = 8'b00011111; // 1780 :  31 - 0x1f
      12'h6F5: dout  = 8'b00011111; // 1781 :  31 - 0x1f
      12'h6F6: dout  = 8'b00001111; // 1782 :  15 - 0xf
      12'h6F7: dout  = 8'b00000111; // 1783 :   7 - 0x7
      12'h6F8: dout  = 8'b00000011; // 1784 :   3 - 0x3 -- plane 1
      12'h6F9: dout  = 8'b01000100; // 1785 :  68 - 0x44
      12'h6FA: dout  = 8'b00101000; // 1786 :  40 - 0x28
      12'h6FB: dout  = 8'b00010000; // 1787 :  16 - 0x10
      12'h6FC: dout  = 8'b00001000; // 1788 :   8 - 0x8
      12'h6FD: dout  = 8'b00000100; // 1789 :   4 - 0x4
      12'h6FE: dout  = 8'b00000011; // 1790 :   3 - 0x3
      12'h6FF: dout  = 8'b00000100; // 1791 :   4 - 0x4
      12'h700: dout  = 8'b00000011; // 1792 :   3 - 0x3 -- Sprite 0x70
      12'h701: dout  = 8'b00000111; // 1793 :   7 - 0x7
      12'h702: dout  = 8'b00001111; // 1794 :  15 - 0xf
      12'h703: dout  = 8'b00011111; // 1795 :  31 - 0x1f
      12'h704: dout  = 8'b00111111; // 1796 :  63 - 0x3f
      12'h705: dout  = 8'b01110111; // 1797 : 119 - 0x77
      12'h706: dout  = 8'b01110111; // 1798 : 119 - 0x77
      12'h707: dout  = 8'b11110101; // 1799 : 245 - 0xf5
      12'h708: dout  = 8'b00000011; // 1800 :   3 - 0x3 -- plane 1
      12'h709: dout  = 8'b00000111; // 1801 :   7 - 0x7
      12'h70A: dout  = 8'b00001111; // 1802 :  15 - 0xf
      12'h70B: dout  = 8'b00011111; // 1803 :  31 - 0x1f
      12'h70C: dout  = 8'b00100111; // 1804 :  39 - 0x27
      12'h70D: dout  = 8'b01111011; // 1805 : 123 - 0x7b
      12'h70E: dout  = 8'b01111000; // 1806 : 120 - 0x78
      12'h70F: dout  = 8'b11111011; // 1807 : 251 - 0xfb
      12'h710: dout  = 8'b11000000; // 1808 : 192 - 0xc0 -- Sprite 0x71
      12'h711: dout  = 8'b11100000; // 1809 : 224 - 0xe0
      12'h712: dout  = 8'b11110000; // 1810 : 240 - 0xf0
      12'h713: dout  = 8'b11111000; // 1811 : 248 - 0xf8
      12'h714: dout  = 8'b11111100; // 1812 : 252 - 0xfc
      12'h715: dout  = 8'b11101110; // 1813 : 238 - 0xee
      12'h716: dout  = 8'b11101110; // 1814 : 238 - 0xee
      12'h717: dout  = 8'b10101111; // 1815 : 175 - 0xaf
      12'h718: dout  = 8'b11000000; // 1816 : 192 - 0xc0 -- plane 1
      12'h719: dout  = 8'b11100000; // 1817 : 224 - 0xe0
      12'h71A: dout  = 8'b11110000; // 1818 : 240 - 0xf0
      12'h71B: dout  = 8'b11111000; // 1819 : 248 - 0xf8
      12'h71C: dout  = 8'b11100100; // 1820 : 228 - 0xe4
      12'h71D: dout  = 8'b11011110; // 1821 : 222 - 0xde
      12'h71E: dout  = 8'b00011110; // 1822 :  30 - 0x1e
      12'h71F: dout  = 8'b11011111; // 1823 : 223 - 0xdf
      12'h720: dout  = 8'b11110001; // 1824 : 241 - 0xf1 -- Sprite 0x72
      12'h721: dout  = 8'b11111111; // 1825 : 255 - 0xff
      12'h722: dout  = 8'b01111000; // 1826 : 120 - 0x78
      12'h723: dout  = 8'b00000000; // 1827 :   0 - 0x0
      12'h724: dout  = 8'b00000000; // 1828 :   0 - 0x0
      12'h725: dout  = 8'b00011000; // 1829 :  24 - 0x18
      12'h726: dout  = 8'b00011100; // 1830 :  28 - 0x1c
      12'h727: dout  = 8'b00001110; // 1831 :  14 - 0xe
      12'h728: dout  = 8'b11111111; // 1832 : 255 - 0xff -- plane 1
      12'h729: dout  = 8'b11111111; // 1833 : 255 - 0xff
      12'h72A: dout  = 8'b01111111; // 1834 : 127 - 0x7f
      12'h72B: dout  = 8'b00001111; // 1835 :  15 - 0xf
      12'h72C: dout  = 8'b00001111; // 1836 :  15 - 0xf
      12'h72D: dout  = 8'b00000111; // 1837 :   7 - 0x7
      12'h72E: dout  = 8'b00000011; // 1838 :   3 - 0x3
      12'h72F: dout  = 8'b00000000; // 1839 :   0 - 0x0
      12'h730: dout  = 8'b10001111; // 1840 : 143 - 0x8f -- Sprite 0x73
      12'h731: dout  = 8'b11111111; // 1841 : 255 - 0xff
      12'h732: dout  = 8'b00011110; // 1842 :  30 - 0x1e
      12'h733: dout  = 8'b00000000; // 1843 :   0 - 0x0
      12'h734: dout  = 8'b00001100; // 1844 :  12 - 0xc
      12'h735: dout  = 8'b00111110; // 1845 :  62 - 0x3e
      12'h736: dout  = 8'b01111110; // 1846 : 126 - 0x7e
      12'h737: dout  = 8'b01111100; // 1847 : 124 - 0x7c
      12'h738: dout  = 8'b11111111; // 1848 : 255 - 0xff -- plane 1
      12'h739: dout  = 8'b11111111; // 1849 : 255 - 0xff
      12'h73A: dout  = 8'b11111110; // 1850 : 254 - 0xfe
      12'h73B: dout  = 8'b11110000; // 1851 : 240 - 0xf0
      12'h73C: dout  = 8'b11110000; // 1852 : 240 - 0xf0
      12'h73D: dout  = 8'b11000000; // 1853 : 192 - 0xc0
      12'h73E: dout  = 8'b10000000; // 1854 : 128 - 0x80
      12'h73F: dout  = 8'b00000000; // 1855 :   0 - 0x0
      12'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0x74
      12'h741: dout  = 8'b00000000; // 1857 :   0 - 0x0
      12'h742: dout  = 8'b00000000; // 1858 :   0 - 0x0
      12'h743: dout  = 8'b00000000; // 1859 :   0 - 0x0
      12'h744: dout  = 8'b00000000; // 1860 :   0 - 0x0
      12'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      12'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      12'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      12'h748: dout  = 8'b00000000; // 1864 :   0 - 0x0 -- plane 1
      12'h749: dout  = 8'b00000000; // 1865 :   0 - 0x0
      12'h74A: dout  = 8'b00011000; // 1866 :  24 - 0x18
      12'h74B: dout  = 8'b00100100; // 1867 :  36 - 0x24
      12'h74C: dout  = 8'b00100100; // 1868 :  36 - 0x24
      12'h74D: dout  = 8'b00011000; // 1869 :  24 - 0x18
      12'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      12'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout  = 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0x75
      12'h751: dout  = 8'b00000010; // 1873 :   2 - 0x2
      12'h752: dout  = 8'b01000001; // 1874 :  65 - 0x41
      12'h753: dout  = 8'b01000001; // 1875 :  65 - 0x41
      12'h754: dout  = 8'b01100001; // 1876 :  97 - 0x61
      12'h755: dout  = 8'b00110011; // 1877 :  51 - 0x33
      12'h756: dout  = 8'b00000110; // 1878 :   6 - 0x6
      12'h757: dout  = 8'b00111100; // 1879 :  60 - 0x3c
      12'h758: dout  = 8'b00111100; // 1880 :  60 - 0x3c -- plane 1
      12'h759: dout  = 8'b01111110; // 1881 : 126 - 0x7e
      12'h75A: dout  = 8'b11111111; // 1882 : 255 - 0xff
      12'h75B: dout  = 8'b11111111; // 1883 : 255 - 0xff
      12'h75C: dout  = 8'b11111111; // 1884 : 255 - 0xff
      12'h75D: dout  = 8'b11111111; // 1885 : 255 - 0xff
      12'h75E: dout  = 8'b01111110; // 1886 : 126 - 0x7e
      12'h75F: dout  = 8'b00111100; // 1887 :  60 - 0x3c
      12'h760: dout  = 8'b00000011; // 1888 :   3 - 0x3 -- Sprite 0x76
      12'h761: dout  = 8'b00000111; // 1889 :   7 - 0x7
      12'h762: dout  = 8'b00001111; // 1890 :  15 - 0xf
      12'h763: dout  = 8'b00011111; // 1891 :  31 - 0x1f
      12'h764: dout  = 8'b00111111; // 1892 :  63 - 0x3f
      12'h765: dout  = 8'b01111111; // 1893 : 127 - 0x7f
      12'h766: dout  = 8'b01111111; // 1894 : 127 - 0x7f
      12'h767: dout  = 8'b11111111; // 1895 : 255 - 0xff
      12'h768: dout  = 8'b00000011; // 1896 :   3 - 0x3 -- plane 1
      12'h769: dout  = 8'b00000111; // 1897 :   7 - 0x7
      12'h76A: dout  = 8'b00001111; // 1898 :  15 - 0xf
      12'h76B: dout  = 8'b00011111; // 1899 :  31 - 0x1f
      12'h76C: dout  = 8'b00111111; // 1900 :  63 - 0x3f
      12'h76D: dout  = 8'b01100011; // 1901 :  99 - 0x63
      12'h76E: dout  = 8'b01000001; // 1902 :  65 - 0x41
      12'h76F: dout  = 8'b11000001; // 1903 : 193 - 0xc1
      12'h770: dout  = 8'b11000000; // 1904 : 192 - 0xc0 -- Sprite 0x77
      12'h771: dout  = 8'b11100000; // 1905 : 224 - 0xe0
      12'h772: dout  = 8'b11110000; // 1906 : 240 - 0xf0
      12'h773: dout  = 8'b11111000; // 1907 : 248 - 0xf8
      12'h774: dout  = 8'b11111100; // 1908 : 252 - 0xfc
      12'h775: dout  = 8'b11111110; // 1909 : 254 - 0xfe
      12'h776: dout  = 8'b11111110; // 1910 : 254 - 0xfe
      12'h777: dout  = 8'b11111111; // 1911 : 255 - 0xff
      12'h778: dout  = 8'b11000000; // 1912 : 192 - 0xc0 -- plane 1
      12'h779: dout  = 8'b10000000; // 1913 : 128 - 0x80
      12'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      12'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      12'h77C: dout  = 8'b10001100; // 1916 : 140 - 0x8c
      12'h77D: dout  = 8'b11111110; // 1917 : 254 - 0xfe
      12'h77E: dout  = 8'b11111110; // 1918 : 254 - 0xfe
      12'h77F: dout  = 8'b11110011; // 1919 : 243 - 0xf3
      12'h780: dout  = 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0x78
      12'h781: dout  = 8'b11111111; // 1921 : 255 - 0xff
      12'h782: dout  = 8'b11111111; // 1922 : 255 - 0xff
      12'h783: dout  = 8'b01111000; // 1923 : 120 - 0x78
      12'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout  = 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout  = 8'b11000001; // 1928 : 193 - 0xc1 -- plane 1
      12'h789: dout  = 8'b11100011; // 1929 : 227 - 0xe3
      12'h78A: dout  = 8'b11111111; // 1930 : 255 - 0xff
      12'h78B: dout  = 8'b01000111; // 1931 :  71 - 0x47
      12'h78C: dout  = 8'b00001111; // 1932 :  15 - 0xf
      12'h78D: dout  = 8'b00001111; // 1933 :  15 - 0xf
      12'h78E: dout  = 8'b00001111; // 1934 :  15 - 0xf
      12'h78F: dout  = 8'b00000111; // 1935 :   7 - 0x7
      12'h790: dout  = 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0x79
      12'h791: dout  = 8'b11111111; // 1937 : 255 - 0xff
      12'h792: dout  = 8'b11111111; // 1938 : 255 - 0xff
      12'h793: dout  = 8'b00011110; // 1939 :  30 - 0x1e
      12'h794: dout  = 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout  = 8'b00100000; // 1941 :  32 - 0x20
      12'h796: dout  = 8'b00100000; // 1942 :  32 - 0x20
      12'h797: dout  = 8'b01000000; // 1943 :  64 - 0x40
      12'h798: dout  = 8'b11110001; // 1944 : 241 - 0xf1 -- plane 1
      12'h799: dout  = 8'b11111001; // 1945 : 249 - 0xf9
      12'h79A: dout  = 8'b11111111; // 1946 : 255 - 0xff
      12'h79B: dout  = 8'b11100010; // 1947 : 226 - 0xe2
      12'h79C: dout  = 8'b11110000; // 1948 : 240 - 0xf0
      12'h79D: dout  = 8'b11110000; // 1949 : 240 - 0xf0
      12'h79E: dout  = 8'b11110000; // 1950 : 240 - 0xf0
      12'h79F: dout  = 8'b11100000; // 1951 : 224 - 0xe0
      12'h7A0: dout  = 8'b00010110; // 1952 :  22 - 0x16 -- Sprite 0x7a
      12'h7A1: dout  = 8'b00011111; // 1953 :  31 - 0x1f
      12'h7A2: dout  = 8'b00111111; // 1954 :  63 - 0x3f
      12'h7A3: dout  = 8'b01111111; // 1955 : 127 - 0x7f
      12'h7A4: dout  = 8'b00111101; // 1956 :  61 - 0x3d
      12'h7A5: dout  = 8'b00011101; // 1957 :  29 - 0x1d
      12'h7A6: dout  = 8'b00111111; // 1958 :  63 - 0x3f
      12'h7A7: dout  = 8'b00011111; // 1959 :  31 - 0x1f
      12'h7A8: dout  = 8'b00010110; // 1960 :  22 - 0x16 -- plane 1
      12'h7A9: dout  = 8'b00011111; // 1961 :  31 - 0x1f
      12'h7AA: dout  = 8'b00000000; // 1962 :   0 - 0x0
      12'h7AB: dout  = 8'b00000000; // 1963 :   0 - 0x0
      12'h7AC: dout  = 8'b00000101; // 1964 :   5 - 0x5
      12'h7AD: dout  = 8'b00001101; // 1965 :  13 - 0xd
      12'h7AE: dout  = 8'b00111111; // 1966 :  63 - 0x3f
      12'h7AF: dout  = 8'b00011111; // 1967 :  31 - 0x1f
      12'h7B0: dout  = 8'b10000000; // 1968 : 128 - 0x80 -- Sprite 0x7b
      12'h7B1: dout  = 8'b10000000; // 1969 : 128 - 0x80
      12'h7B2: dout  = 8'b11000000; // 1970 : 192 - 0xc0
      12'h7B3: dout  = 8'b11100000; // 1971 : 224 - 0xe0
      12'h7B4: dout  = 8'b11110000; // 1972 : 240 - 0xf0
      12'h7B5: dout  = 8'b11110000; // 1973 : 240 - 0xf0
      12'h7B6: dout  = 8'b11110000; // 1974 : 240 - 0xf0
      12'h7B7: dout  = 8'b11111000; // 1975 : 248 - 0xf8
      12'h7B8: dout  = 8'b10000000; // 1976 : 128 - 0x80 -- plane 1
      12'h7B9: dout  = 8'b10000000; // 1977 : 128 - 0x80
      12'h7BA: dout  = 8'b00000000; // 1978 :   0 - 0x0
      12'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout  = 8'b10100000; // 1981 : 160 - 0xa0
      12'h7BE: dout  = 8'b10100000; // 1982 : 160 - 0xa0
      12'h7BF: dout  = 8'b11100000; // 1983 : 224 - 0xe0
      12'h7C0: dout  = 8'b00111100; // 1984 :  60 - 0x3c -- Sprite 0x7c
      12'h7C1: dout  = 8'b11111010; // 1985 : 250 - 0xfa
      12'h7C2: dout  = 8'b10110001; // 1986 : 177 - 0xb1
      12'h7C3: dout  = 8'b01110010; // 1987 : 114 - 0x72
      12'h7C4: dout  = 8'b11110010; // 1988 : 242 - 0xf2
      12'h7C5: dout  = 8'b11011011; // 1989 : 219 - 0xdb
      12'h7C6: dout  = 8'b11011111; // 1990 : 223 - 0xdf
      12'h7C7: dout  = 8'b01011111; // 1991 :  95 - 0x5f
      12'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0 -- plane 1
      12'h7C9: dout  = 8'b00000100; // 1993 :   4 - 0x4
      12'h7CA: dout  = 8'b01001110; // 1994 :  78 - 0x4e
      12'h7CB: dout  = 8'b10001100; // 1995 : 140 - 0x8c
      12'h7CC: dout  = 8'b00001100; // 1996 :  12 - 0xc
      12'h7CD: dout  = 8'b01111111; // 1997 : 127 - 0x7f
      12'h7CE: dout  = 8'b11111111; // 1998 : 255 - 0xff
      12'h7CF: dout  = 8'b11111111; // 1999 : 255 - 0xff
      12'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0x7d
      12'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      12'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      12'h7D3: dout  = 8'b00000001; // 2003 :   1 - 0x1
      12'h7D4: dout  = 8'b00000001; // 2004 :   1 - 0x1
      12'h7D5: dout  = 8'b00000001; // 2005 :   1 - 0x1
      12'h7D6: dout  = 8'b00000110; // 2006 :   6 - 0x6
      12'h7D7: dout  = 8'b00011110; // 2007 :  30 - 0x1e
      12'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0 -- plane 1
      12'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      12'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      12'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      12'h7DC: dout  = 8'b00000000; // 2012 :   0 - 0x0
      12'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      12'h7DE: dout  = 8'b00000001; // 2014 :   1 - 0x1
      12'h7DF: dout  = 8'b00000001; // 2015 :   1 - 0x1
      12'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0x7e
      12'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      12'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      12'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      12'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      12'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      12'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout  = 8'b11111111; // 2024 : 255 - 0xff -- plane 1
      12'h7E9: dout  = 8'b01111111; // 2025 : 127 - 0x7f
      12'h7EA: dout  = 8'b00111111; // 2026 :  63 - 0x3f
      12'h7EB: dout  = 8'b00011111; // 2027 :  31 - 0x1f
      12'h7EC: dout  = 8'b00001111; // 2028 :  15 - 0xf
      12'h7ED: dout  = 8'b00000111; // 2029 :   7 - 0x7
      12'h7EE: dout  = 8'b00000011; // 2030 :   3 - 0x3
      12'h7EF: dout  = 8'b00000001; // 2031 :   1 - 0x1
      12'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0x7f
      12'h7F1: dout  = 8'b01111100; // 2033 : 124 - 0x7c
      12'h7F2: dout  = 8'b11010110; // 2034 : 214 - 0xd6
      12'h7F3: dout  = 8'b10010010; // 2035 : 146 - 0x92
      12'h7F4: dout  = 8'b10111010; // 2036 : 186 - 0xba
      12'h7F5: dout  = 8'b11101110; // 2037 : 238 - 0xee
      12'h7F6: dout  = 8'b11111110; // 2038 : 254 - 0xfe
      12'h7F7: dout  = 8'b00111000; // 2039 :  56 - 0x38
      12'h7F8: dout  = 8'b11111111; // 2040 : 255 - 0xff -- plane 1
      12'h7F9: dout  = 8'b10000011; // 2041 : 131 - 0x83
      12'h7FA: dout  = 8'b00101001; // 2042 :  41 - 0x29
      12'h7FB: dout  = 8'b01101101; // 2043 : 109 - 0x6d
      12'h7FC: dout  = 8'b01000101; // 2044 :  69 - 0x45
      12'h7FD: dout  = 8'b00010001; // 2045 :  17 - 0x11
      12'h7FE: dout  = 8'b00000001; // 2046 :   1 - 0x1
      12'h7FF: dout  = 8'b11000111; // 2047 : 199 - 0xc7
      12'h800: dout  = 8'b00000000; // 2048 :   0 - 0x0 -- Sprite 0x80
      12'h801: dout  = 8'b00010101; // 2049 :  21 - 0x15
      12'h802: dout  = 8'b00111111; // 2050 :  63 - 0x3f
      12'h803: dout  = 8'b01100010; // 2051 :  98 - 0x62
      12'h804: dout  = 8'b01011111; // 2052 :  95 - 0x5f
      12'h805: dout  = 8'b11111111; // 2053 : 255 - 0xff
      12'h806: dout  = 8'b10011111; // 2054 : 159 - 0x9f
      12'h807: dout  = 8'b01111101; // 2055 : 125 - 0x7d
      12'h808: dout  = 8'b00001000; // 2056 :   8 - 0x8 -- plane 1
      12'h809: dout  = 8'b00001000; // 2057 :   8 - 0x8
      12'h80A: dout  = 8'b00000010; // 2058 :   2 - 0x2
      12'h80B: dout  = 8'b00011111; // 2059 :  31 - 0x1f
      12'h80C: dout  = 8'b00100010; // 2060 :  34 - 0x22
      12'h80D: dout  = 8'b00000010; // 2061 :   2 - 0x2
      12'h80E: dout  = 8'b00000010; // 2062 :   2 - 0x2
      12'h80F: dout  = 8'b00000000; // 2063 :   0 - 0x0
      12'h810: dout  = 8'b00000000; // 2064 :   0 - 0x0 -- Sprite 0x81
      12'h811: dout  = 8'b00000000; // 2065 :   0 - 0x0
      12'h812: dout  = 8'b00000000; // 2066 :   0 - 0x0
      12'h813: dout  = 8'b00000000; // 2067 :   0 - 0x0
      12'h814: dout  = 8'b00000000; // 2068 :   0 - 0x0
      12'h815: dout  = 8'b00000000; // 2069 :   0 - 0x0
      12'h816: dout  = 8'b00000000; // 2070 :   0 - 0x0
      12'h817: dout  = 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout  = 8'b00001000; // 2072 :   8 - 0x8 -- plane 1
      12'h819: dout  = 8'b00001000; // 2073 :   8 - 0x8
      12'h81A: dout  = 8'b00001000; // 2074 :   8 - 0x8
      12'h81B: dout  = 8'b00001000; // 2075 :   8 - 0x8
      12'h81C: dout  = 8'b00001000; // 2076 :   8 - 0x8
      12'h81D: dout  = 8'b00001000; // 2077 :   8 - 0x8
      12'h81E: dout  = 8'b00001000; // 2078 :   8 - 0x8
      12'h81F: dout  = 8'b00001000; // 2079 :   8 - 0x8
      12'h820: dout  = 8'b00101111; // 2080 :  47 - 0x2f -- Sprite 0x82
      12'h821: dout  = 8'b00011110; // 2081 :  30 - 0x1e
      12'h822: dout  = 8'b00101111; // 2082 :  47 - 0x2f
      12'h823: dout  = 8'b00101111; // 2083 :  47 - 0x2f
      12'h824: dout  = 8'b00101111; // 2084 :  47 - 0x2f
      12'h825: dout  = 8'b00010101; // 2085 :  21 - 0x15
      12'h826: dout  = 8'b00001101; // 2086 :  13 - 0xd
      12'h827: dout  = 8'b00001110; // 2087 :  14 - 0xe
      12'h828: dout  = 8'b00010000; // 2088 :  16 - 0x10 -- plane 1
      12'h829: dout  = 8'b00011110; // 2089 :  30 - 0x1e
      12'h82A: dout  = 8'b00010000; // 2090 :  16 - 0x10
      12'h82B: dout  = 8'b01010000; // 2091 :  80 - 0x50
      12'h82C: dout  = 8'b00010000; // 2092 :  16 - 0x10
      12'h82D: dout  = 8'b00001000; // 2093 :   8 - 0x8
      12'h82E: dout  = 8'b00000000; // 2094 :   0 - 0x0
      12'h82F: dout  = 8'b00000000; // 2095 :   0 - 0x0
      12'h830: dout  = 8'b00000000; // 2096 :   0 - 0x0 -- Sprite 0x83
      12'h831: dout  = 8'b00000000; // 2097 :   0 - 0x0
      12'h832: dout  = 8'b00000000; // 2098 :   0 - 0x0
      12'h833: dout  = 8'b00000000; // 2099 :   0 - 0x0
      12'h834: dout  = 8'b00000000; // 2100 :   0 - 0x0
      12'h835: dout  = 8'b00000000; // 2101 :   0 - 0x0
      12'h836: dout  = 8'b00000000; // 2102 :   0 - 0x0
      12'h837: dout  = 8'b00000000; // 2103 :   0 - 0x0
      12'h838: dout  = 8'b00000000; // 2104 :   0 - 0x0 -- plane 1
      12'h839: dout  = 8'b00000000; // 2105 :   0 - 0x0
      12'h83A: dout  = 8'b00000000; // 2106 :   0 - 0x0
      12'h83B: dout  = 8'b11111110; // 2107 : 254 - 0xfe
      12'h83C: dout  = 8'b00000000; // 2108 :   0 - 0x0
      12'h83D: dout  = 8'b00000000; // 2109 :   0 - 0x0
      12'h83E: dout  = 8'b00000000; // 2110 :   0 - 0x0
      12'h83F: dout  = 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout  = 8'b00011100; // 2112 :  28 - 0x1c -- Sprite 0x84
      12'h841: dout  = 8'b00111110; // 2113 :  62 - 0x3e
      12'h842: dout  = 8'b01111111; // 2114 : 127 - 0x7f
      12'h843: dout  = 8'b11111111; // 2115 : 255 - 0xff
      12'h844: dout  = 8'b11111111; // 2116 : 255 - 0xff
      12'h845: dout  = 8'b11111110; // 2117 : 254 - 0xfe
      12'h846: dout  = 8'b01111100; // 2118 : 124 - 0x7c
      12'h847: dout  = 8'b00111000; // 2119 :  56 - 0x38
      12'h848: dout  = 8'b00011100; // 2120 :  28 - 0x1c -- plane 1
      12'h849: dout  = 8'b00101010; // 2121 :  42 - 0x2a
      12'h84A: dout  = 8'b01110111; // 2122 : 119 - 0x77
      12'h84B: dout  = 8'b11101110; // 2123 : 238 - 0xee
      12'h84C: dout  = 8'b11011101; // 2124 : 221 - 0xdd
      12'h84D: dout  = 8'b10101010; // 2125 : 170 - 0xaa
      12'h84E: dout  = 8'b01110100; // 2126 : 116 - 0x74
      12'h84F: dout  = 8'b00101000; // 2127 :  40 - 0x28
      12'h850: dout  = 8'b00000000; // 2128 :   0 - 0x0 -- Sprite 0x85
      12'h851: dout  = 8'b11111111; // 2129 : 255 - 0xff
      12'h852: dout  = 8'b11111111; // 2130 : 255 - 0xff
      12'h853: dout  = 8'b11111111; // 2131 : 255 - 0xff
      12'h854: dout  = 8'b11111111; // 2132 : 255 - 0xff
      12'h855: dout  = 8'b11111111; // 2133 : 255 - 0xff
      12'h856: dout  = 8'b11111111; // 2134 : 255 - 0xff
      12'h857: dout  = 8'b11111111; // 2135 : 255 - 0xff
      12'h858: dout  = 8'b11111111; // 2136 : 255 - 0xff -- plane 1
      12'h859: dout  = 8'b11111110; // 2137 : 254 - 0xfe
      12'h85A: dout  = 8'b11111110; // 2138 : 254 - 0xfe
      12'h85B: dout  = 8'b00000000; // 2139 :   0 - 0x0
      12'h85C: dout  = 8'b11101111; // 2140 : 239 - 0xef
      12'h85D: dout  = 8'b11101111; // 2141 : 239 - 0xef
      12'h85E: dout  = 8'b11101111; // 2142 : 239 - 0xef
      12'h85F: dout  = 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout  = 8'b11111111; // 2144 : 255 - 0xff -- Sprite 0x86
      12'h861: dout  = 8'b11111111; // 2145 : 255 - 0xff
      12'h862: dout  = 8'b11111111; // 2146 : 255 - 0xff
      12'h863: dout  = 8'b11111111; // 2147 : 255 - 0xff
      12'h864: dout  = 8'b11111111; // 2148 : 255 - 0xff
      12'h865: dout  = 8'b11111111; // 2149 : 255 - 0xff
      12'h866: dout  = 8'b11111111; // 2150 : 255 - 0xff
      12'h867: dout  = 8'b11111111; // 2151 : 255 - 0xff
      12'h868: dout  = 8'b11111110; // 2152 : 254 - 0xfe -- plane 1
      12'h869: dout  = 8'b11111110; // 2153 : 254 - 0xfe
      12'h86A: dout  = 8'b11111110; // 2154 : 254 - 0xfe
      12'h86B: dout  = 8'b00000000; // 2155 :   0 - 0x0
      12'h86C: dout  = 8'b11101111; // 2156 : 239 - 0xef
      12'h86D: dout  = 8'b11101111; // 2157 : 239 - 0xef
      12'h86E: dout  = 8'b11101111; // 2158 : 239 - 0xef
      12'h86F: dout  = 8'b00000000; // 2159 :   0 - 0x0
      12'h870: dout  = 8'b01111111; // 2160 : 127 - 0x7f -- Sprite 0x87
      12'h871: dout  = 8'b11111111; // 2161 : 255 - 0xff
      12'h872: dout  = 8'b11111111; // 2162 : 255 - 0xff
      12'h873: dout  = 8'b11111111; // 2163 : 255 - 0xff
      12'h874: dout  = 8'b11111111; // 2164 : 255 - 0xff
      12'h875: dout  = 8'b11111111; // 2165 : 255 - 0xff
      12'h876: dout  = 8'b11111111; // 2166 : 255 - 0xff
      12'h877: dout  = 8'b11111111; // 2167 : 255 - 0xff
      12'h878: dout  = 8'b00000000; // 2168 :   0 - 0x0 -- plane 1
      12'h879: dout  = 8'b01111111; // 2169 : 127 - 0x7f
      12'h87A: dout  = 8'b01011111; // 2170 :  95 - 0x5f
      12'h87B: dout  = 8'b01111111; // 2171 : 127 - 0x7f
      12'h87C: dout  = 8'b01111111; // 2172 : 127 - 0x7f
      12'h87D: dout  = 8'b01111111; // 2173 : 127 - 0x7f
      12'h87E: dout  = 8'b01111111; // 2174 : 127 - 0x7f
      12'h87F: dout  = 8'b01111111; // 2175 : 127 - 0x7f
      12'h880: dout  = 8'b01101000; // 2176 : 104 - 0x68 -- Sprite 0x88
      12'h881: dout  = 8'b01001110; // 2177 :  78 - 0x4e
      12'h882: dout  = 8'b11100000; // 2178 : 224 - 0xe0
      12'h883: dout  = 8'b11100000; // 2179 : 224 - 0xe0
      12'h884: dout  = 8'b11100000; // 2180 : 224 - 0xe0
      12'h885: dout  = 8'b11110000; // 2181 : 240 - 0xf0
      12'h886: dout  = 8'b11111000; // 2182 : 248 - 0xf8
      12'h887: dout  = 8'b11111100; // 2183 : 252 - 0xfc
      12'h888: dout  = 8'b10111000; // 2184 : 184 - 0xb8 -- plane 1
      12'h889: dout  = 8'b10011110; // 2185 : 158 - 0x9e
      12'h88A: dout  = 8'b10000000; // 2186 : 128 - 0x80
      12'h88B: dout  = 8'b11000000; // 2187 : 192 - 0xc0
      12'h88C: dout  = 8'b11100000; // 2188 : 224 - 0xe0
      12'h88D: dout  = 8'b11110000; // 2189 : 240 - 0xf0
      12'h88E: dout  = 8'b11111000; // 2190 : 248 - 0xf8
      12'h88F: dout  = 8'b01111100; // 2191 : 124 - 0x7c
      12'h890: dout  = 8'b00111111; // 2192 :  63 - 0x3f -- Sprite 0x89
      12'h891: dout  = 8'b01011100; // 2193 :  92 - 0x5c
      12'h892: dout  = 8'b00111001; // 2194 :  57 - 0x39
      12'h893: dout  = 8'b00111011; // 2195 :  59 - 0x3b
      12'h894: dout  = 8'b10111011; // 2196 : 187 - 0xbb
      12'h895: dout  = 8'b11111001; // 2197 : 249 - 0xf9
      12'h896: dout  = 8'b11111100; // 2198 : 252 - 0xfc
      12'h897: dout  = 8'b11111110; // 2199 : 254 - 0xfe
      12'h898: dout  = 8'b00000000; // 2200 :   0 - 0x0 -- plane 1
      12'h899: dout  = 8'b00100011; // 2201 :  35 - 0x23
      12'h89A: dout  = 8'b01010111; // 2202 :  87 - 0x57
      12'h89B: dout  = 8'b01001111; // 2203 :  79 - 0x4f
      12'h89C: dout  = 8'b01010111; // 2204 :  87 - 0x57
      12'h89D: dout  = 8'b00100111; // 2205 :  39 - 0x27
      12'h89E: dout  = 8'b11000011; // 2206 : 195 - 0xc3
      12'h89F: dout  = 8'b00100001; // 2207 :  33 - 0x21
      12'h8A0: dout  = 8'b11000000; // 2208 : 192 - 0xc0 -- Sprite 0x8a
      12'h8A1: dout  = 8'b11110000; // 2209 : 240 - 0xf0
      12'h8A2: dout  = 8'b11110000; // 2210 : 240 - 0xf0
      12'h8A3: dout  = 8'b11110000; // 2211 : 240 - 0xf0
      12'h8A4: dout  = 8'b11110000; // 2212 : 240 - 0xf0
      12'h8A5: dout  = 8'b11100000; // 2213 : 224 - 0xe0
      12'h8A6: dout  = 8'b11000000; // 2214 : 192 - 0xc0
      12'h8A7: dout  = 8'b00000000; // 2215 :   0 - 0x0
      12'h8A8: dout  = 8'b00000000; // 2216 :   0 - 0x0 -- plane 1
      12'h8A9: dout  = 8'b00110000; // 2217 :  48 - 0x30
      12'h8AA: dout  = 8'b01110000; // 2218 : 112 - 0x70
      12'h8AB: dout  = 8'b01110000; // 2219 : 112 - 0x70
      12'h8AC: dout  = 8'b11110000; // 2220 : 240 - 0xf0
      12'h8AD: dout  = 8'b11100000; // 2221 : 224 - 0xe0
      12'h8AE: dout  = 8'b11000000; // 2222 : 192 - 0xc0
      12'h8AF: dout  = 8'b00000000; // 2223 :   0 - 0x0
      12'h8B0: dout  = 8'b11111110; // 2224 : 254 - 0xfe -- Sprite 0x8b
      12'h8B1: dout  = 8'b11111100; // 2225 : 252 - 0xfc
      12'h8B2: dout  = 8'b01100001; // 2226 :  97 - 0x61
      12'h8B3: dout  = 8'b00001111; // 2227 :  15 - 0xf
      12'h8B4: dout  = 8'b11111111; // 2228 : 255 - 0xff
      12'h8B5: dout  = 8'b11111110; // 2229 : 254 - 0xfe
      12'h8B6: dout  = 8'b11110000; // 2230 : 240 - 0xf0
      12'h8B7: dout  = 8'b11100000; // 2231 : 224 - 0xe0
      12'h8B8: dout  = 8'b00010011; // 2232 :  19 - 0x13 -- plane 1
      12'h8B9: dout  = 8'b00001111; // 2233 :  15 - 0xf
      12'h8BA: dout  = 8'b00011110; // 2234 :  30 - 0x1e
      12'h8BB: dout  = 8'b11110000; // 2235 : 240 - 0xf0
      12'h8BC: dout  = 8'b11111100; // 2236 : 252 - 0xfc
      12'h8BD: dout  = 8'b11111000; // 2237 : 248 - 0xf8
      12'h8BE: dout  = 8'b11110000; // 2238 : 240 - 0xf0
      12'h8BF: dout  = 8'b11100000; // 2239 : 224 - 0xe0
      12'h8C0: dout  = 8'b01101110; // 2240 : 110 - 0x6e -- Sprite 0x8c
      12'h8C1: dout  = 8'b01000000; // 2241 :  64 - 0x40
      12'h8C2: dout  = 8'b11100000; // 2242 : 224 - 0xe0
      12'h8C3: dout  = 8'b11100000; // 2243 : 224 - 0xe0
      12'h8C4: dout  = 8'b11100000; // 2244 : 224 - 0xe0
      12'h8C5: dout  = 8'b11100000; // 2245 : 224 - 0xe0
      12'h8C6: dout  = 8'b11100000; // 2246 : 224 - 0xe0
      12'h8C7: dout  = 8'b11000000; // 2247 : 192 - 0xc0
      12'h8C8: dout  = 8'b10111110; // 2248 : 190 - 0xbe -- plane 1
      12'h8C9: dout  = 8'b10010000; // 2249 : 144 - 0x90
      12'h8CA: dout  = 8'b10000000; // 2250 : 128 - 0x80
      12'h8CB: dout  = 8'b11000000; // 2251 : 192 - 0xc0
      12'h8CC: dout  = 8'b11000000; // 2252 : 192 - 0xc0
      12'h8CD: dout  = 8'b10000000; // 2253 : 128 - 0x80
      12'h8CE: dout  = 8'b00000000; // 2254 :   0 - 0x0
      12'h8CF: dout  = 8'b00000000; // 2255 :   0 - 0x0
      12'h8D0: dout  = 8'b00000001; // 2256 :   1 - 0x1 -- Sprite 0x8d
      12'h8D1: dout  = 8'b00000001; // 2257 :   1 - 0x1
      12'h8D2: dout  = 8'b00000011; // 2258 :   3 - 0x3
      12'h8D3: dout  = 8'b00000011; // 2259 :   3 - 0x3
      12'h8D4: dout  = 8'b00000111; // 2260 :   7 - 0x7
      12'h8D5: dout  = 8'b01111111; // 2261 : 127 - 0x7f
      12'h8D6: dout  = 8'b01111111; // 2262 : 127 - 0x7f
      12'h8D7: dout  = 8'b00111111; // 2263 :  63 - 0x3f
      12'h8D8: dout  = 8'b00000001; // 2264 :   1 - 0x1 -- plane 1
      12'h8D9: dout  = 8'b00000001; // 2265 :   1 - 0x1
      12'h8DA: dout  = 8'b00000011; // 2266 :   3 - 0x3
      12'h8DB: dout  = 8'b00000011; // 2267 :   3 - 0x3
      12'h8DC: dout  = 8'b00000111; // 2268 :   7 - 0x7
      12'h8DD: dout  = 8'b01111111; // 2269 : 127 - 0x7f
      12'h8DE: dout  = 8'b01111101; // 2270 : 125 - 0x7d
      12'h8DF: dout  = 8'b00111101; // 2271 :  61 - 0x3d
      12'h8E0: dout  = 8'b00000110; // 2272 :   6 - 0x6 -- Sprite 0x8e
      12'h8E1: dout  = 8'b00000111; // 2273 :   7 - 0x7
      12'h8E2: dout  = 8'b00111111; // 2274 :  63 - 0x3f
      12'h8E3: dout  = 8'b00111100; // 2275 :  60 - 0x3c
      12'h8E4: dout  = 8'b00011001; // 2276 :  25 - 0x19
      12'h8E5: dout  = 8'b01111011; // 2277 : 123 - 0x7b
      12'h8E6: dout  = 8'b01111111; // 2278 : 127 - 0x7f
      12'h8E7: dout  = 8'b00111111; // 2279 :  63 - 0x3f
      12'h8E8: dout  = 8'b00000110; // 2280 :   6 - 0x6 -- plane 1
      12'h8E9: dout  = 8'b00000100; // 2281 :   4 - 0x4
      12'h8EA: dout  = 8'b00110000; // 2282 :  48 - 0x30
      12'h8EB: dout  = 8'b00100011; // 2283 :  35 - 0x23
      12'h8EC: dout  = 8'b00000110; // 2284 :   6 - 0x6
      12'h8ED: dout  = 8'b01100100; // 2285 : 100 - 0x64
      12'h8EE: dout  = 8'b01100000; // 2286 :  96 - 0x60
      12'h8EF: dout  = 8'b00000000; // 2287 :   0 - 0x0
      12'h8F0: dout  = 8'b00111111; // 2288 :  63 - 0x3f -- Sprite 0x8f
      12'h8F1: dout  = 8'b01111111; // 2289 : 127 - 0x7f
      12'h8F2: dout  = 8'b01111111; // 2290 : 127 - 0x7f
      12'h8F3: dout  = 8'b00011111; // 2291 :  31 - 0x1f
      12'h8F4: dout  = 8'b00111111; // 2292 :  63 - 0x3f
      12'h8F5: dout  = 8'b00111111; // 2293 :  63 - 0x3f
      12'h8F6: dout  = 8'b00000111; // 2294 :   7 - 0x7
      12'h8F7: dout  = 8'b00000110; // 2295 :   6 - 0x6
      12'h8F8: dout  = 8'b00000000; // 2296 :   0 - 0x0 -- plane 1
      12'h8F9: dout  = 8'b01100000; // 2297 :  96 - 0x60
      12'h8FA: dout  = 8'b01100000; // 2298 :  96 - 0x60
      12'h8FB: dout  = 8'b00000000; // 2299 :   0 - 0x0
      12'h8FC: dout  = 8'b00100000; // 2300 :  32 - 0x20
      12'h8FD: dout  = 8'b00110000; // 2301 :  48 - 0x30
      12'h8FE: dout  = 8'b00000100; // 2302 :   4 - 0x4
      12'h8FF: dout  = 8'b00000110; // 2303 :   6 - 0x6
      12'h900: dout  = 8'b00000011; // 2304 :   3 - 0x3 -- Sprite 0x90
      12'h901: dout  = 8'b00000111; // 2305 :   7 - 0x7
      12'h902: dout  = 8'b00001111; // 2306 :  15 - 0xf
      12'h903: dout  = 8'b00001111; // 2307 :  15 - 0xf
      12'h904: dout  = 8'b00001111; // 2308 :  15 - 0xf
      12'h905: dout  = 8'b00001111; // 2309 :  15 - 0xf
      12'h906: dout  = 8'b00000111; // 2310 :   7 - 0x7
      12'h907: dout  = 8'b00000011; // 2311 :   3 - 0x3
      12'h908: dout  = 8'b00000000; // 2312 :   0 - 0x0 -- plane 1
      12'h909: dout  = 8'b00000001; // 2313 :   1 - 0x1
      12'h90A: dout  = 8'b00000001; // 2314 :   1 - 0x1
      12'h90B: dout  = 8'b00000000; // 2315 :   0 - 0x0
      12'h90C: dout  = 8'b00000000; // 2316 :   0 - 0x0
      12'h90D: dout  = 8'b00000000; // 2317 :   0 - 0x0
      12'h90E: dout  = 8'b00000000; // 2318 :   0 - 0x0
      12'h90F: dout  = 8'b00000000; // 2319 :   0 - 0x0
      12'h910: dout  = 8'b11111000; // 2320 : 248 - 0xf8 -- Sprite 0x91
      12'h911: dout  = 8'b11111000; // 2321 : 248 - 0xf8
      12'h912: dout  = 8'b11111000; // 2322 : 248 - 0xf8
      12'h913: dout  = 8'b10100000; // 2323 : 160 - 0xa0
      12'h914: dout  = 8'b11100001; // 2324 : 225 - 0xe1
      12'h915: dout  = 8'b11111111; // 2325 : 255 - 0xff
      12'h916: dout  = 8'b11111111; // 2326 : 255 - 0xff
      12'h917: dout  = 8'b11111111; // 2327 : 255 - 0xff
      12'h918: dout  = 8'b11111110; // 2328 : 254 - 0xfe -- plane 1
      12'h919: dout  = 8'b11111111; // 2329 : 255 - 0xff
      12'h91A: dout  = 8'b11111111; // 2330 : 255 - 0xff
      12'h91B: dout  = 8'b01000000; // 2331 :  64 - 0x40
      12'h91C: dout  = 8'b00000001; // 2332 :   1 - 0x1
      12'h91D: dout  = 8'b00000011; // 2333 :   3 - 0x3
      12'h91E: dout  = 8'b00000011; // 2334 :   3 - 0x3
      12'h91F: dout  = 8'b00000011; // 2335 :   3 - 0x3
      12'h920: dout  = 8'b00001111; // 2336 :  15 - 0xf -- Sprite 0x92
      12'h921: dout  = 8'b00001111; // 2337 :  15 - 0xf
      12'h922: dout  = 8'b00001111; // 2338 :  15 - 0xf
      12'h923: dout  = 8'b00011111; // 2339 :  31 - 0x1f
      12'h924: dout  = 8'b00011111; // 2340 :  31 - 0x1f
      12'h925: dout  = 8'b00011111; // 2341 :  31 - 0x1f
      12'h926: dout  = 8'b00001111; // 2342 :  15 - 0xf
      12'h927: dout  = 8'b00000111; // 2343 :   7 - 0x7
      12'h928: dout  = 8'b00000001; // 2344 :   1 - 0x1 -- plane 1
      12'h929: dout  = 8'b00000001; // 2345 :   1 - 0x1
      12'h92A: dout  = 8'b00000000; // 2346 :   0 - 0x0
      12'h92B: dout  = 8'b00000000; // 2347 :   0 - 0x0
      12'h92C: dout  = 8'b00000000; // 2348 :   0 - 0x0
      12'h92D: dout  = 8'b00000000; // 2349 :   0 - 0x0
      12'h92E: dout  = 8'b00000000; // 2350 :   0 - 0x0
      12'h92F: dout  = 8'b00000000; // 2351 :   0 - 0x0
      12'h930: dout  = 8'b11100000; // 2352 : 224 - 0xe0 -- Sprite 0x93
      12'h931: dout  = 8'b11111000; // 2353 : 248 - 0xf8
      12'h932: dout  = 8'b11111000; // 2354 : 248 - 0xf8
      12'h933: dout  = 8'b11111000; // 2355 : 248 - 0xf8
      12'h934: dout  = 8'b11111111; // 2356 : 255 - 0xff
      12'h935: dout  = 8'b11111110; // 2357 : 254 - 0xfe
      12'h936: dout  = 8'b11110000; // 2358 : 240 - 0xf0
      12'h937: dout  = 8'b11000000; // 2359 : 192 - 0xc0
      12'h938: dout  = 8'b11100000; // 2360 : 224 - 0xe0 -- plane 1
      12'h939: dout  = 8'b11111110; // 2361 : 254 - 0xfe
      12'h93A: dout  = 8'b11111111; // 2362 : 255 - 0xff
      12'h93B: dout  = 8'b01111111; // 2363 : 127 - 0x7f
      12'h93C: dout  = 8'b00000011; // 2364 :   3 - 0x3
      12'h93D: dout  = 8'b00000010; // 2365 :   2 - 0x2
      12'h93E: dout  = 8'b00000000; // 2366 :   0 - 0x0
      12'h93F: dout  = 8'b00000000; // 2367 :   0 - 0x0
      12'h940: dout  = 8'b00000001; // 2368 :   1 - 0x1 -- Sprite 0x94
      12'h941: dout  = 8'b00001111; // 2369 :  15 - 0xf
      12'h942: dout  = 8'b00001111; // 2370 :  15 - 0xf
      12'h943: dout  = 8'b00011111; // 2371 :  31 - 0x1f
      12'h944: dout  = 8'b00111001; // 2372 :  57 - 0x39
      12'h945: dout  = 8'b00110011; // 2373 :  51 - 0x33
      12'h946: dout  = 8'b00110111; // 2374 :  55 - 0x37
      12'h947: dout  = 8'b01111111; // 2375 : 127 - 0x7f
      12'h948: dout  = 8'b00000001; // 2376 :   1 - 0x1 -- plane 1
      12'h949: dout  = 8'b00001101; // 2377 :  13 - 0xd
      12'h94A: dout  = 8'b00001000; // 2378 :   8 - 0x8
      12'h94B: dout  = 8'b00000000; // 2379 :   0 - 0x0
      12'h94C: dout  = 8'b00110110; // 2380 :  54 - 0x36
      12'h94D: dout  = 8'b00101100; // 2381 :  44 - 0x2c
      12'h94E: dout  = 8'b00001000; // 2382 :   8 - 0x8
      12'h94F: dout  = 8'b01100000; // 2383 :  96 - 0x60
      12'h950: dout  = 8'b01111111; // 2384 : 127 - 0x7f -- Sprite 0x95
      12'h951: dout  = 8'b00111111; // 2385 :  63 - 0x3f
      12'h952: dout  = 8'b00111111; // 2386 :  63 - 0x3f
      12'h953: dout  = 8'b00111111; // 2387 :  63 - 0x3f
      12'h954: dout  = 8'b00011111; // 2388 :  31 - 0x1f
      12'h955: dout  = 8'b00001111; // 2389 :  15 - 0xf
      12'h956: dout  = 8'b00001111; // 2390 :  15 - 0xf
      12'h957: dout  = 8'b00000001; // 2391 :   1 - 0x1
      12'h958: dout  = 8'b01100000; // 2392 :  96 - 0x60 -- plane 1
      12'h959: dout  = 8'b00000000; // 2393 :   0 - 0x0
      12'h95A: dout  = 8'b00100000; // 2394 :  32 - 0x20
      12'h95B: dout  = 8'b00110000; // 2395 :  48 - 0x30
      12'h95C: dout  = 8'b00000000; // 2396 :   0 - 0x0
      12'h95D: dout  = 8'b00001000; // 2397 :   8 - 0x8
      12'h95E: dout  = 8'b00001101; // 2398 :  13 - 0xd
      12'h95F: dout  = 8'b00000001; // 2399 :   1 - 0x1
      12'h960: dout  = 8'b00000000; // 2400 :   0 - 0x0 -- Sprite 0x96
      12'h961: dout  = 8'b00000000; // 2401 :   0 - 0x0
      12'h962: dout  = 8'b00000011; // 2402 :   3 - 0x3
      12'h963: dout  = 8'b00000011; // 2403 :   3 - 0x3
      12'h964: dout  = 8'b01000111; // 2404 :  71 - 0x47
      12'h965: dout  = 8'b01100111; // 2405 : 103 - 0x67
      12'h966: dout  = 8'b01110111; // 2406 : 119 - 0x77
      12'h967: dout  = 8'b01110111; // 2407 : 119 - 0x77
      12'h968: dout  = 8'b00000001; // 2408 :   1 - 0x1 -- plane 1
      12'h969: dout  = 8'b00000001; // 2409 :   1 - 0x1
      12'h96A: dout  = 8'b00000011; // 2410 :   3 - 0x3
      12'h96B: dout  = 8'b01000011; // 2411 :  67 - 0x43
      12'h96C: dout  = 8'b01100111; // 2412 : 103 - 0x67
      12'h96D: dout  = 8'b01110111; // 2413 : 119 - 0x77
      12'h96E: dout  = 8'b01111011; // 2414 : 123 - 0x7b
      12'h96F: dout  = 8'b01111000; // 2415 : 120 - 0x78
      12'h970: dout  = 8'b00000000; // 2416 :   0 - 0x0 -- Sprite 0x97
      12'h971: dout  = 8'b00000000; // 2417 :   0 - 0x0
      12'h972: dout  = 8'b00000000; // 2418 :   0 - 0x0
      12'h973: dout  = 8'b00000000; // 2419 :   0 - 0x0
      12'h974: dout  = 8'b10001000; // 2420 : 136 - 0x88
      12'h975: dout  = 8'b10011000; // 2421 : 152 - 0x98
      12'h976: dout  = 8'b11111000; // 2422 : 248 - 0xf8
      12'h977: dout  = 8'b11110000; // 2423 : 240 - 0xf0
      12'h978: dout  = 8'b00000000; // 2424 :   0 - 0x0 -- plane 1
      12'h979: dout  = 8'b00000000; // 2425 :   0 - 0x0
      12'h97A: dout  = 8'b10000000; // 2426 : 128 - 0x80
      12'h97B: dout  = 8'b10000100; // 2427 : 132 - 0x84
      12'h97C: dout  = 8'b11001100; // 2428 : 204 - 0xcc
      12'h97D: dout  = 8'b11011100; // 2429 : 220 - 0xdc
      12'h97E: dout  = 8'b10111100; // 2430 : 188 - 0xbc
      12'h97F: dout  = 8'b00111100; // 2431 :  60 - 0x3c
      12'h980: dout  = 8'b01111110; // 2432 : 126 - 0x7e -- Sprite 0x98
      12'h981: dout  = 8'b01111111; // 2433 : 127 - 0x7f
      12'h982: dout  = 8'b11111111; // 2434 : 255 - 0xff
      12'h983: dout  = 8'b00011111; // 2435 :  31 - 0x1f
      12'h984: dout  = 8'b00000111; // 2436 :   7 - 0x7
      12'h985: dout  = 8'b00110000; // 2437 :  48 - 0x30
      12'h986: dout  = 8'b00011100; // 2438 :  28 - 0x1c
      12'h987: dout  = 8'b00001100; // 2439 :  12 - 0xc
      12'h988: dout  = 8'b00110011; // 2440 :  51 - 0x33 -- plane 1
      12'h989: dout  = 8'b00000111; // 2441 :   7 - 0x7
      12'h98A: dout  = 8'b00000111; // 2442 :   7 - 0x7
      12'h98B: dout  = 8'b11100011; // 2443 : 227 - 0xe3
      12'h98C: dout  = 8'b00111000; // 2444 :  56 - 0x38
      12'h98D: dout  = 8'b00111111; // 2445 :  63 - 0x3f
      12'h98E: dout  = 8'b00011100; // 2446 :  28 - 0x1c
      12'h98F: dout  = 8'b00001100; // 2447 :  12 - 0xc
      12'h990: dout  = 8'b01111110; // 2448 : 126 - 0x7e -- Sprite 0x99
      12'h991: dout  = 8'b00111000; // 2449 :  56 - 0x38
      12'h992: dout  = 8'b11110110; // 2450 : 246 - 0xf6
      12'h993: dout  = 8'b11101101; // 2451 : 237 - 0xed
      12'h994: dout  = 8'b11011111; // 2452 : 223 - 0xdf
      12'h995: dout  = 8'b00111000; // 2453 :  56 - 0x38
      12'h996: dout  = 8'b01110000; // 2454 : 112 - 0x70
      12'h997: dout  = 8'b01100000; // 2455 :  96 - 0x60
      12'h998: dout  = 8'b10011000; // 2456 : 152 - 0x98 -- plane 1
      12'h999: dout  = 8'b11000111; // 2457 : 199 - 0xc7
      12'h99A: dout  = 8'b11001000; // 2458 : 200 - 0xc8
      12'h99B: dout  = 8'b10010010; // 2459 : 146 - 0x92
      12'h99C: dout  = 8'b00110000; // 2460 :  48 - 0x30
      12'h99D: dout  = 8'b11111000; // 2461 : 248 - 0xf8
      12'h99E: dout  = 8'b01110000; // 2462 : 112 - 0x70
      12'h99F: dout  = 8'b01100000; // 2463 :  96 - 0x60
      12'h9A0: dout  = 8'b00000000; // 2464 :   0 - 0x0 -- Sprite 0x9a
      12'h9A1: dout  = 8'b00000000; // 2465 :   0 - 0x0
      12'h9A2: dout  = 8'b00000000; // 2466 :   0 - 0x0
      12'h9A3: dout  = 8'b00000011; // 2467 :   3 - 0x3
      12'h9A4: dout  = 8'b00000011; // 2468 :   3 - 0x3
      12'h9A5: dout  = 8'b01000111; // 2469 :  71 - 0x47
      12'h9A6: dout  = 8'b01100111; // 2470 : 103 - 0x67
      12'h9A7: dout  = 8'b01110111; // 2471 : 119 - 0x77
      12'h9A8: dout  = 8'b00000000; // 2472 :   0 - 0x0 -- plane 1
      12'h9A9: dout  = 8'b00000001; // 2473 :   1 - 0x1
      12'h9AA: dout  = 8'b00000001; // 2474 :   1 - 0x1
      12'h9AB: dout  = 8'b00000011; // 2475 :   3 - 0x3
      12'h9AC: dout  = 8'b01000011; // 2476 :  67 - 0x43
      12'h9AD: dout  = 8'b01100111; // 2477 : 103 - 0x67
      12'h9AE: dout  = 8'b01110111; // 2478 : 119 - 0x77
      12'h9AF: dout  = 8'b01111011; // 2479 : 123 - 0x7b
      12'h9B0: dout  = 8'b00000000; // 2480 :   0 - 0x0 -- Sprite 0x9b
      12'h9B1: dout  = 8'b00000000; // 2481 :   0 - 0x0
      12'h9B2: dout  = 8'b00000000; // 2482 :   0 - 0x0
      12'h9B3: dout  = 8'b00000000; // 2483 :   0 - 0x0
      12'h9B4: dout  = 8'b00000000; // 2484 :   0 - 0x0
      12'h9B5: dout  = 8'b10001000; // 2485 : 136 - 0x88
      12'h9B6: dout  = 8'b10011000; // 2486 : 152 - 0x98
      12'h9B7: dout  = 8'b11111000; // 2487 : 248 - 0xf8
      12'h9B8: dout  = 8'b00000000; // 2488 :   0 - 0x0 -- plane 1
      12'h9B9: dout  = 8'b00000000; // 2489 :   0 - 0x0
      12'h9BA: dout  = 8'b00000000; // 2490 :   0 - 0x0
      12'h9BB: dout  = 8'b10000000; // 2491 : 128 - 0x80
      12'h9BC: dout  = 8'b10000100; // 2492 : 132 - 0x84
      12'h9BD: dout  = 8'b11001100; // 2493 : 204 - 0xcc
      12'h9BE: dout  = 8'b11011100; // 2494 : 220 - 0xdc
      12'h9BF: dout  = 8'b10111100; // 2495 : 188 - 0xbc
      12'h9C0: dout  = 8'b01110111; // 2496 : 119 - 0x77 -- Sprite 0x9c
      12'h9C1: dout  = 8'b01111110; // 2497 : 126 - 0x7e
      12'h9C2: dout  = 8'b01111111; // 2498 : 127 - 0x7f
      12'h9C3: dout  = 8'b11111111; // 2499 : 255 - 0xff
      12'h9C4: dout  = 8'b00011111; // 2500 :  31 - 0x1f
      12'h9C5: dout  = 8'b00000111; // 2501 :   7 - 0x7
      12'h9C6: dout  = 8'b01110000; // 2502 : 112 - 0x70
      12'h9C7: dout  = 8'b11110000; // 2503 : 240 - 0xf0
      12'h9C8: dout  = 8'b01111000; // 2504 : 120 - 0x78 -- plane 1
      12'h9C9: dout  = 8'b00110011; // 2505 :  51 - 0x33
      12'h9CA: dout  = 8'b00000111; // 2506 :   7 - 0x7
      12'h9CB: dout  = 8'b00000111; // 2507 :   7 - 0x7
      12'h9CC: dout  = 8'b11100011; // 2508 : 227 - 0xe3
      12'h9CD: dout  = 8'b00111000; // 2509 :  56 - 0x38
      12'h9CE: dout  = 8'b01111111; // 2510 : 127 - 0x7f
      12'h9CF: dout  = 8'b11110000; // 2511 : 240 - 0xf0
      12'h9D0: dout  = 8'b11110000; // 2512 : 240 - 0xf0 -- Sprite 0x9d
      12'h9D1: dout  = 8'b01111110; // 2513 : 126 - 0x7e
      12'h9D2: dout  = 8'b00111000; // 2514 :  56 - 0x38
      12'h9D3: dout  = 8'b11110110; // 2515 : 246 - 0xf6
      12'h9D4: dout  = 8'b11101101; // 2516 : 237 - 0xed
      12'h9D5: dout  = 8'b11011111; // 2517 : 223 - 0xdf
      12'h9D6: dout  = 8'b00111000; // 2518 :  56 - 0x38
      12'h9D7: dout  = 8'b00111100; // 2519 :  60 - 0x3c
      12'h9D8: dout  = 8'b00111100; // 2520 :  60 - 0x3c -- plane 1
      12'h9D9: dout  = 8'b10011000; // 2521 : 152 - 0x98
      12'h9DA: dout  = 8'b11000111; // 2522 : 199 - 0xc7
      12'h9DB: dout  = 8'b11001000; // 2523 : 200 - 0xc8
      12'h9DC: dout  = 8'b10010010; // 2524 : 146 - 0x92
      12'h9DD: dout  = 8'b00110000; // 2525 :  48 - 0x30
      12'h9DE: dout  = 8'b11111000; // 2526 : 248 - 0xf8
      12'h9DF: dout  = 8'b00111100; // 2527 :  60 - 0x3c
      12'h9E0: dout  = 8'b00000011; // 2528 :   3 - 0x3 -- Sprite 0x9e
      12'h9E1: dout  = 8'b00000111; // 2529 :   7 - 0x7
      12'h9E2: dout  = 8'b00001010; // 2530 :  10 - 0xa
      12'h9E3: dout  = 8'b00011010; // 2531 :  26 - 0x1a
      12'h9E4: dout  = 8'b00011100; // 2532 :  28 - 0x1c
      12'h9E5: dout  = 8'b00011110; // 2533 :  30 - 0x1e
      12'h9E6: dout  = 8'b00001011; // 2534 :  11 - 0xb
      12'h9E7: dout  = 8'b00001000; // 2535 :   8 - 0x8
      12'h9E8: dout  = 8'b00000000; // 2536 :   0 - 0x0 -- plane 1
      12'h9E9: dout  = 8'b00010000; // 2537 :  16 - 0x10
      12'h9EA: dout  = 8'b01111111; // 2538 : 127 - 0x7f
      12'h9EB: dout  = 8'b01111111; // 2539 : 127 - 0x7f
      12'h9EC: dout  = 8'b01111111; // 2540 : 127 - 0x7f
      12'h9ED: dout  = 8'b00011111; // 2541 :  31 - 0x1f
      12'h9EE: dout  = 8'b00001111; // 2542 :  15 - 0xf
      12'h9EF: dout  = 8'b00001111; // 2543 :  15 - 0xf
      12'h9F0: dout  = 8'b00011100; // 2544 :  28 - 0x1c -- Sprite 0x9f
      12'h9F1: dout  = 8'b00111111; // 2545 :  63 - 0x3f
      12'h9F2: dout  = 8'b00111111; // 2546 :  63 - 0x3f
      12'h9F3: dout  = 8'b00111101; // 2547 :  61 - 0x3d
      12'h9F4: dout  = 8'b00111111; // 2548 :  63 - 0x3f
      12'h9F5: dout  = 8'b00011111; // 2549 :  31 - 0x1f
      12'h9F6: dout  = 8'b00000000; // 2550 :   0 - 0x0
      12'h9F7: dout  = 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout  = 8'b00000011; // 2552 :   3 - 0x3 -- plane 1
      12'h9F9: dout  = 8'b00110011; // 2553 :  51 - 0x33
      12'h9FA: dout  = 8'b00111001; // 2554 :  57 - 0x39
      12'h9FB: dout  = 8'b00111010; // 2555 :  58 - 0x3a
      12'h9FC: dout  = 8'b00111000; // 2556 :  56 - 0x38
      12'h9FD: dout  = 8'b00011000; // 2557 :  24 - 0x18
      12'h9FE: dout  = 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout  = 8'b00000000; // 2560 :   0 - 0x0 -- Sprite 0xa0
      12'hA01: dout  = 8'b00000000; // 2561 :   0 - 0x0
      12'hA02: dout  = 8'b00000100; // 2562 :   4 - 0x4
      12'hA03: dout  = 8'b01001100; // 2563 :  76 - 0x4c
      12'hA04: dout  = 8'b01001110; // 2564 :  78 - 0x4e
      12'hA05: dout  = 8'b01001110; // 2565 :  78 - 0x4e
      12'hA06: dout  = 8'b01000110; // 2566 :  70 - 0x46
      12'hA07: dout  = 8'b01101111; // 2567 : 111 - 0x6f
      12'hA08: dout  = 8'b00010000; // 2568 :  16 - 0x10 -- plane 1
      12'hA09: dout  = 8'b00111000; // 2569 :  56 - 0x38
      12'hA0A: dout  = 8'b00111100; // 2570 :  60 - 0x3c
      12'hA0B: dout  = 8'b01110100; // 2571 : 116 - 0x74
      12'hA0C: dout  = 8'b01110110; // 2572 : 118 - 0x76
      12'hA0D: dout  = 8'b01110110; // 2573 : 118 - 0x76
      12'hA0E: dout  = 8'b01111110; // 2574 : 126 - 0x7e
      12'hA0F: dout  = 8'b01111101; // 2575 : 125 - 0x7d
      12'hA10: dout  = 8'b00000000; // 2576 :   0 - 0x0 -- Sprite 0xa1
      12'hA11: dout  = 8'b00011111; // 2577 :  31 - 0x1f
      12'hA12: dout  = 8'b00111111; // 2578 :  63 - 0x3f
      12'hA13: dout  = 8'b00111111; // 2579 :  63 - 0x3f
      12'hA14: dout  = 8'b01001111; // 2580 :  79 - 0x4f
      12'hA15: dout  = 8'b01011111; // 2581 :  95 - 0x5f
      12'hA16: dout  = 8'b01111111; // 2582 : 127 - 0x7f
      12'hA17: dout  = 8'b01111111; // 2583 : 127 - 0x7f
      12'hA18: dout  = 8'b00000000; // 2584 :   0 - 0x0 -- plane 1
      12'hA19: dout  = 8'b00000000; // 2585 :   0 - 0x0
      12'hA1A: dout  = 8'b00010001; // 2586 :  17 - 0x11
      12'hA1B: dout  = 8'b00001010; // 2587 :  10 - 0xa
      12'hA1C: dout  = 8'b00110100; // 2588 :  52 - 0x34
      12'hA1D: dout  = 8'b00101010; // 2589 :  42 - 0x2a
      12'hA1E: dout  = 8'b01010001; // 2590 :  81 - 0x51
      12'hA1F: dout  = 8'b00100000; // 2591 :  32 - 0x20
      12'hA20: dout  = 8'b01111111; // 2592 : 127 - 0x7f -- Sprite 0xa2
      12'hA21: dout  = 8'b01100111; // 2593 : 103 - 0x67
      12'hA22: dout  = 8'b10100011; // 2594 : 163 - 0xa3
      12'hA23: dout  = 8'b10110000; // 2595 : 176 - 0xb0
      12'hA24: dout  = 8'b11011000; // 2596 : 216 - 0xd8
      12'hA25: dout  = 8'b11011110; // 2597 : 222 - 0xde
      12'hA26: dout  = 8'b11011100; // 2598 : 220 - 0xdc
      12'hA27: dout  = 8'b11001000; // 2599 : 200 - 0xc8
      12'hA28: dout  = 8'b01111111; // 2600 : 127 - 0x7f -- plane 1
      12'hA29: dout  = 8'b01100111; // 2601 : 103 - 0x67
      12'hA2A: dout  = 8'b01100011; // 2602 :  99 - 0x63
      12'hA2B: dout  = 8'b01110000; // 2603 : 112 - 0x70
      12'hA2C: dout  = 8'b00111000; // 2604 :  56 - 0x38
      12'hA2D: dout  = 8'b00111110; // 2605 :  62 - 0x3e
      12'hA2E: dout  = 8'b01111100; // 2606 : 124 - 0x7c
      12'hA2F: dout  = 8'b10111000; // 2607 : 184 - 0xb8
      12'hA30: dout  = 8'b01111111; // 2608 : 127 - 0x7f -- Sprite 0xa3
      12'hA31: dout  = 8'b01111111; // 2609 : 127 - 0x7f
      12'hA32: dout  = 8'b01111111; // 2610 : 127 - 0x7f
      12'hA33: dout  = 8'b00011111; // 2611 :  31 - 0x1f
      12'hA34: dout  = 8'b01000111; // 2612 :  71 - 0x47
      12'hA35: dout  = 8'b01110000; // 2613 : 112 - 0x70
      12'hA36: dout  = 8'b01110000; // 2614 : 112 - 0x70
      12'hA37: dout  = 8'b00111001; // 2615 :  57 - 0x39
      12'hA38: dout  = 8'b01010001; // 2616 :  81 - 0x51 -- plane 1
      12'hA39: dout  = 8'b00001010; // 2617 :  10 - 0xa
      12'hA3A: dout  = 8'b00000100; // 2618 :   4 - 0x4
      12'hA3B: dout  = 8'b11101010; // 2619 : 234 - 0xea
      12'hA3C: dout  = 8'b01111001; // 2620 : 121 - 0x79
      12'hA3D: dout  = 8'b01111111; // 2621 : 127 - 0x7f
      12'hA3E: dout  = 8'b01110000; // 2622 : 112 - 0x70
      12'hA3F: dout  = 8'b00111001; // 2623 :  57 - 0x39
      12'hA40: dout  = 8'b11101000; // 2624 : 232 - 0xe8 -- Sprite 0xa4
      12'hA41: dout  = 8'b11101000; // 2625 : 232 - 0xe8
      12'hA42: dout  = 8'b11100000; // 2626 : 224 - 0xe0
      12'hA43: dout  = 8'b11000000; // 2627 : 192 - 0xc0
      12'hA44: dout  = 8'b00010000; // 2628 :  16 - 0x10
      12'hA45: dout  = 8'b01110000; // 2629 : 112 - 0x70
      12'hA46: dout  = 8'b11100000; // 2630 : 224 - 0xe0
      12'hA47: dout  = 8'b11000000; // 2631 : 192 - 0xc0
      12'hA48: dout  = 8'b01011000; // 2632 :  88 - 0x58 -- plane 1
      12'hA49: dout  = 8'b00111000; // 2633 :  56 - 0x38
      12'hA4A: dout  = 8'b00010000; // 2634 :  16 - 0x10
      12'hA4B: dout  = 8'b00110000; // 2635 :  48 - 0x30
      12'hA4C: dout  = 8'b11110000; // 2636 : 240 - 0xf0
      12'hA4D: dout  = 8'b11110000; // 2637 : 240 - 0xf0
      12'hA4E: dout  = 8'b11100000; // 2638 : 224 - 0xe0
      12'hA4F: dout  = 8'b11000000; // 2639 : 192 - 0xc0
      12'hA50: dout  = 8'b00000000; // 2640 :   0 - 0x0 -- Sprite 0xa5
      12'hA51: dout  = 8'b00000000; // 2641 :   0 - 0x0
      12'hA52: dout  = 8'b00000000; // 2642 :   0 - 0x0
      12'hA53: dout  = 8'b00100000; // 2643 :  32 - 0x20
      12'hA54: dout  = 8'b01100110; // 2644 : 102 - 0x66
      12'hA55: dout  = 8'b01100110; // 2645 : 102 - 0x66
      12'hA56: dout  = 8'b01100110; // 2646 : 102 - 0x66
      12'hA57: dout  = 8'b01100010; // 2647 :  98 - 0x62
      12'hA58: dout  = 8'b00000000; // 2648 :   0 - 0x0 -- plane 1
      12'hA59: dout  = 8'b00001000; // 2649 :   8 - 0x8
      12'hA5A: dout  = 8'b00011100; // 2650 :  28 - 0x1c
      12'hA5B: dout  = 8'b00111100; // 2651 :  60 - 0x3c
      12'hA5C: dout  = 8'b01111010; // 2652 : 122 - 0x7a
      12'hA5D: dout  = 8'b01111010; // 2653 : 122 - 0x7a
      12'hA5E: dout  = 8'b01111010; // 2654 : 122 - 0x7a
      12'hA5F: dout  = 8'b01111110; // 2655 : 126 - 0x7e
      12'hA60: dout  = 8'b00000000; // 2656 :   0 - 0x0 -- Sprite 0xa6
      12'hA61: dout  = 8'b00000000; // 2657 :   0 - 0x0
      12'hA62: dout  = 8'b00011111; // 2658 :  31 - 0x1f
      12'hA63: dout  = 8'b00111111; // 2659 :  63 - 0x3f
      12'hA64: dout  = 8'b01111111; // 2660 : 127 - 0x7f
      12'hA65: dout  = 8'b01001111; // 2661 :  79 - 0x4f
      12'hA66: dout  = 8'b01011111; // 2662 :  95 - 0x5f
      12'hA67: dout  = 8'b01111111; // 2663 : 127 - 0x7f
      12'hA68: dout  = 8'b00000000; // 2664 :   0 - 0x0 -- plane 1
      12'hA69: dout  = 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout  = 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout  = 8'b00010001; // 2667 :  17 - 0x11
      12'hA6C: dout  = 8'b00001010; // 2668 :  10 - 0xa
      12'hA6D: dout  = 8'b00110100; // 2669 :  52 - 0x34
      12'hA6E: dout  = 8'b00101010; // 2670 :  42 - 0x2a
      12'hA6F: dout  = 8'b01010001; // 2671 :  81 - 0x51
      12'hA70: dout  = 8'b01110111; // 2672 : 119 - 0x77 -- Sprite 0xa7
      12'hA71: dout  = 8'b01111111; // 2673 : 127 - 0x7f
      12'hA72: dout  = 8'b00111111; // 2674 :  63 - 0x3f
      12'hA73: dout  = 8'b10110111; // 2675 : 183 - 0xb7
      12'hA74: dout  = 8'b10110011; // 2676 : 179 - 0xb3
      12'hA75: dout  = 8'b11011011; // 2677 : 219 - 0xdb
      12'hA76: dout  = 8'b11011010; // 2678 : 218 - 0xda
      12'hA77: dout  = 8'b11011000; // 2679 : 216 - 0xd8
      12'hA78: dout  = 8'b01111111; // 2680 : 127 - 0x7f -- plane 1
      12'hA79: dout  = 8'b01111101; // 2681 : 125 - 0x7d
      12'hA7A: dout  = 8'b00111111; // 2682 :  63 - 0x3f
      12'hA7B: dout  = 8'b00110111; // 2683 :  55 - 0x37
      12'hA7C: dout  = 8'b00110011; // 2684 :  51 - 0x33
      12'hA7D: dout  = 8'b00111011; // 2685 :  59 - 0x3b
      12'hA7E: dout  = 8'b00111010; // 2686 :  58 - 0x3a
      12'hA7F: dout  = 8'b01111000; // 2687 : 120 - 0x78
      12'hA80: dout  = 8'b01111111; // 2688 : 127 - 0x7f -- Sprite 0xa8
      12'hA81: dout  = 8'b01111111; // 2689 : 127 - 0x7f
      12'hA82: dout  = 8'b01111111; // 2690 : 127 - 0x7f
      12'hA83: dout  = 8'b01111111; // 2691 : 127 - 0x7f
      12'hA84: dout  = 8'b00011111; // 2692 :  31 - 0x1f
      12'hA85: dout  = 8'b00000111; // 2693 :   7 - 0x7
      12'hA86: dout  = 8'b01110000; // 2694 : 112 - 0x70
      12'hA87: dout  = 8'b11110000; // 2695 : 240 - 0xf0
      12'hA88: dout  = 8'b00100000; // 2696 :  32 - 0x20 -- plane 1
      12'hA89: dout  = 8'b01010001; // 2697 :  81 - 0x51
      12'hA8A: dout  = 8'b00001010; // 2698 :  10 - 0xa
      12'hA8B: dout  = 8'b00000100; // 2699 :   4 - 0x4
      12'hA8C: dout  = 8'b11101010; // 2700 : 234 - 0xea
      12'hA8D: dout  = 8'b00111001; // 2701 :  57 - 0x39
      12'hA8E: dout  = 8'b01111111; // 2702 : 127 - 0x7f
      12'hA8F: dout  = 8'b11110000; // 2703 : 240 - 0xf0
      12'hA90: dout  = 8'b11001100; // 2704 : 204 - 0xcc -- Sprite 0xa9
      12'hA91: dout  = 8'b11101000; // 2705 : 232 - 0xe8
      12'hA92: dout  = 8'b11101000; // 2706 : 232 - 0xe8
      12'hA93: dout  = 8'b11100000; // 2707 : 224 - 0xe0
      12'hA94: dout  = 8'b11000000; // 2708 : 192 - 0xc0
      12'hA95: dout  = 8'b00011000; // 2709 :  24 - 0x18
      12'hA96: dout  = 8'b01111100; // 2710 : 124 - 0x7c
      12'hA97: dout  = 8'b00111110; // 2711 :  62 - 0x3e
      12'hA98: dout  = 8'b10111100; // 2712 : 188 - 0xbc -- plane 1
      12'hA99: dout  = 8'b01011000; // 2713 :  88 - 0x58
      12'hA9A: dout  = 8'b00111000; // 2714 :  56 - 0x38
      12'hA9B: dout  = 8'b00010000; // 2715 :  16 - 0x10
      12'hA9C: dout  = 8'b00110000; // 2716 :  48 - 0x30
      12'hA9D: dout  = 8'b11111000; // 2717 : 248 - 0xf8
      12'hA9E: dout  = 8'b11111100; // 2718 : 252 - 0xfc
      12'hA9F: dout  = 8'b00111110; // 2719 :  62 - 0x3e
      12'hAA0: dout  = 8'b00000011; // 2720 :   3 - 0x3 -- Sprite 0xaa
      12'hAA1: dout  = 8'b00001111; // 2721 :  15 - 0xf
      12'hAA2: dout  = 8'b00011111; // 2722 :  31 - 0x1f
      12'hAA3: dout  = 8'b00111111; // 2723 :  63 - 0x3f
      12'hAA4: dout  = 8'b00111011; // 2724 :  59 - 0x3b
      12'hAA5: dout  = 8'b00111111; // 2725 :  63 - 0x3f
      12'hAA6: dout  = 8'b01111111; // 2726 : 127 - 0x7f
      12'hAA7: dout  = 8'b01111111; // 2727 : 127 - 0x7f
      12'hAA8: dout  = 8'b00000000; // 2728 :   0 - 0x0 -- plane 1
      12'hAA9: dout  = 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout  = 8'b00000000; // 2730 :   0 - 0x0
      12'hAAB: dout  = 8'b00000110; // 2731 :   6 - 0x6
      12'hAAC: dout  = 8'b00001110; // 2732 :  14 - 0xe
      12'hAAD: dout  = 8'b00001100; // 2733 :  12 - 0xc
      12'hAAE: dout  = 8'b00000000; // 2734 :   0 - 0x0
      12'hAAF: dout  = 8'b00000000; // 2735 :   0 - 0x0
      12'hAB0: dout  = 8'b10000000; // 2736 : 128 - 0x80 -- Sprite 0xab
      12'hAB1: dout  = 8'b11110000; // 2737 : 240 - 0xf0
      12'hAB2: dout  = 8'b11111000; // 2738 : 248 - 0xf8
      12'hAB3: dout  = 8'b11111100; // 2739 : 252 - 0xfc
      12'hAB4: dout  = 8'b11111110; // 2740 : 254 - 0xfe
      12'hAB5: dout  = 8'b11111110; // 2741 : 254 - 0xfe
      12'hAB6: dout  = 8'b11111111; // 2742 : 255 - 0xff
      12'hAB7: dout  = 8'b11111110; // 2743 : 254 - 0xfe
      12'hAB8: dout  = 8'b00000000; // 2744 :   0 - 0x0 -- plane 1
      12'hAB9: dout  = 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout  = 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout  = 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout  = 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout  = 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout  = 8'b00001111; // 2750 :  15 - 0xf
      12'hABF: dout  = 8'b00011000; // 2751 :  24 - 0x18
      12'hAC0: dout  = 8'b01111111; // 2752 : 127 - 0x7f -- Sprite 0xac
      12'hAC1: dout  = 8'b01111111; // 2753 : 127 - 0x7f
      12'hAC2: dout  = 8'b01111111; // 2754 : 127 - 0x7f
      12'hAC3: dout  = 8'b01111111; // 2755 : 127 - 0x7f
      12'hAC4: dout  = 8'b11111111; // 2756 : 255 - 0xff
      12'hAC5: dout  = 8'b00001111; // 2757 :  15 - 0xf
      12'hAC6: dout  = 8'b00000011; // 2758 :   3 - 0x3
      12'hAC7: dout  = 8'b00000000; // 2759 :   0 - 0x0
      12'hAC8: dout  = 8'b00000000; // 2760 :   0 - 0x0 -- plane 1
      12'hAC9: dout  = 8'b00000000; // 2761 :   0 - 0x0
      12'hACA: dout  = 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout  = 8'b00000000; // 2763 :   0 - 0x0
      12'hACC: dout  = 8'b11111000; // 2764 : 248 - 0xf8
      12'hACD: dout  = 8'b00111110; // 2765 :  62 - 0x3e
      12'hACE: dout  = 8'b00111011; // 2766 :  59 - 0x3b
      12'hACF: dout  = 8'b00011000; // 2767 :  24 - 0x18
      12'hAD0: dout  = 8'b11111110; // 2768 : 254 - 0xfe -- Sprite 0xad
      12'hAD1: dout  = 8'b11111011; // 2769 : 251 - 0xfb
      12'hAD2: dout  = 8'b11111111; // 2770 : 255 - 0xff
      12'hAD3: dout  = 8'b11111111; // 2771 : 255 - 0xff
      12'hAD4: dout  = 8'b11110110; // 2772 : 246 - 0xf6
      12'hAD5: dout  = 8'b11100000; // 2773 : 224 - 0xe0
      12'hAD6: dout  = 8'b11000000; // 2774 : 192 - 0xc0
      12'hAD7: dout  = 8'b00000000; // 2775 :   0 - 0x0
      12'hAD8: dout  = 8'b00010000; // 2776 :  16 - 0x10 -- plane 1
      12'hAD9: dout  = 8'b00010100; // 2777 :  20 - 0x14
      12'hADA: dout  = 8'b00010000; // 2778 :  16 - 0x10
      12'hADB: dout  = 8'b00010000; // 2779 :  16 - 0x10
      12'hADC: dout  = 8'b00111000; // 2780 :  56 - 0x38
      12'hADD: dout  = 8'b01111000; // 2781 : 120 - 0x78
      12'hADE: dout  = 8'b11111000; // 2782 : 248 - 0xf8
      12'hADF: dout  = 8'b00110000; // 2783 :  48 - 0x30
      12'hAE0: dout  = 8'b00000000; // 2784 :   0 - 0x0 -- Sprite 0xae
      12'hAE1: dout  = 8'b00000011; // 2785 :   3 - 0x3
      12'hAE2: dout  = 8'b00001111; // 2786 :  15 - 0xf
      12'hAE3: dout  = 8'b00011111; // 2787 :  31 - 0x1f
      12'hAE4: dout  = 8'b00111111; // 2788 :  63 - 0x3f
      12'hAE5: dout  = 8'b00111011; // 2789 :  59 - 0x3b
      12'hAE6: dout  = 8'b00111111; // 2790 :  63 - 0x3f
      12'hAE7: dout  = 8'b01111111; // 2791 : 127 - 0x7f
      12'hAE8: dout  = 8'b00000000; // 2792 :   0 - 0x0 -- plane 1
      12'hAE9: dout  = 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout  = 8'b00000000; // 2794 :   0 - 0x0
      12'hAEB: dout  = 8'b00000000; // 2795 :   0 - 0x0
      12'hAEC: dout  = 8'b00000110; // 2796 :   6 - 0x6
      12'hAED: dout  = 8'b00001110; // 2797 :  14 - 0xe
      12'hAEE: dout  = 8'b00001100; // 2798 :  12 - 0xc
      12'hAEF: dout  = 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout  = 8'b00000000; // 2800 :   0 - 0x0 -- Sprite 0xaf
      12'hAF1: dout  = 8'b11000000; // 2801 : 192 - 0xc0
      12'hAF2: dout  = 8'b11110000; // 2802 : 240 - 0xf0
      12'hAF3: dout  = 8'b11111000; // 2803 : 248 - 0xf8
      12'hAF4: dout  = 8'b11111100; // 2804 : 252 - 0xfc
      12'hAF5: dout  = 8'b11111110; // 2805 : 254 - 0xfe
      12'hAF6: dout  = 8'b11111110; // 2806 : 254 - 0xfe
      12'hAF7: dout  = 8'b11111111; // 2807 : 255 - 0xff
      12'hAF8: dout  = 8'b00000000; // 2808 :   0 - 0x0 -- plane 1
      12'hAF9: dout  = 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout  = 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout  = 8'b00000000; // 2811 :   0 - 0x0
      12'hAFC: dout  = 8'b00000000; // 2812 :   0 - 0x0
      12'hAFD: dout  = 8'b00000000; // 2813 :   0 - 0x0
      12'hAFE: dout  = 8'b00000000; // 2814 :   0 - 0x0
      12'hAFF: dout  = 8'b00001111; // 2815 :  15 - 0xf
      12'hB00: dout  = 8'b01111111; // 2816 : 127 - 0x7f -- Sprite 0xb0
      12'hB01: dout  = 8'b01111111; // 2817 : 127 - 0x7f
      12'hB02: dout  = 8'b01111111; // 2818 : 127 - 0x7f
      12'hB03: dout  = 8'b01111111; // 2819 : 127 - 0x7f
      12'hB04: dout  = 8'b01111111; // 2820 : 127 - 0x7f
      12'hB05: dout  = 8'b11111111; // 2821 : 255 - 0xff
      12'hB06: dout  = 8'b00001111; // 2822 :  15 - 0xf
      12'hB07: dout  = 8'b00000011; // 2823 :   3 - 0x3
      12'hB08: dout  = 8'b00000000; // 2824 :   0 - 0x0 -- plane 1
      12'hB09: dout  = 8'b00000000; // 2825 :   0 - 0x0
      12'hB0A: dout  = 8'b00000000; // 2826 :   0 - 0x0
      12'hB0B: dout  = 8'b00000000; // 2827 :   0 - 0x0
      12'hB0C: dout  = 8'b00000000; // 2828 :   0 - 0x0
      12'hB0D: dout  = 8'b11111000; // 2829 : 248 - 0xf8
      12'hB0E: dout  = 8'b01111110; // 2830 : 126 - 0x7e
      12'hB0F: dout  = 8'b11110011; // 2831 : 243 - 0xf3
      12'hB10: dout  = 8'b11111110; // 2832 : 254 - 0xfe -- Sprite 0xb1
      12'hB11: dout  = 8'b11111110; // 2833 : 254 - 0xfe
      12'hB12: dout  = 8'b11111011; // 2834 : 251 - 0xfb
      12'hB13: dout  = 8'b11111111; // 2835 : 255 - 0xff
      12'hB14: dout  = 8'b11111111; // 2836 : 255 - 0xff
      12'hB15: dout  = 8'b11110110; // 2837 : 246 - 0xf6
      12'hB16: dout  = 8'b11100000; // 2838 : 224 - 0xe0
      12'hB17: dout  = 8'b11000000; // 2839 : 192 - 0xc0
      12'hB18: dout  = 8'b00011000; // 2840 :  24 - 0x18 -- plane 1
      12'hB19: dout  = 8'b00010000; // 2841 :  16 - 0x10
      12'hB1A: dout  = 8'b00010100; // 2842 :  20 - 0x14
      12'hB1B: dout  = 8'b00010000; // 2843 :  16 - 0x10
      12'hB1C: dout  = 8'b00010000; // 2844 :  16 - 0x10
      12'hB1D: dout  = 8'b00111000; // 2845 :  56 - 0x38
      12'hB1E: dout  = 8'b01111100; // 2846 : 124 - 0x7c
      12'hB1F: dout  = 8'b11011110; // 2847 : 222 - 0xde
      12'hB20: dout  = 8'b00000000; // 2848 :   0 - 0x0 -- Sprite 0xb2
      12'hB21: dout  = 8'b00000001; // 2849 :   1 - 0x1
      12'hB22: dout  = 8'b00000001; // 2850 :   1 - 0x1
      12'hB23: dout  = 8'b00000001; // 2851 :   1 - 0x1
      12'hB24: dout  = 8'b00000001; // 2852 :   1 - 0x1
      12'hB25: dout  = 8'b00000000; // 2853 :   0 - 0x0
      12'hB26: dout  = 8'b00000000; // 2854 :   0 - 0x0
      12'hB27: dout  = 8'b00001000; // 2855 :   8 - 0x8
      12'hB28: dout  = 8'b00000000; // 2856 :   0 - 0x0 -- plane 1
      12'hB29: dout  = 8'b00001101; // 2857 :  13 - 0xd
      12'hB2A: dout  = 8'b00011110; // 2858 :  30 - 0x1e
      12'hB2B: dout  = 8'b00011110; // 2859 :  30 - 0x1e
      12'hB2C: dout  = 8'b00011110; // 2860 :  30 - 0x1e
      12'hB2D: dout  = 8'b00011111; // 2861 :  31 - 0x1f
      12'hB2E: dout  = 8'b00001111; // 2862 :  15 - 0xf
      12'hB2F: dout  = 8'b00000111; // 2863 :   7 - 0x7
      12'hB30: dout  = 8'b01111000; // 2864 : 120 - 0x78 -- Sprite 0xb3
      12'hB31: dout  = 8'b11110000; // 2865 : 240 - 0xf0
      12'hB32: dout  = 8'b11111000; // 2866 : 248 - 0xf8
      12'hB33: dout  = 8'b11100100; // 2867 : 228 - 0xe4
      12'hB34: dout  = 8'b11000000; // 2868 : 192 - 0xc0
      12'hB35: dout  = 8'b11001010; // 2869 : 202 - 0xca
      12'hB36: dout  = 8'b11001010; // 2870 : 202 - 0xca
      12'hB37: dout  = 8'b11000000; // 2871 : 192 - 0xc0
      12'hB38: dout  = 8'b01111000; // 2872 : 120 - 0x78 -- plane 1
      12'hB39: dout  = 8'b11110000; // 2873 : 240 - 0xf0
      12'hB3A: dout  = 8'b00000000; // 2874 :   0 - 0x0
      12'hB3B: dout  = 8'b00011010; // 2875 :  26 - 0x1a
      12'hB3C: dout  = 8'b00111111; // 2876 :  63 - 0x3f
      12'hB3D: dout  = 8'b00110101; // 2877 :  53 - 0x35
      12'hB3E: dout  = 8'b00110101; // 2878 :  53 - 0x35
      12'hB3F: dout  = 8'b00111111; // 2879 :  63 - 0x3f
      12'hB40: dout  = 8'b00001111; // 2880 :  15 - 0xf -- Sprite 0xb4
      12'hB41: dout  = 8'b00011111; // 2881 :  31 - 0x1f
      12'hB42: dout  = 8'b10011111; // 2882 : 159 - 0x9f
      12'hB43: dout  = 8'b11111111; // 2883 : 255 - 0xff
      12'hB44: dout  = 8'b11111111; // 2884 : 255 - 0xff
      12'hB45: dout  = 8'b01111111; // 2885 : 127 - 0x7f
      12'hB46: dout  = 8'b01110100; // 2886 : 116 - 0x74
      12'hB47: dout  = 8'b00100000; // 2887 :  32 - 0x20
      12'hB48: dout  = 8'b00000000; // 2888 :   0 - 0x0 -- plane 1
      12'hB49: dout  = 8'b00000000; // 2889 :   0 - 0x0
      12'hB4A: dout  = 8'b10000000; // 2890 : 128 - 0x80
      12'hB4B: dout  = 8'b11100000; // 2891 : 224 - 0xe0
      12'hB4C: dout  = 8'b11100000; // 2892 : 224 - 0xe0
      12'hB4D: dout  = 8'b01110000; // 2893 : 112 - 0x70
      12'hB4E: dout  = 8'b01110011; // 2894 : 115 - 0x73
      12'hB4F: dout  = 8'b00100001; // 2895 :  33 - 0x21
      12'hB50: dout  = 8'b11100100; // 2896 : 228 - 0xe4 -- Sprite 0xb5
      12'hB51: dout  = 8'b11111111; // 2897 : 255 - 0xff
      12'hB52: dout  = 8'b11111110; // 2898 : 254 - 0xfe
      12'hB53: dout  = 8'b11111100; // 2899 : 252 - 0xfc
      12'hB54: dout  = 8'b10011100; // 2900 : 156 - 0x9c
      12'hB55: dout  = 8'b00011110; // 2901 :  30 - 0x1e
      12'hB56: dout  = 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout  = 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout  = 8'b00011010; // 2904 :  26 - 0x1a -- plane 1
      12'hB59: dout  = 8'b00000111; // 2905 :   7 - 0x7
      12'hB5A: dout  = 8'b00001100; // 2906 :  12 - 0xc
      12'hB5B: dout  = 8'b00011000; // 2907 :  24 - 0x18
      12'hB5C: dout  = 8'b01111000; // 2908 : 120 - 0x78
      12'hB5D: dout  = 8'b11111110; // 2909 : 254 - 0xfe
      12'hB5E: dout  = 8'b11111100; // 2910 : 252 - 0xfc
      12'hB5F: dout  = 8'b11110000; // 2911 : 240 - 0xf0
      12'hB60: dout  = 8'b00000000; // 2912 :   0 - 0x0 -- Sprite 0xb6
      12'hB61: dout  = 8'b00000001; // 2913 :   1 - 0x1
      12'hB62: dout  = 8'b00000011; // 2914 :   3 - 0x3
      12'hB63: dout  = 8'b00000011; // 2915 :   3 - 0x3
      12'hB64: dout  = 8'b00000111; // 2916 :   7 - 0x7
      12'hB65: dout  = 8'b00000011; // 2917 :   3 - 0x3
      12'hB66: dout  = 8'b00000001; // 2918 :   1 - 0x1
      12'hB67: dout  = 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout  = 8'b00000000; // 2920 :   0 - 0x0 -- plane 1
      12'hB69: dout  = 8'b00000001; // 2921 :   1 - 0x1
      12'hB6A: dout  = 8'b00000010; // 2922 :   2 - 0x2
      12'hB6B: dout  = 8'b00000000; // 2923 :   0 - 0x0
      12'hB6C: dout  = 8'b00111000; // 2924 :  56 - 0x38
      12'hB6D: dout  = 8'b01111100; // 2925 : 124 - 0x7c
      12'hB6E: dout  = 8'b01111110; // 2926 : 126 - 0x7e
      12'hB6F: dout  = 8'b00111111; // 2927 :  63 - 0x3f
      12'hB70: dout  = 8'b00000000; // 2928 :   0 - 0x0 -- Sprite 0xb7
      12'hB71: dout  = 8'b01011111; // 2929 :  95 - 0x5f
      12'hB72: dout  = 8'b01111111; // 2930 : 127 - 0x7f
      12'hB73: dout  = 8'b01111111; // 2931 : 127 - 0x7f
      12'hB74: dout  = 8'b00111111; // 2932 :  63 - 0x3f
      12'hB75: dout  = 8'b00111111; // 2933 :  63 - 0x3f
      12'hB76: dout  = 8'b00010100; // 2934 :  20 - 0x14
      12'hB77: dout  = 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout  = 8'b00111111; // 2936 :  63 - 0x3f -- plane 1
      12'hB79: dout  = 8'b01000000; // 2937 :  64 - 0x40
      12'hB7A: dout  = 8'b01100000; // 2938 :  96 - 0x60
      12'hB7B: dout  = 8'b01100000; // 2939 :  96 - 0x60
      12'hB7C: dout  = 8'b00100000; // 2940 :  32 - 0x20
      12'hB7D: dout  = 8'b00110000; // 2941 :  48 - 0x30
      12'hB7E: dout  = 8'b00010011; // 2942 :  19 - 0x13
      12'hB7F: dout  = 8'b00000001; // 2943 :   1 - 0x1
      12'hB80: dout  = 8'b11000000; // 2944 : 192 - 0xc0 -- Sprite 0xb8
      12'hB81: dout  = 8'b11100000; // 2945 : 224 - 0xe0
      12'hB82: dout  = 8'b11110000; // 2946 : 240 - 0xf0
      12'hB83: dout  = 8'b00110000; // 2947 :  48 - 0x30
      12'hB84: dout  = 8'b00111000; // 2948 :  56 - 0x38
      12'hB85: dout  = 8'b00111100; // 2949 :  60 - 0x3c
      12'hB86: dout  = 8'b00111100; // 2950 :  60 - 0x3c
      12'hB87: dout  = 8'b11111100; // 2951 : 252 - 0xfc
      12'hB88: dout  = 8'b11000000; // 2952 : 192 - 0xc0 -- plane 1
      12'hB89: dout  = 8'b11100000; // 2953 : 224 - 0xe0
      12'hB8A: dout  = 8'b00110000; // 2954 :  48 - 0x30
      12'hB8B: dout  = 8'b11010000; // 2955 : 208 - 0xd0
      12'hB8C: dout  = 8'b11010000; // 2956 : 208 - 0xd0
      12'hB8D: dout  = 8'b11010000; // 2957 : 208 - 0xd0
      12'hB8E: dout  = 8'b11010000; // 2958 : 208 - 0xd0
      12'hB8F: dout  = 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout  = 8'b00000111; // 2960 :   7 - 0x7 -- Sprite 0xb9
      12'hB91: dout  = 8'b00001111; // 2961 :  15 - 0xf
      12'hB92: dout  = 8'b00011111; // 2962 :  31 - 0x1f
      12'hB93: dout  = 8'b00100010; // 2963 :  34 - 0x22
      12'hB94: dout  = 8'b00100000; // 2964 :  32 - 0x20
      12'hB95: dout  = 8'b00100101; // 2965 :  37 - 0x25
      12'hB96: dout  = 8'b00100101; // 2966 :  37 - 0x25
      12'hB97: dout  = 8'b00011111; // 2967 :  31 - 0x1f
      12'hB98: dout  = 8'b00000111; // 2968 :   7 - 0x7 -- plane 1
      12'hB99: dout  = 8'b00001111; // 2969 :  15 - 0xf
      12'hB9A: dout  = 8'b00000010; // 2970 :   2 - 0x2
      12'hB9B: dout  = 8'b00011101; // 2971 :  29 - 0x1d
      12'hB9C: dout  = 8'b00011111; // 2972 :  31 - 0x1f
      12'hB9D: dout  = 8'b00011010; // 2973 :  26 - 0x1a
      12'hB9E: dout  = 8'b00011010; // 2974 :  26 - 0x1a
      12'hB9F: dout  = 8'b00000010; // 2975 :   2 - 0x2
      12'hBA0: dout  = 8'b11111110; // 2976 : 254 - 0xfe -- Sprite 0xba
      12'hBA1: dout  = 8'b11111110; // 2977 : 254 - 0xfe
      12'hBA2: dout  = 8'b01111110; // 2978 : 126 - 0x7e
      12'hBA3: dout  = 8'b00111010; // 2979 :  58 - 0x3a
      12'hBA4: dout  = 8'b00000010; // 2980 :   2 - 0x2
      12'hBA5: dout  = 8'b00000001; // 2981 :   1 - 0x1
      12'hBA6: dout  = 8'b01000001; // 2982 :  65 - 0x41
      12'hBA7: dout  = 8'b01000001; // 2983 :  65 - 0x41
      12'hBA8: dout  = 8'b00111000; // 2984 :  56 - 0x38 -- plane 1
      12'hBA9: dout  = 8'b01111100; // 2985 : 124 - 0x7c
      12'hBAA: dout  = 8'b11111100; // 2986 : 252 - 0xfc
      12'hBAB: dout  = 8'b11111100; // 2987 : 252 - 0xfc
      12'hBAC: dout  = 8'b11111100; // 2988 : 252 - 0xfc
      12'hBAD: dout  = 8'b11111110; // 2989 : 254 - 0xfe
      12'hBAE: dout  = 8'b10111110; // 2990 : 190 - 0xbe
      12'hBAF: dout  = 8'b10111110; // 2991 : 190 - 0xbe
      12'hBB0: dout  = 8'b00011111; // 2992 :  31 - 0x1f -- Sprite 0xbb
      12'hBB1: dout  = 8'b00111111; // 2993 :  63 - 0x3f
      12'hBB2: dout  = 8'b01111110; // 2994 : 126 - 0x7e
      12'hBB3: dout  = 8'b01011100; // 2995 :  92 - 0x5c
      12'hBB4: dout  = 8'b01000000; // 2996 :  64 - 0x40
      12'hBB5: dout  = 8'b10000000; // 2997 : 128 - 0x80
      12'hBB6: dout  = 8'b10000010; // 2998 : 130 - 0x82
      12'hBB7: dout  = 8'b10000010; // 2999 : 130 - 0x82
      12'hBB8: dout  = 8'b00011100; // 3000 :  28 - 0x1c -- plane 1
      12'hBB9: dout  = 8'b00111110; // 3001 :  62 - 0x3e
      12'hBBA: dout  = 8'b00111111; // 3002 :  63 - 0x3f
      12'hBBB: dout  = 8'b00111111; // 3003 :  63 - 0x3f
      12'hBBC: dout  = 8'b00111111; // 3004 :  63 - 0x3f
      12'hBBD: dout  = 8'b01111111; // 3005 : 127 - 0x7f
      12'hBBE: dout  = 8'b01111101; // 3006 : 125 - 0x7d
      12'hBBF: dout  = 8'b01111101; // 3007 : 125 - 0x7d
      12'hBC0: dout  = 8'b10000010; // 3008 : 130 - 0x82 -- Sprite 0xbc
      12'hBC1: dout  = 8'b10000000; // 3009 : 128 - 0x80
      12'hBC2: dout  = 8'b10100000; // 3010 : 160 - 0xa0
      12'hBC3: dout  = 8'b01000100; // 3011 :  68 - 0x44
      12'hBC4: dout  = 8'b01000011; // 3012 :  67 - 0x43
      12'hBC5: dout  = 8'b01000000; // 3013 :  64 - 0x40
      12'hBC6: dout  = 8'b00100001; // 3014 :  33 - 0x21
      12'hBC7: dout  = 8'b00011110; // 3015 :  30 - 0x1e
      12'hBC8: dout  = 8'b01111101; // 3016 : 125 - 0x7d -- plane 1
      12'hBC9: dout  = 8'b01111111; // 3017 : 127 - 0x7f
      12'hBCA: dout  = 8'b01011111; // 3018 :  95 - 0x5f
      12'hBCB: dout  = 8'b00111011; // 3019 :  59 - 0x3b
      12'hBCC: dout  = 8'b00111100; // 3020 :  60 - 0x3c
      12'hBCD: dout  = 8'b00111111; // 3021 :  63 - 0x3f
      12'hBCE: dout  = 8'b00011110; // 3022 :  30 - 0x1e
      12'hBCF: dout  = 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout  = 8'b00011100; // 3024 :  28 - 0x1c -- Sprite 0xbd
      12'hBD1: dout  = 8'b00111111; // 3025 :  63 - 0x3f
      12'hBD2: dout  = 8'b00111110; // 3026 :  62 - 0x3e
      12'hBD3: dout  = 8'b00111100; // 3027 :  60 - 0x3c
      12'hBD4: dout  = 8'b01000000; // 3028 :  64 - 0x40
      12'hBD5: dout  = 8'b10000000; // 3029 : 128 - 0x80
      12'hBD6: dout  = 8'b10000010; // 3030 : 130 - 0x82
      12'hBD7: dout  = 8'b10000010; // 3031 : 130 - 0x82
      12'hBD8: dout  = 8'b00011100; // 3032 :  28 - 0x1c -- plane 1
      12'hBD9: dout  = 8'b00111110; // 3033 :  62 - 0x3e
      12'hBDA: dout  = 8'b00111111; // 3034 :  63 - 0x3f
      12'hBDB: dout  = 8'b00011111; // 3035 :  31 - 0x1f
      12'hBDC: dout  = 8'b00111111; // 3036 :  63 - 0x3f
      12'hBDD: dout  = 8'b01111111; // 3037 : 127 - 0x7f
      12'hBDE: dout  = 8'b01111101; // 3038 : 125 - 0x7d
      12'hBDF: dout  = 8'b01111101; // 3039 : 125 - 0x7d
      12'hBE0: dout  = 8'b00000000; // 3040 :   0 - 0x0 -- Sprite 0xbe
      12'hBE1: dout  = 8'b00000000; // 3041 :   0 - 0x0
      12'hBE2: dout  = 8'b10000000; // 3042 : 128 - 0x80
      12'hBE3: dout  = 8'b10000000; // 3043 : 128 - 0x80
      12'hBE4: dout  = 8'b10010010; // 3044 : 146 - 0x92
      12'hBE5: dout  = 8'b10011101; // 3045 : 157 - 0x9d
      12'hBE6: dout  = 8'b11000111; // 3046 : 199 - 0xc7
      12'hBE7: dout  = 8'b11101111; // 3047 : 239 - 0xef
      12'hBE8: dout  = 8'b00000000; // 3048 :   0 - 0x0 -- plane 1
      12'hBE9: dout  = 8'b00000000; // 3049 :   0 - 0x0
      12'hBEA: dout  = 8'b00000000; // 3050 :   0 - 0x0
      12'hBEB: dout  = 8'b01100000; // 3051 :  96 - 0x60
      12'hBEC: dout  = 8'b01100010; // 3052 :  98 - 0x62
      12'hBED: dout  = 8'b01100101; // 3053 : 101 - 0x65
      12'hBEE: dout  = 8'b00111111; // 3054 :  63 - 0x3f
      12'hBEF: dout  = 8'b00011111; // 3055 :  31 - 0x1f
      12'hBF0: dout  = 8'b00000000; // 3056 :   0 - 0x0 -- Sprite 0xbf
      12'hBF1: dout  = 8'b00100011; // 3057 :  35 - 0x23
      12'hBF2: dout  = 8'b00110011; // 3058 :  51 - 0x33
      12'hBF3: dout  = 8'b00111111; // 3059 :  63 - 0x3f
      12'hBF4: dout  = 8'b00111111; // 3060 :  63 - 0x3f
      12'hBF5: dout  = 8'b01111111; // 3061 : 127 - 0x7f
      12'hBF6: dout  = 8'b01111111; // 3062 : 127 - 0x7f
      12'hBF7: dout  = 8'b01111111; // 3063 : 127 - 0x7f
      12'hBF8: dout  = 8'b01110000; // 3064 : 112 - 0x70 -- plane 1
      12'hBF9: dout  = 8'b00111100; // 3065 :  60 - 0x3c
      12'hBFA: dout  = 8'b00111100; // 3066 :  60 - 0x3c
      12'hBFB: dout  = 8'b00011000; // 3067 :  24 - 0x18
      12'hBFC: dout  = 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout  = 8'b00000000; // 3069 :   0 - 0x0
      12'hBFE: dout  = 8'b00000010; // 3070 :   2 - 0x2
      12'hBFF: dout  = 8'b00000111; // 3071 :   7 - 0x7
      12'hC00: dout  = 8'b11111110; // 3072 : 254 - 0xfe -- Sprite 0xc0
      12'hC01: dout  = 8'b11111000; // 3073 : 248 - 0xf8
      12'hC02: dout  = 8'b10100000; // 3074 : 160 - 0xa0
      12'hC03: dout  = 8'b00000000; // 3075 :   0 - 0x0
      12'hC04: dout  = 8'b00000000; // 3076 :   0 - 0x0
      12'hC05: dout  = 8'b00000000; // 3077 :   0 - 0x0
      12'hC06: dout  = 8'b10000000; // 3078 : 128 - 0x80
      12'hC07: dout  = 8'b10000000; // 3079 : 128 - 0x80
      12'hC08: dout  = 8'b11001111; // 3080 : 207 - 0xcf -- plane 1
      12'hC09: dout  = 8'b01111010; // 3081 : 122 - 0x7a
      12'hC0A: dout  = 8'b01011010; // 3082 :  90 - 0x5a
      12'hC0B: dout  = 8'b00010000; // 3083 :  16 - 0x10
      12'hC0C: dout  = 8'b00000000; // 3084 :   0 - 0x0
      12'hC0D: dout  = 8'b00000000; // 3085 :   0 - 0x0
      12'hC0E: dout  = 8'b11000000; // 3086 : 192 - 0xc0
      12'hC0F: dout  = 8'b10000000; // 3087 : 128 - 0x80
      12'hC10: dout  = 8'b01111110; // 3088 : 126 - 0x7e -- Sprite 0xc1
      12'hC11: dout  = 8'b01111111; // 3089 : 127 - 0x7f
      12'hC12: dout  = 8'b01111101; // 3090 : 125 - 0x7d
      12'hC13: dout  = 8'b00111111; // 3091 :  63 - 0x3f
      12'hC14: dout  = 8'b00011110; // 3092 :  30 - 0x1e
      12'hC15: dout  = 8'b10001111; // 3093 : 143 - 0x8f
      12'hC16: dout  = 8'b10001111; // 3094 : 143 - 0x8f
      12'hC17: dout  = 8'b00011001; // 3095 :  25 - 0x19
      12'hC18: dout  = 8'b10000101; // 3096 : 133 - 0x85 -- plane 1
      12'hC19: dout  = 8'b10000100; // 3097 : 132 - 0x84
      12'hC1A: dout  = 8'b10000110; // 3098 : 134 - 0x86
      12'hC1B: dout  = 8'b11000110; // 3099 : 198 - 0xc6
      12'hC1C: dout  = 8'b11100111; // 3100 : 231 - 0xe7
      12'hC1D: dout  = 8'b01110011; // 3101 : 115 - 0x73
      12'hC1E: dout  = 8'b01110011; // 3102 : 115 - 0x73
      12'hC1F: dout  = 8'b11100001; // 3103 : 225 - 0xe1
      12'hC20: dout  = 8'b11100000; // 3104 : 224 - 0xe0 -- Sprite 0xc2
      12'hC21: dout  = 8'b00001110; // 3105 :  14 - 0xe
      12'hC22: dout  = 8'b01110011; // 3106 : 115 - 0x73
      12'hC23: dout  = 8'b11110011; // 3107 : 243 - 0xf3
      12'hC24: dout  = 8'b11111001; // 3108 : 249 - 0xf9
      12'hC25: dout  = 8'b11111001; // 3109 : 249 - 0xf9
      12'hC26: dout  = 8'b11111000; // 3110 : 248 - 0xf8
      12'hC27: dout  = 8'b01110000; // 3111 : 112 - 0x70
      12'hC28: dout  = 8'b10000000; // 3112 : 128 - 0x80 -- plane 1
      12'hC29: dout  = 8'b01001110; // 3113 :  78 - 0x4e
      12'hC2A: dout  = 8'b01110111; // 3114 : 119 - 0x77
      12'hC2B: dout  = 8'b11110011; // 3115 : 243 - 0xf3
      12'hC2C: dout  = 8'b11111011; // 3116 : 251 - 0xfb
      12'hC2D: dout  = 8'b11111001; // 3117 : 249 - 0xf9
      12'hC2E: dout  = 8'b11111010; // 3118 : 250 - 0xfa
      12'hC2F: dout  = 8'b01111000; // 3119 : 120 - 0x78
      12'hC30: dout  = 8'b00001110; // 3120 :  14 - 0xe -- Sprite 0xc3
      12'hC31: dout  = 8'b01100110; // 3121 : 102 - 0x66
      12'hC32: dout  = 8'b11100010; // 3122 : 226 - 0xe2
      12'hC33: dout  = 8'b11110110; // 3123 : 246 - 0xf6
      12'hC34: dout  = 8'b11111111; // 3124 : 255 - 0xff
      12'hC35: dout  = 8'b11111111; // 3125 : 255 - 0xff
      12'hC36: dout  = 8'b00011111; // 3126 :  31 - 0x1f
      12'hC37: dout  = 8'b10011000; // 3127 : 152 - 0x98
      12'hC38: dout  = 8'b00010001; // 3128 :  17 - 0x11 -- plane 1
      12'hC39: dout  = 8'b00111001; // 3129 :  57 - 0x39
      12'hC3A: dout  = 8'b01111101; // 3130 : 125 - 0x7d
      12'hC3B: dout  = 8'b00111001; // 3131 :  57 - 0x39
      12'hC3C: dout  = 8'b00000000; // 3132 :   0 - 0x0
      12'hC3D: dout  = 8'b00000000; // 3133 :   0 - 0x0
      12'hC3E: dout  = 8'b11100000; // 3134 : 224 - 0xe0
      12'hC3F: dout  = 8'b11100111; // 3135 : 231 - 0xe7
      12'hC40: dout  = 8'b00000000; // 3136 :   0 - 0x0 -- Sprite 0xc4
      12'hC41: dout  = 8'b00000000; // 3137 :   0 - 0x0
      12'hC42: dout  = 8'b00000000; // 3138 :   0 - 0x0
      12'hC43: dout  = 8'b00000100; // 3139 :   4 - 0x4
      12'hC44: dout  = 8'b00001111; // 3140 :  15 - 0xf
      12'hC45: dout  = 8'b00001111; // 3141 :  15 - 0xf
      12'hC46: dout  = 8'b00011111; // 3142 :  31 - 0x1f
      12'hC47: dout  = 8'b00000111; // 3143 :   7 - 0x7
      12'hC48: dout  = 8'b00000000; // 3144 :   0 - 0x0 -- plane 1
      12'hC49: dout  = 8'b00000000; // 3145 :   0 - 0x0
      12'hC4A: dout  = 8'b00000111; // 3146 :   7 - 0x7
      12'hC4B: dout  = 8'b00000111; // 3147 :   7 - 0x7
      12'hC4C: dout  = 8'b00010110; // 3148 :  22 - 0x16
      12'hC4D: dout  = 8'b00010000; // 3149 :  16 - 0x10
      12'hC4E: dout  = 8'b00000000; // 3150 :   0 - 0x0
      12'hC4F: dout  = 8'b00111000; // 3151 :  56 - 0x38
      12'hC50: dout  = 8'b11110011; // 3152 : 243 - 0xf3 -- Sprite 0xc5
      12'hC51: dout  = 8'b11100111; // 3153 : 231 - 0xe7
      12'hC52: dout  = 8'b11101110; // 3154 : 238 - 0xee
      12'hC53: dout  = 8'b11101100; // 3155 : 236 - 0xec
      12'hC54: dout  = 8'b11001101; // 3156 : 205 - 0xcd
      12'hC55: dout  = 8'b11001111; // 3157 : 207 - 0xcf
      12'hC56: dout  = 8'b11001111; // 3158 : 207 - 0xcf
      12'hC57: dout  = 8'b11011111; // 3159 : 223 - 0xdf
      12'hC58: dout  = 8'b11001111; // 3160 : 207 - 0xcf -- plane 1
      12'hC59: dout  = 8'b00011111; // 3161 :  31 - 0x1f
      12'hC5A: dout  = 8'b00010111; // 3162 :  23 - 0x17
      12'hC5B: dout  = 8'b00010000; // 3163 :  16 - 0x10
      12'hC5C: dout  = 8'b00110011; // 3164 :  51 - 0x33
      12'hC5D: dout  = 8'b00110000; // 3165 :  48 - 0x30
      12'hC5E: dout  = 8'b00110000; // 3166 :  48 - 0x30
      12'hC5F: dout  = 8'b00100000; // 3167 :  32 - 0x20
      12'hC60: dout  = 8'b00100111; // 3168 :  39 - 0x27 -- Sprite 0xc6
      12'hC61: dout  = 8'b00111111; // 3169 :  63 - 0x3f
      12'hC62: dout  = 8'b00111111; // 3170 :  63 - 0x3f
      12'hC63: dout  = 8'b01111000; // 3171 : 120 - 0x78
      12'hC64: dout  = 8'b00111100; // 3172 :  60 - 0x3c
      12'hC65: dout  = 8'b00011111; // 3173 :  31 - 0x1f
      12'hC66: dout  = 8'b00011111; // 3174 :  31 - 0x1f
      12'hC67: dout  = 8'b01110011; // 3175 : 115 - 0x73
      12'hC68: dout  = 8'b00111000; // 3176 :  56 - 0x38 -- plane 1
      12'hC69: dout  = 8'b00110000; // 3177 :  48 - 0x30
      12'hC6A: dout  = 8'b01000000; // 3178 :  64 - 0x40
      12'hC6B: dout  = 8'b11000111; // 3179 : 199 - 0xc7
      12'hC6C: dout  = 8'b00000111; // 3180 :   7 - 0x7
      12'hC6D: dout  = 8'b01100110; // 3181 : 102 - 0x66
      12'hC6E: dout  = 8'b11100000; // 3182 : 224 - 0xe0
      12'hC6F: dout  = 8'b01101100; // 3183 : 108 - 0x6c
      12'hC70: dout  = 8'b10011111; // 3184 : 159 - 0x9f -- Sprite 0xc7
      12'hC71: dout  = 8'b00111110; // 3185 :  62 - 0x3e
      12'hC72: dout  = 8'b01111100; // 3186 : 124 - 0x7c
      12'hC73: dout  = 8'b11111100; // 3187 : 252 - 0xfc
      12'hC74: dout  = 8'b11111000; // 3188 : 248 - 0xf8
      12'hC75: dout  = 8'b11111000; // 3189 : 248 - 0xf8
      12'hC76: dout  = 8'b11000000; // 3190 : 192 - 0xc0
      12'hC77: dout  = 8'b01000000; // 3191 :  64 - 0x40
      12'hC78: dout  = 8'b01100000; // 3192 :  96 - 0x60 -- plane 1
      12'hC79: dout  = 8'b11000000; // 3193 : 192 - 0xc0
      12'hC7A: dout  = 8'b10000000; // 3194 : 128 - 0x80
      12'hC7B: dout  = 8'b00000100; // 3195 :   4 - 0x4
      12'hC7C: dout  = 8'b10011110; // 3196 : 158 - 0x9e
      12'hC7D: dout  = 8'b11111111; // 3197 : 255 - 0xff
      12'hC7E: dout  = 8'b11110000; // 3198 : 240 - 0xf0
      12'hC7F: dout  = 8'b11111000; // 3199 : 248 - 0xf8
      12'hC80: dout  = 8'b01111111; // 3200 : 127 - 0x7f -- Sprite 0xc8
      12'hC81: dout  = 8'b01111110; // 3201 : 126 - 0x7e
      12'hC82: dout  = 8'b01111000; // 3202 : 120 - 0x78
      12'hC83: dout  = 8'b00000001; // 3203 :   1 - 0x1
      12'hC84: dout  = 8'b00000111; // 3204 :   7 - 0x7
      12'hC85: dout  = 8'b00011111; // 3205 :  31 - 0x1f
      12'hC86: dout  = 8'b00111100; // 3206 :  60 - 0x3c
      12'hC87: dout  = 8'b01111100; // 3207 : 124 - 0x7c
      12'hC88: dout  = 8'b00100100; // 3208 :  36 - 0x24 -- plane 1
      12'hC89: dout  = 8'b00000001; // 3209 :   1 - 0x1
      12'hC8A: dout  = 8'b00000111; // 3210 :   7 - 0x7
      12'hC8B: dout  = 8'b11111110; // 3211 : 254 - 0xfe
      12'hC8C: dout  = 8'b11111111; // 3212 : 255 - 0xff
      12'hC8D: dout  = 8'b01111111; // 3213 : 127 - 0x7f
      12'hC8E: dout  = 8'b00111111; // 3214 :  63 - 0x3f
      12'hC8F: dout  = 8'b01111111; // 3215 : 127 - 0x7f
      12'hC90: dout  = 8'b11111100; // 3216 : 252 - 0xfc -- Sprite 0xc9
      12'hC91: dout  = 8'b11111000; // 3217 : 248 - 0xf8
      12'hC92: dout  = 8'b10100000; // 3218 : 160 - 0xa0
      12'hC93: dout  = 8'b11111110; // 3219 : 254 - 0xfe
      12'hC94: dout  = 8'b11111100; // 3220 : 252 - 0xfc
      12'hC95: dout  = 8'b11110000; // 3221 : 240 - 0xf0
      12'hC96: dout  = 8'b10000000; // 3222 : 128 - 0x80
      12'hC97: dout  = 8'b00000000; // 3223 :   0 - 0x0
      12'hC98: dout  = 8'b11001111; // 3224 : 207 - 0xcf -- plane 1
      12'hC99: dout  = 8'b01111010; // 3225 : 122 - 0x7a
      12'hC9A: dout  = 8'b00001010; // 3226 :  10 - 0xa
      12'hC9B: dout  = 8'b11111110; // 3227 : 254 - 0xfe
      12'hC9C: dout  = 8'b11111100; // 3228 : 252 - 0xfc
      12'hC9D: dout  = 8'b00000000; // 3229 :   0 - 0x0
      12'hC9E: dout  = 8'b00000000; // 3230 :   0 - 0x0
      12'hC9F: dout  = 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout  = 8'b01111110; // 3232 : 126 - 0x7e -- Sprite 0xca
      12'hCA1: dout  = 8'b01111111; // 3233 : 127 - 0x7f
      12'hCA2: dout  = 8'b01111111; // 3234 : 127 - 0x7f
      12'hCA3: dout  = 8'b00111111; // 3235 :  63 - 0x3f
      12'hCA4: dout  = 8'b00011111; // 3236 :  31 - 0x1f
      12'hCA5: dout  = 8'b10001111; // 3237 : 143 - 0x8f
      12'hCA6: dout  = 8'b10001111; // 3238 : 143 - 0x8f
      12'hCA7: dout  = 8'b00011000; // 3239 :  24 - 0x18
      12'hCA8: dout  = 8'b10000101; // 3240 : 133 - 0x85 -- plane 1
      12'hCA9: dout  = 8'b10000110; // 3241 : 134 - 0x86
      12'hCAA: dout  = 8'b10000011; // 3242 : 131 - 0x83
      12'hCAB: dout  = 8'b11000011; // 3243 : 195 - 0xc3
      12'hCAC: dout  = 8'b11100001; // 3244 : 225 - 0xe1
      12'hCAD: dout  = 8'b01110000; // 3245 : 112 - 0x70
      12'hCAE: dout  = 8'b01110000; // 3246 : 112 - 0x70
      12'hCAF: dout  = 8'b11100000; // 3247 : 224 - 0xe0
      12'hCB0: dout  = 8'b10011111; // 3248 : 159 - 0x9f -- Sprite 0xcb
      12'hCB1: dout  = 8'b00111110; // 3249 :  62 - 0x3e
      12'hCB2: dout  = 8'b01111100; // 3250 : 124 - 0x7c
      12'hCB3: dout  = 8'b11111000; // 3251 : 248 - 0xf8
      12'hCB4: dout  = 8'b11111000; // 3252 : 248 - 0xf8
      12'hCB5: dout  = 8'b00111100; // 3253 :  60 - 0x3c
      12'hCB6: dout  = 8'b00011000; // 3254 :  24 - 0x18
      12'hCB7: dout  = 8'b11111000; // 3255 : 248 - 0xf8
      12'hCB8: dout  = 8'b01100000; // 3256 :  96 - 0x60 -- plane 1
      12'hCB9: dout  = 8'b11000000; // 3257 : 192 - 0xc0
      12'hCBA: dout  = 8'b10000000; // 3258 : 128 - 0x80
      12'hCBB: dout  = 8'b00000000; // 3259 :   0 - 0x0
      12'hCBC: dout  = 8'b10011000; // 3260 : 152 - 0x98
      12'hCBD: dout  = 8'b11111100; // 3261 : 252 - 0xfc
      12'hCBE: dout  = 8'b11111110; // 3262 : 254 - 0xfe
      12'hCBF: dout  = 8'b11111111; // 3263 : 255 - 0xff
      12'hCC0: dout  = 8'b01111111; // 3264 : 127 - 0x7f -- Sprite 0xcc
      12'hCC1: dout  = 8'b01111111; // 3265 : 127 - 0x7f
      12'hCC2: dout  = 8'b01111000; // 3266 : 120 - 0x78
      12'hCC3: dout  = 8'b00000001; // 3267 :   1 - 0x1
      12'hCC4: dout  = 8'b00000111; // 3268 :   7 - 0x7
      12'hCC5: dout  = 8'b00010011; // 3269 :  19 - 0x13
      12'hCC6: dout  = 8'b11110001; // 3270 : 241 - 0xf1
      12'hCC7: dout  = 8'b00000011; // 3271 :   3 - 0x3
      12'hCC8: dout  = 8'b00100100; // 3272 :  36 - 0x24 -- plane 1
      12'hCC9: dout  = 8'b00000000; // 3273 :   0 - 0x0
      12'hCCA: dout  = 8'b00000111; // 3274 :   7 - 0x7
      12'hCCB: dout  = 8'b11111110; // 3275 : 254 - 0xfe
      12'hCCC: dout  = 8'b11111111; // 3276 : 255 - 0xff
      12'hCCD: dout  = 8'b01111111; // 3277 : 127 - 0x7f
      12'hCCE: dout  = 8'b11111111; // 3278 : 255 - 0xff
      12'hCCF: dout  = 8'b00000011; // 3279 :   3 - 0x3
      12'hCD0: dout  = 8'b00000000; // 3280 :   0 - 0x0 -- Sprite 0xcd
      12'hCD1: dout  = 8'b00000000; // 3281 :   0 - 0x0
      12'hCD2: dout  = 8'b00011100; // 3282 :  28 - 0x1c
      12'hCD3: dout  = 8'b00011101; // 3283 :  29 - 0x1d
      12'hCD4: dout  = 8'b00011011; // 3284 :  27 - 0x1b
      12'hCD5: dout  = 8'b11000011; // 3285 : 195 - 0xc3
      12'hCD6: dout  = 8'b11100011; // 3286 : 227 - 0xe3
      12'hCD7: dout  = 8'b11100001; // 3287 : 225 - 0xe1
      12'hCD8: dout  = 8'b00000011; // 3288 :   3 - 0x3 -- plane 1
      12'hCD9: dout  = 8'b00001111; // 3289 :  15 - 0xf
      12'hCDA: dout  = 8'b00100011; // 3290 :  35 - 0x23
      12'hCDB: dout  = 8'b01100010; // 3291 :  98 - 0x62
      12'hCDC: dout  = 8'b01100100; // 3292 : 100 - 0x64
      12'hCDD: dout  = 8'b00111100; // 3293 :  60 - 0x3c
      12'hCDE: dout  = 8'b00011100; // 3294 :  28 - 0x1c
      12'hCDF: dout  = 8'b00011110; // 3295 :  30 - 0x1e
      12'hCE0: dout  = 8'b11100000; // 3296 : 224 - 0xe0 -- Sprite 0xce
      12'hCE1: dout  = 8'b11001101; // 3297 : 205 - 0xcd
      12'hCE2: dout  = 8'b00011101; // 3298 :  29 - 0x1d
      12'hCE3: dout  = 8'b01001111; // 3299 :  79 - 0x4f
      12'hCE4: dout  = 8'b11101110; // 3300 : 238 - 0xee
      12'hCE5: dout  = 8'b11111111; // 3301 : 255 - 0xff
      12'hCE6: dout  = 8'b00111111; // 3302 :  63 - 0x3f
      12'hCE7: dout  = 8'b00111111; // 3303 :  63 - 0x3f
      12'hCE8: dout  = 8'b00011111; // 3304 :  31 - 0x1f -- plane 1
      12'hCE9: dout  = 8'b00111101; // 3305 :  61 - 0x3d
      12'hCEA: dout  = 8'b01101101; // 3306 : 109 - 0x6d
      12'hCEB: dout  = 8'b01001111; // 3307 :  79 - 0x4f
      12'hCEC: dout  = 8'b11101110; // 3308 : 238 - 0xee
      12'hCED: dout  = 8'b11110011; // 3309 : 243 - 0xf3
      12'hCEE: dout  = 8'b00100000; // 3310 :  32 - 0x20
      12'hCEF: dout  = 8'b00000011; // 3311 :   3 - 0x3
      12'hCF0: dout  = 8'b00111111; // 3312 :  63 - 0x3f -- Sprite 0xcf
      12'hCF1: dout  = 8'b00111111; // 3313 :  63 - 0x3f
      12'hCF2: dout  = 8'b00000000; // 3314 :   0 - 0x0
      12'hCF3: dout  = 8'b00000000; // 3315 :   0 - 0x0
      12'hCF4: dout  = 8'b01110000; // 3316 : 112 - 0x70
      12'hCF5: dout  = 8'b10111000; // 3317 : 184 - 0xb8
      12'hCF6: dout  = 8'b11111100; // 3318 : 252 - 0xfc
      12'hCF7: dout  = 8'b11111100; // 3319 : 252 - 0xfc
      12'hCF8: dout  = 8'b00000111; // 3320 :   7 - 0x7 -- plane 1
      12'hCF9: dout  = 8'b00000111; // 3321 :   7 - 0x7
      12'hCFA: dout  = 8'b00011111; // 3322 :  31 - 0x1f
      12'hCFB: dout  = 8'b00111111; // 3323 :  63 - 0x3f
      12'hCFC: dout  = 8'b00001111; // 3324 :  15 - 0xf
      12'hCFD: dout  = 8'b01000111; // 3325 :  71 - 0x47
      12'hCFE: dout  = 8'b00000011; // 3326 :   3 - 0x3
      12'hCFF: dout  = 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout  = 8'b00000111; // 3328 :   7 - 0x7 -- Sprite 0xd0
      12'hD01: dout  = 8'b00001111; // 3329 :  15 - 0xf
      12'hD02: dout  = 8'b00011111; // 3330 :  31 - 0x1f
      12'hD03: dout  = 8'b00111111; // 3331 :  63 - 0x3f
      12'hD04: dout  = 8'b00111110; // 3332 :  62 - 0x3e
      12'hD05: dout  = 8'b01111100; // 3333 : 124 - 0x7c
      12'hD06: dout  = 8'b01111000; // 3334 : 120 - 0x78
      12'hD07: dout  = 8'b01111000; // 3335 : 120 - 0x78
      12'hD08: dout  = 8'b00000000; // 3336 :   0 - 0x0 -- plane 1
      12'hD09: dout  = 8'b00000000; // 3337 :   0 - 0x0
      12'hD0A: dout  = 8'b00000011; // 3338 :   3 - 0x3
      12'hD0B: dout  = 8'b00000111; // 3339 :   7 - 0x7
      12'hD0C: dout  = 8'b00001111; // 3340 :  15 - 0xf
      12'hD0D: dout  = 8'b00001111; // 3341 :  15 - 0xf
      12'hD0E: dout  = 8'b00011111; // 3342 :  31 - 0x1f
      12'hD0F: dout  = 8'b00011111; // 3343 :  31 - 0x1f
      12'hD10: dout  = 8'b00111111; // 3344 :  63 - 0x3f -- Sprite 0xd1
      12'hD11: dout  = 8'b01011100; // 3345 :  92 - 0x5c
      12'hD12: dout  = 8'b00111001; // 3346 :  57 - 0x39
      12'hD13: dout  = 8'b00111011; // 3347 :  59 - 0x3b
      12'hD14: dout  = 8'b10111111; // 3348 : 191 - 0xbf
      12'hD15: dout  = 8'b11111111; // 3349 : 255 - 0xff
      12'hD16: dout  = 8'b11111110; // 3350 : 254 - 0xfe
      12'hD17: dout  = 8'b11111110; // 3351 : 254 - 0xfe
      12'hD18: dout  = 8'b00000000; // 3352 :   0 - 0x0 -- plane 1
      12'hD19: dout  = 8'b00100011; // 3353 :  35 - 0x23
      12'hD1A: dout  = 8'b01010111; // 3354 :  87 - 0x57
      12'hD1B: dout  = 8'b01001111; // 3355 :  79 - 0x4f
      12'hD1C: dout  = 8'b01010111; // 3356 :  87 - 0x57
      12'hD1D: dout  = 8'b00101111; // 3357 :  47 - 0x2f
      12'hD1E: dout  = 8'b11011111; // 3358 : 223 - 0xdf
      12'hD1F: dout  = 8'b00100001; // 3359 :  33 - 0x21
      12'hD20: dout  = 8'b11000000; // 3360 : 192 - 0xc0 -- Sprite 0xd2
      12'hD21: dout  = 8'b11000000; // 3361 : 192 - 0xc0
      12'hD22: dout  = 8'b10000000; // 3362 : 128 - 0x80
      12'hD23: dout  = 8'b10000000; // 3363 : 128 - 0x80
      12'hD24: dout  = 8'b10000000; // 3364 : 128 - 0x80
      12'hD25: dout  = 8'b10000000; // 3365 : 128 - 0x80
      12'hD26: dout  = 8'b00000000; // 3366 :   0 - 0x0
      12'hD27: dout  = 8'b00000000; // 3367 :   0 - 0x0
      12'hD28: dout  = 8'b00000000; // 3368 :   0 - 0x0 -- plane 1
      12'hD29: dout  = 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout  = 8'b00000000; // 3370 :   0 - 0x0
      12'hD2B: dout  = 8'b00000000; // 3371 :   0 - 0x0
      12'hD2C: dout  = 8'b10000000; // 3372 : 128 - 0x80
      12'hD2D: dout  = 8'b10000000; // 3373 : 128 - 0x80
      12'hD2E: dout  = 8'b00000000; // 3374 :   0 - 0x0
      12'hD2F: dout  = 8'b00000000; // 3375 :   0 - 0x0
      12'hD30: dout  = 8'b11111110; // 3376 : 254 - 0xfe -- Sprite 0xd3
      12'hD31: dout  = 8'b11111100; // 3377 : 252 - 0xfc
      12'hD32: dout  = 8'b01100001; // 3378 :  97 - 0x61
      12'hD33: dout  = 8'b00001111; // 3379 :  15 - 0xf
      12'hD34: dout  = 8'b01111111; // 3380 : 127 - 0x7f
      12'hD35: dout  = 8'b00111111; // 3381 :  63 - 0x3f
      12'hD36: dout  = 8'b00011111; // 3382 :  31 - 0x1f
      12'hD37: dout  = 8'b00011110; // 3383 :  30 - 0x1e
      12'hD38: dout  = 8'b00100011; // 3384 :  35 - 0x23 -- plane 1
      12'hD39: dout  = 8'b00001111; // 3385 :  15 - 0xf
      12'hD3A: dout  = 8'b00011110; // 3386 :  30 - 0x1e
      12'hD3B: dout  = 8'b11110000; // 3387 : 240 - 0xf0
      12'hD3C: dout  = 8'b00011100; // 3388 :  28 - 0x1c
      12'hD3D: dout  = 8'b00111111; // 3389 :  63 - 0x3f
      12'hD3E: dout  = 8'b00011111; // 3390 :  31 - 0x1f
      12'hD3F: dout  = 8'b00011110; // 3391 :  30 - 0x1e
      12'hD40: dout  = 8'b11110000; // 3392 : 240 - 0xf0 -- Sprite 0xd4
      12'hD41: dout  = 8'b01111000; // 3393 : 120 - 0x78
      12'hD42: dout  = 8'b11100100; // 3394 : 228 - 0xe4
      12'hD43: dout  = 8'b11001000; // 3395 : 200 - 0xc8
      12'hD44: dout  = 8'b11001100; // 3396 : 204 - 0xcc
      12'hD45: dout  = 8'b10111110; // 3397 : 190 - 0xbe
      12'hD46: dout  = 8'b10111110; // 3398 : 190 - 0xbe
      12'hD47: dout  = 8'b00111110; // 3399 :  62 - 0x3e
      12'hD48: dout  = 8'b00000000; // 3400 :   0 - 0x0 -- plane 1
      12'hD49: dout  = 8'b10000000; // 3401 : 128 - 0x80
      12'hD4A: dout  = 8'b00011000; // 3402 :  24 - 0x18
      12'hD4B: dout  = 8'b00110000; // 3403 :  48 - 0x30
      12'hD4C: dout  = 8'b00110100; // 3404 :  52 - 0x34
      12'hD4D: dout  = 8'b11111110; // 3405 : 254 - 0xfe
      12'hD4E: dout  = 8'b11111110; // 3406 : 254 - 0xfe
      12'hD4F: dout  = 8'b11111110; // 3407 : 254 - 0xfe
      12'hD50: dout  = 8'b00000000; // 3408 :   0 - 0x0 -- Sprite 0xd5
      12'hD51: dout  = 8'b00000001; // 3409 :   1 - 0x1
      12'hD52: dout  = 8'b00000000; // 3410 :   0 - 0x0
      12'hD53: dout  = 8'b00000111; // 3411 :   7 - 0x7
      12'hD54: dout  = 8'b00000111; // 3412 :   7 - 0x7
      12'hD55: dout  = 8'b00000111; // 3413 :   7 - 0x7
      12'hD56: dout  = 8'b00000111; // 3414 :   7 - 0x7
      12'hD57: dout  = 8'b00011111; // 3415 :  31 - 0x1f
      12'hD58: dout  = 8'b00000000; // 3416 :   0 - 0x0 -- plane 1
      12'hD59: dout  = 8'b00000000; // 3417 :   0 - 0x0
      12'hD5A: dout  = 8'b00000001; // 3418 :   1 - 0x1
      12'hD5B: dout  = 8'b00000100; // 3419 :   4 - 0x4
      12'hD5C: dout  = 8'b00000110; // 3420 :   6 - 0x6
      12'hD5D: dout  = 8'b00000110; // 3421 :   6 - 0x6
      12'hD5E: dout  = 8'b00000111; // 3422 :   7 - 0x7
      12'hD5F: dout  = 8'b00000111; // 3423 :   7 - 0x7
      12'hD60: dout  = 8'b00000000; // 3424 :   0 - 0x0 -- Sprite 0xd6
      12'hD61: dout  = 8'b00000000; // 3425 :   0 - 0x0
      12'hD62: dout  = 8'b00001111; // 3426 :  15 - 0xf
      12'hD63: dout  = 8'b00111111; // 3427 :  63 - 0x3f
      12'hD64: dout  = 8'b00111111; // 3428 :  63 - 0x3f
      12'hD65: dout  = 8'b00001111; // 3429 :  15 - 0xf
      12'hD66: dout  = 8'b00000000; // 3430 :   0 - 0x0
      12'hD67: dout  = 8'b00000000; // 3431 :   0 - 0x0
      12'hD68: dout  = 8'b00001111; // 3432 :  15 - 0xf -- plane 1
      12'hD69: dout  = 8'b00111111; // 3433 :  63 - 0x3f
      12'hD6A: dout  = 8'b01111111; // 3434 : 127 - 0x7f
      12'hD6B: dout  = 8'b11111000; // 3435 : 248 - 0xf8
      12'hD6C: dout  = 8'b11111000; // 3436 : 248 - 0xf8
      12'hD6D: dout  = 8'b01111111; // 3437 : 127 - 0x7f
      12'hD6E: dout  = 8'b00111111; // 3438 :  63 - 0x3f
      12'hD6F: dout  = 8'b00001111; // 3439 :  15 - 0xf
      12'hD70: dout  = 8'b01111000; // 3440 : 120 - 0x78 -- Sprite 0xd7
      12'hD71: dout  = 8'b01111100; // 3441 : 124 - 0x7c
      12'hD72: dout  = 8'b01111110; // 3442 : 126 - 0x7e
      12'hD73: dout  = 8'b01111111; // 3443 : 127 - 0x7f
      12'hD74: dout  = 8'b00111111; // 3444 :  63 - 0x3f
      12'hD75: dout  = 8'b00111111; // 3445 :  63 - 0x3f
      12'hD76: dout  = 8'b00011011; // 3446 :  27 - 0x1b
      12'hD77: dout  = 8'b00001001; // 3447 :   9 - 0x9
      12'hD78: dout  = 8'b00011111; // 3448 :  31 - 0x1f -- plane 1
      12'hD79: dout  = 8'b00011111; // 3449 :  31 - 0x1f
      12'hD7A: dout  = 8'b00011111; // 3450 :  31 - 0x1f
      12'hD7B: dout  = 8'b00001011; // 3451 :  11 - 0xb
      12'hD7C: dout  = 8'b00000001; // 3452 :   1 - 0x1
      12'hD7D: dout  = 8'b00000001; // 3453 :   1 - 0x1
      12'hD7E: dout  = 8'b00000000; // 3454 :   0 - 0x0
      12'hD7F: dout  = 8'b00000000; // 3455 :   0 - 0x0
      12'hD80: dout  = 8'b00001100; // 3456 :  12 - 0xc -- Sprite 0xd8
      12'hD81: dout  = 8'b00000000; // 3457 :   0 - 0x0
      12'hD82: dout  = 8'b00000000; // 3458 :   0 - 0x0
      12'hD83: dout  = 8'b00000000; // 3459 :   0 - 0x0
      12'hD84: dout  = 8'b00000111; // 3460 :   7 - 0x7
      12'hD85: dout  = 8'b01111111; // 3461 : 127 - 0x7f
      12'hD86: dout  = 8'b01111100; // 3462 : 124 - 0x7c
      12'hD87: dout  = 8'b00000000; // 3463 :   0 - 0x0
      12'hD88: dout  = 8'b00000011; // 3464 :   3 - 0x3 -- plane 1
      12'hD89: dout  = 8'b00011111; // 3465 :  31 - 0x1f
      12'hD8A: dout  = 8'b00111111; // 3466 :  63 - 0x3f
      12'hD8B: dout  = 8'b00111111; // 3467 :  63 - 0x3f
      12'hD8C: dout  = 8'b01111000; // 3468 : 120 - 0x78
      12'hD8D: dout  = 8'b00000000; // 3469 :   0 - 0x0
      12'hD8E: dout  = 8'b00000011; // 3470 :   3 - 0x3
      12'hD8F: dout  = 8'b11111111; // 3471 : 255 - 0xff
      12'hD90: dout  = 8'b00000001; // 3472 :   1 - 0x1 -- Sprite 0xd9
      12'hD91: dout  = 8'b11100001; // 3473 : 225 - 0xe1
      12'hD92: dout  = 8'b01110001; // 3474 : 113 - 0x71
      12'hD93: dout  = 8'b01111001; // 3475 : 121 - 0x79
      12'hD94: dout  = 8'b00111101; // 3476 :  61 - 0x3d
      12'hD95: dout  = 8'b00111101; // 3477 :  61 - 0x3d
      12'hD96: dout  = 8'b00011111; // 3478 :  31 - 0x1f
      12'hD97: dout  = 8'b00000011; // 3479 :   3 - 0x3
      12'hD98: dout  = 8'b00000000; // 3480 :   0 - 0x0 -- plane 1
      12'hD99: dout  = 8'b00000000; // 3481 :   0 - 0x0
      12'hD9A: dout  = 8'b00000000; // 3482 :   0 - 0x0
      12'hD9B: dout  = 8'b00000000; // 3483 :   0 - 0x0
      12'hD9C: dout  = 8'b00000000; // 3484 :   0 - 0x0
      12'hD9D: dout  = 8'b00000000; // 3485 :   0 - 0x0
      12'hD9E: dout  = 8'b00000000; // 3486 :   0 - 0x0
      12'hD9F: dout  = 8'b00000000; // 3487 :   0 - 0x0
      12'hDA0: dout  = 8'b00111111; // 3488 :  63 - 0x3f -- Sprite 0xda
      12'hDA1: dout  = 8'b00111111; // 3489 :  63 - 0x3f
      12'hDA2: dout  = 8'b00011111; // 3490 :  31 - 0x1f
      12'hDA3: dout  = 8'b00011011; // 3491 :  27 - 0x1b
      12'hDA4: dout  = 8'b00110110; // 3492 :  54 - 0x36
      12'hDA5: dout  = 8'b00110000; // 3493 :  48 - 0x30
      12'hDA6: dout  = 8'b01111111; // 3494 : 127 - 0x7f
      12'hDA7: dout  = 8'b00111111; // 3495 :  63 - 0x3f
      12'hDA8: dout  = 8'b00100011; // 3496 :  35 - 0x23 -- plane 1
      12'hDA9: dout  = 8'b00100111; // 3497 :  39 - 0x27
      12'hDAA: dout  = 8'b00011111; // 3498 :  31 - 0x1f
      12'hDAB: dout  = 8'b00000111; // 3499 :   7 - 0x7
      12'hDAC: dout  = 8'b00001111; // 3500 :  15 - 0xf
      12'hDAD: dout  = 8'b00011111; // 3501 :  31 - 0x1f
      12'hDAE: dout  = 8'b01111111; // 3502 : 127 - 0x7f
      12'hDAF: dout  = 8'b00111111; // 3503 :  63 - 0x3f
      12'hDB0: dout  = 8'b11111000; // 3504 : 248 - 0xf8 -- Sprite 0xdb
      12'hDB1: dout  = 8'b11111000; // 3505 : 248 - 0xf8
      12'hDB2: dout  = 8'b11111000; // 3506 : 248 - 0xf8
      12'hDB3: dout  = 8'b10111000; // 3507 : 184 - 0xb8
      12'hDB4: dout  = 8'b00011000; // 3508 :  24 - 0x18
      12'hDB5: dout  = 8'b11011000; // 3509 : 216 - 0xd8
      12'hDB6: dout  = 8'b11011000; // 3510 : 216 - 0xd8
      12'hDB7: dout  = 8'b10111000; // 3511 : 184 - 0xb8
      12'hDB8: dout  = 8'b11100000; // 3512 : 224 - 0xe0 -- plane 1
      12'hDB9: dout  = 8'b10000000; // 3513 : 128 - 0x80
      12'hDBA: dout  = 8'b10000000; // 3514 : 128 - 0x80
      12'hDBB: dout  = 8'b01000000; // 3515 :  64 - 0x40
      12'hDBC: dout  = 8'b11100000; // 3516 : 224 - 0xe0
      12'hDBD: dout  = 8'b11100000; // 3517 : 224 - 0xe0
      12'hDBE: dout  = 8'b11100000; // 3518 : 224 - 0xe0
      12'hDBF: dout  = 8'b11000000; // 3519 : 192 - 0xc0
      12'hDC0: dout  = 8'b00000001; // 3520 :   1 - 0x1 -- Sprite 0xdc
      12'hDC1: dout  = 8'b00000010; // 3521 :   2 - 0x2
      12'hDC2: dout  = 8'b00000100; // 3522 :   4 - 0x4
      12'hDC3: dout  = 8'b00000100; // 3523 :   4 - 0x4
      12'hDC4: dout  = 8'b00001000; // 3524 :   8 - 0x8
      12'hDC5: dout  = 8'b00001000; // 3525 :   8 - 0x8
      12'hDC6: dout  = 8'b00010000; // 3526 :  16 - 0x10
      12'hDC7: dout  = 8'b00010000; // 3527 :  16 - 0x10
      12'hDC8: dout  = 8'b00000011; // 3528 :   3 - 0x3 -- plane 1
      12'hDC9: dout  = 8'b00000111; // 3529 :   7 - 0x7
      12'hDCA: dout  = 8'b00001111; // 3530 :  15 - 0xf
      12'hDCB: dout  = 8'b00011111; // 3531 :  31 - 0x1f
      12'hDCC: dout  = 8'b00111111; // 3532 :  63 - 0x3f
      12'hDCD: dout  = 8'b01111111; // 3533 : 127 - 0x7f
      12'hDCE: dout  = 8'b11111111; // 3534 : 255 - 0xff
      12'hDCF: dout  = 8'b00011111; // 3535 :  31 - 0x1f
      12'hDD0: dout  = 8'b00000000; // 3536 :   0 - 0x0 -- Sprite 0xdd
      12'hDD1: dout  = 8'b00001111; // 3537 :  15 - 0xf
      12'hDD2: dout  = 8'b00010011; // 3538 :  19 - 0x13
      12'hDD3: dout  = 8'b00001101; // 3539 :  13 - 0xd
      12'hDD4: dout  = 8'b00001101; // 3540 :  13 - 0xd
      12'hDD5: dout  = 8'b00010011; // 3541 :  19 - 0x13
      12'hDD6: dout  = 8'b00001100; // 3542 :  12 - 0xc
      12'hDD7: dout  = 8'b00100000; // 3543 :  32 - 0x20
      12'hDD8: dout  = 8'b00011111; // 3544 :  31 - 0x1f -- plane 1
      12'hDD9: dout  = 8'b00010000; // 3545 :  16 - 0x10
      12'hDDA: dout  = 8'b00001100; // 3546 :  12 - 0xc
      12'hDDB: dout  = 8'b00010010; // 3547 :  18 - 0x12
      12'hDDC: dout  = 8'b00010010; // 3548 :  18 - 0x12
      12'hDDD: dout  = 8'b00101100; // 3549 :  44 - 0x2c
      12'hDDE: dout  = 8'b00111111; // 3550 :  63 - 0x3f
      12'hDDF: dout  = 8'b00111111; // 3551 :  63 - 0x3f
      12'hDE0: dout  = 8'b00000000; // 3552 :   0 - 0x0 -- Sprite 0xde
      12'hDE1: dout  = 8'b00100100; // 3553 :  36 - 0x24
      12'hDE2: dout  = 8'b00000000; // 3554 :   0 - 0x0
      12'hDE3: dout  = 8'b00100100; // 3555 :  36 - 0x24
      12'hDE4: dout  = 8'b00000000; // 3556 :   0 - 0x0
      12'hDE5: dout  = 8'b00000100; // 3557 :   4 - 0x4
      12'hDE6: dout  = 8'b00000000; // 3558 :   0 - 0x0
      12'hDE7: dout  = 8'b00000000; // 3559 :   0 - 0x0
      12'hDE8: dout  = 8'b00110111; // 3560 :  55 - 0x37 -- plane 1
      12'hDE9: dout  = 8'b00110110; // 3561 :  54 - 0x36
      12'hDEA: dout  = 8'b00110110; // 3562 :  54 - 0x36
      12'hDEB: dout  = 8'b00110110; // 3563 :  54 - 0x36
      12'hDEC: dout  = 8'b00010110; // 3564 :  22 - 0x16
      12'hDED: dout  = 8'b00010110; // 3565 :  22 - 0x16
      12'hDEE: dout  = 8'b00010010; // 3566 :  18 - 0x12
      12'hDEF: dout  = 8'b00000010; // 3567 :   2 - 0x2
      12'hDF0: dout  = 8'b00001111; // 3568 :  15 - 0xf -- Sprite 0xdf
      12'hDF1: dout  = 8'b01000001; // 3569 :  65 - 0x41
      12'hDF2: dout  = 8'b00000000; // 3570 :   0 - 0x0
      12'hDF3: dout  = 8'b10001000; // 3571 : 136 - 0x88
      12'hDF4: dout  = 8'b00000000; // 3572 :   0 - 0x0
      12'hDF5: dout  = 8'b01000100; // 3573 :  68 - 0x44
      12'hDF6: dout  = 8'b00000000; // 3574 :   0 - 0x0
      12'hDF7: dout  = 8'b00000000; // 3575 :   0 - 0x0
      12'hDF8: dout  = 8'b00010000; // 3576 :  16 - 0x10 -- plane 1
      12'hDF9: dout  = 8'b01111110; // 3577 : 126 - 0x7e
      12'hDFA: dout  = 8'b11111111; // 3578 : 255 - 0xff
      12'hDFB: dout  = 8'b11111111; // 3579 : 255 - 0xff
      12'hDFC: dout  = 8'b11110110; // 3580 : 246 - 0xf6
      12'hDFD: dout  = 8'b01110110; // 3581 : 118 - 0x76
      12'hDFE: dout  = 8'b00111010; // 3582 :  58 - 0x3a
      12'hDFF: dout  = 8'b00011010; // 3583 :  26 - 0x1a
      12'hE00: dout  = 8'b00111000; // 3584 :  56 - 0x38 -- Sprite 0xe0
      12'hE01: dout  = 8'b01111100; // 3585 : 124 - 0x7c
      12'hE02: dout  = 8'b11111110; // 3586 : 254 - 0xfe
      12'hE03: dout  = 8'b11111110; // 3587 : 254 - 0xfe
      12'hE04: dout  = 8'b00111011; // 3588 :  59 - 0x3b
      12'hE05: dout  = 8'b00000011; // 3589 :   3 - 0x3
      12'hE06: dout  = 8'b00000011; // 3590 :   3 - 0x3
      12'hE07: dout  = 8'b00000011; // 3591 :   3 - 0x3
      12'hE08: dout  = 8'b00000000; // 3592 :   0 - 0x0 -- plane 1
      12'hE09: dout  = 8'b00000000; // 3593 :   0 - 0x0
      12'hE0A: dout  = 8'b00111000; // 3594 :  56 - 0x38
      12'hE0B: dout  = 8'b00000100; // 3595 :   4 - 0x4
      12'hE0C: dout  = 8'b00000000; // 3596 :   0 - 0x0
      12'hE0D: dout  = 8'b00000000; // 3597 :   0 - 0x0
      12'hE0E: dout  = 8'b00000000; // 3598 :   0 - 0x0
      12'hE0F: dout  = 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout  = 8'b00000011; // 3600 :   3 - 0x3 -- Sprite 0xe1
      12'hE11: dout  = 8'b00110011; // 3601 :  51 - 0x33
      12'hE12: dout  = 8'b01111011; // 3602 : 123 - 0x7b
      12'hE13: dout  = 8'b01111111; // 3603 : 127 - 0x7f
      12'hE14: dout  = 8'b11111111; // 3604 : 255 - 0xff
      12'hE15: dout  = 8'b11111011; // 3605 : 251 - 0xfb
      12'hE16: dout  = 8'b00000011; // 3606 :   3 - 0x3
      12'hE17: dout  = 8'b00000011; // 3607 :   3 - 0x3
      12'hE18: dout  = 8'b00000000; // 3608 :   0 - 0x0 -- plane 1
      12'hE19: dout  = 8'b00000000; // 3609 :   0 - 0x0
      12'hE1A: dout  = 8'b00000000; // 3610 :   0 - 0x0
      12'hE1B: dout  = 8'b00111000; // 3611 :  56 - 0x38
      12'hE1C: dout  = 8'b01000000; // 3612 :  64 - 0x40
      12'hE1D: dout  = 8'b00000000; // 3613 :   0 - 0x0
      12'hE1E: dout  = 8'b00000000; // 3614 :   0 - 0x0
      12'hE1F: dout  = 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout  = 8'b11011100; // 3616 : 220 - 0xdc -- Sprite 0xe2
      12'hE21: dout  = 8'b11000000; // 3617 : 192 - 0xc0
      12'hE22: dout  = 8'b11100000; // 3618 : 224 - 0xe0
      12'hE23: dout  = 8'b11100000; // 3619 : 224 - 0xe0
      12'hE24: dout  = 8'b11100000; // 3620 : 224 - 0xe0
      12'hE25: dout  = 8'b11100000; // 3621 : 224 - 0xe0
      12'hE26: dout  = 8'b11100000; // 3622 : 224 - 0xe0
      12'hE27: dout  = 8'b11000000; // 3623 : 192 - 0xc0
      12'hE28: dout  = 8'b11111100; // 3624 : 252 - 0xfc -- plane 1
      12'hE29: dout  = 8'b10100000; // 3625 : 160 - 0xa0
      12'hE2A: dout  = 8'b10000000; // 3626 : 128 - 0x80
      12'hE2B: dout  = 8'b10000000; // 3627 : 128 - 0x80
      12'hE2C: dout  = 8'b00000000; // 3628 :   0 - 0x0
      12'hE2D: dout  = 8'b00000000; // 3629 :   0 - 0x0
      12'hE2E: dout  = 8'b00000000; // 3630 :   0 - 0x0
      12'hE2F: dout  = 8'b00000000; // 3631 :   0 - 0x0
      12'hE30: dout  = 8'b00111111; // 3632 :  63 - 0x3f -- Sprite 0xe3
      12'hE31: dout  = 8'b01011111; // 3633 :  95 - 0x5f
      12'hE32: dout  = 8'b00111111; // 3634 :  63 - 0x3f
      12'hE33: dout  = 8'b00111111; // 3635 :  63 - 0x3f
      12'hE34: dout  = 8'b10111011; // 3636 : 187 - 0xbb
      12'hE35: dout  = 8'b11111000; // 3637 : 248 - 0xf8
      12'hE36: dout  = 8'b11111110; // 3638 : 254 - 0xfe
      12'hE37: dout  = 8'b11111110; // 3639 : 254 - 0xfe
      12'hE38: dout  = 8'b00000111; // 3640 :   7 - 0x7 -- plane 1
      12'hE39: dout  = 8'b00100111; // 3641 :  39 - 0x27
      12'hE3A: dout  = 8'b01010111; // 3642 :  87 - 0x57
      12'hE3B: dout  = 8'b01001111; // 3643 :  79 - 0x4f
      12'hE3C: dout  = 8'b01010111; // 3644 :  87 - 0x57
      12'hE3D: dout  = 8'b00100111; // 3645 :  39 - 0x27
      12'hE3E: dout  = 8'b11000001; // 3646 : 193 - 0xc1
      12'hE3F: dout  = 8'b00100001; // 3647 :  33 - 0x21
      12'hE40: dout  = 8'b00011111; // 3648 :  31 - 0x1f -- Sprite 0xe4
      12'hE41: dout  = 8'b00001111; // 3649 :  15 - 0xf
      12'hE42: dout  = 8'b00001111; // 3650 :  15 - 0xf
      12'hE43: dout  = 8'b00011111; // 3651 :  31 - 0x1f
      12'hE44: dout  = 8'b00011111; // 3652 :  31 - 0x1f
      12'hE45: dout  = 8'b00011110; // 3653 :  30 - 0x1e
      12'hE46: dout  = 8'b00111000; // 3654 :  56 - 0x38
      12'hE47: dout  = 8'b00110000; // 3655 :  48 - 0x30
      12'hE48: dout  = 8'b00011101; // 3656 :  29 - 0x1d -- plane 1
      12'hE49: dout  = 8'b00001111; // 3657 :  15 - 0xf
      12'hE4A: dout  = 8'b00001111; // 3658 :  15 - 0xf
      12'hE4B: dout  = 8'b00011111; // 3659 :  31 - 0x1f
      12'hE4C: dout  = 8'b00011111; // 3660 :  31 - 0x1f
      12'hE4D: dout  = 8'b00011110; // 3661 :  30 - 0x1e
      12'hE4E: dout  = 8'b00111000; // 3662 :  56 - 0x38
      12'hE4F: dout  = 8'b00110000; // 3663 :  48 - 0x30
      12'hE50: dout  = 8'b00000000; // 3664 :   0 - 0x0 -- Sprite 0xe5
      12'hE51: dout  = 8'b00100000; // 3665 :  32 - 0x20
      12'hE52: dout  = 8'b01100000; // 3666 :  96 - 0x60
      12'hE53: dout  = 8'b01100000; // 3667 :  96 - 0x60
      12'hE54: dout  = 8'b01110000; // 3668 : 112 - 0x70
      12'hE55: dout  = 8'b11110000; // 3669 : 240 - 0xf0
      12'hE56: dout  = 8'b11111000; // 3670 : 248 - 0xf8
      12'hE57: dout  = 8'b11111000; // 3671 : 248 - 0xf8
      12'hE58: dout  = 8'b00000000; // 3672 :   0 - 0x0 -- plane 1
      12'hE59: dout  = 8'b00000000; // 3673 :   0 - 0x0
      12'hE5A: dout  = 8'b00111000; // 3674 :  56 - 0x38
      12'hE5B: dout  = 8'b00010000; // 3675 :  16 - 0x10
      12'hE5C: dout  = 8'b01001100; // 3676 :  76 - 0x4c
      12'hE5D: dout  = 8'b00011000; // 3677 :  24 - 0x18
      12'hE5E: dout  = 8'b10000110; // 3678 : 134 - 0x86
      12'hE5F: dout  = 8'b00100100; // 3679 :  36 - 0x24
      12'hE60: dout  = 8'b11111000; // 3680 : 248 - 0xf8 -- Sprite 0xe6
      12'hE61: dout  = 8'b11111100; // 3681 : 252 - 0xfc
      12'hE62: dout  = 8'b11111100; // 3682 : 252 - 0xfc
      12'hE63: dout  = 8'b01111110; // 3683 : 126 - 0x7e
      12'hE64: dout  = 8'b01111110; // 3684 : 126 - 0x7e
      12'hE65: dout  = 8'b00111110; // 3685 :  62 - 0x3e
      12'hE66: dout  = 8'b00011111; // 3686 :  31 - 0x1f
      12'hE67: dout  = 8'b00000111; // 3687 :   7 - 0x7
      12'hE68: dout  = 8'b00000000; // 3688 :   0 - 0x0 -- plane 1
      12'hE69: dout  = 8'b01000010; // 3689 :  66 - 0x42
      12'hE6A: dout  = 8'b00001010; // 3690 :  10 - 0xa
      12'hE6B: dout  = 8'b01000000; // 3691 :  64 - 0x40
      12'hE6C: dout  = 8'b00010000; // 3692 :  16 - 0x10
      12'hE6D: dout  = 8'b00000010; // 3693 :   2 - 0x2
      12'hE6E: dout  = 8'b00001000; // 3694 :   8 - 0x8
      12'hE6F: dout  = 8'b00000010; // 3695 :   2 - 0x2
      12'hE70: dout  = 8'b00000000; // 3696 :   0 - 0x0 -- Sprite 0xe7
      12'hE71: dout  = 8'b11000000; // 3697 : 192 - 0xc0
      12'hE72: dout  = 8'b01110000; // 3698 : 112 - 0x70
      12'hE73: dout  = 8'b10111000; // 3699 : 184 - 0xb8
      12'hE74: dout  = 8'b11110100; // 3700 : 244 - 0xf4
      12'hE75: dout  = 8'b11110010; // 3701 : 242 - 0xf2
      12'hE76: dout  = 8'b11110101; // 3702 : 245 - 0xf5
      12'hE77: dout  = 8'b01111011; // 3703 : 123 - 0x7b
      12'hE78: dout  = 8'b00000000; // 3704 :   0 - 0x0 -- plane 1
      12'hE79: dout  = 8'b00000000; // 3705 :   0 - 0x0
      12'hE7A: dout  = 8'b10000000; // 3706 : 128 - 0x80
      12'hE7B: dout  = 8'b01000000; // 3707 :  64 - 0x40
      12'hE7C: dout  = 8'b00001000; // 3708 :   8 - 0x8
      12'hE7D: dout  = 8'b00001100; // 3709 :  12 - 0xc
      12'hE7E: dout  = 8'b00001010; // 3710 :  10 - 0xa
      12'hE7F: dout  = 8'b10000100; // 3711 : 132 - 0x84
      12'hE80: dout  = 8'b00000000; // 3712 :   0 - 0x0 -- Sprite 0xe8
      12'hE81: dout  = 8'b11011111; // 3713 : 223 - 0xdf
      12'hE82: dout  = 8'b00010000; // 3714 :  16 - 0x10
      12'hE83: dout  = 8'b11111111; // 3715 : 255 - 0xff
      12'hE84: dout  = 8'b11011111; // 3716 : 223 - 0xdf
      12'hE85: dout  = 8'b11111111; // 3717 : 255 - 0xff
      12'hE86: dout  = 8'b11111111; // 3718 : 255 - 0xff
      12'hE87: dout  = 8'b11111001; // 3719 : 249 - 0xf9
      12'hE88: dout  = 8'b00000000; // 3720 :   0 - 0x0 -- plane 1
      12'hE89: dout  = 8'b00000000; // 3721 :   0 - 0x0
      12'hE8A: dout  = 8'b11001111; // 3722 : 207 - 0xcf
      12'hE8B: dout  = 8'b00100000; // 3723 :  32 - 0x20
      12'hE8C: dout  = 8'b00100000; // 3724 :  32 - 0x20
      12'hE8D: dout  = 8'b00100000; // 3725 :  32 - 0x20
      12'hE8E: dout  = 8'b00100110; // 3726 :  38 - 0x26
      12'hE8F: dout  = 8'b00101110; // 3727 :  46 - 0x2e
      12'hE90: dout  = 8'b00011111; // 3728 :  31 - 0x1f -- Sprite 0xe9
      12'hE91: dout  = 8'b00011111; // 3729 :  31 - 0x1f
      12'hE92: dout  = 8'b00111110; // 3730 :  62 - 0x3e
      12'hE93: dout  = 8'b11111100; // 3731 : 252 - 0xfc
      12'hE94: dout  = 8'b11111000; // 3732 : 248 - 0xf8
      12'hE95: dout  = 8'b11110000; // 3733 : 240 - 0xf0
      12'hE96: dout  = 8'b11000000; // 3734 : 192 - 0xc0
      12'hE97: dout  = 8'b00000000; // 3735 :   0 - 0x0
      12'hE98: dout  = 8'b11100000; // 3736 : 224 - 0xe0 -- plane 1
      12'hE99: dout  = 8'b11100000; // 3737 : 224 - 0xe0
      12'hE9A: dout  = 8'b11000000; // 3738 : 192 - 0xc0
      12'hE9B: dout  = 8'b00000000; // 3739 :   0 - 0x0
      12'hE9C: dout  = 8'b00000000; // 3740 :   0 - 0x0
      12'hE9D: dout  = 8'b00000000; // 3741 :   0 - 0x0
      12'hE9E: dout  = 8'b00000000; // 3742 :   0 - 0x0
      12'hE9F: dout  = 8'b00000000; // 3743 :   0 - 0x0
      12'hEA0: dout  = 8'b11111000; // 3744 : 248 - 0xf8 -- Sprite 0xea
      12'hEA1: dout  = 8'b11111100; // 3745 : 252 - 0xfc
      12'hEA2: dout  = 8'b11111110; // 3746 : 254 - 0xfe
      12'hEA3: dout  = 8'b11111111; // 3747 : 255 - 0xff
      12'hEA4: dout  = 8'b11111111; // 3748 : 255 - 0xff
      12'hEA5: dout  = 8'b11011111; // 3749 : 223 - 0xdf
      12'hEA6: dout  = 8'b11011111; // 3750 : 223 - 0xdf
      12'hEA7: dout  = 8'b00000000; // 3751 :   0 - 0x0
      12'hEA8: dout  = 8'b00101111; // 3752 :  47 - 0x2f -- plane 1
      12'hEA9: dout  = 8'b00100011; // 3753 :  35 - 0x23
      12'hEAA: dout  = 8'b00100001; // 3754 :  33 - 0x21
      12'hEAB: dout  = 8'b00100000; // 3755 :  32 - 0x20
      12'hEAC: dout  = 8'b00100000; // 3756 :  32 - 0x20
      12'hEAD: dout  = 8'b00000000; // 3757 :   0 - 0x0
      12'hEAE: dout  = 8'b00000000; // 3758 :   0 - 0x0
      12'hEAF: dout  = 8'b00000000; // 3759 :   0 - 0x0
      12'hEB0: dout  = 8'b11000001; // 3760 : 193 - 0xc1 -- Sprite 0xeb
      12'hEB1: dout  = 8'b11110001; // 3761 : 241 - 0xf1
      12'hEB2: dout  = 8'b01111001; // 3762 : 121 - 0x79
      12'hEB3: dout  = 8'b01111101; // 3763 : 125 - 0x7d
      12'hEB4: dout  = 8'b00111101; // 3764 :  61 - 0x3d
      12'hEB5: dout  = 8'b00111111; // 3765 :  63 - 0x3f
      12'hEB6: dout  = 8'b00011111; // 3766 :  31 - 0x1f
      12'hEB7: dout  = 8'b00000011; // 3767 :   3 - 0x3
      12'hEB8: dout  = 8'b11000001; // 3768 : 193 - 0xc1 -- plane 1
      12'hEB9: dout  = 8'b10110001; // 3769 : 177 - 0xb1
      12'hEBA: dout  = 8'b01011001; // 3770 :  89 - 0x59
      12'hEBB: dout  = 8'b01101101; // 3771 : 109 - 0x6d
      12'hEBC: dout  = 8'b00110101; // 3772 :  53 - 0x35
      12'hEBD: dout  = 8'b00111011; // 3773 :  59 - 0x3b
      12'hEBE: dout  = 8'b00011111; // 3774 :  31 - 0x1f
      12'hEBF: dout  = 8'b00000011; // 3775 :   3 - 0x3
      12'hEC0: dout  = 8'b00000010; // 3776 :   2 - 0x2 -- Sprite 0xec
      12'hEC1: dout  = 8'b00000110; // 3777 :   6 - 0x6
      12'hEC2: dout  = 8'b00001110; // 3778 :  14 - 0xe
      12'hEC3: dout  = 8'b00001110; // 3779 :  14 - 0xe
      12'hEC4: dout  = 8'b00011110; // 3780 :  30 - 0x1e
      12'hEC5: dout  = 8'b00011110; // 3781 :  30 - 0x1e
      12'hEC6: dout  = 8'b00111110; // 3782 :  62 - 0x3e
      12'hEC7: dout  = 8'b00111110; // 3783 :  62 - 0x3e
      12'hEC8: dout  = 8'b00000000; // 3784 :   0 - 0x0 -- plane 1
      12'hEC9: dout  = 8'b00000010; // 3785 :   2 - 0x2
      12'hECA: dout  = 8'b00000000; // 3786 :   0 - 0x0
      12'hECB: dout  = 8'b00001000; // 3787 :   8 - 0x8
      12'hECC: dout  = 8'b00000010; // 3788 :   2 - 0x2
      12'hECD: dout  = 8'b00000000; // 3789 :   0 - 0x0
      12'hECE: dout  = 8'b00101000; // 3790 :  40 - 0x28
      12'hECF: dout  = 8'b00000000; // 3791 :   0 - 0x0
      12'hED0: dout  = 8'b00111110; // 3792 :  62 - 0x3e -- Sprite 0xed
      12'hED1: dout  = 8'b00111110; // 3793 :  62 - 0x3e
      12'hED2: dout  = 8'b00111110; // 3794 :  62 - 0x3e
      12'hED3: dout  = 8'b00111110; // 3795 :  62 - 0x3e
      12'hED4: dout  = 8'b00011110; // 3796 :  30 - 0x1e
      12'hED5: dout  = 8'b00011110; // 3797 :  30 - 0x1e
      12'hED6: dout  = 8'b00001110; // 3798 :  14 - 0xe
      12'hED7: dout  = 8'b00000010; // 3799 :   2 - 0x2
      12'hED8: dout  = 8'b00000100; // 3800 :   4 - 0x4 -- plane 1
      12'hED9: dout  = 8'b00010000; // 3801 :  16 - 0x10
      12'hEDA: dout  = 8'b00000010; // 3802 :   2 - 0x2
      12'hEDB: dout  = 8'b00010000; // 3803 :  16 - 0x10
      12'hEDC: dout  = 8'b00000100; // 3804 :   4 - 0x4
      12'hEDD: dout  = 8'b00000000; // 3805 :   0 - 0x0
      12'hEDE: dout  = 8'b00001010; // 3806 :  10 - 0xa
      12'hEDF: dout  = 8'b00000000; // 3807 :   0 - 0x0
      12'hEE0: dout  = 8'b11000001; // 3808 : 193 - 0xc1 -- Sprite 0xee
      12'hEE1: dout  = 8'b11110001; // 3809 : 241 - 0xf1
      12'hEE2: dout  = 8'b01111001; // 3810 : 121 - 0x79
      12'hEE3: dout  = 8'b01111101; // 3811 : 125 - 0x7d
      12'hEE4: dout  = 8'b00111101; // 3812 :  61 - 0x3d
      12'hEE5: dout  = 8'b00111111; // 3813 :  63 - 0x3f
      12'hEE6: dout  = 8'b00011111; // 3814 :  31 - 0x1f
      12'hEE7: dout  = 8'b00000011; // 3815 :   3 - 0x3
      12'hEE8: dout  = 8'b11000001; // 3816 : 193 - 0xc1 -- plane 1
      12'hEE9: dout  = 8'b10110001; // 3817 : 177 - 0xb1
      12'hEEA: dout  = 8'b01011001; // 3818 :  89 - 0x59
      12'hEEB: dout  = 8'b01101101; // 3819 : 109 - 0x6d
      12'hEEC: dout  = 8'b00110101; // 3820 :  53 - 0x35
      12'hEED: dout  = 8'b00111011; // 3821 :  59 - 0x3b
      12'hEEE: dout  = 8'b00011111; // 3822 :  31 - 0x1f
      12'hEEF: dout  = 8'b00000011; // 3823 :   3 - 0x3
      12'hEF0: dout  = 8'b01111100; // 3824 : 124 - 0x7c -- Sprite 0xef
      12'hEF1: dout  = 8'b00000000; // 3825 :   0 - 0x0
      12'hEF2: dout  = 8'b00000000; // 3826 :   0 - 0x0
      12'hEF3: dout  = 8'b11111111; // 3827 : 255 - 0xff
      12'hEF4: dout  = 8'b11000011; // 3828 : 195 - 0xc3
      12'hEF5: dout  = 8'b01111111; // 3829 : 127 - 0x7f
      12'hEF6: dout  = 8'b00011111; // 3830 :  31 - 0x1f
      12'hEF7: dout  = 8'b00000011; // 3831 :   3 - 0x3
      12'hEF8: dout  = 8'b00000000; // 3832 :   0 - 0x0 -- plane 1
      12'hEF9: dout  = 8'b00001111; // 3833 :  15 - 0xf
      12'hEFA: dout  = 8'b00011111; // 3834 :  31 - 0x1f
      12'hEFB: dout  = 8'b11111111; // 3835 : 255 - 0xff
      12'hEFC: dout  = 8'b11111100; // 3836 : 252 - 0xfc
      12'hEFD: dout  = 8'b01100011; // 3837 :  99 - 0x63
      12'hEFE: dout  = 8'b00011111; // 3838 :  31 - 0x1f
      12'hEFF: dout  = 8'b00000011; // 3839 :   3 - 0x3
      12'hF00: dout  = 8'b11111111; // 3840 : 255 - 0xff -- Sprite 0xf0
      12'hF01: dout  = 8'b11111111; // 3841 : 255 - 0xff
      12'hF02: dout  = 8'b01111100; // 3842 : 124 - 0x7c
      12'hF03: dout  = 8'b00000000; // 3843 :   0 - 0x0
      12'hF04: dout  = 8'b00000000; // 3844 :   0 - 0x0
      12'hF05: dout  = 8'b01111100; // 3845 : 124 - 0x7c
      12'hF06: dout  = 8'b11111111; // 3846 : 255 - 0xff
      12'hF07: dout  = 8'b11111111; // 3847 : 255 - 0xff
      12'hF08: dout  = 8'b00000000; // 3848 :   0 - 0x0 -- plane 1
      12'hF09: dout  = 8'b00000000; // 3849 :   0 - 0x0
      12'hF0A: dout  = 8'b11111110; // 3850 : 254 - 0xfe
      12'hF0B: dout  = 8'b11000110; // 3851 : 198 - 0xc6
      12'hF0C: dout  = 8'b11000110; // 3852 : 198 - 0xc6
      12'hF0D: dout  = 8'b11111110; // 3853 : 254 - 0xfe
      12'hF0E: dout  = 8'b00000000; // 3854 :   0 - 0x0
      12'hF0F: dout  = 8'b00000000; // 3855 :   0 - 0x0
      12'hF10: dout  = 8'b11111111; // 3856 : 255 - 0xff -- Sprite 0xf1
      12'hF11: dout  = 8'b11111111; // 3857 : 255 - 0xff
      12'hF12: dout  = 8'b00000000; // 3858 :   0 - 0x0
      12'hF13: dout  = 8'b00000100; // 3859 :   4 - 0x4
      12'hF14: dout  = 8'b00001100; // 3860 :  12 - 0xc
      12'hF15: dout  = 8'b00011000; // 3861 :  24 - 0x18
      12'hF16: dout  = 8'b00110000; // 3862 :  48 - 0x30
      12'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout  = 8'b00000000; // 3864 :   0 - 0x0 -- plane 1
      12'hF19: dout  = 8'b00000000; // 3865 :   0 - 0x0
      12'hF1A: dout  = 8'b00000110; // 3866 :   6 - 0x6
      12'hF1B: dout  = 8'b00000110; // 3867 :   6 - 0x6
      12'hF1C: dout  = 8'b00001100; // 3868 :  12 - 0xc
      12'hF1D: dout  = 8'b00011000; // 3869 :  24 - 0x18
      12'hF1E: dout  = 8'b01110000; // 3870 : 112 - 0x70
      12'hF1F: dout  = 8'b01100000; // 3871 :  96 - 0x60
      12'hF20: dout  = 8'b11111111; // 3872 : 255 - 0xff -- Sprite 0xf2
      12'hF21: dout  = 8'b11111111; // 3873 : 255 - 0xff
      12'hF22: dout  = 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout  = 8'b00000100; // 3875 :   4 - 0x4
      12'hF24: dout  = 8'b00000100; // 3876 :   4 - 0x4
      12'hF25: dout  = 8'b00000100; // 3877 :   4 - 0x4
      12'hF26: dout  = 8'b00001000; // 3878 :   8 - 0x8
      12'hF27: dout  = 8'b00001000; // 3879 :   8 - 0x8
      12'hF28: dout  = 8'b00000000; // 3880 :   0 - 0x0 -- plane 1
      12'hF29: dout  = 8'b00000000; // 3881 :   0 - 0x0
      12'hF2A: dout  = 8'b00000110; // 3882 :   6 - 0x6
      12'hF2B: dout  = 8'b00000110; // 3883 :   6 - 0x6
      12'hF2C: dout  = 8'b00000100; // 3884 :   4 - 0x4
      12'hF2D: dout  = 8'b00000100; // 3885 :   4 - 0x4
      12'hF2E: dout  = 8'b00001000; // 3886 :   8 - 0x8
      12'hF2F: dout  = 8'b00001000; // 3887 :   8 - 0x8
      12'hF30: dout  = 8'b00001000; // 3888 :   8 - 0x8 -- Sprite 0xf3
      12'hF31: dout  = 8'b00010000; // 3889 :  16 - 0x10
      12'hF32: dout  = 8'b00010000; // 3890 :  16 - 0x10
      12'hF33: dout  = 8'b00000000; // 3891 :   0 - 0x0
      12'hF34: dout  = 8'b00000000; // 3892 :   0 - 0x0
      12'hF35: dout  = 8'b00010000; // 3893 :  16 - 0x10
      12'hF36: dout  = 8'b00010000; // 3894 :  16 - 0x10
      12'hF37: dout  = 8'b00001000; // 3895 :   8 - 0x8
      12'hF38: dout  = 8'b00001000; // 3896 :   8 - 0x8 -- plane 1
      12'hF39: dout  = 8'b00010000; // 3897 :  16 - 0x10
      12'hF3A: dout  = 8'b00110000; // 3898 :  48 - 0x30
      12'hF3B: dout  = 8'b00110000; // 3899 :  48 - 0x30
      12'hF3C: dout  = 8'b00110000; // 3900 :  48 - 0x30
      12'hF3D: dout  = 8'b00110000; // 3901 :  48 - 0x30
      12'hF3E: dout  = 8'b00010000; // 3902 :  16 - 0x10
      12'hF3F: dout  = 8'b00001000; // 3903 :   8 - 0x8
      12'hF40: dout  = 8'b01111111; // 3904 : 127 - 0x7f -- Sprite 0xf4
      12'hF41: dout  = 8'b00111111; // 3905 :  63 - 0x3f
      12'hF42: dout  = 8'b00111111; // 3906 :  63 - 0x3f
      12'hF43: dout  = 8'b00111110; // 3907 :  62 - 0x3e
      12'hF44: dout  = 8'b00011111; // 3908 :  31 - 0x1f
      12'hF45: dout  = 8'b00001111; // 3909 :  15 - 0xf
      12'hF46: dout  = 8'b00000011; // 3910 :   3 - 0x3
      12'hF47: dout  = 8'b00000000; // 3911 :   0 - 0x0
      12'hF48: dout  = 8'b00000000; // 3912 :   0 - 0x0 -- plane 1
      12'hF49: dout  = 8'b00000000; // 3913 :   0 - 0x0
      12'hF4A: dout  = 8'b00000001; // 3914 :   1 - 0x1
      12'hF4B: dout  = 8'b00000011; // 3915 :   3 - 0x3
      12'hF4C: dout  = 8'b00000001; // 3916 :   1 - 0x1
      12'hF4D: dout  = 8'b00000000; // 3917 :   0 - 0x0
      12'hF4E: dout  = 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout  = 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout  = 8'b00000011; // 3920 :   3 - 0x3 -- Sprite 0xf5
      12'hF51: dout  = 8'b00001111; // 3921 :  15 - 0xf
      12'hF52: dout  = 8'b11111111; // 3922 : 255 - 0xff
      12'hF53: dout  = 8'b01111111; // 3923 : 127 - 0x7f
      12'hF54: dout  = 8'b01111111; // 3924 : 127 - 0x7f
      12'hF55: dout  = 8'b01111111; // 3925 : 127 - 0x7f
      12'hF56: dout  = 8'b01111111; // 3926 : 127 - 0x7f
      12'hF57: dout  = 8'b01111111; // 3927 : 127 - 0x7f
      12'hF58: dout  = 8'b00000011; // 3928 :   3 - 0x3 -- plane 1
      12'hF59: dout  = 8'b00001110; // 3929 :  14 - 0xe
      12'hF5A: dout  = 8'b11111000; // 3930 : 248 - 0xf8
      12'hF5B: dout  = 8'b00000000; // 3931 :   0 - 0x0
      12'hF5C: dout  = 8'b00000000; // 3932 :   0 - 0x0
      12'hF5D: dout  = 8'b00000000; // 3933 :   0 - 0x0
      12'hF5E: dout  = 8'b00000000; // 3934 :   0 - 0x0
      12'hF5F: dout  = 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout  = 8'b00000000; // 3936 :   0 - 0x0 -- Sprite 0xf6
      12'hF61: dout  = 8'b00000000; // 3937 :   0 - 0x0
      12'hF62: dout  = 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout  = 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout  = 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout  = 8'b00000000; // 3941 :   0 - 0x0
      12'hF66: dout  = 8'b00000000; // 3942 :   0 - 0x0
      12'hF67: dout  = 8'b00000000; // 3943 :   0 - 0x0
      12'hF68: dout  = 8'b00100010; // 3944 :  34 - 0x22 -- plane 1
      12'hF69: dout  = 8'b01100101; // 3945 : 101 - 0x65
      12'hF6A: dout  = 8'b00100101; // 3946 :  37 - 0x25
      12'hF6B: dout  = 8'b00100101; // 3947 :  37 - 0x25
      12'hF6C: dout  = 8'b00100101; // 3948 :  37 - 0x25
      12'hF6D: dout  = 8'b00100101; // 3949 :  37 - 0x25
      12'hF6E: dout  = 8'b01110111; // 3950 : 119 - 0x77
      12'hF6F: dout  = 8'b01110010; // 3951 : 114 - 0x72
      12'hF70: dout  = 8'b00000000; // 3952 :   0 - 0x0 -- Sprite 0xf7
      12'hF71: dout  = 8'b00000000; // 3953 :   0 - 0x0
      12'hF72: dout  = 8'b00000000; // 3954 :   0 - 0x0
      12'hF73: dout  = 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout  = 8'b00000000; // 3956 :   0 - 0x0
      12'hF75: dout  = 8'b00000000; // 3957 :   0 - 0x0
      12'hF76: dout  = 8'b00000000; // 3958 :   0 - 0x0
      12'hF77: dout  = 8'b00000000; // 3959 :   0 - 0x0
      12'hF78: dout  = 8'b01100010; // 3960 :  98 - 0x62 -- plane 1
      12'hF79: dout  = 8'b10010101; // 3961 : 149 - 0x95
      12'hF7A: dout  = 8'b00010101; // 3962 :  21 - 0x15
      12'hF7B: dout  = 8'b00100101; // 3963 :  37 - 0x25
      12'hF7C: dout  = 8'b01000101; // 3964 :  69 - 0x45
      12'hF7D: dout  = 8'b10000101; // 3965 : 133 - 0x85
      12'hF7E: dout  = 8'b11110111; // 3966 : 247 - 0xf7
      12'hF7F: dout  = 8'b11110010; // 3967 : 242 - 0xf2
      12'hF80: dout  = 8'b00000000; // 3968 :   0 - 0x0 -- Sprite 0xf8
      12'hF81: dout  = 8'b00000000; // 3969 :   0 - 0x0
      12'hF82: dout  = 8'b00000000; // 3970 :   0 - 0x0
      12'hF83: dout  = 8'b00000000; // 3971 :   0 - 0x0
      12'hF84: dout  = 8'b00000000; // 3972 :   0 - 0x0
      12'hF85: dout  = 8'b00000000; // 3973 :   0 - 0x0
      12'hF86: dout  = 8'b00000000; // 3974 :   0 - 0x0
      12'hF87: dout  = 8'b00000000; // 3975 :   0 - 0x0
      12'hF88: dout  = 8'b10100010; // 3976 : 162 - 0xa2 -- plane 1
      12'hF89: dout  = 8'b10100101; // 3977 : 165 - 0xa5
      12'hF8A: dout  = 8'b10100101; // 3978 : 165 - 0xa5
      12'hF8B: dout  = 8'b10100101; // 3979 : 165 - 0xa5
      12'hF8C: dout  = 8'b11110101; // 3980 : 245 - 0xf5
      12'hF8D: dout  = 8'b11110101; // 3981 : 245 - 0xf5
      12'hF8E: dout  = 8'b00100111; // 3982 :  39 - 0x27
      12'hF8F: dout  = 8'b00100010; // 3983 :  34 - 0x22
      12'hF90: dout  = 8'b00000000; // 3984 :   0 - 0x0 -- Sprite 0xf9
      12'hF91: dout  = 8'b00000000; // 3985 :   0 - 0x0
      12'hF92: dout  = 8'b00000000; // 3986 :   0 - 0x0
      12'hF93: dout  = 8'b00000000; // 3987 :   0 - 0x0
      12'hF94: dout  = 8'b00000000; // 3988 :   0 - 0x0
      12'hF95: dout  = 8'b00000000; // 3989 :   0 - 0x0
      12'hF96: dout  = 8'b00000000; // 3990 :   0 - 0x0
      12'hF97: dout  = 8'b00000000; // 3991 :   0 - 0x0
      12'hF98: dout  = 8'b11110010; // 3992 : 242 - 0xf2 -- plane 1
      12'hF99: dout  = 8'b10000101; // 3993 : 133 - 0x85
      12'hF9A: dout  = 8'b10000101; // 3994 : 133 - 0x85
      12'hF9B: dout  = 8'b11100101; // 3995 : 229 - 0xe5
      12'hF9C: dout  = 8'b00010101; // 3996 :  21 - 0x15
      12'hF9D: dout  = 8'b00010101; // 3997 :  21 - 0x15
      12'hF9E: dout  = 8'b11110111; // 3998 : 247 - 0xf7
      12'hF9F: dout  = 8'b11100010; // 3999 : 226 - 0xe2
      12'hFA0: dout  = 8'b00000000; // 4000 :   0 - 0x0 -- Sprite 0xfa
      12'hFA1: dout  = 8'b00000000; // 4001 :   0 - 0x0
      12'hFA2: dout  = 8'b00000000; // 4002 :   0 - 0x0
      12'hFA3: dout  = 8'b00000000; // 4003 :   0 - 0x0
      12'hFA4: dout  = 8'b00000000; // 4004 :   0 - 0x0
      12'hFA5: dout  = 8'b00000000; // 4005 :   0 - 0x0
      12'hFA6: dout  = 8'b00000000; // 4006 :   0 - 0x0
      12'hFA7: dout  = 8'b00000000; // 4007 :   0 - 0x0
      12'hFA8: dout  = 8'b01100010; // 4008 :  98 - 0x62 -- plane 1
      12'hFA9: dout  = 8'b10010101; // 4009 : 149 - 0x95
      12'hFAA: dout  = 8'b01010101; // 4010 :  85 - 0x55
      12'hFAB: dout  = 8'b01100101; // 4011 : 101 - 0x65
      12'hFAC: dout  = 8'b10110101; // 4012 : 181 - 0xb5
      12'hFAD: dout  = 8'b10010101; // 4013 : 149 - 0x95
      12'hFAE: dout  = 8'b10010111; // 4014 : 151 - 0x97
      12'hFAF: dout  = 8'b01100010; // 4015 :  98 - 0x62
      12'hFB0: dout  = 8'b00000000; // 4016 :   0 - 0x0 -- Sprite 0xfb
      12'hFB1: dout  = 8'b00000000; // 4017 :   0 - 0x0
      12'hFB2: dout  = 8'b00000000; // 4018 :   0 - 0x0
      12'hFB3: dout  = 8'b00000000; // 4019 :   0 - 0x0
      12'hFB4: dout  = 8'b00000000; // 4020 :   0 - 0x0
      12'hFB5: dout  = 8'b00000000; // 4021 :   0 - 0x0
      12'hFB6: dout  = 8'b00000000; // 4022 :   0 - 0x0
      12'hFB7: dout  = 8'b00000000; // 4023 :   0 - 0x0
      12'hFB8: dout  = 8'b00100000; // 4024 :  32 - 0x20 -- plane 1
      12'hFB9: dout  = 8'b01010000; // 4025 :  80 - 0x50
      12'hFBA: dout  = 8'b01010000; // 4026 :  80 - 0x50
      12'hFBB: dout  = 8'b01010000; // 4027 :  80 - 0x50
      12'hFBC: dout  = 8'b01010000; // 4028 :  80 - 0x50
      12'hFBD: dout  = 8'b01010000; // 4029 :  80 - 0x50
      12'hFBE: dout  = 8'b01110000; // 4030 : 112 - 0x70
      12'hFBF: dout  = 8'b00100000; // 4031 :  32 - 0x20
      12'hFC0: dout  = 8'b00000000; // 4032 :   0 - 0x0 -- Sprite 0xfc
      12'hFC1: dout  = 8'b00000000; // 4033 :   0 - 0x0
      12'hFC2: dout  = 8'b00000000; // 4034 :   0 - 0x0
      12'hFC3: dout  = 8'b00000000; // 4035 :   0 - 0x0
      12'hFC4: dout  = 8'b00000000; // 4036 :   0 - 0x0
      12'hFC5: dout  = 8'b00000000; // 4037 :   0 - 0x0
      12'hFC6: dout  = 8'b00000000; // 4038 :   0 - 0x0
      12'hFC7: dout  = 8'b00000000; // 4039 :   0 - 0x0
      12'hFC8: dout  = 8'b00000000; // 4040 :   0 - 0x0 -- plane 1
      12'hFC9: dout  = 8'b00000000; // 4041 :   0 - 0x0
      12'hFCA: dout  = 8'b00000000; // 4042 :   0 - 0x0
      12'hFCB: dout  = 8'b00000000; // 4043 :   0 - 0x0
      12'hFCC: dout  = 8'b00000000; // 4044 :   0 - 0x0
      12'hFCD: dout  = 8'b00000000; // 4045 :   0 - 0x0
      12'hFCE: dout  = 8'b00000000; // 4046 :   0 - 0x0
      12'hFCF: dout  = 8'b00000000; // 4047 :   0 - 0x0
      12'hFD0: dout  = 8'b00000000; // 4048 :   0 - 0x0 -- Sprite 0xfd
      12'hFD1: dout  = 8'b00000000; // 4049 :   0 - 0x0
      12'hFD2: dout  = 8'b00000000; // 4050 :   0 - 0x0
      12'hFD3: dout  = 8'b00000000; // 4051 :   0 - 0x0
      12'hFD4: dout  = 8'b00000000; // 4052 :   0 - 0x0
      12'hFD5: dout  = 8'b00000000; // 4053 :   0 - 0x0
      12'hFD6: dout  = 8'b00000000; // 4054 :   0 - 0x0
      12'hFD7: dout  = 8'b00000000; // 4055 :   0 - 0x0
      12'hFD8: dout  = 8'b01100110; // 4056 : 102 - 0x66 -- plane 1
      12'hFD9: dout  = 8'b11100110; // 4057 : 230 - 0xe6
      12'hFDA: dout  = 8'b01100110; // 4058 : 102 - 0x66
      12'hFDB: dout  = 8'b01100110; // 4059 : 102 - 0x66
      12'hFDC: dout  = 8'b01100110; // 4060 : 102 - 0x66
      12'hFDD: dout  = 8'b01100111; // 4061 : 103 - 0x67
      12'hFDE: dout  = 8'b11110011; // 4062 : 243 - 0xf3
      12'hFDF: dout  = 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout  = 8'b00000000; // 4064 :   0 - 0x0 -- Sprite 0xfe
      12'hFE1: dout  = 8'b00000000; // 4065 :   0 - 0x0
      12'hFE2: dout  = 8'b00000000; // 4066 :   0 - 0x0
      12'hFE3: dout  = 8'b00000000; // 4067 :   0 - 0x0
      12'hFE4: dout  = 8'b00000000; // 4068 :   0 - 0x0
      12'hFE5: dout  = 8'b00000000; // 4069 :   0 - 0x0
      12'hFE6: dout  = 8'b00000000; // 4070 :   0 - 0x0
      12'hFE7: dout  = 8'b00000000; // 4071 :   0 - 0x0
      12'hFE8: dout  = 8'b01011110; // 4072 :  94 - 0x5e -- plane 1
      12'hFE9: dout  = 8'b01011001; // 4073 :  89 - 0x59
      12'hFEA: dout  = 8'b01011001; // 4074 :  89 - 0x59
      12'hFEB: dout  = 8'b01011001; // 4075 :  89 - 0x59
      12'hFEC: dout  = 8'b01011110; // 4076 :  94 - 0x5e
      12'hFED: dout  = 8'b11011000; // 4077 : 216 - 0xd8
      12'hFEE: dout  = 8'b10011000; // 4078 : 152 - 0x98
      12'hFEF: dout  = 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout  = 8'b00000000; // 4080 :   0 - 0x0 -- Sprite 0xff
      12'hFF1: dout  = 8'b00000000; // 4081 :   0 - 0x0
      12'hFF2: dout  = 8'b00000000; // 4082 :   0 - 0x0
      12'hFF3: dout  = 8'b00000000; // 4083 :   0 - 0x0
      12'hFF4: dout  = 8'b00000000; // 4084 :   0 - 0x0
      12'hFF5: dout  = 8'b01111100; // 4085 : 124 - 0x7c
      12'hFF6: dout  = 8'b00111000; // 4086 :  56 - 0x38
      12'hFF7: dout  = 8'b00000000; // 4087 :   0 - 0x0
      12'hFF8: dout  = 8'b00000000; // 4088 :   0 - 0x0 -- plane 1
      12'hFF9: dout  = 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout  = 8'b00000000; // 4090 :   0 - 0x0
      12'hFFB: dout  = 8'b00000000; // 4091 :   0 - 0x0
      12'hFFC: dout  = 8'b00000000; // 4092 :   0 - 0x0
      12'hFFD: dout  = 8'b00000100; // 4093 :   4 - 0x4
      12'hFFE: dout  = 8'b00001000; // 4094 :   8 - 0x8
      12'hFFF: dout  = 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
