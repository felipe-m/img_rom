//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: pacman_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_PACMAN_color0
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout <= 8'b00000000; //    1 :   0 - 0x0
      12'h2: dout <= 8'b00000000; //    2 :   0 - 0x0
      12'h3: dout <= 8'b00000000; //    3 :   0 - 0x0
      12'h4: dout <= 8'b00000000; //    4 :   0 - 0x0
      12'h5: dout <= 8'b00000000; //    5 :   0 - 0x0
      12'h6: dout <= 8'b00000000; //    6 :   0 - 0x0
      12'h7: dout <= 8'b00000000; //    7 :   0 - 0x0
      12'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      12'h9: dout <= 8'b00111000; //    9 :  56 - 0x38
      12'hA: dout <= 8'b01111100; //   10 : 124 - 0x7c
      12'hB: dout <= 8'b11111110; //   11 : 254 - 0xfe
      12'hC: dout <= 8'b11111110; //   12 : 254 - 0xfe
      12'hD: dout <= 8'b11111110; //   13 : 254 - 0xfe
      12'hE: dout <= 8'b01111100; //   14 : 124 - 0x7c
      12'hF: dout <= 8'b00111000; //   15 :  56 - 0x38
      12'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x2
      12'h11: dout <= 8'b00000000; //   17 :   0 - 0x0
      12'h12: dout <= 8'b00000000; //   18 :   0 - 0x0
      12'h13: dout <= 8'b00000000; //   19 :   0 - 0x0
      12'h14: dout <= 8'b00000000; //   20 :   0 - 0x0
      12'h15: dout <= 8'b00000000; //   21 :   0 - 0x0
      12'h16: dout <= 8'b00000000; //   22 :   0 - 0x0
      12'h17: dout <= 8'b00000000; //   23 :   0 - 0x0
      12'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- Sprite 0x3
      12'h19: dout <= 8'b00000000; //   25 :   0 - 0x0
      12'h1A: dout <= 8'b00000000; //   26 :   0 - 0x0
      12'h1B: dout <= 8'b00011000; //   27 :  24 - 0x18
      12'h1C: dout <= 8'b00011000; //   28 :  24 - 0x18
      12'h1D: dout <= 8'b00000000; //   29 :   0 - 0x0
      12'h1E: dout <= 8'b00000000; //   30 :   0 - 0x0
      12'h1F: dout <= 8'b00000000; //   31 :   0 - 0x0
      12'h20: dout <= 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x4
      12'h21: dout <= 8'b00000000; //   33 :   0 - 0x0
      12'h22: dout <= 8'b00000000; //   34 :   0 - 0x0
      12'h23: dout <= 8'b00000000; //   35 :   0 - 0x0
      12'h24: dout <= 8'b00000000; //   36 :   0 - 0x0
      12'h25: dout <= 8'b00000000; //   37 :   0 - 0x0
      12'h26: dout <= 8'b00000000; //   38 :   0 - 0x0
      12'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout <= 8'b00000000; //   40 :   0 - 0x0 -- Sprite 0x5
      12'h29: dout <= 8'b00000000; //   41 :   0 - 0x0
      12'h2A: dout <= 8'b00000000; //   42 :   0 - 0x0
      12'h2B: dout <= 8'b00000000; //   43 :   0 - 0x0
      12'h2C: dout <= 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout <= 8'b00000000; //   45 :   0 - 0x0
      12'h2E: dout <= 8'b00000000; //   46 :   0 - 0x0
      12'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout <= 8'b00000000; //   48 :   0 - 0x0 -- Sprite 0x6
      12'h31: dout <= 8'b00000000; //   49 :   0 - 0x0
      12'h32: dout <= 8'b00000000; //   50 :   0 - 0x0
      12'h33: dout <= 8'b00000000; //   51 :   0 - 0x0
      12'h34: dout <= 8'b00000000; //   52 :   0 - 0x0
      12'h35: dout <= 8'b00000000; //   53 :   0 - 0x0
      12'h36: dout <= 8'b00000000; //   54 :   0 - 0x0
      12'h37: dout <= 8'b00000000; //   55 :   0 - 0x0
      12'h38: dout <= 8'b00000000; //   56 :   0 - 0x0 -- Sprite 0x7
      12'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      12'h3A: dout <= 8'b00000000; //   58 :   0 - 0x0
      12'h3B: dout <= 8'b00000000; //   59 :   0 - 0x0
      12'h3C: dout <= 8'b00000000; //   60 :   0 - 0x0
      12'h3D: dout <= 8'b00000000; //   61 :   0 - 0x0
      12'h3E: dout <= 8'b00000000; //   62 :   0 - 0x0
      12'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout <= 8'b00000000; //   64 :   0 - 0x0 -- Sprite 0x8
      12'h41: dout <= 8'b00000000; //   65 :   0 - 0x0
      12'h42: dout <= 8'b00000000; //   66 :   0 - 0x0
      12'h43: dout <= 8'b00000000; //   67 :   0 - 0x0
      12'h44: dout <= 8'b00000000; //   68 :   0 - 0x0
      12'h45: dout <= 8'b00000000; //   69 :   0 - 0x0
      12'h46: dout <= 8'b00000000; //   70 :   0 - 0x0
      12'h47: dout <= 8'b00000000; //   71 :   0 - 0x0
      12'h48: dout <= 8'b00000000; //   72 :   0 - 0x0 -- Sprite 0x9
      12'h49: dout <= 8'b00000000; //   73 :   0 - 0x0
      12'h4A: dout <= 8'b00000000; //   74 :   0 - 0x0
      12'h4B: dout <= 8'b00011000; //   75 :  24 - 0x18
      12'h4C: dout <= 8'b00011000; //   76 :  24 - 0x18
      12'h4D: dout <= 8'b00000000; //   77 :   0 - 0x0
      12'h4E: dout <= 8'b00000000; //   78 :   0 - 0x0
      12'h4F: dout <= 8'b00000000; //   79 :   0 - 0x0
      12'h50: dout <= 8'b00000000; //   80 :   0 - 0x0 -- Sprite 0xa
      12'h51: dout <= 8'b00000000; //   81 :   0 - 0x0
      12'h52: dout <= 8'b00000000; //   82 :   0 - 0x0
      12'h53: dout <= 8'b00000000; //   83 :   0 - 0x0
      12'h54: dout <= 8'b00000000; //   84 :   0 - 0x0
      12'h55: dout <= 8'b00000000; //   85 :   0 - 0x0
      12'h56: dout <= 8'b00000000; //   86 :   0 - 0x0
      12'h57: dout <= 8'b00000000; //   87 :   0 - 0x0
      12'h58: dout <= 8'b00000000; //   88 :   0 - 0x0 -- Sprite 0xb
      12'h59: dout <= 8'b00000000; //   89 :   0 - 0x0
      12'h5A: dout <= 8'b00000000; //   90 :   0 - 0x0
      12'h5B: dout <= 8'b00000000; //   91 :   0 - 0x0
      12'h5C: dout <= 8'b00000000; //   92 :   0 - 0x0
      12'h5D: dout <= 8'b00000000; //   93 :   0 - 0x0
      12'h5E: dout <= 8'b00000000; //   94 :   0 - 0x0
      12'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0xc
      12'h61: dout <= 8'b00000000; //   97 :   0 - 0x0
      12'h62: dout <= 8'b00000000; //   98 :   0 - 0x0
      12'h63: dout <= 8'b00000000; //   99 :   0 - 0x0
      12'h64: dout <= 8'b00000000; //  100 :   0 - 0x0
      12'h65: dout <= 8'b00000000; //  101 :   0 - 0x0
      12'h66: dout <= 8'b00000000; //  102 :   0 - 0x0
      12'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      12'h68: dout <= 8'b00000000; //  104 :   0 - 0x0 -- Sprite 0xd
      12'h69: dout <= 8'b00000000; //  105 :   0 - 0x0
      12'h6A: dout <= 8'b00000000; //  106 :   0 - 0x0
      12'h6B: dout <= 8'b00000000; //  107 :   0 - 0x0
      12'h6C: dout <= 8'b00000000; //  108 :   0 - 0x0
      12'h6D: dout <= 8'b00000000; //  109 :   0 - 0x0
      12'h6E: dout <= 8'b00000000; //  110 :   0 - 0x0
      12'h6F: dout <= 8'b00000000; //  111 :   0 - 0x0
      12'h70: dout <= 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0xe
      12'h71: dout <= 8'b00000000; //  113 :   0 - 0x0
      12'h72: dout <= 8'b00000000; //  114 :   0 - 0x0
      12'h73: dout <= 8'b00000000; //  115 :   0 - 0x0
      12'h74: dout <= 8'b00000000; //  116 :   0 - 0x0
      12'h75: dout <= 8'b00000000; //  117 :   0 - 0x0
      12'h76: dout <= 8'b00000000; //  118 :   0 - 0x0
      12'h77: dout <= 8'b00000000; //  119 :   0 - 0x0
      12'h78: dout <= 8'b00000000; //  120 :   0 - 0x0 -- Sprite 0xf
      12'h79: dout <= 8'b00000000; //  121 :   0 - 0x0
      12'h7A: dout <= 8'b00000000; //  122 :   0 - 0x0
      12'h7B: dout <= 8'b00000000; //  123 :   0 - 0x0
      12'h7C: dout <= 8'b00000000; //  124 :   0 - 0x0
      12'h7D: dout <= 8'b00000000; //  125 :   0 - 0x0
      12'h7E: dout <= 8'b00000000; //  126 :   0 - 0x0
      12'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout <= 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      12'h81: dout <= 8'b00000000; //  129 :   0 - 0x0
      12'h82: dout <= 8'b11111111; //  130 : 255 - 0xff
      12'h83: dout <= 8'b00000000; //  131 :   0 - 0x0
      12'h84: dout <= 8'b00000000; //  132 :   0 - 0x0
      12'h85: dout <= 8'b11111111; //  133 : 255 - 0xff
      12'h86: dout <= 8'b00000000; //  134 :   0 - 0x0
      12'h87: dout <= 8'b00000000; //  135 :   0 - 0x0
      12'h88: dout <= 8'b00100100; //  136 :  36 - 0x24 -- Sprite 0x11
      12'h89: dout <= 8'b00100100; //  137 :  36 - 0x24
      12'h8A: dout <= 8'b00100100; //  138 :  36 - 0x24
      12'h8B: dout <= 8'b00100100; //  139 :  36 - 0x24
      12'h8C: dout <= 8'b00100100; //  140 :  36 - 0x24
      12'h8D: dout <= 8'b00100100; //  141 :  36 - 0x24
      12'h8E: dout <= 8'b00100100; //  142 :  36 - 0x24
      12'h8F: dout <= 8'b00100100; //  143 :  36 - 0x24
      12'h90: dout <= 8'b00100100; //  144 :  36 - 0x24 -- Sprite 0x12
      12'h91: dout <= 8'b00100100; //  145 :  36 - 0x24
      12'h92: dout <= 8'b11000011; //  146 : 195 - 0xc3
      12'h93: dout <= 8'b00000000; //  147 :   0 - 0x0
      12'h94: dout <= 8'b00000000; //  148 :   0 - 0x0
      12'h95: dout <= 8'b11111111; //  149 : 255 - 0xff
      12'h96: dout <= 8'b00000000; //  150 :   0 - 0x0
      12'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      12'h98: dout <= 8'b00000000; //  152 :   0 - 0x0 -- Sprite 0x13
      12'h99: dout <= 8'b00000000; //  153 :   0 - 0x0
      12'h9A: dout <= 8'b11111111; //  154 : 255 - 0xff
      12'h9B: dout <= 8'b00000000; //  155 :   0 - 0x0
      12'h9C: dout <= 8'b00000000; //  156 :   0 - 0x0
      12'h9D: dout <= 8'b11000011; //  157 : 195 - 0xc3
      12'h9E: dout <= 8'b00100100; //  158 :  36 - 0x24
      12'h9F: dout <= 8'b00100100; //  159 :  36 - 0x24
      12'hA0: dout <= 8'b00100100; //  160 :  36 - 0x24 -- Sprite 0x14
      12'hA1: dout <= 8'b00100100; //  161 :  36 - 0x24
      12'hA2: dout <= 8'b11000100; //  162 : 196 - 0xc4
      12'hA3: dout <= 8'b00000100; //  163 :   4 - 0x4
      12'hA4: dout <= 8'b00000100; //  164 :   4 - 0x4
      12'hA5: dout <= 8'b11000100; //  165 : 196 - 0xc4
      12'hA6: dout <= 8'b00100100; //  166 :  36 - 0x24
      12'hA7: dout <= 8'b00100100; //  167 :  36 - 0x24
      12'hA8: dout <= 8'b00100100; //  168 :  36 - 0x24 -- Sprite 0x15
      12'hA9: dout <= 8'b00100100; //  169 :  36 - 0x24
      12'hAA: dout <= 8'b00100011; //  170 :  35 - 0x23
      12'hAB: dout <= 8'b00100000; //  171 :  32 - 0x20
      12'hAC: dout <= 8'b00100000; //  172 :  32 - 0x20
      12'hAD: dout <= 8'b00100011; //  173 :  35 - 0x23
      12'hAE: dout <= 8'b00100100; //  174 :  36 - 0x24
      12'hAF: dout <= 8'b00100100; //  175 :  36 - 0x24
      12'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0x16
      12'hB1: dout <= 8'b00000000; //  177 :   0 - 0x0
      12'hB2: dout <= 8'b00001111; //  178 :  15 - 0xf
      12'hB3: dout <= 8'b00010000; //  179 :  16 - 0x10
      12'hB4: dout <= 8'b11110000; //  180 : 240 - 0xf0
      12'hB5: dout <= 8'b00001111; //  181 :  15 - 0xf
      12'hB6: dout <= 8'b00000000; //  182 :   0 - 0x0
      12'hB7: dout <= 8'b00000000; //  183 :   0 - 0x0
      12'hB8: dout <= 8'b00000000; //  184 :   0 - 0x0 -- Sprite 0x17
      12'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      12'hBA: dout <= 8'b11110000; //  186 : 240 - 0xf0
      12'hBB: dout <= 8'b00001000; //  187 :   8 - 0x8
      12'hBC: dout <= 8'b00001111; //  188 :  15 - 0xf
      12'hBD: dout <= 8'b11110000; //  189 : 240 - 0xf0
      12'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      12'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0x18
      12'hC1: dout <= 8'b00000000; //  193 :   0 - 0x0
      12'hC2: dout <= 8'b11110000; //  194 : 240 - 0xf0
      12'hC3: dout <= 8'b00001000; //  195 :   8 - 0x8
      12'hC4: dout <= 8'b00001000; //  196 :   8 - 0x8
      12'hC5: dout <= 8'b11110000; //  197 : 240 - 0xf0
      12'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      12'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      12'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0 -- Sprite 0x19
      12'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      12'hCA: dout <= 8'b00001111; //  202 :  15 - 0xf
      12'hCB: dout <= 8'b00010000; //  203 :  16 - 0x10
      12'hCC: dout <= 8'b00010000; //  204 :  16 - 0x10
      12'hCD: dout <= 8'b00001111; //  205 :  15 - 0xf
      12'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      12'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      12'hD0: dout <= 8'b00100100; //  208 :  36 - 0x24 -- Sprite 0x1a
      12'hD1: dout <= 8'b00100100; //  209 :  36 - 0x24
      12'hD2: dout <= 8'b00100100; //  210 :  36 - 0x24
      12'hD3: dout <= 8'b00100100; //  211 :  36 - 0x24
      12'hD4: dout <= 8'b00011000; //  212 :  24 - 0x18
      12'hD5: dout <= 8'b00000000; //  213 :   0 - 0x0
      12'hD6: dout <= 8'b00000000; //  214 :   0 - 0x0
      12'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      12'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x1b
      12'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      12'hDA: dout <= 8'b00000000; //  218 :   0 - 0x0
      12'hDB: dout <= 8'b00011000; //  219 :  24 - 0x18
      12'hDC: dout <= 8'b00100100; //  220 :  36 - 0x24
      12'hDD: dout <= 8'b00100100; //  221 :  36 - 0x24
      12'hDE: dout <= 8'b00100100; //  222 :  36 - 0x24
      12'hDF: dout <= 8'b00100100; //  223 :  36 - 0x24
      12'hE0: dout <= 8'b00100100; //  224 :  36 - 0x24 -- Sprite 0x1c
      12'hE1: dout <= 8'b00100100; //  225 :  36 - 0x24
      12'hE2: dout <= 8'b11000100; //  226 : 196 - 0xc4
      12'hE3: dout <= 8'b00000100; //  227 :   4 - 0x4
      12'hE4: dout <= 8'b00001000; //  228 :   8 - 0x8
      12'hE5: dout <= 8'b11110000; //  229 : 240 - 0xf0
      12'hE6: dout <= 8'b00000000; //  230 :   0 - 0x0
      12'hE7: dout <= 8'b00000000; //  231 :   0 - 0x0
      12'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0 -- Sprite 0x1d
      12'hE9: dout <= 8'b00000000; //  233 :   0 - 0x0
      12'hEA: dout <= 8'b11110000; //  234 : 240 - 0xf0
      12'hEB: dout <= 8'b00001000; //  235 :   8 - 0x8
      12'hEC: dout <= 8'b00000100; //  236 :   4 - 0x4
      12'hED: dout <= 8'b11000100; //  237 : 196 - 0xc4
      12'hEE: dout <= 8'b00100100; //  238 :  36 - 0x24
      12'hEF: dout <= 8'b00100100; //  239 :  36 - 0x24
      12'hF0: dout <= 8'b00100100; //  240 :  36 - 0x24 -- Sprite 0x1e
      12'hF1: dout <= 8'b00100100; //  241 :  36 - 0x24
      12'hF2: dout <= 8'b00100011; //  242 :  35 - 0x23
      12'hF3: dout <= 8'b00100000; //  243 :  32 - 0x20
      12'hF4: dout <= 8'b00010000; //  244 :  16 - 0x10
      12'hF5: dout <= 8'b00001111; //  245 :  15 - 0xf
      12'hF6: dout <= 8'b00000000; //  246 :   0 - 0x0
      12'hF7: dout <= 8'b00000000; //  247 :   0 - 0x0
      12'hF8: dout <= 8'b00000000; //  248 :   0 - 0x0 -- Sprite 0x1f
      12'hF9: dout <= 8'b00000000; //  249 :   0 - 0x0
      12'hFA: dout <= 8'b00001111; //  250 :  15 - 0xf
      12'hFB: dout <= 8'b00010000; //  251 :  16 - 0x10
      12'hFC: dout <= 8'b00100000; //  252 :  32 - 0x20
      12'hFD: dout <= 8'b00100011; //  253 :  35 - 0x23
      12'hFE: dout <= 8'b00100100; //  254 :  36 - 0x24
      12'hFF: dout <= 8'b00100100; //  255 :  36 - 0x24
      12'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      12'h101: dout <= 8'b00000000; //  257 :   0 - 0x0
      12'h102: dout <= 8'b00000000; //  258 :   0 - 0x0
      12'h103: dout <= 8'b00000000; //  259 :   0 - 0x0
      12'h104: dout <= 8'b00000000; //  260 :   0 - 0x0
      12'h105: dout <= 8'b00000000; //  261 :   0 - 0x0
      12'h106: dout <= 8'b00000000; //  262 :   0 - 0x0
      12'h107: dout <= 8'b00000000; //  263 :   0 - 0x0
      12'h108: dout <= 8'b00000000; //  264 :   0 - 0x0 -- Sprite 0x21
      12'h109: dout <= 8'b00000000; //  265 :   0 - 0x0
      12'h10A: dout <= 8'b11110000; //  266 : 240 - 0xf0
      12'h10B: dout <= 8'b00001000; //  267 :   8 - 0x8
      12'h10C: dout <= 8'b00001000; //  268 :   8 - 0x8
      12'h10D: dout <= 8'b11110000; //  269 : 240 - 0xf0
      12'h10E: dout <= 8'b00000000; //  270 :   0 - 0x0
      12'h10F: dout <= 8'b00000000; //  271 :   0 - 0x0
      12'h110: dout <= 8'b00000000; //  272 :   0 - 0x0 -- Sprite 0x22
      12'h111: dout <= 8'b00000000; //  273 :   0 - 0x0
      12'h112: dout <= 8'b00001111; //  274 :  15 - 0xf
      12'h113: dout <= 8'b00010000; //  275 :  16 - 0x10
      12'h114: dout <= 8'b00010000; //  276 :  16 - 0x10
      12'h115: dout <= 8'b00001111; //  277 :  15 - 0xf
      12'h116: dout <= 8'b00000000; //  278 :   0 - 0x0
      12'h117: dout <= 8'b00000000; //  279 :   0 - 0x0
      12'h118: dout <= 8'b11111111; //  280 : 255 - 0xff -- Sprite 0x23
      12'h119: dout <= 8'b11111111; //  281 : 255 - 0xff
      12'h11A: dout <= 8'b11100001; //  282 : 225 - 0xe1
      12'h11B: dout <= 8'b11100001; //  283 : 225 - 0xe1
      12'h11C: dout <= 8'b11100001; //  284 : 225 - 0xe1
      12'h11D: dout <= 8'b11100001; //  285 : 225 - 0xe1
      12'h11E: dout <= 8'b11100001; //  286 : 225 - 0xe1
      12'h11F: dout <= 8'b11100001; //  287 : 225 - 0xe1
      12'h120: dout <= 8'b10000111; //  288 : 135 - 0x87 -- Sprite 0x24
      12'h121: dout <= 8'b11000111; //  289 : 199 - 0xc7
      12'h122: dout <= 8'b11000000; //  290 : 192 - 0xc0
      12'h123: dout <= 8'b11000111; //  291 : 199 - 0xc7
      12'h124: dout <= 8'b11001111; //  292 : 207 - 0xcf
      12'h125: dout <= 8'b11001110; //  293 : 206 - 0xce
      12'h126: dout <= 8'b11001111; //  294 : 207 - 0xcf
      12'h127: dout <= 8'b11000111; //  295 : 199 - 0xc7
      12'h128: dout <= 8'b11111000; //  296 : 248 - 0xf8 -- Sprite 0x25
      12'h129: dout <= 8'b11111100; //  297 : 252 - 0xfc
      12'h12A: dout <= 8'b00011100; //  298 :  28 - 0x1c
      12'h12B: dout <= 8'b11111100; //  299 : 252 - 0xfc
      12'h12C: dout <= 8'b11111100; //  300 : 252 - 0xfc
      12'h12D: dout <= 8'b00011100; //  301 :  28 - 0x1c
      12'h12E: dout <= 8'b11111100; //  302 : 252 - 0xfc
      12'h12F: dout <= 8'b11111100; //  303 : 252 - 0xfc
      12'h130: dout <= 8'b11111111; //  304 : 255 - 0xff -- Sprite 0x26
      12'h131: dout <= 8'b11111111; //  305 : 255 - 0xff
      12'h132: dout <= 8'b11100111; //  306 : 231 - 0xe7
      12'h133: dout <= 8'b11100111; //  307 : 231 - 0xe7
      12'h134: dout <= 8'b11100111; //  308 : 231 - 0xe7
      12'h135: dout <= 8'b11100111; //  309 : 231 - 0xe7
      12'h136: dout <= 8'b11100111; //  310 : 231 - 0xe7
      12'h137: dout <= 8'b11100111; //  311 : 231 - 0xe7
      12'h138: dout <= 8'b11110000; //  312 : 240 - 0xf0 -- Sprite 0x27
      12'h139: dout <= 8'b11111001; //  313 : 249 - 0xf9
      12'h13A: dout <= 8'b00111001; //  314 :  57 - 0x39
      12'h13B: dout <= 8'b00111001; //  315 :  57 - 0x39
      12'h13C: dout <= 8'b00111001; //  316 :  57 - 0x39
      12'h13D: dout <= 8'b00111001; //  317 :  57 - 0x39
      12'h13E: dout <= 8'b00111001; //  318 :  57 - 0x39
      12'h13F: dout <= 8'b00111000; //  319 :  56 - 0x38
      12'h140: dout <= 8'b11111111; //  320 : 255 - 0xff -- Sprite 0x28
      12'h141: dout <= 8'b11111111; //  321 : 255 - 0xff
      12'h142: dout <= 8'b11000000; //  322 : 192 - 0xc0
      12'h143: dout <= 8'b11000000; //  323 : 192 - 0xc0
      12'h144: dout <= 8'b11000000; //  324 : 192 - 0xc0
      12'h145: dout <= 8'b11000000; //  325 : 192 - 0xc0
      12'h146: dout <= 8'b11111111; //  326 : 255 - 0xff
      12'h147: dout <= 8'b11111111; //  327 : 255 - 0xff
      12'h148: dout <= 8'b00011111; //  328 :  31 - 0x1f -- Sprite 0x29
      12'h149: dout <= 8'b00111111; //  329 :  63 - 0x3f
      12'h14A: dout <= 8'b00110000; //  330 :  48 - 0x30
      12'h14B: dout <= 8'b00110000; //  331 :  48 - 0x30
      12'h14C: dout <= 8'b00110000; //  332 :  48 - 0x30
      12'h14D: dout <= 8'b00110000; //  333 :  48 - 0x30
      12'h14E: dout <= 8'b00111111; //  334 :  63 - 0x3f
      12'h14F: dout <= 8'b00011111; //  335 :  31 - 0x1f
      12'h150: dout <= 8'b11100011; //  336 : 227 - 0xe3 -- Sprite 0x2a
      12'h151: dout <= 8'b11110011; //  337 : 243 - 0xf3
      12'h152: dout <= 8'b01110000; //  338 : 112 - 0x70
      12'h153: dout <= 8'b01110000; //  339 : 112 - 0x70
      12'h154: dout <= 8'b01110000; //  340 : 112 - 0x70
      12'h155: dout <= 8'b01110000; //  341 : 112 - 0x70
      12'h156: dout <= 8'b11110000; //  342 : 240 - 0xf0
      12'h157: dout <= 8'b11100000; //  343 : 224 - 0xe0
      12'h158: dout <= 8'b11111110; //  344 : 254 - 0xfe -- Sprite 0x2b
      12'h159: dout <= 8'b11111110; //  345 : 254 - 0xfe
      12'h15A: dout <= 8'b01110000; //  346 : 112 - 0x70
      12'h15B: dout <= 8'b01110000; //  347 : 112 - 0x70
      12'h15C: dout <= 8'b01110000; //  348 : 112 - 0x70
      12'h15D: dout <= 8'b01110000; //  349 : 112 - 0x70
      12'h15E: dout <= 8'b01110000; //  350 : 112 - 0x70
      12'h15F: dout <= 8'b01110000; //  351 : 112 - 0x70
      12'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x2c
      12'h161: dout <= 8'b00000000; //  353 :   0 - 0x0
      12'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      12'h163: dout <= 8'b00000000; //  355 :   0 - 0x0
      12'h164: dout <= 8'b11111111; //  356 : 255 - 0xff
      12'h165: dout <= 8'b00000000; //  357 :   0 - 0x0
      12'h166: dout <= 8'b00000000; //  358 :   0 - 0x0
      12'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout <= 8'b00000000; //  360 :   0 - 0x0 -- Sprite 0x2d
      12'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      12'h16A: dout <= 8'b00000000; //  362 :   0 - 0x0
      12'h16B: dout <= 8'b00000000; //  363 :   0 - 0x0
      12'h16C: dout <= 8'b00000000; //  364 :   0 - 0x0
      12'h16D: dout <= 8'b00000000; //  365 :   0 - 0x0
      12'h16E: dout <= 8'b00000000; //  366 :   0 - 0x0
      12'h16F: dout <= 8'b00000000; //  367 :   0 - 0x0
      12'h170: dout <= 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x2e
      12'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      12'h172: dout <= 8'b00000000; //  370 :   0 - 0x0
      12'h173: dout <= 8'b00011000; //  371 :  24 - 0x18
      12'h174: dout <= 8'b00011000; //  372 :  24 - 0x18
      12'h175: dout <= 8'b00000000; //  373 :   0 - 0x0
      12'h176: dout <= 8'b00000000; //  374 :   0 - 0x0
      12'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      12'h178: dout <= 8'b00000000; //  376 :   0 - 0x0 -- Sprite 0x2f
      12'h179: dout <= 8'b00000000; //  377 :   0 - 0x0
      12'h17A: dout <= 8'b00000000; //  378 :   0 - 0x0
      12'h17B: dout <= 8'b00000000; //  379 :   0 - 0x0
      12'h17C: dout <= 8'b00000000; //  380 :   0 - 0x0
      12'h17D: dout <= 8'b00000000; //  381 :   0 - 0x0
      12'h17E: dout <= 8'b00000000; //  382 :   0 - 0x0
      12'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      12'h180: dout <= 8'b00011100; //  384 :  28 - 0x1c -- Sprite 0x30
      12'h181: dout <= 8'b00100110; //  385 :  38 - 0x26
      12'h182: dout <= 8'b01100011; //  386 :  99 - 0x63
      12'h183: dout <= 8'b01100011; //  387 :  99 - 0x63
      12'h184: dout <= 8'b01100011; //  388 :  99 - 0x63
      12'h185: dout <= 8'b00110010; //  389 :  50 - 0x32
      12'h186: dout <= 8'b00011100; //  390 :  28 - 0x1c
      12'h187: dout <= 8'b00000000; //  391 :   0 - 0x0
      12'h188: dout <= 8'b00001100; //  392 :  12 - 0xc -- Sprite 0x31
      12'h189: dout <= 8'b00011100; //  393 :  28 - 0x1c
      12'h18A: dout <= 8'b00001100; //  394 :  12 - 0xc
      12'h18B: dout <= 8'b00001100; //  395 :  12 - 0xc
      12'h18C: dout <= 8'b00001100; //  396 :  12 - 0xc
      12'h18D: dout <= 8'b00001100; //  397 :  12 - 0xc
      12'h18E: dout <= 8'b00111111; //  398 :  63 - 0x3f
      12'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      12'h190: dout <= 8'b00111110; //  400 :  62 - 0x3e -- Sprite 0x32
      12'h191: dout <= 8'b01100011; //  401 :  99 - 0x63
      12'h192: dout <= 8'b00000111; //  402 :   7 - 0x7
      12'h193: dout <= 8'b00011110; //  403 :  30 - 0x1e
      12'h194: dout <= 8'b00111100; //  404 :  60 - 0x3c
      12'h195: dout <= 8'b01110000; //  405 : 112 - 0x70
      12'h196: dout <= 8'b01111111; //  406 : 127 - 0x7f
      12'h197: dout <= 8'b00000000; //  407 :   0 - 0x0
      12'h198: dout <= 8'b00111111; //  408 :  63 - 0x3f -- Sprite 0x33
      12'h199: dout <= 8'b00000110; //  409 :   6 - 0x6
      12'h19A: dout <= 8'b00001100; //  410 :  12 - 0xc
      12'h19B: dout <= 8'b00011110; //  411 :  30 - 0x1e
      12'h19C: dout <= 8'b00000011; //  412 :   3 - 0x3
      12'h19D: dout <= 8'b01100011; //  413 :  99 - 0x63
      12'h19E: dout <= 8'b00111110; //  414 :  62 - 0x3e
      12'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout <= 8'b00001110; //  416 :  14 - 0xe -- Sprite 0x34
      12'h1A1: dout <= 8'b00011110; //  417 :  30 - 0x1e
      12'h1A2: dout <= 8'b00110110; //  418 :  54 - 0x36
      12'h1A3: dout <= 8'b01100110; //  419 : 102 - 0x66
      12'h1A4: dout <= 8'b01111111; //  420 : 127 - 0x7f
      12'h1A5: dout <= 8'b00000110; //  421 :   6 - 0x6
      12'h1A6: dout <= 8'b00000110; //  422 :   6 - 0x6
      12'h1A7: dout <= 8'b00000000; //  423 :   0 - 0x0
      12'h1A8: dout <= 8'b01111110; //  424 : 126 - 0x7e -- Sprite 0x35
      12'h1A9: dout <= 8'b01100000; //  425 :  96 - 0x60
      12'h1AA: dout <= 8'b01111110; //  426 : 126 - 0x7e
      12'h1AB: dout <= 8'b00000011; //  427 :   3 - 0x3
      12'h1AC: dout <= 8'b00000011; //  428 :   3 - 0x3
      12'h1AD: dout <= 8'b01100011; //  429 :  99 - 0x63
      12'h1AE: dout <= 8'b00111110; //  430 :  62 - 0x3e
      12'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      12'h1B0: dout <= 8'b00011110; //  432 :  30 - 0x1e -- Sprite 0x36
      12'h1B1: dout <= 8'b00110000; //  433 :  48 - 0x30
      12'h1B2: dout <= 8'b01100000; //  434 :  96 - 0x60
      12'h1B3: dout <= 8'b01111110; //  435 : 126 - 0x7e
      12'h1B4: dout <= 8'b01100011; //  436 :  99 - 0x63
      12'h1B5: dout <= 8'b01100011; //  437 :  99 - 0x63
      12'h1B6: dout <= 8'b00111110; //  438 :  62 - 0x3e
      12'h1B7: dout <= 8'b00000000; //  439 :   0 - 0x0
      12'h1B8: dout <= 8'b01111111; //  440 : 127 - 0x7f -- Sprite 0x37
      12'h1B9: dout <= 8'b01100011; //  441 :  99 - 0x63
      12'h1BA: dout <= 8'b00000110; //  442 :   6 - 0x6
      12'h1BB: dout <= 8'b00001100; //  443 :  12 - 0xc
      12'h1BC: dout <= 8'b00011000; //  444 :  24 - 0x18
      12'h1BD: dout <= 8'b00011000; //  445 :  24 - 0x18
      12'h1BE: dout <= 8'b00011000; //  446 :  24 - 0x18
      12'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout <= 8'b00111100; //  448 :  60 - 0x3c -- Sprite 0x38
      12'h1C1: dout <= 8'b01100010; //  449 :  98 - 0x62
      12'h1C2: dout <= 8'b01110010; //  450 : 114 - 0x72
      12'h1C3: dout <= 8'b00111100; //  451 :  60 - 0x3c
      12'h1C4: dout <= 8'b01001111; //  452 :  79 - 0x4f
      12'h1C5: dout <= 8'b01000011; //  453 :  67 - 0x43
      12'h1C6: dout <= 8'b00111110; //  454 :  62 - 0x3e
      12'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      12'h1C8: dout <= 8'b00111110; //  456 :  62 - 0x3e -- Sprite 0x39
      12'h1C9: dout <= 8'b01100011; //  457 :  99 - 0x63
      12'h1CA: dout <= 8'b01100011; //  458 :  99 - 0x63
      12'h1CB: dout <= 8'b00111111; //  459 :  63 - 0x3f
      12'h1CC: dout <= 8'b00000011; //  460 :   3 - 0x3
      12'h1CD: dout <= 8'b00000110; //  461 :   6 - 0x6
      12'h1CE: dout <= 8'b00111100; //  462 :  60 - 0x3c
      12'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      12'h1D1: dout <= 8'b00000000; //  465 :   0 - 0x0
      12'h1D2: dout <= 8'b00000000; //  466 :   0 - 0x0
      12'h1D3: dout <= 8'b01111110; //  467 : 126 - 0x7e
      12'h1D4: dout <= 8'b00000000; //  468 :   0 - 0x0
      12'h1D5: dout <= 8'b00000000; //  469 :   0 - 0x0
      12'h1D6: dout <= 8'b00000000; //  470 :   0 - 0x0
      12'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      12'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0 -- Sprite 0x3b
      12'h1D9: dout <= 8'b00000010; //  473 :   2 - 0x2
      12'h1DA: dout <= 8'b00000100; //  474 :   4 - 0x4
      12'h1DB: dout <= 8'b00001000; //  475 :   8 - 0x8
      12'h1DC: dout <= 8'b00010000; //  476 :  16 - 0x10
      12'h1DD: dout <= 8'b00100000; //  477 :  32 - 0x20
      12'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      12'h1E1: dout <= 8'b00000111; //  481 :   7 - 0x7
      12'h1E2: dout <= 8'b00011111; //  482 :  31 - 0x1f
      12'h1E3: dout <= 8'b00111111; //  483 :  63 - 0x3f
      12'h1E4: dout <= 8'b00111111; //  484 :  63 - 0x3f
      12'h1E5: dout <= 8'b00001111; //  485 :  15 - 0xf
      12'h1E6: dout <= 8'b00000011; //  486 :   3 - 0x3
      12'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      12'h1E9: dout <= 8'b11000000; //  489 : 192 - 0xc0
      12'h1EA: dout <= 8'b11110000; //  490 : 240 - 0xf0
      12'h1EB: dout <= 8'b11111000; //  491 : 248 - 0xf8
      12'h1EC: dout <= 8'b11111000; //  492 : 248 - 0xf8
      12'h1ED: dout <= 8'b11111100; //  493 : 252 - 0xfc
      12'h1EE: dout <= 8'b11111100; //  494 : 252 - 0xfc
      12'h1EF: dout <= 8'b11111100; //  495 : 252 - 0xfc
      12'h1F0: dout <= 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      12'h1F1: dout <= 8'b00000011; //  497 :   3 - 0x3
      12'h1F2: dout <= 8'b00001111; //  498 :  15 - 0xf
      12'h1F3: dout <= 8'b00111111; //  499 :  63 - 0x3f
      12'h1F4: dout <= 8'b00111111; //  500 :  63 - 0x3f
      12'h1F5: dout <= 8'b00011111; //  501 :  31 - 0x1f
      12'h1F6: dout <= 8'b00000111; //  502 :   7 - 0x7
      12'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      12'h1F8: dout <= 8'b11111100; //  504 : 252 - 0xfc -- Sprite 0x3f
      12'h1F9: dout <= 8'b11111100; //  505 : 252 - 0xfc
      12'h1FA: dout <= 8'b11111100; //  506 : 252 - 0xfc
      12'h1FB: dout <= 8'b11111000; //  507 : 248 - 0xf8
      12'h1FC: dout <= 8'b11111000; //  508 : 248 - 0xf8
      12'h1FD: dout <= 8'b11110000; //  509 : 240 - 0xf0
      12'h1FE: dout <= 8'b11000000; //  510 : 192 - 0xc0
      12'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout <= 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x40
      12'h201: dout <= 8'b00000000; //  513 :   0 - 0x0
      12'h202: dout <= 8'b00000000; //  514 :   0 - 0x0
      12'h203: dout <= 8'b00000000; //  515 :   0 - 0x0
      12'h204: dout <= 8'b00000000; //  516 :   0 - 0x0
      12'h205: dout <= 8'b00000000; //  517 :   0 - 0x0
      12'h206: dout <= 8'b00000000; //  518 :   0 - 0x0
      12'h207: dout <= 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout <= 8'b00011100; //  520 :  28 - 0x1c -- Sprite 0x41
      12'h209: dout <= 8'b00110110; //  521 :  54 - 0x36
      12'h20A: dout <= 8'b01100011; //  522 :  99 - 0x63
      12'h20B: dout <= 8'b01100011; //  523 :  99 - 0x63
      12'h20C: dout <= 8'b01111111; //  524 : 127 - 0x7f
      12'h20D: dout <= 8'b01100011; //  525 :  99 - 0x63
      12'h20E: dout <= 8'b01100011; //  526 :  99 - 0x63
      12'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout <= 8'b01111110; //  528 : 126 - 0x7e -- Sprite 0x42
      12'h211: dout <= 8'b01100011; //  529 :  99 - 0x63
      12'h212: dout <= 8'b01100011; //  530 :  99 - 0x63
      12'h213: dout <= 8'b01111110; //  531 : 126 - 0x7e
      12'h214: dout <= 8'b01100011; //  532 :  99 - 0x63
      12'h215: dout <= 8'b01100011; //  533 :  99 - 0x63
      12'h216: dout <= 8'b01111110; //  534 : 126 - 0x7e
      12'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      12'h218: dout <= 8'b00011110; //  536 :  30 - 0x1e -- Sprite 0x43
      12'h219: dout <= 8'b00110011; //  537 :  51 - 0x33
      12'h21A: dout <= 8'b01100000; //  538 :  96 - 0x60
      12'h21B: dout <= 8'b01100000; //  539 :  96 - 0x60
      12'h21C: dout <= 8'b01100000; //  540 :  96 - 0x60
      12'h21D: dout <= 8'b00110011; //  541 :  51 - 0x33
      12'h21E: dout <= 8'b00011110; //  542 :  30 - 0x1e
      12'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout <= 8'b01111100; //  544 : 124 - 0x7c -- Sprite 0x44
      12'h221: dout <= 8'b01100110; //  545 : 102 - 0x66
      12'h222: dout <= 8'b01100011; //  546 :  99 - 0x63
      12'h223: dout <= 8'b01100011; //  547 :  99 - 0x63
      12'h224: dout <= 8'b01100011; //  548 :  99 - 0x63
      12'h225: dout <= 8'b01100110; //  549 : 102 - 0x66
      12'h226: dout <= 8'b01111100; //  550 : 124 - 0x7c
      12'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      12'h228: dout <= 8'b01111111; //  552 : 127 - 0x7f -- Sprite 0x45
      12'h229: dout <= 8'b01100000; //  553 :  96 - 0x60
      12'h22A: dout <= 8'b01100000; //  554 :  96 - 0x60
      12'h22B: dout <= 8'b01111110; //  555 : 126 - 0x7e
      12'h22C: dout <= 8'b01100000; //  556 :  96 - 0x60
      12'h22D: dout <= 8'b01100000; //  557 :  96 - 0x60
      12'h22E: dout <= 8'b01111111; //  558 : 127 - 0x7f
      12'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout <= 8'b01111111; //  560 : 127 - 0x7f -- Sprite 0x46
      12'h231: dout <= 8'b01100000; //  561 :  96 - 0x60
      12'h232: dout <= 8'b01100000; //  562 :  96 - 0x60
      12'h233: dout <= 8'b01111110; //  563 : 126 - 0x7e
      12'h234: dout <= 8'b01100000; //  564 :  96 - 0x60
      12'h235: dout <= 8'b01100000; //  565 :  96 - 0x60
      12'h236: dout <= 8'b01100000; //  566 :  96 - 0x60
      12'h237: dout <= 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout <= 8'b00011111; //  568 :  31 - 0x1f -- Sprite 0x47
      12'h239: dout <= 8'b00110000; //  569 :  48 - 0x30
      12'h23A: dout <= 8'b01100000; //  570 :  96 - 0x60
      12'h23B: dout <= 8'b01100111; //  571 : 103 - 0x67
      12'h23C: dout <= 8'b01100011; //  572 :  99 - 0x63
      12'h23D: dout <= 8'b00110011; //  573 :  51 - 0x33
      12'h23E: dout <= 8'b00011111; //  574 :  31 - 0x1f
      12'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout <= 8'b01100011; //  576 :  99 - 0x63 -- Sprite 0x48
      12'h241: dout <= 8'b01100011; //  577 :  99 - 0x63
      12'h242: dout <= 8'b01100011; //  578 :  99 - 0x63
      12'h243: dout <= 8'b01111111; //  579 : 127 - 0x7f
      12'h244: dout <= 8'b01100011; //  580 :  99 - 0x63
      12'h245: dout <= 8'b01100011; //  581 :  99 - 0x63
      12'h246: dout <= 8'b01100011; //  582 :  99 - 0x63
      12'h247: dout <= 8'b00000000; //  583 :   0 - 0x0
      12'h248: dout <= 8'b00111111; //  584 :  63 - 0x3f -- Sprite 0x49
      12'h249: dout <= 8'b00001100; //  585 :  12 - 0xc
      12'h24A: dout <= 8'b00001100; //  586 :  12 - 0xc
      12'h24B: dout <= 8'b00001100; //  587 :  12 - 0xc
      12'h24C: dout <= 8'b00001100; //  588 :  12 - 0xc
      12'h24D: dout <= 8'b00001100; //  589 :  12 - 0xc
      12'h24E: dout <= 8'b00111111; //  590 :  63 - 0x3f
      12'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout <= 8'b00000011; //  592 :   3 - 0x3 -- Sprite 0x4a
      12'h251: dout <= 8'b00000011; //  593 :   3 - 0x3
      12'h252: dout <= 8'b00000011; //  594 :   3 - 0x3
      12'h253: dout <= 8'b00000011; //  595 :   3 - 0x3
      12'h254: dout <= 8'b00000011; //  596 :   3 - 0x3
      12'h255: dout <= 8'b01100011; //  597 :  99 - 0x63
      12'h256: dout <= 8'b00111110; //  598 :  62 - 0x3e
      12'h257: dout <= 8'b00000000; //  599 :   0 - 0x0
      12'h258: dout <= 8'b01100011; //  600 :  99 - 0x63 -- Sprite 0x4b
      12'h259: dout <= 8'b01100110; //  601 : 102 - 0x66
      12'h25A: dout <= 8'b01101100; //  602 : 108 - 0x6c
      12'h25B: dout <= 8'b01111000; //  603 : 120 - 0x78
      12'h25C: dout <= 8'b01111100; //  604 : 124 - 0x7c
      12'h25D: dout <= 8'b01100110; //  605 : 102 - 0x66
      12'h25E: dout <= 8'b01100011; //  606 :  99 - 0x63
      12'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout <= 8'b01100000; //  608 :  96 - 0x60 -- Sprite 0x4c
      12'h261: dout <= 8'b01100000; //  609 :  96 - 0x60
      12'h262: dout <= 8'b01100000; //  610 :  96 - 0x60
      12'h263: dout <= 8'b01100000; //  611 :  96 - 0x60
      12'h264: dout <= 8'b01100000; //  612 :  96 - 0x60
      12'h265: dout <= 8'b01100000; //  613 :  96 - 0x60
      12'h266: dout <= 8'b01111111; //  614 : 127 - 0x7f
      12'h267: dout <= 8'b00000000; //  615 :   0 - 0x0
      12'h268: dout <= 8'b01100011; //  616 :  99 - 0x63 -- Sprite 0x4d
      12'h269: dout <= 8'b01110111; //  617 : 119 - 0x77
      12'h26A: dout <= 8'b01111111; //  618 : 127 - 0x7f
      12'h26B: dout <= 8'b01111111; //  619 : 127 - 0x7f
      12'h26C: dout <= 8'b01101011; //  620 : 107 - 0x6b
      12'h26D: dout <= 8'b01100011; //  621 :  99 - 0x63
      12'h26E: dout <= 8'b01100011; //  622 :  99 - 0x63
      12'h26F: dout <= 8'b00000000; //  623 :   0 - 0x0
      12'h270: dout <= 8'b01100011; //  624 :  99 - 0x63 -- Sprite 0x4e
      12'h271: dout <= 8'b01110011; //  625 : 115 - 0x73
      12'h272: dout <= 8'b01111011; //  626 : 123 - 0x7b
      12'h273: dout <= 8'b01111111; //  627 : 127 - 0x7f
      12'h274: dout <= 8'b01101111; //  628 : 111 - 0x6f
      12'h275: dout <= 8'b01100111; //  629 : 103 - 0x67
      12'h276: dout <= 8'b01100011; //  630 :  99 - 0x63
      12'h277: dout <= 8'b00000000; //  631 :   0 - 0x0
      12'h278: dout <= 8'b00111110; //  632 :  62 - 0x3e -- Sprite 0x4f
      12'h279: dout <= 8'b01100011; //  633 :  99 - 0x63
      12'h27A: dout <= 8'b01100011; //  634 :  99 - 0x63
      12'h27B: dout <= 8'b01100011; //  635 :  99 - 0x63
      12'h27C: dout <= 8'b01100011; //  636 :  99 - 0x63
      12'h27D: dout <= 8'b01100011; //  637 :  99 - 0x63
      12'h27E: dout <= 8'b00111110; //  638 :  62 - 0x3e
      12'h27F: dout <= 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout <= 8'b01111110; //  640 : 126 - 0x7e -- Sprite 0x50
      12'h281: dout <= 8'b01100011; //  641 :  99 - 0x63
      12'h282: dout <= 8'b01100011; //  642 :  99 - 0x63
      12'h283: dout <= 8'b01100011; //  643 :  99 - 0x63
      12'h284: dout <= 8'b01111110; //  644 : 126 - 0x7e
      12'h285: dout <= 8'b01100000; //  645 :  96 - 0x60
      12'h286: dout <= 8'b01100000; //  646 :  96 - 0x60
      12'h287: dout <= 8'b00000000; //  647 :   0 - 0x0
      12'h288: dout <= 8'b00111110; //  648 :  62 - 0x3e -- Sprite 0x51
      12'h289: dout <= 8'b01100011; //  649 :  99 - 0x63
      12'h28A: dout <= 8'b01100011; //  650 :  99 - 0x63
      12'h28B: dout <= 8'b01100011; //  651 :  99 - 0x63
      12'h28C: dout <= 8'b01101111; //  652 : 111 - 0x6f
      12'h28D: dout <= 8'b01100110; //  653 : 102 - 0x66
      12'h28E: dout <= 8'b00111101; //  654 :  61 - 0x3d
      12'h28F: dout <= 8'b00000000; //  655 :   0 - 0x0
      12'h290: dout <= 8'b01111110; //  656 : 126 - 0x7e -- Sprite 0x52
      12'h291: dout <= 8'b01100011; //  657 :  99 - 0x63
      12'h292: dout <= 8'b01100011; //  658 :  99 - 0x63
      12'h293: dout <= 8'b01100111; //  659 : 103 - 0x67
      12'h294: dout <= 8'b01111100; //  660 : 124 - 0x7c
      12'h295: dout <= 8'b01101110; //  661 : 110 - 0x6e
      12'h296: dout <= 8'b01100111; //  662 : 103 - 0x67
      12'h297: dout <= 8'b00000000; //  663 :   0 - 0x0
      12'h298: dout <= 8'b00111100; //  664 :  60 - 0x3c -- Sprite 0x53
      12'h299: dout <= 8'b01100110; //  665 : 102 - 0x66
      12'h29A: dout <= 8'b01100000; //  666 :  96 - 0x60
      12'h29B: dout <= 8'b00111110; //  667 :  62 - 0x3e
      12'h29C: dout <= 8'b00000011; //  668 :   3 - 0x3
      12'h29D: dout <= 8'b01100011; //  669 :  99 - 0x63
      12'h29E: dout <= 8'b00111110; //  670 :  62 - 0x3e
      12'h29F: dout <= 8'b00000000; //  671 :   0 - 0x0
      12'h2A0: dout <= 8'b00111111; //  672 :  63 - 0x3f -- Sprite 0x54
      12'h2A1: dout <= 8'b00001100; //  673 :  12 - 0xc
      12'h2A2: dout <= 8'b00001100; //  674 :  12 - 0xc
      12'h2A3: dout <= 8'b00001100; //  675 :  12 - 0xc
      12'h2A4: dout <= 8'b00001100; //  676 :  12 - 0xc
      12'h2A5: dout <= 8'b00001100; //  677 :  12 - 0xc
      12'h2A6: dout <= 8'b00001100; //  678 :  12 - 0xc
      12'h2A7: dout <= 8'b00000000; //  679 :   0 - 0x0
      12'h2A8: dout <= 8'b01100011; //  680 :  99 - 0x63 -- Sprite 0x55
      12'h2A9: dout <= 8'b01100011; //  681 :  99 - 0x63
      12'h2AA: dout <= 8'b01100011; //  682 :  99 - 0x63
      12'h2AB: dout <= 8'b01100011; //  683 :  99 - 0x63
      12'h2AC: dout <= 8'b01100011; //  684 :  99 - 0x63
      12'h2AD: dout <= 8'b01100011; //  685 :  99 - 0x63
      12'h2AE: dout <= 8'b00111110; //  686 :  62 - 0x3e
      12'h2AF: dout <= 8'b00000000; //  687 :   0 - 0x0
      12'h2B0: dout <= 8'b01100011; //  688 :  99 - 0x63 -- Sprite 0x56
      12'h2B1: dout <= 8'b01100011; //  689 :  99 - 0x63
      12'h2B2: dout <= 8'b01100011; //  690 :  99 - 0x63
      12'h2B3: dout <= 8'b01110111; //  691 : 119 - 0x77
      12'h2B4: dout <= 8'b00111110; //  692 :  62 - 0x3e
      12'h2B5: dout <= 8'b00011100; //  693 :  28 - 0x1c
      12'h2B6: dout <= 8'b00001000; //  694 :   8 - 0x8
      12'h2B7: dout <= 8'b00000000; //  695 :   0 - 0x0
      12'h2B8: dout <= 8'b01100011; //  696 :  99 - 0x63 -- Sprite 0x57
      12'h2B9: dout <= 8'b01100011; //  697 :  99 - 0x63
      12'h2BA: dout <= 8'b01101011; //  698 : 107 - 0x6b
      12'h2BB: dout <= 8'b01111111; //  699 : 127 - 0x7f
      12'h2BC: dout <= 8'b01111111; //  700 : 127 - 0x7f
      12'h2BD: dout <= 8'b01110111; //  701 : 119 - 0x77
      12'h2BE: dout <= 8'b01100011; //  702 :  99 - 0x63
      12'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout <= 8'b01100011; //  704 :  99 - 0x63 -- Sprite 0x58
      12'h2C1: dout <= 8'b01110111; //  705 : 119 - 0x77
      12'h2C2: dout <= 8'b00111110; //  706 :  62 - 0x3e
      12'h2C3: dout <= 8'b00011100; //  707 :  28 - 0x1c
      12'h2C4: dout <= 8'b00111110; //  708 :  62 - 0x3e
      12'h2C5: dout <= 8'b01110111; //  709 : 119 - 0x77
      12'h2C6: dout <= 8'b01100011; //  710 :  99 - 0x63
      12'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout <= 8'b00110011; //  712 :  51 - 0x33 -- Sprite 0x59
      12'h2C9: dout <= 8'b00110011; //  713 :  51 - 0x33
      12'h2CA: dout <= 8'b00110011; //  714 :  51 - 0x33
      12'h2CB: dout <= 8'b00011110; //  715 :  30 - 0x1e
      12'h2CC: dout <= 8'b00001100; //  716 :  12 - 0xc
      12'h2CD: dout <= 8'b00001100; //  717 :  12 - 0xc
      12'h2CE: dout <= 8'b00001100; //  718 :  12 - 0xc
      12'h2CF: dout <= 8'b00000000; //  719 :   0 - 0x0
      12'h2D0: dout <= 8'b01111111; //  720 : 127 - 0x7f -- Sprite 0x5a
      12'h2D1: dout <= 8'b00000111; //  721 :   7 - 0x7
      12'h2D2: dout <= 8'b00001110; //  722 :  14 - 0xe
      12'h2D3: dout <= 8'b00011100; //  723 :  28 - 0x1c
      12'h2D4: dout <= 8'b00111000; //  724 :  56 - 0x38
      12'h2D5: dout <= 8'b01110000; //  725 : 112 - 0x70
      12'h2D6: dout <= 8'b01111111; //  726 : 127 - 0x7f
      12'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      12'h2D8: dout <= 8'b00000000; //  728 :   0 - 0x0 -- Sprite 0x5b
      12'h2D9: dout <= 8'b00000000; //  729 :   0 - 0x0
      12'h2DA: dout <= 8'b00000000; //  730 :   0 - 0x0
      12'h2DB: dout <= 8'b00000000; //  731 :   0 - 0x0
      12'h2DC: dout <= 8'b00000000; //  732 :   0 - 0x0
      12'h2DD: dout <= 8'b00110000; //  733 :  48 - 0x30
      12'h2DE: dout <= 8'b00110000; //  734 :  48 - 0x30
      12'h2DF: dout <= 8'b00000000; //  735 :   0 - 0x0
      12'h2E0: dout <= 8'b11000000; //  736 : 192 - 0xc0 -- Sprite 0x5c
      12'h2E1: dout <= 8'b11110000; //  737 : 240 - 0xf0
      12'h2E2: dout <= 8'b11111100; //  738 : 252 - 0xfc
      12'h2E3: dout <= 8'b11111111; //  739 : 255 - 0xff
      12'h2E4: dout <= 8'b11111100; //  740 : 252 - 0xfc
      12'h2E5: dout <= 8'b11110000; //  741 : 240 - 0xf0
      12'h2E6: dout <= 8'b11000000; //  742 : 192 - 0xc0
      12'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout <= 8'b00111100; //  744 :  60 - 0x3c -- Sprite 0x5d
      12'h2E9: dout <= 8'b01000010; //  745 :  66 - 0x42
      12'h2EA: dout <= 8'b10011001; //  746 : 153 - 0x99
      12'h2EB: dout <= 8'b10100001; //  747 : 161 - 0xa1
      12'h2EC: dout <= 8'b10100001; //  748 : 161 - 0xa1
      12'h2ED: dout <= 8'b10011001; //  749 : 153 - 0x99
      12'h2EE: dout <= 8'b01000010; //  750 :  66 - 0x42
      12'h2EF: dout <= 8'b00111100; //  751 :  60 - 0x3c
      12'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x5e
      12'h2F1: dout <= 8'b00000000; //  753 :   0 - 0x0
      12'h2F2: dout <= 8'b00010000; //  754 :  16 - 0x10
      12'h2F3: dout <= 8'b00010000; //  755 :  16 - 0x10
      12'h2F4: dout <= 8'b00010000; //  756 :  16 - 0x10
      12'h2F5: dout <= 8'b00010000; //  757 :  16 - 0x10
      12'h2F6: dout <= 8'b00000000; //  758 :   0 - 0x0
      12'h2F7: dout <= 8'b00000000; //  759 :   0 - 0x0
      12'h2F8: dout <= 8'b00110110; //  760 :  54 - 0x36 -- Sprite 0x5f
      12'h2F9: dout <= 8'b00110110; //  761 :  54 - 0x36
      12'h2FA: dout <= 8'b00010010; //  762 :  18 - 0x12
      12'h2FB: dout <= 8'b00000000; //  763 :   0 - 0x0
      12'h2FC: dout <= 8'b00000000; //  764 :   0 - 0x0
      12'h2FD: dout <= 8'b00000000; //  765 :   0 - 0x0
      12'h2FE: dout <= 8'b00000000; //  766 :   0 - 0x0
      12'h2FF: dout <= 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout <= 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      12'h301: dout <= 8'b00000000; //  769 :   0 - 0x0
      12'h302: dout <= 8'b00000000; //  770 :   0 - 0x0
      12'h303: dout <= 8'b00000000; //  771 :   0 - 0x0
      12'h304: dout <= 8'b00000000; //  772 :   0 - 0x0
      12'h305: dout <= 8'b00000001; //  773 :   1 - 0x1
      12'h306: dout <= 8'b00011110; //  774 :  30 - 0x1e
      12'h307: dout <= 8'b00111011; //  775 :  59 - 0x3b
      12'h308: dout <= 8'b00000000; //  776 :   0 - 0x0 -- Sprite 0x61
      12'h309: dout <= 8'b00000000; //  777 :   0 - 0x0
      12'h30A: dout <= 8'b00001100; //  778 :  12 - 0xc
      12'h30B: dout <= 8'b00111100; //  779 :  60 - 0x3c
      12'h30C: dout <= 8'b11010000; //  780 : 208 - 0xd0
      12'h30D: dout <= 8'b00010000; //  781 :  16 - 0x10
      12'h30E: dout <= 8'b00100000; //  782 :  32 - 0x20
      12'h30F: dout <= 8'b01000000; //  783 :  64 - 0x40
      12'h310: dout <= 8'b00111110; //  784 :  62 - 0x3e -- Sprite 0x62
      12'h311: dout <= 8'b00101101; //  785 :  45 - 0x2d
      12'h312: dout <= 8'b00110101; //  786 :  53 - 0x35
      12'h313: dout <= 8'b00011101; //  787 :  29 - 0x1d
      12'h314: dout <= 8'b00000001; //  788 :   1 - 0x1
      12'h315: dout <= 8'b00000000; //  789 :   0 - 0x0
      12'h316: dout <= 8'b00000000; //  790 :   0 - 0x0
      12'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout <= 8'b10110000; //  792 : 176 - 0xb0 -- Sprite 0x63
      12'h319: dout <= 8'b10111000; //  793 : 184 - 0xb8
      12'h31A: dout <= 8'b11111000; //  794 : 248 - 0xf8
      12'h31B: dout <= 8'b01111000; //  795 : 120 - 0x78
      12'h31C: dout <= 8'b10011000; //  796 : 152 - 0x98
      12'h31D: dout <= 8'b11110000; //  797 : 240 - 0xf0
      12'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      12'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout <= 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x64
      12'h321: dout <= 8'b00000000; //  801 :   0 - 0x0
      12'h322: dout <= 8'b00000111; //  802 :   7 - 0x7
      12'h323: dout <= 8'b00000011; //  803 :   3 - 0x3
      12'h324: dout <= 8'b00001101; //  804 :  13 - 0xd
      12'h325: dout <= 8'b00011110; //  805 :  30 - 0x1e
      12'h326: dout <= 8'b00010111; //  806 :  23 - 0x17
      12'h327: dout <= 8'b00011101; //  807 :  29 - 0x1d
      12'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- Sprite 0x65
      12'h329: dout <= 8'b10000000; //  809 : 128 - 0x80
      12'h32A: dout <= 8'b01110000; //  810 : 112 - 0x70
      12'h32B: dout <= 8'b11100000; //  811 : 224 - 0xe0
      12'h32C: dout <= 8'b11011000; //  812 : 216 - 0xd8
      12'h32D: dout <= 8'b10111100; //  813 : 188 - 0xbc
      12'h32E: dout <= 8'b01110100; //  814 : 116 - 0x74
      12'h32F: dout <= 8'b11011100; //  815 : 220 - 0xdc
      12'h330: dout <= 8'b00011111; //  816 :  31 - 0x1f -- Sprite 0x66
      12'h331: dout <= 8'b00001011; //  817 :  11 - 0xb
      12'h332: dout <= 8'b00001111; //  818 :  15 - 0xf
      12'h333: dout <= 8'b00000101; //  819 :   5 - 0x5
      12'h334: dout <= 8'b00000011; //  820 :   3 - 0x3
      12'h335: dout <= 8'b00000001; //  821 :   1 - 0x1
      12'h336: dout <= 8'b00000000; //  822 :   0 - 0x0
      12'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      12'h338: dout <= 8'b11111100; //  824 : 252 - 0xfc -- Sprite 0x67
      12'h339: dout <= 8'b01101000; //  825 : 104 - 0x68
      12'h33A: dout <= 8'b11111000; //  826 : 248 - 0xf8
      12'h33B: dout <= 8'b10110000; //  827 : 176 - 0xb0
      12'h33C: dout <= 8'b11100000; //  828 : 224 - 0xe0
      12'h33D: dout <= 8'b10000000; //  829 : 128 - 0x80
      12'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      12'h341: dout <= 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout <= 8'b00000000; //  834 :   0 - 0x0
      12'h343: dout <= 8'b00000000; //  835 :   0 - 0x0
      12'h344: dout <= 8'b00000000; //  836 :   0 - 0x0
      12'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      12'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout <= 8'b00000000; //  840 :   0 - 0x0 -- Sprite 0x69
      12'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout <= 8'b00000000; //  842 :   0 - 0x0
      12'h34B: dout <= 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout <= 8'b00000000; //  844 :   0 - 0x0
      12'h34D: dout <= 8'b00000000; //  845 :   0 - 0x0
      12'h34E: dout <= 8'b00000000; //  846 :   0 - 0x0
      12'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      12'h351: dout <= 8'b00000000; //  849 :   0 - 0x0
      12'h352: dout <= 8'b00000000; //  850 :   0 - 0x0
      12'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      12'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      12'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout <= 8'b00000000; //  856 :   0 - 0x0 -- Sprite 0x6b
      12'h359: dout <= 8'b00000000; //  857 :   0 - 0x0
      12'h35A: dout <= 8'b00000000; //  858 :   0 - 0x0
      12'h35B: dout <= 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout <= 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x6c
      12'h361: dout <= 8'b00000000; //  865 :   0 - 0x0
      12'h362: dout <= 8'b00000001; //  866 :   1 - 0x1
      12'h363: dout <= 8'b00011101; //  867 :  29 - 0x1d
      12'h364: dout <= 8'b00111110; //  868 :  62 - 0x3e
      12'h365: dout <= 8'b00111111; //  869 :  63 - 0x3f
      12'h366: dout <= 8'b00111111; //  870 :  63 - 0x3f
      12'h367: dout <= 8'b00111111; //  871 :  63 - 0x3f
      12'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      12'h369: dout <= 8'b10000000; //  873 : 128 - 0x80
      12'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout <= 8'b01110000; //  875 : 112 - 0x70
      12'h36C: dout <= 8'b11111000; //  876 : 248 - 0xf8
      12'h36D: dout <= 8'b11111100; //  877 : 252 - 0xfc
      12'h36E: dout <= 8'b11111100; //  878 : 252 - 0xfc
      12'h36F: dout <= 8'b11111100; //  879 : 252 - 0xfc
      12'h370: dout <= 8'b00111111; //  880 :  63 - 0x3f -- Sprite 0x6e
      12'h371: dout <= 8'b00111111; //  881 :  63 - 0x3f
      12'h372: dout <= 8'b00011111; //  882 :  31 - 0x1f
      12'h373: dout <= 8'b00011111; //  883 :  31 - 0x1f
      12'h374: dout <= 8'b00001111; //  884 :  15 - 0xf
      12'h375: dout <= 8'b00000110; //  885 :   6 - 0x6
      12'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout <= 8'b11101100; //  888 : 236 - 0xec -- Sprite 0x6f
      12'h379: dout <= 8'b11101100; //  889 : 236 - 0xec
      12'h37A: dout <= 8'b11011000; //  890 : 216 - 0xd8
      12'h37B: dout <= 8'b11111000; //  891 : 248 - 0xf8
      12'h37C: dout <= 8'b11110000; //  892 : 240 - 0xf0
      12'h37D: dout <= 8'b11100000; //  893 : 224 - 0xe0
      12'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x70
      12'h381: dout <= 8'b00000100; //  897 :   4 - 0x4
      12'h382: dout <= 8'b00000011; //  898 :   3 - 0x3
      12'h383: dout <= 8'b00000000; //  899 :   0 - 0x0
      12'h384: dout <= 8'b00000001; //  900 :   1 - 0x1
      12'h385: dout <= 8'b00000111; //  901 :   7 - 0x7
      12'h386: dout <= 8'b00001111; //  902 :  15 - 0xf
      12'h387: dout <= 8'b00001100; //  903 :  12 - 0xc
      12'h388: dout <= 8'b00000000; //  904 :   0 - 0x0 -- Sprite 0x71
      12'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout <= 8'b11100000; //  906 : 224 - 0xe0
      12'h38B: dout <= 8'b10000000; //  907 : 128 - 0x80
      12'h38C: dout <= 8'b01000000; //  908 :  64 - 0x40
      12'h38D: dout <= 8'b11110000; //  909 : 240 - 0xf0
      12'h38E: dout <= 8'b10011000; //  910 : 152 - 0x98
      12'h38F: dout <= 8'b11111000; //  911 : 248 - 0xf8
      12'h390: dout <= 8'b00011111; //  912 :  31 - 0x1f -- Sprite 0x72
      12'h391: dout <= 8'b00010011; //  913 :  19 - 0x13
      12'h392: dout <= 8'b00011111; //  914 :  31 - 0x1f
      12'h393: dout <= 8'b00001111; //  915 :  15 - 0xf
      12'h394: dout <= 8'b00001001; //  916 :   9 - 0x9
      12'h395: dout <= 8'b00000111; //  917 :   7 - 0x7
      12'h396: dout <= 8'b00000001; //  918 :   1 - 0x1
      12'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout <= 8'b11100100; //  920 : 228 - 0xe4 -- Sprite 0x73
      12'h399: dout <= 8'b00111100; //  921 :  60 - 0x3c
      12'h39A: dout <= 8'b11100100; //  922 : 228 - 0xe4
      12'h39B: dout <= 8'b00111000; //  923 :  56 - 0x38
      12'h39C: dout <= 8'b11111000; //  924 : 248 - 0xf8
      12'h39D: dout <= 8'b11110000; //  925 : 240 - 0xf0
      12'h39E: dout <= 8'b11000000; //  926 : 192 - 0xc0
      12'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x74
      12'h3A1: dout <= 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout <= 8'b00000000; //  930 :   0 - 0x0
      12'h3A3: dout <= 8'b00000000; //  931 :   0 - 0x0
      12'h3A4: dout <= 8'b00000000; //  932 :   0 - 0x0
      12'h3A5: dout <= 8'b00000000; //  933 :   0 - 0x0
      12'h3A6: dout <= 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0 -- Sprite 0x75
      12'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout <= 8'b00000000; //  938 :   0 - 0x0
      12'h3AB: dout <= 8'b00000000; //  939 :   0 - 0x0
      12'h3AC: dout <= 8'b00000000; //  940 :   0 - 0x0
      12'h3AD: dout <= 8'b00000000; //  941 :   0 - 0x0
      12'h3AE: dout <= 8'b00000000; //  942 :   0 - 0x0
      12'h3AF: dout <= 8'b00000000; //  943 :   0 - 0x0
      12'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x76
      12'h3B1: dout <= 8'b00000000; //  945 :   0 - 0x0
      12'h3B2: dout <= 8'b00000000; //  946 :   0 - 0x0
      12'h3B3: dout <= 8'b00000000; //  947 :   0 - 0x0
      12'h3B4: dout <= 8'b00000000; //  948 :   0 - 0x0
      12'h3B5: dout <= 8'b00000000; //  949 :   0 - 0x0
      12'h3B6: dout <= 8'b00000000; //  950 :   0 - 0x0
      12'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout <= 8'b00000000; //  952 :   0 - 0x0 -- Sprite 0x77
      12'h3B9: dout <= 8'b00000000; //  953 :   0 - 0x0
      12'h3BA: dout <= 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout <= 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout <= 8'b00000000; //  956 :   0 - 0x0
      12'h3BD: dout <= 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout <= 8'b00000000; //  958 :   0 - 0x0
      12'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x78
      12'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      12'h3C4: dout <= 8'b00000000; //  964 :   0 - 0x0
      12'h3C5: dout <= 8'b00000000; //  965 :   0 - 0x0
      12'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- Sprite 0x79
      12'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x7a
      12'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      12'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      12'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0 -- Sprite 0x7b
      12'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      12'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      12'h3E1: dout <= 8'b00000001; //  993 :   1 - 0x1
      12'h3E2: dout <= 8'b00000110; //  994 :   6 - 0x6
      12'h3E3: dout <= 8'b00000111; //  995 :   7 - 0x7
      12'h3E4: dout <= 8'b00000111; //  996 :   7 - 0x7
      12'h3E5: dout <= 8'b00000111; //  997 :   7 - 0x7
      12'h3E6: dout <= 8'b00000001; //  998 :   1 - 0x1
      12'h3E7: dout <= 8'b00000011; //  999 :   3 - 0x3
      12'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0 -- Sprite 0x7d
      12'h3E9: dout <= 8'b11000000; // 1001 : 192 - 0xc0
      12'h3EA: dout <= 8'b00110000; // 1002 :  48 - 0x30
      12'h3EB: dout <= 8'b11110000; // 1003 : 240 - 0xf0
      12'h3EC: dout <= 8'b11110000; // 1004 : 240 - 0xf0
      12'h3ED: dout <= 8'b11110000; // 1005 : 240 - 0xf0
      12'h3EE: dout <= 8'b01000000; // 1006 :  64 - 0x40
      12'h3EF: dout <= 8'b01000000; // 1007 :  64 - 0x40
      12'h3F0: dout <= 8'b00000001; // 1008 :   1 - 0x1 -- Sprite 0x7e
      12'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout <= 8'b00000001; // 1010 :   1 - 0x1
      12'h3F3: dout <= 8'b00000011; // 1011 :   3 - 0x3
      12'h3F4: dout <= 8'b00000001; // 1012 :   1 - 0x1
      12'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout <= 8'b01000000; // 1016 :  64 - 0x40 -- Sprite 0x7f
      12'h3F9: dout <= 8'b01000000; // 1017 :  64 - 0x40
      12'h3FA: dout <= 8'b01000000; // 1018 :  64 - 0x40
      12'h3FB: dout <= 8'b01000000; // 1019 :  64 - 0x40
      12'h3FC: dout <= 8'b01000000; // 1020 :  64 - 0x40
      12'h3FD: dout <= 8'b10000000; // 1021 : 128 - 0x80
      12'h3FE: dout <= 8'b00000000; // 1022 :   0 - 0x0
      12'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout <= 8'b11111111; // 1024 : 255 - 0xff -- Sprite 0x80
      12'h401: dout <= 8'b11111111; // 1025 : 255 - 0xff
      12'h402: dout <= 8'b11111111; // 1026 : 255 - 0xff
      12'h403: dout <= 8'b11111111; // 1027 : 255 - 0xff
      12'h404: dout <= 8'b11000000; // 1028 : 192 - 0xc0
      12'h405: dout <= 8'b11000000; // 1029 : 192 - 0xc0
      12'h406: dout <= 8'b11000000; // 1030 : 192 - 0xc0
      12'h407: dout <= 8'b11000111; // 1031 : 199 - 0xc7
      12'h408: dout <= 8'b11111111; // 1032 : 255 - 0xff -- Sprite 0x81
      12'h409: dout <= 8'b11111111; // 1033 : 255 - 0xff
      12'h40A: dout <= 8'b11111111; // 1034 : 255 - 0xff
      12'h40B: dout <= 8'b11111111; // 1035 : 255 - 0xff
      12'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      12'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      12'h40F: dout <= 8'b11111111; // 1039 : 255 - 0xff
      12'h410: dout <= 8'b11111111; // 1040 : 255 - 0xff -- Sprite 0x82
      12'h411: dout <= 8'b11111111; // 1041 : 255 - 0xff
      12'h412: dout <= 8'b11111111; // 1042 : 255 - 0xff
      12'h413: dout <= 8'b11111111; // 1043 : 255 - 0xff
      12'h414: dout <= 8'b01111111; // 1044 : 127 - 0x7f
      12'h415: dout <= 8'b00111111; // 1045 :  63 - 0x3f
      12'h416: dout <= 8'b00011111; // 1046 :  31 - 0x1f
      12'h417: dout <= 8'b11001111; // 1047 : 207 - 0xcf
      12'h418: dout <= 8'b11111111; // 1048 : 255 - 0xff -- Sprite 0x83
      12'h419: dout <= 8'b11111111; // 1049 : 255 - 0xff
      12'h41A: dout <= 8'b11111111; // 1050 : 255 - 0xff
      12'h41B: dout <= 8'b11110111; // 1051 : 247 - 0xf7
      12'h41C: dout <= 8'b11110111; // 1052 : 247 - 0xf7
      12'h41D: dout <= 8'b11100010; // 1053 : 226 - 0xe2
      12'h41E: dout <= 8'b11100000; // 1054 : 224 - 0xe0
      12'h41F: dout <= 8'b11000110; // 1055 : 198 - 0xc6
      12'h420: dout <= 8'b11111111; // 1056 : 255 - 0xff -- Sprite 0x84
      12'h421: dout <= 8'b11111111; // 1057 : 255 - 0xff
      12'h422: dout <= 8'b11111111; // 1058 : 255 - 0xff
      12'h423: dout <= 8'b11111111; // 1059 : 255 - 0xff
      12'h424: dout <= 8'b10111111; // 1060 : 191 - 0xbf
      12'h425: dout <= 8'b10111111; // 1061 : 191 - 0xbf
      12'h426: dout <= 8'b00011111; // 1062 :  31 - 0x1f
      12'h427: dout <= 8'b00011111; // 1063 :  31 - 0x1f
      12'h428: dout <= 8'b11111111; // 1064 : 255 - 0xff -- Sprite 0x85
      12'h429: dout <= 8'b11111111; // 1065 : 255 - 0xff
      12'h42A: dout <= 8'b11111111; // 1066 : 255 - 0xff
      12'h42B: dout <= 8'b11111111; // 1067 : 255 - 0xff
      12'h42C: dout <= 8'b11111110; // 1068 : 254 - 0xfe
      12'h42D: dout <= 8'b11111000; // 1069 : 248 - 0xf8
      12'h42E: dout <= 8'b11100000; // 1070 : 224 - 0xe0
      12'h42F: dout <= 8'b11000000; // 1071 : 192 - 0xc0
      12'h430: dout <= 8'b11111111; // 1072 : 255 - 0xff -- Sprite 0x86
      12'h431: dout <= 8'b11111111; // 1073 : 255 - 0xff
      12'h432: dout <= 8'b11111111; // 1074 : 255 - 0xff
      12'h433: dout <= 8'b11111111; // 1075 : 255 - 0xff
      12'h434: dout <= 8'b00000111; // 1076 :   7 - 0x7
      12'h435: dout <= 8'b00000000; // 1077 :   0 - 0x0
      12'h436: dout <= 8'b00111111; // 1078 :  63 - 0x3f
      12'h437: dout <= 8'b11111111; // 1079 : 255 - 0xff
      12'h438: dout <= 8'b11111111; // 1080 : 255 - 0xff -- Sprite 0x87
      12'h439: dout <= 8'b11111111; // 1081 : 255 - 0xff
      12'h43A: dout <= 8'b11111111; // 1082 : 255 - 0xff
      12'h43B: dout <= 8'b11111111; // 1083 : 255 - 0xff
      12'h43C: dout <= 8'b11111111; // 1084 : 255 - 0xff
      12'h43D: dout <= 8'b11111111; // 1085 : 255 - 0xff
      12'h43E: dout <= 8'b00111111; // 1086 :  63 - 0x3f
      12'h43F: dout <= 8'b11001111; // 1087 : 207 - 0xcf
      12'h440: dout <= 8'b11111111; // 1088 : 255 - 0xff -- Sprite 0x88
      12'h441: dout <= 8'b11111111; // 1089 : 255 - 0xff
      12'h442: dout <= 8'b11111111; // 1090 : 255 - 0xff
      12'h443: dout <= 8'b11111111; // 1091 : 255 - 0xff
      12'h444: dout <= 8'b11111111; // 1092 : 255 - 0xff
      12'h445: dout <= 8'b11111111; // 1093 : 255 - 0xff
      12'h446: dout <= 8'b11111111; // 1094 : 255 - 0xff
      12'h447: dout <= 8'b11111111; // 1095 : 255 - 0xff
      12'h448: dout <= 8'b11111111; // 1096 : 255 - 0xff -- Sprite 0x89
      12'h449: dout <= 8'b11111111; // 1097 : 255 - 0xff
      12'h44A: dout <= 8'b11111111; // 1098 : 255 - 0xff
      12'h44B: dout <= 8'b01110111; // 1099 : 119 - 0x77
      12'h44C: dout <= 8'b00010011; // 1100 :  19 - 0x13
      12'h44D: dout <= 8'b00000001; // 1101 :   1 - 0x1
      12'h44E: dout <= 8'b00010000; // 1102 :  16 - 0x10
      12'h44F: dout <= 8'b00011000; // 1103 :  24 - 0x18
      12'h450: dout <= 8'b11111111; // 1104 : 255 - 0xff -- Sprite 0x8a
      12'h451: dout <= 8'b11111111; // 1105 : 255 - 0xff
      12'h452: dout <= 8'b11111111; // 1106 : 255 - 0xff
      12'h453: dout <= 8'b11111111; // 1107 : 255 - 0xff
      12'h454: dout <= 8'b11111111; // 1108 : 255 - 0xff
      12'h455: dout <= 8'b11111111; // 1109 : 255 - 0xff
      12'h456: dout <= 8'b11111111; // 1110 : 255 - 0xff
      12'h457: dout <= 8'b01111111; // 1111 : 127 - 0x7f
      12'h458: dout <= 8'b11111111; // 1112 : 255 - 0xff -- Sprite 0x8b
      12'h459: dout <= 8'b11111111; // 1113 : 255 - 0xff
      12'h45A: dout <= 8'b11111111; // 1114 : 255 - 0xff
      12'h45B: dout <= 8'b11110111; // 1115 : 247 - 0xf7
      12'h45C: dout <= 8'b11100101; // 1116 : 229 - 0xe5
      12'h45D: dout <= 8'b11000001; // 1117 : 193 - 0xc1
      12'h45E: dout <= 8'b10000100; // 1118 : 132 - 0x84
      12'h45F: dout <= 8'b00001100; // 1119 :  12 - 0xc
      12'h460: dout <= 8'b11111111; // 1120 : 255 - 0xff -- Sprite 0x8c
      12'h461: dout <= 8'b11111111; // 1121 : 255 - 0xff
      12'h462: dout <= 8'b11111111; // 1122 : 255 - 0xff
      12'h463: dout <= 8'b11111111; // 1123 : 255 - 0xff
      12'h464: dout <= 8'b11111111; // 1124 : 255 - 0xff
      12'h465: dout <= 8'b01111111; // 1125 : 127 - 0x7f
      12'h466: dout <= 8'b01111110; // 1126 : 126 - 0x7e
      12'h467: dout <= 8'b01111110; // 1127 : 126 - 0x7e
      12'h468: dout <= 8'b11111111; // 1128 : 255 - 0xff -- Sprite 0x8d
      12'h469: dout <= 8'b11111111; // 1129 : 255 - 0xff
      12'h46A: dout <= 8'b10111111; // 1130 : 191 - 0xbf
      12'h46B: dout <= 8'b10110111; // 1131 : 183 - 0xb7
      12'h46C: dout <= 8'b00010111; // 1132 :  23 - 0x17
      12'h46D: dout <= 8'b00000011; // 1133 :   3 - 0x3
      12'h46E: dout <= 8'b00100011; // 1134 :  35 - 0x23
      12'h46F: dout <= 8'b00100001; // 1135 :  33 - 0x21
      12'h470: dout <= 8'b11111111; // 1136 : 255 - 0xff -- Sprite 0x8e
      12'h471: dout <= 8'b11111111; // 1137 : 255 - 0xff
      12'h472: dout <= 8'b11111011; // 1138 : 251 - 0xfb
      12'h473: dout <= 8'b11111001; // 1139 : 249 - 0xf9
      12'h474: dout <= 8'b11111000; // 1140 : 248 - 0xf8
      12'h475: dout <= 8'b11111000; // 1141 : 248 - 0xf8
      12'h476: dout <= 8'b11111000; // 1142 : 248 - 0xf8
      12'h477: dout <= 8'b11111000; // 1143 : 248 - 0xf8
      12'h478: dout <= 8'b11111111; // 1144 : 255 - 0xff -- Sprite 0x8f
      12'h479: dout <= 8'b11111111; // 1145 : 255 - 0xff
      12'h47A: dout <= 8'b01111000; // 1146 : 120 - 0x78
      12'h47B: dout <= 8'b00111000; // 1147 :  56 - 0x38
      12'h47C: dout <= 8'b00011000; // 1148 :  24 - 0x18
      12'h47D: dout <= 8'b00001000; // 1149 :   8 - 0x8
      12'h47E: dout <= 8'b10000000; // 1150 : 128 - 0x80
      12'h47F: dout <= 8'b11000000; // 1151 : 192 - 0xc0
      12'h480: dout <= 8'b11111111; // 1152 : 255 - 0xff -- Sprite 0x90
      12'h481: dout <= 8'b11111111; // 1153 : 255 - 0xff
      12'h482: dout <= 8'b00000001; // 1154 :   1 - 0x1
      12'h483: dout <= 8'b00000001; // 1155 :   1 - 0x1
      12'h484: dout <= 8'b00000001; // 1156 :   1 - 0x1
      12'h485: dout <= 8'b00000000; // 1157 :   0 - 0x0
      12'h486: dout <= 8'b11111111; // 1158 : 255 - 0xff
      12'h487: dout <= 8'b11111111; // 1159 : 255 - 0xff
      12'h488: dout <= 8'b11111111; // 1160 : 255 - 0xff -- Sprite 0x91
      12'h489: dout <= 8'b11111111; // 1161 : 255 - 0xff
      12'h48A: dout <= 8'b11111111; // 1162 : 255 - 0xff
      12'h48B: dout <= 8'b11111111; // 1163 : 255 - 0xff
      12'h48C: dout <= 8'b11111111; // 1164 : 255 - 0xff
      12'h48D: dout <= 8'b11111111; // 1165 : 255 - 0xff
      12'h48E: dout <= 8'b01111111; // 1166 : 127 - 0x7f
      12'h48F: dout <= 8'b00111111; // 1167 :  63 - 0x3f
      12'h490: dout <= 8'b11000111; // 1168 : 199 - 0xc7 -- Sprite 0x92
      12'h491: dout <= 8'b11000111; // 1169 : 199 - 0xc7
      12'h492: dout <= 8'b11000111; // 1170 : 199 - 0xc7
      12'h493: dout <= 8'b11000111; // 1171 : 199 - 0xc7
      12'h494: dout <= 8'b11000111; // 1172 : 199 - 0xc7
      12'h495: dout <= 8'b11000111; // 1173 : 199 - 0xc7
      12'h496: dout <= 8'b11000111; // 1174 : 199 - 0xc7
      12'h497: dout <= 8'b11000111; // 1175 : 199 - 0xc7
      12'h498: dout <= 8'b11111111; // 1176 : 255 - 0xff -- Sprite 0x93
      12'h499: dout <= 8'b11111111; // 1177 : 255 - 0xff
      12'h49A: dout <= 8'b11111111; // 1178 : 255 - 0xff
      12'h49B: dout <= 8'b11111111; // 1179 : 255 - 0xff
      12'h49C: dout <= 8'b11111001; // 1180 : 249 - 0xf9
      12'h49D: dout <= 8'b11111001; // 1181 : 249 - 0xf9
      12'h49E: dout <= 8'b11111111; // 1182 : 255 - 0xff
      12'h49F: dout <= 8'b11111111; // 1183 : 255 - 0xff
      12'h4A0: dout <= 8'b11110111; // 1184 : 247 - 0xf7 -- Sprite 0x94
      12'h4A1: dout <= 8'b11111011; // 1185 : 251 - 0xfb
      12'h4A2: dout <= 8'b11111011; // 1186 : 251 - 0xfb
      12'h4A3: dout <= 8'b11111101; // 1187 : 253 - 0xfd
      12'h4A4: dout <= 8'b11111100; // 1188 : 252 - 0xfc
      12'h4A5: dout <= 8'b11111100; // 1189 : 252 - 0xfc
      12'h4A6: dout <= 8'b01111100; // 1190 : 124 - 0x7c
      12'h4A7: dout <= 8'b01111100; // 1191 : 124 - 0x7c
      12'h4A8: dout <= 8'b11000111; // 1192 : 199 - 0xc7 -- Sprite 0x95
      12'h4A9: dout <= 8'b10001111; // 1193 : 143 - 0x8f
      12'h4AA: dout <= 8'b10001111; // 1194 : 143 - 0x8f
      12'h4AB: dout <= 8'b00011111; // 1195 :  31 - 0x1f
      12'h4AC: dout <= 8'b00011111; // 1196 :  31 - 0x1f
      12'h4AD: dout <= 8'b00111111; // 1197 :  63 - 0x3f
      12'h4AE: dout <= 8'b00111111; // 1198 :  63 - 0x3f
      12'h4AF: dout <= 8'b01111111; // 1199 : 127 - 0x7f
      12'h4B0: dout <= 8'b00001111; // 1200 :  15 - 0xf -- Sprite 0x96
      12'h4B1: dout <= 8'b00001111; // 1201 :  15 - 0xf
      12'h4B2: dout <= 8'b10000111; // 1202 : 135 - 0x87
      12'h4B3: dout <= 8'b10000111; // 1203 : 135 - 0x87
      12'h4B4: dout <= 8'b11000010; // 1204 : 194 - 0xc2
      12'h4B5: dout <= 8'b11000010; // 1205 : 194 - 0xc2
      12'h4B6: dout <= 8'b11100000; // 1206 : 224 - 0xe0
      12'h4B7: dout <= 8'b11100000; // 1207 : 224 - 0xe0
      12'h4B8: dout <= 8'b10000011; // 1208 : 131 - 0x83 -- Sprite 0x97
      12'h4B9: dout <= 8'b10001111; // 1209 : 143 - 0x8f
      12'h4BA: dout <= 8'b00001111; // 1210 :  15 - 0xf
      12'h4BB: dout <= 8'b00011111; // 1211 :  31 - 0x1f
      12'h4BC: dout <= 8'b00011111; // 1212 :  31 - 0x1f
      12'h4BD: dout <= 8'b00111111; // 1213 :  63 - 0x3f
      12'h4BE: dout <= 8'b00111111; // 1214 :  63 - 0x3f
      12'h4BF: dout <= 8'b00111111; // 1215 :  63 - 0x3f
      12'h4C0: dout <= 8'b11111111; // 1216 : 255 - 0xff -- Sprite 0x98
      12'h4C1: dout <= 8'b11111111; // 1217 : 255 - 0xff
      12'h4C2: dout <= 8'b11111111; // 1218 : 255 - 0xff
      12'h4C3: dout <= 8'b11111110; // 1219 : 254 - 0xfe
      12'h4C4: dout <= 8'b11111001; // 1220 : 249 - 0xf9
      12'h4C5: dout <= 8'b11100111; // 1221 : 231 - 0xe7
      12'h4C6: dout <= 8'b11111100; // 1222 : 252 - 0xfc
      12'h4C7: dout <= 8'b11110000; // 1223 : 240 - 0xf0
      12'h4C8: dout <= 8'b11110111; // 1224 : 247 - 0xf7 -- Sprite 0x99
      12'h4C9: dout <= 8'b11111011; // 1225 : 251 - 0xfb
      12'h4CA: dout <= 8'b11111011; // 1226 : 251 - 0xfb
      12'h4CB: dout <= 8'b01110011; // 1227 : 115 - 0x73
      12'h4CC: dout <= 8'b11000001; // 1228 : 193 - 0xc1
      12'h4CD: dout <= 8'b00000011; // 1229 :   3 - 0x3
      12'h4CE: dout <= 8'b00001111; // 1230 :  15 - 0xf
      12'h4CF: dout <= 8'b00111111; // 1231 :  63 - 0x3f
      12'h4D0: dout <= 8'b11111111; // 1232 : 255 - 0xff -- Sprite 0x9a
      12'h4D1: dout <= 8'b11111111; // 1233 : 255 - 0xff
      12'h4D2: dout <= 8'b11111111; // 1234 : 255 - 0xff
      12'h4D3: dout <= 8'b10000000; // 1235 : 128 - 0x80
      12'h4D4: dout <= 8'b10000000; // 1236 : 128 - 0x80
      12'h4D5: dout <= 8'b10000000; // 1237 : 128 - 0x80
      12'h4D6: dout <= 8'b10001111; // 1238 : 143 - 0x8f
      12'h4D7: dout <= 8'b10001111; // 1239 : 143 - 0x8f
      12'h4D8: dout <= 8'b11111111; // 1240 : 255 - 0xff -- Sprite 0x9b
      12'h4D9: dout <= 8'b11111111; // 1241 : 255 - 0xff
      12'h4DA: dout <= 8'b11111111; // 1242 : 255 - 0xff
      12'h4DB: dout <= 8'b00001111; // 1243 :  15 - 0xf
      12'h4DC: dout <= 8'b00001111; // 1244 :  15 - 0xf
      12'h4DD: dout <= 8'b00000111; // 1245 :   7 - 0x7
      12'h4DE: dout <= 8'b11110111; // 1246 : 247 - 0xf7
      12'h4DF: dout <= 8'b11110001; // 1247 : 241 - 0xf1
      12'h4E0: dout <= 8'b00011100; // 1248 :  28 - 0x1c -- Sprite 0x9c
      12'h4E1: dout <= 8'b00011110; // 1249 :  30 - 0x1e
      12'h4E2: dout <= 8'b00011111; // 1250 :  31 - 0x1f
      12'h4E3: dout <= 8'b00011111; // 1251 :  31 - 0x1f
      12'h4E4: dout <= 8'b00011111; // 1252 :  31 - 0x1f
      12'h4E5: dout <= 8'b00011111; // 1253 :  31 - 0x1f
      12'h4E6: dout <= 8'b00011111; // 1254 :  31 - 0x1f
      12'h4E7: dout <= 8'b00011111; // 1255 :  31 - 0x1f
      12'h4E8: dout <= 8'b00111110; // 1256 :  62 - 0x3e -- Sprite 0x9d
      12'h4E9: dout <= 8'b00011100; // 1257 :  28 - 0x1c
      12'h4EA: dout <= 8'b00001000; // 1258 :   8 - 0x8
      12'h4EB: dout <= 8'b10000000; // 1259 : 128 - 0x80
      12'h4EC: dout <= 8'b11000001; // 1260 : 193 - 0xc1
      12'h4ED: dout <= 8'b11100011; // 1261 : 227 - 0xe3
      12'h4EE: dout <= 8'b11110111; // 1262 : 247 - 0xf7
      12'h4EF: dout <= 8'b11111111; // 1263 : 255 - 0xff
      12'h4F0: dout <= 8'b00011100; // 1264 :  28 - 0x1c -- Sprite 0x9e
      12'h4F1: dout <= 8'b00111100; // 1265 :  60 - 0x3c
      12'h4F2: dout <= 8'b01111100; // 1266 : 124 - 0x7c
      12'h4F3: dout <= 8'b11111100; // 1267 : 252 - 0xfc
      12'h4F4: dout <= 8'b11111100; // 1268 : 252 - 0xfc
      12'h4F5: dout <= 8'b11111100; // 1269 : 252 - 0xfc
      12'h4F6: dout <= 8'b11111100; // 1270 : 252 - 0xfc
      12'h4F7: dout <= 8'b11111100; // 1271 : 252 - 0xfc
      12'h4F8: dout <= 8'b01111100; // 1272 : 124 - 0x7c -- Sprite 0x9f
      12'h4F9: dout <= 8'b01111100; // 1273 : 124 - 0x7c
      12'h4FA: dout <= 8'b01111000; // 1274 : 120 - 0x78
      12'h4FB: dout <= 8'b01111000; // 1275 : 120 - 0x78
      12'h4FC: dout <= 8'b01110001; // 1276 : 113 - 0x71
      12'h4FD: dout <= 8'b01110001; // 1277 : 113 - 0x71
      12'h4FE: dout <= 8'b01100011; // 1278 :  99 - 0x63
      12'h4FF: dout <= 8'b01100011; // 1279 :  99 - 0x63
      12'h500: dout <= 8'b01110001; // 1280 : 113 - 0x71 -- Sprite 0xa0
      12'h501: dout <= 8'b01110000; // 1281 : 112 - 0x70
      12'h502: dout <= 8'b11111000; // 1282 : 248 - 0xf8
      12'h503: dout <= 8'b11111000; // 1283 : 248 - 0xf8
      12'h504: dout <= 8'b11111100; // 1284 : 252 - 0xfc
      12'h505: dout <= 8'b11111100; // 1285 : 252 - 0xfc
      12'h506: dout <= 8'b11111110; // 1286 : 254 - 0xfe
      12'h507: dout <= 8'b11111110; // 1287 : 254 - 0xfe
      12'h508: dout <= 8'b11111000; // 1288 : 248 - 0xf8 -- Sprite 0xa1
      12'h509: dout <= 8'b11111000; // 1289 : 248 - 0xf8
      12'h50A: dout <= 8'b11111000; // 1290 : 248 - 0xf8
      12'h50B: dout <= 8'b01111000; // 1291 : 120 - 0x78
      12'h50C: dout <= 8'b01111000; // 1292 : 120 - 0x78
      12'h50D: dout <= 8'b00111000; // 1293 :  56 - 0x38
      12'h50E: dout <= 8'b00111000; // 1294 :  56 - 0x38
      12'h50F: dout <= 8'b00011000; // 1295 :  24 - 0x18
      12'h510: dout <= 8'b11100000; // 1296 : 224 - 0xe0 -- Sprite 0xa2
      12'h511: dout <= 8'b11110000; // 1297 : 240 - 0xf0
      12'h512: dout <= 8'b11111000; // 1298 : 248 - 0xf8
      12'h513: dout <= 8'b11111000; // 1299 : 248 - 0xf8
      12'h514: dout <= 8'b11111100; // 1300 : 252 - 0xfc
      12'h515: dout <= 8'b11111100; // 1301 : 252 - 0xfc
      12'h516: dout <= 8'b11111110; // 1302 : 254 - 0xfe
      12'h517: dout <= 8'b11111111; // 1303 : 255 - 0xff
      12'h518: dout <= 8'b11111111; // 1304 : 255 - 0xff -- Sprite 0xa3
      12'h519: dout <= 8'b11111111; // 1305 : 255 - 0xff
      12'h51A: dout <= 8'b11111111; // 1306 : 255 - 0xff
      12'h51B: dout <= 8'b11111111; // 1307 : 255 - 0xff
      12'h51C: dout <= 8'b11111111; // 1308 : 255 - 0xff
      12'h51D: dout <= 8'b11111111; // 1309 : 255 - 0xff
      12'h51E: dout <= 8'b11111111; // 1310 : 255 - 0xff
      12'h51F: dout <= 8'b11111111; // 1311 : 255 - 0xff
      12'h520: dout <= 8'b00011111; // 1312 :  31 - 0x1f -- Sprite 0xa4
      12'h521: dout <= 8'b00011111; // 1313 :  31 - 0x1f
      12'h522: dout <= 8'b00011111; // 1314 :  31 - 0x1f
      12'h523: dout <= 8'b00011111; // 1315 :  31 - 0x1f
      12'h524: dout <= 8'b00011111; // 1316 :  31 - 0x1f
      12'h525: dout <= 8'b00011111; // 1317 :  31 - 0x1f
      12'h526: dout <= 8'b00011111; // 1318 :  31 - 0x1f
      12'h527: dout <= 8'b00011111; // 1319 :  31 - 0x1f
      12'h528: dout <= 8'b11111000; // 1320 : 248 - 0xf8 -- Sprite 0xa5
      12'h529: dout <= 8'b11111111; // 1321 : 255 - 0xff
      12'h52A: dout <= 8'b11111111; // 1322 : 255 - 0xff
      12'h52B: dout <= 8'b11111000; // 1323 : 248 - 0xf8
      12'h52C: dout <= 8'b11111000; // 1324 : 248 - 0xf8
      12'h52D: dout <= 8'b11111000; // 1325 : 248 - 0xf8
      12'h52E: dout <= 8'b11111000; // 1326 : 248 - 0xf8
      12'h52F: dout <= 8'b11111000; // 1327 : 248 - 0xf8
      12'h530: dout <= 8'b11111100; // 1328 : 252 - 0xfc -- Sprite 0xa6
      12'h531: dout <= 8'b11111000; // 1329 : 248 - 0xf8
      12'h532: dout <= 8'b11110000; // 1330 : 240 - 0xf0
      12'h533: dout <= 8'b00000001; // 1331 :   1 - 0x1
      12'h534: dout <= 8'b00000001; // 1332 :   1 - 0x1
      12'h535: dout <= 8'b00000011; // 1333 :   3 - 0x3
      12'h536: dout <= 8'b11000011; // 1334 : 195 - 0xc3
      12'h537: dout <= 8'b10000111; // 1335 : 135 - 0x87
      12'h538: dout <= 8'b01111111; // 1336 : 127 - 0x7f -- Sprite 0xa7
      12'h539: dout <= 8'b11111001; // 1337 : 249 - 0xf9
      12'h53A: dout <= 8'b11111001; // 1338 : 249 - 0xf9
      12'h53B: dout <= 8'b11111111; // 1339 : 255 - 0xff
      12'h53C: dout <= 8'b11111110; // 1340 : 254 - 0xfe
      12'h53D: dout <= 8'b11111100; // 1341 : 252 - 0xfc
      12'h53E: dout <= 8'b11111111; // 1342 : 255 - 0xff
      12'h53F: dout <= 8'b11111111; // 1343 : 255 - 0xff
      12'h540: dout <= 8'b11110000; // 1344 : 240 - 0xf0 -- Sprite 0xa8
      12'h541: dout <= 8'b11110000; // 1345 : 240 - 0xf0
      12'h542: dout <= 8'b11111000; // 1346 : 248 - 0xf8
      12'h543: dout <= 8'b01111000; // 1347 : 120 - 0x78
      12'h544: dout <= 8'b11111100; // 1348 : 252 - 0xfc
      12'h545: dout <= 8'b11110100; // 1349 : 244 - 0xf4
      12'h546: dout <= 8'b11110110; // 1350 : 246 - 0xf6
      12'h547: dout <= 8'b11111010; // 1351 : 250 - 0xfa
      12'h548: dout <= 8'b00111111; // 1352 :  63 - 0x3f -- Sprite 0xa9
      12'h549: dout <= 8'b00111111; // 1353 :  63 - 0x3f
      12'h54A: dout <= 8'b00111111; // 1354 :  63 - 0x3f
      12'h54B: dout <= 8'b00111111; // 1355 :  63 - 0x3f
      12'h54C: dout <= 8'b00111111; // 1356 :  63 - 0x3f
      12'h54D: dout <= 8'b00011111; // 1357 :  31 - 0x1f
      12'h54E: dout <= 8'b00001111; // 1358 :  15 - 0xf
      12'h54F: dout <= 8'b00000111; // 1359 :   7 - 0x7
      12'h550: dout <= 8'b11100000; // 1360 : 224 - 0xe0 -- Sprite 0xaa
      12'h551: dout <= 8'b11111000; // 1361 : 248 - 0xf8
      12'h552: dout <= 8'b11111111; // 1362 : 255 - 0xff
      12'h553: dout <= 8'b11110011; // 1363 : 243 - 0xf3
      12'h554: dout <= 8'b11111100; // 1364 : 252 - 0xfc
      12'h555: dout <= 8'b11111111; // 1365 : 255 - 0xff
      12'h556: dout <= 8'b11111111; // 1366 : 255 - 0xff
      12'h557: dout <= 8'b11111111; // 1367 : 255 - 0xff
      12'h558: dout <= 8'b11111111; // 1368 : 255 - 0xff -- Sprite 0xab
      12'h559: dout <= 8'b11111111; // 1369 : 255 - 0xff
      12'h55A: dout <= 8'b00111111; // 1370 :  63 - 0x3f
      12'h55B: dout <= 8'b11001111; // 1371 : 207 - 0xcf
      12'h55C: dout <= 8'b11110011; // 1372 : 243 - 0xf3
      12'h55D: dout <= 8'b00111101; // 1373 :  61 - 0x3d
      12'h55E: dout <= 8'b11011000; // 1374 : 216 - 0xd8
      12'h55F: dout <= 8'b10110000; // 1375 : 176 - 0xb0
      12'h560: dout <= 8'b10001111; // 1376 : 143 - 0x8f -- Sprite 0xac
      12'h561: dout <= 8'b11101111; // 1377 : 239 - 0xef
      12'h562: dout <= 8'b11100000; // 1378 : 224 - 0xe0
      12'h563: dout <= 8'b11111000; // 1379 : 248 - 0xf8
      12'h564: dout <= 8'b11111000; // 1380 : 248 - 0xf8
      12'h565: dout <= 8'b11111111; // 1381 : 255 - 0xff
      12'h566: dout <= 8'b11111111; // 1382 : 255 - 0xff
      12'h567: dout <= 8'b11111111; // 1383 : 255 - 0xff
      12'h568: dout <= 8'b11110001; // 1384 : 241 - 0xf1 -- Sprite 0xad
      12'h569: dout <= 8'b11110001; // 1385 : 241 - 0xf1
      12'h56A: dout <= 8'b00000001; // 1386 :   1 - 0x1
      12'h56B: dout <= 8'b00000001; // 1387 :   1 - 0x1
      12'h56C: dout <= 8'b00000001; // 1388 :   1 - 0x1
      12'h56D: dout <= 8'b11111111; // 1389 : 255 - 0xff
      12'h56E: dout <= 8'b11111111; // 1390 : 255 - 0xff
      12'h56F: dout <= 8'b11111111; // 1391 : 255 - 0xff
      12'h570: dout <= 8'b00011111; // 1392 :  31 - 0x1f -- Sprite 0xae
      12'h571: dout <= 8'b00011111; // 1393 :  31 - 0x1f
      12'h572: dout <= 8'b00011111; // 1394 :  31 - 0x1f
      12'h573: dout <= 8'b00011111; // 1395 :  31 - 0x1f
      12'h574: dout <= 8'b00011111; // 1396 :  31 - 0x1f
      12'h575: dout <= 8'b00011111; // 1397 :  31 - 0x1f
      12'h576: dout <= 8'b00011111; // 1398 :  31 - 0x1f
      12'h577: dout <= 8'b00011111; // 1399 :  31 - 0x1f
      12'h578: dout <= 8'b11111100; // 1400 : 252 - 0xfc -- Sprite 0xaf
      12'h579: dout <= 8'b11111100; // 1401 : 252 - 0xfc
      12'h57A: dout <= 8'b11111100; // 1402 : 252 - 0xfc
      12'h57B: dout <= 8'b11111100; // 1403 : 252 - 0xfc
      12'h57C: dout <= 8'b11110100; // 1404 : 244 - 0xf4
      12'h57D: dout <= 8'b11110100; // 1405 : 244 - 0xf4
      12'h57E: dout <= 8'b11110100; // 1406 : 244 - 0xf4
      12'h57F: dout <= 8'b11110100; // 1407 : 244 - 0xf4
      12'h580: dout <= 8'b00001100; // 1408 :  12 - 0xc -- Sprite 0xb0
      12'h581: dout <= 8'b00011100; // 1409 :  28 - 0x1c
      12'h582: dout <= 8'b00001100; // 1410 :  12 - 0xc
      12'h583: dout <= 8'b00001100; // 1411 :  12 - 0xc
      12'h584: dout <= 8'b00001100; // 1412 :  12 - 0xc
      12'h585: dout <= 8'b00001100; // 1413 :  12 - 0xc
      12'h586: dout <= 8'b00111111; // 1414 :  63 - 0x3f
      12'h587: dout <= 8'b00000000; // 1415 :   0 - 0x0
      12'h588: dout <= 8'b00111110; // 1416 :  62 - 0x3e -- Sprite 0xb1
      12'h589: dout <= 8'b01100011; // 1417 :  99 - 0x63
      12'h58A: dout <= 8'b00000111; // 1418 :   7 - 0x7
      12'h58B: dout <= 8'b00011110; // 1419 :  30 - 0x1e
      12'h58C: dout <= 8'b00111100; // 1420 :  60 - 0x3c
      12'h58D: dout <= 8'b01110000; // 1421 : 112 - 0x70
      12'h58E: dout <= 8'b01111111; // 1422 : 127 - 0x7f
      12'h58F: dout <= 8'b00000000; // 1423 :   0 - 0x0
      12'h590: dout <= 8'b01111110; // 1424 : 126 - 0x7e -- Sprite 0xb2
      12'h591: dout <= 8'b01100011; // 1425 :  99 - 0x63
      12'h592: dout <= 8'b01100011; // 1426 :  99 - 0x63
      12'h593: dout <= 8'b01100011; // 1427 :  99 - 0x63
      12'h594: dout <= 8'b01111110; // 1428 : 126 - 0x7e
      12'h595: dout <= 8'b01100000; // 1429 :  96 - 0x60
      12'h596: dout <= 8'b01100000; // 1430 :  96 - 0x60
      12'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      12'h598: dout <= 8'b01100011; // 1432 :  99 - 0x63 -- Sprite 0xb3
      12'h599: dout <= 8'b01100011; // 1433 :  99 - 0x63
      12'h59A: dout <= 8'b01100011; // 1434 :  99 - 0x63
      12'h59B: dout <= 8'b01100011; // 1435 :  99 - 0x63
      12'h59C: dout <= 8'b01100011; // 1436 :  99 - 0x63
      12'h59D: dout <= 8'b01100011; // 1437 :  99 - 0x63
      12'h59E: dout <= 8'b00111110; // 1438 :  62 - 0x3e
      12'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout <= 8'b01100011; // 1440 :  99 - 0x63 -- Sprite 0xb4
      12'h5A1: dout <= 8'b01100011; // 1441 :  99 - 0x63
      12'h5A2: dout <= 8'b01100011; // 1442 :  99 - 0x63
      12'h5A3: dout <= 8'b01111111; // 1443 : 127 - 0x7f
      12'h5A4: dout <= 8'b01100011; // 1444 :  99 - 0x63
      12'h5A5: dout <= 8'b01100011; // 1445 :  99 - 0x63
      12'h5A6: dout <= 8'b01100011; // 1446 :  99 - 0x63
      12'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      12'h5A8: dout <= 8'b00111111; // 1448 :  63 - 0x3f -- Sprite 0xb5
      12'h5A9: dout <= 8'b00001100; // 1449 :  12 - 0xc
      12'h5AA: dout <= 8'b00001100; // 1450 :  12 - 0xc
      12'h5AB: dout <= 8'b00001100; // 1451 :  12 - 0xc
      12'h5AC: dout <= 8'b00001100; // 1452 :  12 - 0xc
      12'h5AD: dout <= 8'b00001100; // 1453 :  12 - 0xc
      12'h5AE: dout <= 8'b00111111; // 1454 :  63 - 0x3f
      12'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      12'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0xb6
      12'h5B1: dout <= 8'b00000000; // 1457 :   0 - 0x0
      12'h5B2: dout <= 8'b00000000; // 1458 :   0 - 0x0
      12'h5B3: dout <= 8'b01111110; // 1459 : 126 - 0x7e
      12'h5B4: dout <= 8'b00000000; // 1460 :   0 - 0x0
      12'h5B5: dout <= 8'b00000000; // 1461 :   0 - 0x0
      12'h5B6: dout <= 8'b00000000; // 1462 :   0 - 0x0
      12'h5B7: dout <= 8'b00000000; // 1463 :   0 - 0x0
      12'h5B8: dout <= 8'b00111100; // 1464 :  60 - 0x3c -- Sprite 0xb7
      12'h5B9: dout <= 8'b01100110; // 1465 : 102 - 0x66
      12'h5BA: dout <= 8'b01100000; // 1466 :  96 - 0x60
      12'h5BB: dout <= 8'b00111110; // 1467 :  62 - 0x3e
      12'h5BC: dout <= 8'b00000011; // 1468 :   3 - 0x3
      12'h5BD: dout <= 8'b01100011; // 1469 :  99 - 0x63
      12'h5BE: dout <= 8'b00111110; // 1470 :  62 - 0x3e
      12'h5BF: dout <= 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout <= 8'b00011110; // 1472 :  30 - 0x1e -- Sprite 0xb8
      12'h5C1: dout <= 8'b00110011; // 1473 :  51 - 0x33
      12'h5C2: dout <= 8'b01100000; // 1474 :  96 - 0x60
      12'h5C3: dout <= 8'b01100000; // 1475 :  96 - 0x60
      12'h5C4: dout <= 8'b01100000; // 1476 :  96 - 0x60
      12'h5C5: dout <= 8'b00110011; // 1477 :  51 - 0x33
      12'h5C6: dout <= 8'b00011110; // 1478 :  30 - 0x1e
      12'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout <= 8'b00111110; // 1480 :  62 - 0x3e -- Sprite 0xb9
      12'h5C9: dout <= 8'b01100011; // 1481 :  99 - 0x63
      12'h5CA: dout <= 8'b01100011; // 1482 :  99 - 0x63
      12'h5CB: dout <= 8'b01100011; // 1483 :  99 - 0x63
      12'h5CC: dout <= 8'b01100011; // 1484 :  99 - 0x63
      12'h5CD: dout <= 8'b01100011; // 1485 :  99 - 0x63
      12'h5CE: dout <= 8'b00111110; // 1486 :  62 - 0x3e
      12'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout <= 8'b01111110; // 1488 : 126 - 0x7e -- Sprite 0xba
      12'h5D1: dout <= 8'b01100011; // 1489 :  99 - 0x63
      12'h5D2: dout <= 8'b01100011; // 1490 :  99 - 0x63
      12'h5D3: dout <= 8'b01100111; // 1491 : 103 - 0x67
      12'h5D4: dout <= 8'b01111100; // 1492 : 124 - 0x7c
      12'h5D5: dout <= 8'b01101110; // 1493 : 110 - 0x6e
      12'h5D6: dout <= 8'b01100111; // 1494 : 103 - 0x67
      12'h5D7: dout <= 8'b00000000; // 1495 :   0 - 0x0
      12'h5D8: dout <= 8'b01111111; // 1496 : 127 - 0x7f -- Sprite 0xbb
      12'h5D9: dout <= 8'b01100000; // 1497 :  96 - 0x60
      12'h5DA: dout <= 8'b01100000; // 1498 :  96 - 0x60
      12'h5DB: dout <= 8'b01111110; // 1499 : 126 - 0x7e
      12'h5DC: dout <= 8'b01100000; // 1500 :  96 - 0x60
      12'h5DD: dout <= 8'b01100000; // 1501 :  96 - 0x60
      12'h5DE: dout <= 8'b01111111; // 1502 : 127 - 0x7f
      12'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0xbc
      12'h5E1: dout <= 8'b00100010; // 1505 :  34 - 0x22
      12'h5E2: dout <= 8'b01100101; // 1506 : 101 - 0x65
      12'h5E3: dout <= 8'b00100101; // 1507 :  37 - 0x25
      12'h5E4: dout <= 8'b00100101; // 1508 :  37 - 0x25
      12'h5E5: dout <= 8'b01110010; // 1509 : 114 - 0x72
      12'h5E6: dout <= 8'b00000000; // 1510 :   0 - 0x0
      12'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0 -- Sprite 0xbd
      12'h5E9: dout <= 8'b01110010; // 1513 : 114 - 0x72
      12'h5EA: dout <= 8'b01000101; // 1514 :  69 - 0x45
      12'h5EB: dout <= 8'b01100101; // 1515 : 101 - 0x65
      12'h5EC: dout <= 8'b00010101; // 1516 :  21 - 0x15
      12'h5ED: dout <= 8'b01100010; // 1517 :  98 - 0x62
      12'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      12'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout <= 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      12'h5F1: dout <= 8'b01100111; // 1521 : 103 - 0x67
      12'h5F2: dout <= 8'b01010010; // 1522 :  82 - 0x52
      12'h5F3: dout <= 8'b01100010; // 1523 :  98 - 0x62
      12'h5F4: dout <= 8'b01000010; // 1524 :  66 - 0x42
      12'h5F5: dout <= 8'b01000010; // 1525 :  66 - 0x42
      12'h5F6: dout <= 8'b00000000; // 1526 :   0 - 0x0
      12'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      12'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      12'h5F9: dout <= 8'b01100000; // 1529 :  96 - 0x60
      12'h5FA: dout <= 8'b10000000; // 1530 : 128 - 0x80
      12'h5FB: dout <= 8'b01000000; // 1531 :  64 - 0x40
      12'h5FC: dout <= 8'b00100000; // 1532 :  32 - 0x20
      12'h5FD: dout <= 8'b11000110; // 1533 : 198 - 0xc6
      12'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      12'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout <= 8'b01100011; // 1536 :  99 - 0x63 -- Sprite 0xc0
      12'h601: dout <= 8'b01100110; // 1537 : 102 - 0x66
      12'h602: dout <= 8'b01101100; // 1538 : 108 - 0x6c
      12'h603: dout <= 8'b01111000; // 1539 : 120 - 0x78
      12'h604: dout <= 8'b01111100; // 1540 : 124 - 0x7c
      12'h605: dout <= 8'b01100110; // 1541 : 102 - 0x66
      12'h606: dout <= 8'b01100011; // 1542 :  99 - 0x63
      12'h607: dout <= 8'b00000000; // 1543 :   0 - 0x0
      12'h608: dout <= 8'b00111111; // 1544 :  63 - 0x3f -- Sprite 0xc1
      12'h609: dout <= 8'b00001100; // 1545 :  12 - 0xc
      12'h60A: dout <= 8'b00001100; // 1546 :  12 - 0xc
      12'h60B: dout <= 8'b00001100; // 1547 :  12 - 0xc
      12'h60C: dout <= 8'b00001100; // 1548 :  12 - 0xc
      12'h60D: dout <= 8'b00001100; // 1549 :  12 - 0xc
      12'h60E: dout <= 8'b00111111; // 1550 :  63 - 0x3f
      12'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout <= 8'b01100011; // 1552 :  99 - 0x63 -- Sprite 0xc2
      12'h611: dout <= 8'b01110111; // 1553 : 119 - 0x77
      12'h612: dout <= 8'b01111111; // 1554 : 127 - 0x7f
      12'h613: dout <= 8'b01111111; // 1555 : 127 - 0x7f
      12'h614: dout <= 8'b01101011; // 1556 : 107 - 0x6b
      12'h615: dout <= 8'b01100011; // 1557 :  99 - 0x63
      12'h616: dout <= 8'b01100011; // 1558 :  99 - 0x63
      12'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      12'h618: dout <= 8'b00011100; // 1560 :  28 - 0x1c -- Sprite 0xc3
      12'h619: dout <= 8'b00110110; // 1561 :  54 - 0x36
      12'h61A: dout <= 8'b01100011; // 1562 :  99 - 0x63
      12'h61B: dout <= 8'b01100011; // 1563 :  99 - 0x63
      12'h61C: dout <= 8'b01111111; // 1564 : 127 - 0x7f
      12'h61D: dout <= 8'b01100011; // 1565 :  99 - 0x63
      12'h61E: dout <= 8'b01100011; // 1566 :  99 - 0x63
      12'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout <= 8'b00011111; // 1568 :  31 - 0x1f -- Sprite 0xc4
      12'h621: dout <= 8'b00110000; // 1569 :  48 - 0x30
      12'h622: dout <= 8'b01100000; // 1570 :  96 - 0x60
      12'h623: dout <= 8'b01100111; // 1571 : 103 - 0x67
      12'h624: dout <= 8'b01100011; // 1572 :  99 - 0x63
      12'h625: dout <= 8'b00110011; // 1573 :  51 - 0x33
      12'h626: dout <= 8'b00011111; // 1574 :  31 - 0x1f
      12'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout <= 8'b01100011; // 1576 :  99 - 0x63 -- Sprite 0xc5
      12'h629: dout <= 8'b01100011; // 1577 :  99 - 0x63
      12'h62A: dout <= 8'b01100011; // 1578 :  99 - 0x63
      12'h62B: dout <= 8'b01100011; // 1579 :  99 - 0x63
      12'h62C: dout <= 8'b01100011; // 1580 :  99 - 0x63
      12'h62D: dout <= 8'b01100011; // 1581 :  99 - 0x63
      12'h62E: dout <= 8'b00111110; // 1582 :  62 - 0x3e
      12'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout <= 8'b01111110; // 1584 : 126 - 0x7e -- Sprite 0xc6
      12'h631: dout <= 8'b01100011; // 1585 :  99 - 0x63
      12'h632: dout <= 8'b01100011; // 1586 :  99 - 0x63
      12'h633: dout <= 8'b01100111; // 1587 : 103 - 0x67
      12'h634: dout <= 8'b01111100; // 1588 : 124 - 0x7c
      12'h635: dout <= 8'b01101110; // 1589 : 110 - 0x6e
      12'h636: dout <= 8'b01100111; // 1590 : 103 - 0x67
      12'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      12'h638: dout <= 8'b01111111; // 1592 : 127 - 0x7f -- Sprite 0xc7
      12'h639: dout <= 8'b01100000; // 1593 :  96 - 0x60
      12'h63A: dout <= 8'b01100000; // 1594 :  96 - 0x60
      12'h63B: dout <= 8'b01111110; // 1595 : 126 - 0x7e
      12'h63C: dout <= 8'b01100000; // 1596 :  96 - 0x60
      12'h63D: dout <= 8'b01100000; // 1597 :  96 - 0x60
      12'h63E: dout <= 8'b01111111; // 1598 : 127 - 0x7f
      12'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout <= 8'b00110110; // 1600 :  54 - 0x36 -- Sprite 0xc8
      12'h641: dout <= 8'b00110110; // 1601 :  54 - 0x36
      12'h642: dout <= 8'b00010010; // 1602 :  18 - 0x12
      12'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      12'h644: dout <= 8'b00000000; // 1604 :   0 - 0x0
      12'h645: dout <= 8'b00000000; // 1605 :   0 - 0x0
      12'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      12'h647: dout <= 8'b00000000; // 1607 :   0 - 0x0
      12'h648: dout <= 8'b00111110; // 1608 :  62 - 0x3e -- Sprite 0xc9
      12'h649: dout <= 8'b01100011; // 1609 :  99 - 0x63
      12'h64A: dout <= 8'b01100011; // 1610 :  99 - 0x63
      12'h64B: dout <= 8'b01100011; // 1611 :  99 - 0x63
      12'h64C: dout <= 8'b01100011; // 1612 :  99 - 0x63
      12'h64D: dout <= 8'b01100011; // 1613 :  99 - 0x63
      12'h64E: dout <= 8'b00111110; // 1614 :  62 - 0x3e
      12'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout <= 8'b00111100; // 1616 :  60 - 0x3c -- Sprite 0xca
      12'h651: dout <= 8'b01100110; // 1617 : 102 - 0x66
      12'h652: dout <= 8'b01100000; // 1618 :  96 - 0x60
      12'h653: dout <= 8'b00111110; // 1619 :  62 - 0x3e
      12'h654: dout <= 8'b00000011; // 1620 :   3 - 0x3
      12'h655: dout <= 8'b01100011; // 1621 :  99 - 0x63
      12'h656: dout <= 8'b00111110; // 1622 :  62 - 0x3e
      12'h657: dout <= 8'b00000000; // 1623 :   0 - 0x0
      12'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- Sprite 0xcb
      12'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      12'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      12'h65C: dout <= 8'b00000000; // 1628 :   0 - 0x0
      12'h65D: dout <= 8'b00000000; // 1629 :   0 - 0x0
      12'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout <= 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0xcc
      12'h661: dout <= 8'b00000000; // 1633 :   0 - 0x0
      12'h662: dout <= 8'b00000000; // 1634 :   0 - 0x0
      12'h663: dout <= 8'b00000000; // 1635 :   0 - 0x0
      12'h664: dout <= 8'b00000000; // 1636 :   0 - 0x0
      12'h665: dout <= 8'b00000000; // 1637 :   0 - 0x0
      12'h666: dout <= 8'b00000000; // 1638 :   0 - 0x0
      12'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      12'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- Sprite 0xcd
      12'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout <= 8'b00000000; // 1643 :   0 - 0x0
      12'h66C: dout <= 8'b00000000; // 1644 :   0 - 0x0
      12'h66D: dout <= 8'b00000000; // 1645 :   0 - 0x0
      12'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      12'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      12'h670: dout <= 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      12'h671: dout <= 8'b00000000; // 1649 :   0 - 0x0
      12'h672: dout <= 8'b00000000; // 1650 :   0 - 0x0
      12'h673: dout <= 8'b00000000; // 1651 :   0 - 0x0
      12'h674: dout <= 8'b00000000; // 1652 :   0 - 0x0
      12'h675: dout <= 8'b00000000; // 1653 :   0 - 0x0
      12'h676: dout <= 8'b00000000; // 1654 :   0 - 0x0
      12'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      12'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- Sprite 0xcf
      12'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      12'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      12'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      12'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout <= 8'b01000111; // 1664 :  71 - 0x47 -- Sprite 0xd0
      12'h681: dout <= 8'b01000111; // 1665 :  71 - 0x47
      12'h682: dout <= 8'b00001111; // 1666 :  15 - 0xf
      12'h683: dout <= 8'b00001111; // 1667 :  15 - 0xf
      12'h684: dout <= 8'b00011111; // 1668 :  31 - 0x1f
      12'h685: dout <= 8'b00011111; // 1669 :  31 - 0x1f
      12'h686: dout <= 8'b00111111; // 1670 :  63 - 0x3f
      12'h687: dout <= 8'b00111111; // 1671 :  63 - 0x3f
      12'h688: dout <= 8'b11111111; // 1672 : 255 - 0xff -- Sprite 0xd1
      12'h689: dout <= 8'b11001111; // 1673 : 207 - 0xcf
      12'h68A: dout <= 8'b11001111; // 1674 : 207 - 0xcf
      12'h68B: dout <= 8'b11111011; // 1675 : 251 - 0xfb
      12'h68C: dout <= 8'b11110111; // 1676 : 247 - 0xf7
      12'h68D: dout <= 8'b11100111; // 1677 : 231 - 0xe7
      12'h68E: dout <= 8'b11111111; // 1678 : 255 - 0xff
      12'h68F: dout <= 8'b11111111; // 1679 : 255 - 0xff
      12'h690: dout <= 8'b00011000; // 1680 :  24 - 0x18 -- Sprite 0xd2
      12'h691: dout <= 8'b00001000; // 1681 :   8 - 0x8
      12'h692: dout <= 8'b10001000; // 1682 : 136 - 0x88
      12'h693: dout <= 8'b10000000; // 1683 : 128 - 0x80
      12'h694: dout <= 8'b01000000; // 1684 :  64 - 0x40
      12'h695: dout <= 8'b01000000; // 1685 :  64 - 0x40
      12'h696: dout <= 8'b10100000; // 1686 : 160 - 0xa0
      12'h697: dout <= 8'b10100000; // 1687 : 160 - 0xa0
      12'h698: dout <= 8'b11111111; // 1688 : 255 - 0xff -- Sprite 0xd3
      12'h699: dout <= 8'b11111111; // 1689 : 255 - 0xff
      12'h69A: dout <= 8'b11111111; // 1690 : 255 - 0xff
      12'h69B: dout <= 8'b11111111; // 1691 : 255 - 0xff
      12'h69C: dout <= 8'b11111101; // 1692 : 253 - 0xfd
      12'h69D: dout <= 8'b11111101; // 1693 : 253 - 0xfd
      12'h69E: dout <= 8'b11111101; // 1694 : 253 - 0xfd
      12'h69F: dout <= 8'b11111101; // 1695 : 253 - 0xfd
      12'h6A0: dout <= 8'b11000111; // 1696 : 199 - 0xc7 -- Sprite 0xd4
      12'h6A1: dout <= 8'b11110111; // 1697 : 247 - 0xf7
      12'h6A2: dout <= 8'b11110000; // 1698 : 240 - 0xf0
      12'h6A3: dout <= 8'b11111000; // 1699 : 248 - 0xf8
      12'h6A4: dout <= 8'b11111000; // 1700 : 248 - 0xf8
      12'h6A5: dout <= 8'b11111111; // 1701 : 255 - 0xff
      12'h6A6: dout <= 8'b11111111; // 1702 : 255 - 0xff
      12'h6A7: dout <= 8'b11111111; // 1703 : 255 - 0xff
      12'h6A8: dout <= 8'b11111000; // 1704 : 248 - 0xf8 -- Sprite 0xd5
      12'h6A9: dout <= 8'b11111000; // 1705 : 248 - 0xf8
      12'h6AA: dout <= 8'b00000000; // 1706 :   0 - 0x0
      12'h6AB: dout <= 8'b00000000; // 1707 :   0 - 0x0
      12'h6AC: dout <= 8'b00000000; // 1708 :   0 - 0x0
      12'h6AD: dout <= 8'b11111111; // 1709 : 255 - 0xff
      12'h6AE: dout <= 8'b11111111; // 1710 : 255 - 0xff
      12'h6AF: dout <= 8'b11111111; // 1711 : 255 - 0xff
      12'h6B0: dout <= 8'b10001111; // 1712 : 143 - 0x8f -- Sprite 0xd6
      12'h6B1: dout <= 8'b11101111; // 1713 : 239 - 0xef
      12'h6B2: dout <= 8'b11000000; // 1714 : 192 - 0xc0
      12'h6B3: dout <= 8'b11110000; // 1715 : 240 - 0xf0
      12'h6B4: dout <= 8'b11100000; // 1716 : 224 - 0xe0
      12'h6B5: dout <= 8'b11111111; // 1717 : 255 - 0xff
      12'h6B6: dout <= 8'b11111111; // 1718 : 255 - 0xff
      12'h6B7: dout <= 8'b11111111; // 1719 : 255 - 0xff
      12'h6B8: dout <= 8'b11111111; // 1720 : 255 - 0xff -- Sprite 0xd7
      12'h6B9: dout <= 8'b11111111; // 1721 : 255 - 0xff
      12'h6BA: dout <= 8'b00000000; // 1722 :   0 - 0x0
      12'h6BB: dout <= 8'b00000000; // 1723 :   0 - 0x0
      12'h6BC: dout <= 8'b00000000; // 1724 :   0 - 0x0
      12'h6BD: dout <= 8'b11111111; // 1725 : 255 - 0xff
      12'h6BE: dout <= 8'b11111111; // 1726 : 255 - 0xff
      12'h6BF: dout <= 8'b11111111; // 1727 : 255 - 0xff
      12'h6C0: dout <= 8'b11000011; // 1728 : 195 - 0xc3 -- Sprite 0xd8
      12'h6C1: dout <= 8'b11111111; // 1729 : 255 - 0xff
      12'h6C2: dout <= 8'b00000000; // 1730 :   0 - 0x0
      12'h6C3: dout <= 8'b00000000; // 1731 :   0 - 0x0
      12'h6C4: dout <= 8'b00000000; // 1732 :   0 - 0x0
      12'h6C5: dout <= 8'b11111111; // 1733 : 255 - 0xff
      12'h6C6: dout <= 8'b11111111; // 1734 : 255 - 0xff
      12'h6C7: dout <= 8'b11111111; // 1735 : 255 - 0xff
      12'h6C8: dout <= 8'b00000011; // 1736 :   3 - 0x3 -- Sprite 0xd9
      12'h6C9: dout <= 8'b10000001; // 1737 : 129 - 0x81
      12'h6CA: dout <= 8'b00000000; // 1738 :   0 - 0x0
      12'h6CB: dout <= 8'b00000000; // 1739 :   0 - 0x0
      12'h6CC: dout <= 8'b00000011; // 1740 :   3 - 0x3
      12'h6CD: dout <= 8'b11111111; // 1741 : 255 - 0xff
      12'h6CE: dout <= 8'b11111111; // 1742 : 255 - 0xff
      12'h6CF: dout <= 8'b11111111; // 1743 : 255 - 0xff
      12'h6D0: dout <= 8'b11111111; // 1744 : 255 - 0xff -- Sprite 0xda
      12'h6D1: dout <= 8'b11111111; // 1745 : 255 - 0xff
      12'h6D2: dout <= 8'b01111110; // 1746 : 126 - 0x7e
      12'h6D3: dout <= 8'b00000000; // 1747 :   0 - 0x0
      12'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      12'h6D5: dout <= 8'b11100000; // 1749 : 224 - 0xe0
      12'h6D6: dout <= 8'b11111111; // 1750 : 255 - 0xff
      12'h6D7: dout <= 8'b11111111; // 1751 : 255 - 0xff
      12'h6D8: dout <= 8'b01100001; // 1752 :  97 - 0x61 -- Sprite 0xdb
      12'h6D9: dout <= 8'b11000011; // 1753 : 195 - 0xc3
      12'h6DA: dout <= 8'b00000111; // 1754 :   7 - 0x7
      12'h6DB: dout <= 8'b00001111; // 1755 :  15 - 0xf
      12'h6DC: dout <= 8'b00011111; // 1756 :  31 - 0x1f
      12'h6DD: dout <= 8'b01111111; // 1757 : 127 - 0x7f
      12'h6DE: dout <= 8'b11111111; // 1758 : 255 - 0xff
      12'h6DF: dout <= 8'b11111111; // 1759 : 255 - 0xff
      12'h6E0: dout <= 8'b00011111; // 1760 :  31 - 0x1f -- Sprite 0xdc
      12'h6E1: dout <= 8'b11011111; // 1761 : 223 - 0xdf
      12'h6E2: dout <= 8'b11000000; // 1762 : 192 - 0xc0
      12'h6E3: dout <= 8'b11110000; // 1763 : 240 - 0xf0
      12'h6E4: dout <= 8'b11110000; // 1764 : 240 - 0xf0
      12'h6E5: dout <= 8'b11111111; // 1765 : 255 - 0xff
      12'h6E6: dout <= 8'b11111111; // 1766 : 255 - 0xff
      12'h6E7: dout <= 8'b11111111; // 1767 : 255 - 0xff
      12'h6E8: dout <= 8'b10000100; // 1768 : 132 - 0x84 -- Sprite 0xdd
      12'h6E9: dout <= 8'b11111100; // 1769 : 252 - 0xfc
      12'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      12'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      12'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      12'h6ED: dout <= 8'b11111111; // 1773 : 255 - 0xff
      12'h6EE: dout <= 8'b11111111; // 1774 : 255 - 0xff
      12'h6EF: dout <= 8'b11111111; // 1775 : 255 - 0xff
      12'h6F0: dout <= 8'b01111111; // 1776 : 127 - 0x7f -- Sprite 0xde
      12'h6F1: dout <= 8'b01111111; // 1777 : 127 - 0x7f
      12'h6F2: dout <= 8'b00000000; // 1778 :   0 - 0x0
      12'h6F3: dout <= 8'b00000000; // 1779 :   0 - 0x0
      12'h6F4: dout <= 8'b00000000; // 1780 :   0 - 0x0
      12'h6F5: dout <= 8'b11111111; // 1781 : 255 - 0xff
      12'h6F6: dout <= 8'b11111111; // 1782 : 255 - 0xff
      12'h6F7: dout <= 8'b11111111; // 1783 : 255 - 0xff
      12'h6F8: dout <= 8'b11111100; // 1784 : 252 - 0xfc -- Sprite 0xdf
      12'h6F9: dout <= 8'b11111111; // 1785 : 255 - 0xff
      12'h6FA: dout <= 8'b00000000; // 1786 :   0 - 0x0
      12'h6FB: dout <= 8'b00000000; // 1787 :   0 - 0x0
      12'h6FC: dout <= 8'b00000000; // 1788 :   0 - 0x0
      12'h6FD: dout <= 8'b11111111; // 1789 : 255 - 0xff
      12'h6FE: dout <= 8'b11111111; // 1790 : 255 - 0xff
      12'h6FF: dout <= 8'b11111111; // 1791 : 255 - 0xff
      12'h700: dout <= 8'b00110000; // 1792 :  48 - 0x30 -- Sprite 0xe0
      12'h701: dout <= 8'b11110000; // 1793 : 240 - 0xf0
      12'h702: dout <= 8'b00000000; // 1794 :   0 - 0x0
      12'h703: dout <= 8'b00000000; // 1795 :   0 - 0x0
      12'h704: dout <= 8'b00000000; // 1796 :   0 - 0x0
      12'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      12'h706: dout <= 8'b11111111; // 1798 : 255 - 0xff
      12'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      12'h708: dout <= 8'b11111111; // 1800 : 255 - 0xff -- Sprite 0xe1
      12'h709: dout <= 8'b11111111; // 1801 : 255 - 0xff
      12'h70A: dout <= 8'b00000000; // 1802 :   0 - 0x0
      12'h70B: dout <= 8'b00000000; // 1803 :   0 - 0x0
      12'h70C: dout <= 8'b00000000; // 1804 :   0 - 0x0
      12'h70D: dout <= 8'b11111111; // 1805 : 255 - 0xff
      12'h70E: dout <= 8'b11111111; // 1806 : 255 - 0xff
      12'h70F: dout <= 8'b11111111; // 1807 : 255 - 0xff
      12'h710: dout <= 8'b11100001; // 1808 : 225 - 0xe1 -- Sprite 0xe2
      12'h711: dout <= 8'b11111111; // 1809 : 255 - 0xff
      12'h712: dout <= 8'b00000000; // 1810 :   0 - 0x0
      12'h713: dout <= 8'b00000000; // 1811 :   0 - 0x0
      12'h714: dout <= 8'b00000000; // 1812 :   0 - 0x0
      12'h715: dout <= 8'b11111111; // 1813 : 255 - 0xff
      12'h716: dout <= 8'b11111111; // 1814 : 255 - 0xff
      12'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      12'h718: dout <= 8'b00011111; // 1816 :  31 - 0x1f -- Sprite 0xe3
      12'h719: dout <= 8'b00011111; // 1817 :  31 - 0x1f
      12'h71A: dout <= 8'b00011111; // 1818 :  31 - 0x1f
      12'h71B: dout <= 8'b00011111; // 1819 :  31 - 0x1f
      12'h71C: dout <= 8'b00011111; // 1820 :  31 - 0x1f
      12'h71D: dout <= 8'b11111111; // 1821 : 255 - 0xff
      12'h71E: dout <= 8'b11111111; // 1822 : 255 - 0xff
      12'h71F: dout <= 8'b11111111; // 1823 : 255 - 0xff
      12'h720: dout <= 8'b00000000; // 1824 :   0 - 0x0 -- Sprite 0xe4
      12'h721: dout <= 8'b00011111; // 1825 :  31 - 0x1f
      12'h722: dout <= 8'b00111111; // 1826 :  63 - 0x3f
      12'h723: dout <= 8'b01111000; // 1827 : 120 - 0x78
      12'h724: dout <= 8'b01110111; // 1828 : 119 - 0x77
      12'h725: dout <= 8'b01101111; // 1829 : 111 - 0x6f
      12'h726: dout <= 8'b01101111; // 1830 : 111 - 0x6f
      12'h727: dout <= 8'b01101111; // 1831 : 111 - 0x6f
      12'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0 -- Sprite 0xe5
      12'h729: dout <= 8'b11111000; // 1833 : 248 - 0xf8
      12'h72A: dout <= 8'b11111100; // 1834 : 252 - 0xfc
      12'h72B: dout <= 8'b00011110; // 1835 :  30 - 0x1e
      12'h72C: dout <= 8'b11101110; // 1836 : 238 - 0xee
      12'h72D: dout <= 8'b11110110; // 1837 : 246 - 0xf6
      12'h72E: dout <= 8'b11110110; // 1838 : 246 - 0xf6
      12'h72F: dout <= 8'b11110110; // 1839 : 246 - 0xf6
      12'h730: dout <= 8'b11110110; // 1840 : 246 - 0xf6 -- Sprite 0xe6
      12'h731: dout <= 8'b11110110; // 1841 : 246 - 0xf6
      12'h732: dout <= 8'b11110110; // 1842 : 246 - 0xf6
      12'h733: dout <= 8'b11101110; // 1843 : 238 - 0xee
      12'h734: dout <= 8'b00011110; // 1844 :  30 - 0x1e
      12'h735: dout <= 8'b11111100; // 1845 : 252 - 0xfc
      12'h736: dout <= 8'b11111000; // 1846 : 248 - 0xf8
      12'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      12'h738: dout <= 8'b01101111; // 1848 : 111 - 0x6f -- Sprite 0xe7
      12'h739: dout <= 8'b01101111; // 1849 : 111 - 0x6f
      12'h73A: dout <= 8'b01101111; // 1850 : 111 - 0x6f
      12'h73B: dout <= 8'b01110111; // 1851 : 119 - 0x77
      12'h73C: dout <= 8'b01111000; // 1852 : 120 - 0x78
      12'h73D: dout <= 8'b00111111; // 1853 :  63 - 0x3f
      12'h73E: dout <= 8'b00011111; // 1854 :  31 - 0x1f
      12'h73F: dout <= 8'b00000000; // 1855 :   0 - 0x0
      12'h740: dout <= 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0xe8
      12'h741: dout <= 8'b11111111; // 1857 : 255 - 0xff
      12'h742: dout <= 8'b11111111; // 1858 : 255 - 0xff
      12'h743: dout <= 8'b00000000; // 1859 :   0 - 0x0
      12'h744: dout <= 8'b11111111; // 1860 : 255 - 0xff
      12'h745: dout <= 8'b11111111; // 1861 : 255 - 0xff
      12'h746: dout <= 8'b11111111; // 1862 : 255 - 0xff
      12'h747: dout <= 8'b11111111; // 1863 : 255 - 0xff
      12'h748: dout <= 8'b11110110; // 1864 : 246 - 0xf6 -- Sprite 0xe9
      12'h749: dout <= 8'b11110110; // 1865 : 246 - 0xf6
      12'h74A: dout <= 8'b11110110; // 1866 : 246 - 0xf6
      12'h74B: dout <= 8'b11110110; // 1867 : 246 - 0xf6
      12'h74C: dout <= 8'b11110110; // 1868 : 246 - 0xf6
      12'h74D: dout <= 8'b11110110; // 1869 : 246 - 0xf6
      12'h74E: dout <= 8'b11110110; // 1870 : 246 - 0xf6
      12'h74F: dout <= 8'b11110110; // 1871 : 246 - 0xf6
      12'h750: dout <= 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0xea
      12'h751: dout <= 8'b11111111; // 1873 : 255 - 0xff
      12'h752: dout <= 8'b11111111; // 1874 : 255 - 0xff
      12'h753: dout <= 8'b11111111; // 1875 : 255 - 0xff
      12'h754: dout <= 8'b00000000; // 1876 :   0 - 0x0
      12'h755: dout <= 8'b11111111; // 1877 : 255 - 0xff
      12'h756: dout <= 8'b11111111; // 1878 : 255 - 0xff
      12'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout <= 8'b01101111; // 1880 : 111 - 0x6f -- Sprite 0xeb
      12'h759: dout <= 8'b01101111; // 1881 : 111 - 0x6f
      12'h75A: dout <= 8'b01101111; // 1882 : 111 - 0x6f
      12'h75B: dout <= 8'b01101111; // 1883 : 111 - 0x6f
      12'h75C: dout <= 8'b01101111; // 1884 : 111 - 0x6f
      12'h75D: dout <= 8'b01101111; // 1885 : 111 - 0x6f
      12'h75E: dout <= 8'b01101111; // 1886 : 111 - 0x6f
      12'h75F: dout <= 8'b01101111; // 1887 : 111 - 0x6f
      12'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      12'h761: dout <= 8'b00000000; // 1889 :   0 - 0x0
      12'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      12'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      12'h765: dout <= 8'b00000000; // 1893 :   0 - 0x0
      12'h766: dout <= 8'b00000000; // 1894 :   0 - 0x0
      12'h767: dout <= 8'b00000000; // 1895 :   0 - 0x0
      12'h768: dout <= 8'b00000000; // 1896 :   0 - 0x0 -- Sprite 0xed
      12'h769: dout <= 8'b00000000; // 1897 :   0 - 0x0
      12'h76A: dout <= 8'b00000000; // 1898 :   0 - 0x0
      12'h76B: dout <= 8'b00000000; // 1899 :   0 - 0x0
      12'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      12'h76D: dout <= 8'b00000000; // 1901 :   0 - 0x0
      12'h76E: dout <= 8'b00000000; // 1902 :   0 - 0x0
      12'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      12'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0xee
      12'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout <= 8'b00000000; // 1906 :   0 - 0x0
      12'h773: dout <= 8'b00000000; // 1907 :   0 - 0x0
      12'h774: dout <= 8'b00000000; // 1908 :   0 - 0x0
      12'h775: dout <= 8'b00000000; // 1909 :   0 - 0x0
      12'h776: dout <= 8'b00000000; // 1910 :   0 - 0x0
      12'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      12'h778: dout <= 8'b00000000; // 1912 :   0 - 0x0 -- Sprite 0xef
      12'h779: dout <= 8'b00000000; // 1913 :   0 - 0x0
      12'h77A: dout <= 8'b00000000; // 1914 :   0 - 0x0
      12'h77B: dout <= 8'b00000000; // 1915 :   0 - 0x0
      12'h77C: dout <= 8'b00000000; // 1916 :   0 - 0x0
      12'h77D: dout <= 8'b00000000; // 1917 :   0 - 0x0
      12'h77E: dout <= 8'b00000000; // 1918 :   0 - 0x0
      12'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      12'h780: dout <= 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0xf0
      12'h781: dout <= 8'b11111111; // 1921 : 255 - 0xff
      12'h782: dout <= 8'b11111111; // 1922 : 255 - 0xff
      12'h783: dout <= 8'b11111111; // 1923 : 255 - 0xff
      12'h784: dout <= 8'b11111111; // 1924 : 255 - 0xff
      12'h785: dout <= 8'b11111111; // 1925 : 255 - 0xff
      12'h786: dout <= 8'b11111111; // 1926 : 255 - 0xff
      12'h787: dout <= 8'b11111111; // 1927 : 255 - 0xff
      12'h788: dout <= 8'b11111111; // 1928 : 255 - 0xff -- Sprite 0xf1
      12'h789: dout <= 8'b11111111; // 1929 : 255 - 0xff
      12'h78A: dout <= 8'b11111111; // 1930 : 255 - 0xff
      12'h78B: dout <= 8'b11111111; // 1931 : 255 - 0xff
      12'h78C: dout <= 8'b11111111; // 1932 : 255 - 0xff
      12'h78D: dout <= 8'b11111111; // 1933 : 255 - 0xff
      12'h78E: dout <= 8'b11111111; // 1934 : 255 - 0xff
      12'h78F: dout <= 8'b11111111; // 1935 : 255 - 0xff
      12'h790: dout <= 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0xf2
      12'h791: dout <= 8'b11111111; // 1937 : 255 - 0xff
      12'h792: dout <= 8'b11111111; // 1938 : 255 - 0xff
      12'h793: dout <= 8'b11111111; // 1939 : 255 - 0xff
      12'h794: dout <= 8'b11111111; // 1940 : 255 - 0xff
      12'h795: dout <= 8'b11111111; // 1941 : 255 - 0xff
      12'h796: dout <= 8'b11111111; // 1942 : 255 - 0xff
      12'h797: dout <= 8'b11111111; // 1943 : 255 - 0xff
      12'h798: dout <= 8'b11111111; // 1944 : 255 - 0xff -- Sprite 0xf3
      12'h799: dout <= 8'b11111111; // 1945 : 255 - 0xff
      12'h79A: dout <= 8'b11111111; // 1946 : 255 - 0xff
      12'h79B: dout <= 8'b11111111; // 1947 : 255 - 0xff
      12'h79C: dout <= 8'b11111111; // 1948 : 255 - 0xff
      12'h79D: dout <= 8'b11111111; // 1949 : 255 - 0xff
      12'h79E: dout <= 8'b11111111; // 1950 : 255 - 0xff
      12'h79F: dout <= 8'b11111111; // 1951 : 255 - 0xff
      12'h7A0: dout <= 8'b11111111; // 1952 : 255 - 0xff -- Sprite 0xf4
      12'h7A1: dout <= 8'b11111111; // 1953 : 255 - 0xff
      12'h7A2: dout <= 8'b11111111; // 1954 : 255 - 0xff
      12'h7A3: dout <= 8'b11111111; // 1955 : 255 - 0xff
      12'h7A4: dout <= 8'b11111111; // 1956 : 255 - 0xff
      12'h7A5: dout <= 8'b11111111; // 1957 : 255 - 0xff
      12'h7A6: dout <= 8'b11111111; // 1958 : 255 - 0xff
      12'h7A7: dout <= 8'b11111111; // 1959 : 255 - 0xff
      12'h7A8: dout <= 8'b11111111; // 1960 : 255 - 0xff -- Sprite 0xf5
      12'h7A9: dout <= 8'b11111111; // 1961 : 255 - 0xff
      12'h7AA: dout <= 8'b11111111; // 1962 : 255 - 0xff
      12'h7AB: dout <= 8'b11111111; // 1963 : 255 - 0xff
      12'h7AC: dout <= 8'b11111111; // 1964 : 255 - 0xff
      12'h7AD: dout <= 8'b11111111; // 1965 : 255 - 0xff
      12'h7AE: dout <= 8'b11111111; // 1966 : 255 - 0xff
      12'h7AF: dout <= 8'b11111111; // 1967 : 255 - 0xff
      12'h7B0: dout <= 8'b11111111; // 1968 : 255 - 0xff -- Sprite 0xf6
      12'h7B1: dout <= 8'b11111111; // 1969 : 255 - 0xff
      12'h7B2: dout <= 8'b11111111; // 1970 : 255 - 0xff
      12'h7B3: dout <= 8'b11111111; // 1971 : 255 - 0xff
      12'h7B4: dout <= 8'b11111111; // 1972 : 255 - 0xff
      12'h7B5: dout <= 8'b11111111; // 1973 : 255 - 0xff
      12'h7B6: dout <= 8'b11111111; // 1974 : 255 - 0xff
      12'h7B7: dout <= 8'b11111111; // 1975 : 255 - 0xff
      12'h7B8: dout <= 8'b11111111; // 1976 : 255 - 0xff -- Sprite 0xf7
      12'h7B9: dout <= 8'b11111111; // 1977 : 255 - 0xff
      12'h7BA: dout <= 8'b11111111; // 1978 : 255 - 0xff
      12'h7BB: dout <= 8'b11111111; // 1979 : 255 - 0xff
      12'h7BC: dout <= 8'b11111111; // 1980 : 255 - 0xff
      12'h7BD: dout <= 8'b11111111; // 1981 : 255 - 0xff
      12'h7BE: dout <= 8'b11111111; // 1982 : 255 - 0xff
      12'h7BF: dout <= 8'b11111111; // 1983 : 255 - 0xff
      12'h7C0: dout <= 8'b11111111; // 1984 : 255 - 0xff -- Sprite 0xf8
      12'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      12'h7C2: dout <= 8'b11111111; // 1986 : 255 - 0xff
      12'h7C3: dout <= 8'b11111111; // 1987 : 255 - 0xff
      12'h7C4: dout <= 8'b11111111; // 1988 : 255 - 0xff
      12'h7C5: dout <= 8'b11111111; // 1989 : 255 - 0xff
      12'h7C6: dout <= 8'b11111111; // 1990 : 255 - 0xff
      12'h7C7: dout <= 8'b11111111; // 1991 : 255 - 0xff
      12'h7C8: dout <= 8'b11111111; // 1992 : 255 - 0xff -- Sprite 0xf9
      12'h7C9: dout <= 8'b11111111; // 1993 : 255 - 0xff
      12'h7CA: dout <= 8'b11111111; // 1994 : 255 - 0xff
      12'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      12'h7CC: dout <= 8'b11111111; // 1996 : 255 - 0xff
      12'h7CD: dout <= 8'b11111111; // 1997 : 255 - 0xff
      12'h7CE: dout <= 8'b11111111; // 1998 : 255 - 0xff
      12'h7CF: dout <= 8'b11111111; // 1999 : 255 - 0xff
      12'h7D0: dout <= 8'b11111111; // 2000 : 255 - 0xff -- Sprite 0xfa
      12'h7D1: dout <= 8'b11111111; // 2001 : 255 - 0xff
      12'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      12'h7D3: dout <= 8'b11111111; // 2003 : 255 - 0xff
      12'h7D4: dout <= 8'b11111111; // 2004 : 255 - 0xff
      12'h7D5: dout <= 8'b11111111; // 2005 : 255 - 0xff
      12'h7D6: dout <= 8'b11111111; // 2006 : 255 - 0xff
      12'h7D7: dout <= 8'b11111111; // 2007 : 255 - 0xff
      12'h7D8: dout <= 8'b11111111; // 2008 : 255 - 0xff -- Sprite 0xfb
      12'h7D9: dout <= 8'b11111111; // 2009 : 255 - 0xff
      12'h7DA: dout <= 8'b11111111; // 2010 : 255 - 0xff
      12'h7DB: dout <= 8'b11111111; // 2011 : 255 - 0xff
      12'h7DC: dout <= 8'b11111111; // 2012 : 255 - 0xff
      12'h7DD: dout <= 8'b11111111; // 2013 : 255 - 0xff
      12'h7DE: dout <= 8'b11111111; // 2014 : 255 - 0xff
      12'h7DF: dout <= 8'b11111111; // 2015 : 255 - 0xff
      12'h7E0: dout <= 8'b11111111; // 2016 : 255 - 0xff -- Sprite 0xfc
      12'h7E1: dout <= 8'b11111111; // 2017 : 255 - 0xff
      12'h7E2: dout <= 8'b11111111; // 2018 : 255 - 0xff
      12'h7E3: dout <= 8'b11111111; // 2019 : 255 - 0xff
      12'h7E4: dout <= 8'b11111111; // 2020 : 255 - 0xff
      12'h7E5: dout <= 8'b11111111; // 2021 : 255 - 0xff
      12'h7E6: dout <= 8'b11111111; // 2022 : 255 - 0xff
      12'h7E7: dout <= 8'b11111111; // 2023 : 255 - 0xff
      12'h7E8: dout <= 8'b11111111; // 2024 : 255 - 0xff -- Sprite 0xfd
      12'h7E9: dout <= 8'b11111111; // 2025 : 255 - 0xff
      12'h7EA: dout <= 8'b11111111; // 2026 : 255 - 0xff
      12'h7EB: dout <= 8'b11111111; // 2027 : 255 - 0xff
      12'h7EC: dout <= 8'b11111111; // 2028 : 255 - 0xff
      12'h7ED: dout <= 8'b11111111; // 2029 : 255 - 0xff
      12'h7EE: dout <= 8'b11111111; // 2030 : 255 - 0xff
      12'h7EF: dout <= 8'b11111111; // 2031 : 255 - 0xff
      12'h7F0: dout <= 8'b11111111; // 2032 : 255 - 0xff -- Sprite 0xfe
      12'h7F1: dout <= 8'b11111111; // 2033 : 255 - 0xff
      12'h7F2: dout <= 8'b11111111; // 2034 : 255 - 0xff
      12'h7F3: dout <= 8'b11111111; // 2035 : 255 - 0xff
      12'h7F4: dout <= 8'b11111111; // 2036 : 255 - 0xff
      12'h7F5: dout <= 8'b11111111; // 2037 : 255 - 0xff
      12'h7F6: dout <= 8'b11111111; // 2038 : 255 - 0xff
      12'h7F7: dout <= 8'b11111111; // 2039 : 255 - 0xff
      12'h7F8: dout <= 8'b11111111; // 2040 : 255 - 0xff -- Sprite 0xff
      12'h7F9: dout <= 8'b11111111; // 2041 : 255 - 0xff
      12'h7FA: dout <= 8'b11111111; // 2042 : 255 - 0xff
      12'h7FB: dout <= 8'b11111111; // 2043 : 255 - 0xff
      12'h7FC: dout <= 8'b11111111; // 2044 : 255 - 0xff
      12'h7FD: dout <= 8'b11111111; // 2045 : 255 - 0xff
      12'h7FE: dout <= 8'b11111111; // 2046 : 255 - 0xff
      12'h7FF: dout <= 8'b11111111; // 2047 : 255 - 0xff
          // Background pattern Table
      12'h800: dout <= 8'b00000000; // 2048 :   0 - 0x0 -- Background 0x0
      12'h801: dout <= 8'b00000011; // 2049 :   3 - 0x3
      12'h802: dout <= 8'b00001111; // 2050 :  15 - 0xf
      12'h803: dout <= 8'b00011111; // 2051 :  31 - 0x1f
      12'h804: dout <= 8'b00111111; // 2052 :  63 - 0x3f
      12'h805: dout <= 8'b00111111; // 2053 :  63 - 0x3f
      12'h806: dout <= 8'b01111111; // 2054 : 127 - 0x7f
      12'h807: dout <= 8'b01111111; // 2055 : 127 - 0x7f
      12'h808: dout <= 8'b00000000; // 2056 :   0 - 0x0 -- Background 0x1
      12'h809: dout <= 8'b11000000; // 2057 : 192 - 0xc0
      12'h80A: dout <= 8'b11110000; // 2058 : 240 - 0xf0
      12'h80B: dout <= 8'b11111000; // 2059 : 248 - 0xf8
      12'h80C: dout <= 8'b11111000; // 2060 : 248 - 0xf8
      12'h80D: dout <= 8'b11111100; // 2061 : 252 - 0xfc
      12'h80E: dout <= 8'b11111100; // 2062 : 252 - 0xfc
      12'h80F: dout <= 8'b11111100; // 2063 : 252 - 0xfc
      12'h810: dout <= 8'b00000000; // 2064 :   0 - 0x0 -- Background 0x2
      12'h811: dout <= 8'b00000111; // 2065 :   7 - 0x7
      12'h812: dout <= 8'b00011111; // 2066 :  31 - 0x1f
      12'h813: dout <= 8'b00111111; // 2067 :  63 - 0x3f
      12'h814: dout <= 8'b00111111; // 2068 :  63 - 0x3f
      12'h815: dout <= 8'b00001111; // 2069 :  15 - 0xf
      12'h816: dout <= 8'b00000011; // 2070 :   3 - 0x3
      12'h817: dout <= 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout <= 8'b00000000; // 2072 :   0 - 0x0 -- Background 0x3
      12'h819: dout <= 8'b00000000; // 2073 :   0 - 0x0
      12'h81A: dout <= 8'b00000111; // 2074 :   7 - 0x7
      12'h81B: dout <= 8'b00011111; // 2075 :  31 - 0x1f
      12'h81C: dout <= 8'b00111111; // 2076 :  63 - 0x3f
      12'h81D: dout <= 8'b00111111; // 2077 :  63 - 0x3f
      12'h81E: dout <= 8'b01111111; // 2078 : 127 - 0x7f
      12'h81F: dout <= 8'b01111111; // 2079 : 127 - 0x7f
      12'h820: dout <= 8'b01111110; // 2080 : 126 - 0x7e -- Background 0x4
      12'h821: dout <= 8'b01111110; // 2081 : 126 - 0x7e
      12'h822: dout <= 8'b01111100; // 2082 : 124 - 0x7c
      12'h823: dout <= 8'b00111100; // 2083 :  60 - 0x3c
      12'h824: dout <= 8'b00111000; // 2084 :  56 - 0x38
      12'h825: dout <= 8'b00011000; // 2085 :  24 - 0x18
      12'h826: dout <= 8'b00000000; // 2086 :   0 - 0x0
      12'h827: dout <= 8'b00000000; // 2087 :   0 - 0x0
      12'h828: dout <= 8'b00000000; // 2088 :   0 - 0x0 -- Background 0x5
      12'h829: dout <= 8'b11000000; // 2089 : 192 - 0xc0
      12'h82A: dout <= 8'b11110000; // 2090 : 240 - 0xf0
      12'h82B: dout <= 8'b11111000; // 2091 : 248 - 0xf8
      12'h82C: dout <= 8'b11111000; // 2092 : 248 - 0xf8
      12'h82D: dout <= 8'b11111100; // 2093 : 252 - 0xfc
      12'h82E: dout <= 8'b01111100; // 2094 : 124 - 0x7c
      12'h82F: dout <= 8'b00111100; // 2095 :  60 - 0x3c
      12'h830: dout <= 8'b00000000; // 2096 :   0 - 0x0 -- Background 0x6
      12'h831: dout <= 8'b00000111; // 2097 :   7 - 0x7
      12'h832: dout <= 8'b00000111; // 2098 :   7 - 0x7
      12'h833: dout <= 8'b00000011; // 2099 :   3 - 0x3
      12'h834: dout <= 8'b00000001; // 2100 :   1 - 0x1
      12'h835: dout <= 8'b00000000; // 2101 :   0 - 0x0
      12'h836: dout <= 8'b00000000; // 2102 :   0 - 0x0
      12'h837: dout <= 8'b00000000; // 2103 :   0 - 0x0
      12'h838: dout <= 8'b00000000; // 2104 :   0 - 0x0 -- Background 0x7
      12'h839: dout <= 8'b00000000; // 2105 :   0 - 0x0
      12'h83A: dout <= 8'b00000111; // 2106 :   7 - 0x7
      12'h83B: dout <= 8'b00011111; // 2107 :  31 - 0x1f
      12'h83C: dout <= 8'b00111111; // 2108 :  63 - 0x3f
      12'h83D: dout <= 8'b00111111; // 2109 :  63 - 0x3f
      12'h83E: dout <= 8'b01111110; // 2110 : 126 - 0x7e
      12'h83F: dout <= 8'b01111100; // 2111 : 124 - 0x7c
      12'h840: dout <= 8'b01111000; // 2112 : 120 - 0x78 -- Background 0x8
      12'h841: dout <= 8'b01110000; // 2113 : 112 - 0x70
      12'h842: dout <= 8'b01100000; // 2114 :  96 - 0x60
      12'h843: dout <= 8'b00000000; // 2115 :   0 - 0x0
      12'h844: dout <= 8'b00000000; // 2116 :   0 - 0x0
      12'h845: dout <= 8'b00000000; // 2117 :   0 - 0x0
      12'h846: dout <= 8'b00000000; // 2118 :   0 - 0x0
      12'h847: dout <= 8'b00000000; // 2119 :   0 - 0x0
      12'h848: dout <= 8'b00000000; // 2120 :   0 - 0x0 -- Background 0x9
      12'h849: dout <= 8'b00000000; // 2121 :   0 - 0x0
      12'h84A: dout <= 8'b00000000; // 2122 :   0 - 0x0
      12'h84B: dout <= 8'b00000000; // 2123 :   0 - 0x0
      12'h84C: dout <= 8'b00000000; // 2124 :   0 - 0x0
      12'h84D: dout <= 8'b01000000; // 2125 :  64 - 0x40
      12'h84E: dout <= 8'b11110000; // 2126 : 240 - 0xf0
      12'h84F: dout <= 8'b11111000; // 2127 : 248 - 0xf8
      12'h850: dout <= 8'b11111110; // 2128 : 254 - 0xfe -- Background 0xa
      12'h851: dout <= 8'b01111111; // 2129 : 127 - 0x7f
      12'h852: dout <= 8'b01111111; // 2130 : 127 - 0x7f
      12'h853: dout <= 8'b00111111; // 2131 :  63 - 0x3f
      12'h854: dout <= 8'b00001110; // 2132 :  14 - 0xe
      12'h855: dout <= 8'b00000000; // 2133 :   0 - 0x0
      12'h856: dout <= 8'b00000000; // 2134 :   0 - 0x0
      12'h857: dout <= 8'b00000000; // 2135 :   0 - 0x0
      12'h858: dout <= 8'b00000000; // 2136 :   0 - 0x0 -- Background 0xb
      12'h859: dout <= 8'b00000000; // 2137 :   0 - 0x0
      12'h85A: dout <= 8'b00000000; // 2138 :   0 - 0x0
      12'h85B: dout <= 8'b00000000; // 2139 :   0 - 0x0
      12'h85C: dout <= 8'b00000000; // 2140 :   0 - 0x0
      12'h85D: dout <= 8'b00000000; // 2141 :   0 - 0x0
      12'h85E: dout <= 8'b00000000; // 2142 :   0 - 0x0
      12'h85F: dout <= 8'b11100000; // 2143 : 224 - 0xe0
      12'h860: dout <= 8'b11111100; // 2144 : 252 - 0xfc -- Background 0xc
      12'h861: dout <= 8'b11111111; // 2145 : 255 - 0xff
      12'h862: dout <= 8'b01111111; // 2146 : 127 - 0x7f
      12'h863: dout <= 8'b00111111; // 2147 :  63 - 0x3f
      12'h864: dout <= 8'b00001110; // 2148 :  14 - 0xe
      12'h865: dout <= 8'b00000000; // 2149 :   0 - 0x0
      12'h866: dout <= 8'b00000000; // 2150 :   0 - 0x0
      12'h867: dout <= 8'b00000000; // 2151 :   0 - 0x0
      12'h868: dout <= 8'b11110000; // 2152 : 240 - 0xf0 -- Background 0xd
      12'h869: dout <= 8'b11111111; // 2153 : 255 - 0xff
      12'h86A: dout <= 8'b11111111; // 2154 : 255 - 0xff
      12'h86B: dout <= 8'b01111111; // 2155 : 127 - 0x7f
      12'h86C: dout <= 8'b00011110; // 2156 :  30 - 0x1e
      12'h86D: dout <= 8'b00000000; // 2157 :   0 - 0x0
      12'h86E: dout <= 8'b00000000; // 2158 :   0 - 0x0
      12'h86F: dout <= 8'b00000000; // 2159 :   0 - 0x0
      12'h870: dout <= 8'b00000000; // 2160 :   0 - 0x0 -- Background 0xe
      12'h871: dout <= 8'b00001111; // 2161 :  15 - 0xf
      12'h872: dout <= 8'b11111111; // 2162 : 255 - 0xff
      12'h873: dout <= 8'b11111111; // 2163 : 255 - 0xff
      12'h874: dout <= 8'b01111111; // 2164 : 127 - 0x7f
      12'h875: dout <= 8'b00011110; // 2165 :  30 - 0x1e
      12'h876: dout <= 8'b00000000; // 2166 :   0 - 0x0
      12'h877: dout <= 8'b00000000; // 2167 :   0 - 0x0
      12'h878: dout <= 8'b00000000; // 2168 :   0 - 0x0 -- Background 0xf
      12'h879: dout <= 8'b00000011; // 2169 :   3 - 0x3
      12'h87A: dout <= 8'b00001111; // 2170 :  15 - 0xf
      12'h87B: dout <= 8'b01111111; // 2171 : 127 - 0x7f
      12'h87C: dout <= 8'b11111111; // 2172 : 255 - 0xff
      12'h87D: dout <= 8'b01111110; // 2173 : 126 - 0x7e
      12'h87E: dout <= 8'b00011100; // 2174 :  28 - 0x1c
      12'h87F: dout <= 8'b00000000; // 2175 :   0 - 0x0
      12'h880: dout <= 8'b00000000; // 2176 :   0 - 0x0 -- Background 0x10
      12'h881: dout <= 8'b00000001; // 2177 :   1 - 0x1
      12'h882: dout <= 8'b00000011; // 2178 :   3 - 0x3
      12'h883: dout <= 8'b00001111; // 2179 :  15 - 0xf
      12'h884: dout <= 8'b00011111; // 2180 :  31 - 0x1f
      12'h885: dout <= 8'b01111111; // 2181 : 127 - 0x7f
      12'h886: dout <= 8'b01111110; // 2182 : 126 - 0x7e
      12'h887: dout <= 8'b00111100; // 2183 :  60 - 0x3c
      12'h888: dout <= 8'b00000000; // 2184 :   0 - 0x0 -- Background 0x11
      12'h889: dout <= 8'b00000001; // 2185 :   1 - 0x1
      12'h88A: dout <= 8'b00000011; // 2186 :   3 - 0x3
      12'h88B: dout <= 8'b00000111; // 2187 :   7 - 0x7
      12'h88C: dout <= 8'b00000111; // 2188 :   7 - 0x7
      12'h88D: dout <= 8'b00001111; // 2189 :  15 - 0xf
      12'h88E: dout <= 8'b00011111; // 2190 :  31 - 0x1f
      12'h88F: dout <= 8'b00001110; // 2191 :  14 - 0xe
      12'h890: dout <= 8'b00000000; // 2192 :   0 - 0x0 -- Background 0x12
      12'h891: dout <= 8'b00000000; // 2193 :   0 - 0x0
      12'h892: dout <= 8'b00000001; // 2194 :   1 - 0x1
      12'h893: dout <= 8'b00000011; // 2195 :   3 - 0x3
      12'h894: dout <= 8'b00000011; // 2196 :   3 - 0x3
      12'h895: dout <= 8'b00000011; // 2197 :   3 - 0x3
      12'h896: dout <= 8'b00000111; // 2198 :   7 - 0x7
      12'h897: dout <= 8'b00000010; // 2199 :   2 - 0x2
      12'h898: dout <= 8'b00000000; // 2200 :   0 - 0x0 -- Background 0x13
      12'h899: dout <= 8'b00000000; // 2201 :   0 - 0x0
      12'h89A: dout <= 8'b00000001; // 2202 :   1 - 0x1
      12'h89B: dout <= 8'b00000001; // 2203 :   1 - 0x1
      12'h89C: dout <= 8'b00000001; // 2204 :   1 - 0x1
      12'h89D: dout <= 8'b00000001; // 2205 :   1 - 0x1
      12'h89E: dout <= 8'b00000001; // 2206 :   1 - 0x1
      12'h89F: dout <= 8'b00000001; // 2207 :   1 - 0x1
      12'h8A0: dout <= 8'b00000000; // 2208 :   0 - 0x0 -- Background 0x14
      12'h8A1: dout <= 8'b00000000; // 2209 :   0 - 0x0
      12'h8A2: dout <= 8'b00000000; // 2210 :   0 - 0x0
      12'h8A3: dout <= 8'b00000000; // 2211 :   0 - 0x0
      12'h8A4: dout <= 8'b00000000; // 2212 :   0 - 0x0
      12'h8A5: dout <= 8'b00000000; // 2213 :   0 - 0x0
      12'h8A6: dout <= 8'b00000100; // 2214 :   4 - 0x4
      12'h8A7: dout <= 8'b00000010; // 2215 :   2 - 0x2
      12'h8A8: dout <= 8'b00000000; // 2216 :   0 - 0x0 -- Background 0x15
      12'h8A9: dout <= 8'b00000000; // 2217 :   0 - 0x0
      12'h8AA: dout <= 8'b00000000; // 2218 :   0 - 0x0
      12'h8AB: dout <= 8'b00000000; // 2219 :   0 - 0x0
      12'h8AC: dout <= 8'b00000000; // 2220 :   0 - 0x0
      12'h8AD: dout <= 8'b00000000; // 2221 :   0 - 0x0
      12'h8AE: dout <= 8'b00100000; // 2222 :  32 - 0x20
      12'h8AF: dout <= 8'b01001000; // 2223 :  72 - 0x48
      12'h8B0: dout <= 8'b00010000; // 2224 :  16 - 0x10 -- Background 0x16
      12'h8B1: dout <= 8'b00001000; // 2225 :   8 - 0x8
      12'h8B2: dout <= 8'b00000000; // 2226 :   0 - 0x0
      12'h8B3: dout <= 8'b00110000; // 2227 :  48 - 0x30
      12'h8B4: dout <= 8'b00000000; // 2228 :   0 - 0x0
      12'h8B5: dout <= 8'b00001000; // 2229 :   8 - 0x8
      12'h8B6: dout <= 8'b00010010; // 2230 :  18 - 0x12
      12'h8B7: dout <= 8'b00000100; // 2231 :   4 - 0x4
      12'h8B8: dout <= 8'b00010000; // 2232 :  16 - 0x10 -- Background 0x17
      12'h8B9: dout <= 8'b00000000; // 2233 :   0 - 0x0
      12'h8BA: dout <= 8'b00001100; // 2234 :  12 - 0xc
      12'h8BB: dout <= 8'b00000000; // 2235 :   0 - 0x0
      12'h8BC: dout <= 8'b00010000; // 2236 :  16 - 0x10
      12'h8BD: dout <= 8'b00001000; // 2237 :   8 - 0x8
      12'h8BE: dout <= 8'b01000000; // 2238 :  64 - 0x40
      12'h8BF: dout <= 8'b00100000; // 2239 :  32 - 0x20
      12'h8C0: dout <= 8'b00000000; // 2240 :   0 - 0x0 -- Background 0x18
      12'h8C1: dout <= 8'b00000000; // 2241 :   0 - 0x0
      12'h8C2: dout <= 8'b00000011; // 2242 :   3 - 0x3
      12'h8C3: dout <= 8'b00000011; // 2243 :   3 - 0x3
      12'h8C4: dout <= 8'b00000001; // 2244 :   1 - 0x1
      12'h8C5: dout <= 8'b00100001; // 2245 :  33 - 0x21
      12'h8C6: dout <= 8'b00100001; // 2246 :  33 - 0x21
      12'h8C7: dout <= 8'b01110011; // 2247 : 115 - 0x73
      12'h8C8: dout <= 8'b01111111; // 2248 : 127 - 0x7f -- Background 0x19
      12'h8C9: dout <= 8'b01111111; // 2249 : 127 - 0x7f
      12'h8CA: dout <= 8'b01111111; // 2250 : 127 - 0x7f
      12'h8CB: dout <= 8'b01111111; // 2251 : 127 - 0x7f
      12'h8CC: dout <= 8'b01101110; // 2252 : 110 - 0x6e
      12'h8CD: dout <= 8'b01000110; // 2253 :  70 - 0x46
      12'h8CE: dout <= 8'b00000000; // 2254 :   0 - 0x0
      12'h8CF: dout <= 8'b00000000; // 2255 :   0 - 0x0
      12'h8D0: dout <= 8'b01111111; // 2256 : 127 - 0x7f -- Background 0x1a
      12'h8D1: dout <= 8'b01111111; // 2257 : 127 - 0x7f
      12'h8D2: dout <= 8'b01111111; // 2258 : 127 - 0x7f
      12'h8D3: dout <= 8'b01111111; // 2259 : 127 - 0x7f
      12'h8D4: dout <= 8'b01111011; // 2260 : 123 - 0x7b
      12'h8D5: dout <= 8'b00110001; // 2261 :  49 - 0x31
      12'h8D6: dout <= 8'b00000000; // 2262 :   0 - 0x0
      12'h8D7: dout <= 8'b00000000; // 2263 :   0 - 0x0
      12'h8D8: dout <= 8'b00000000; // 2264 :   0 - 0x0 -- Background 0x1b
      12'h8D9: dout <= 8'b00000011; // 2265 :   3 - 0x3
      12'h8DA: dout <= 8'b00001111; // 2266 :  15 - 0xf
      12'h8DB: dout <= 8'b00011111; // 2267 :  31 - 0x1f
      12'h8DC: dout <= 8'b00100111; // 2268 :  39 - 0x27
      12'h8DD: dout <= 8'b00000011; // 2269 :   3 - 0x3
      12'h8DE: dout <= 8'b00000011; // 2270 :   3 - 0x3
      12'h8DF: dout <= 8'b01000011; // 2271 :  67 - 0x43
      12'h8E0: dout <= 8'b00000000; // 2272 :   0 - 0x0 -- Background 0x1c
      12'h8E1: dout <= 8'b11000000; // 2273 : 192 - 0xc0
      12'h8E2: dout <= 8'b11110000; // 2274 : 240 - 0xf0
      12'h8E3: dout <= 8'b11111000; // 2275 : 248 - 0xf8
      12'h8E4: dout <= 8'b10011100; // 2276 : 156 - 0x9c
      12'h8E5: dout <= 8'b00001100; // 2277 :  12 - 0xc
      12'h8E6: dout <= 8'b00001100; // 2278 :  12 - 0xc
      12'h8E7: dout <= 8'b00001110; // 2279 :  14 - 0xe
      12'h8E8: dout <= 8'b01100111; // 2280 : 103 - 0x67 -- Background 0x1d
      12'h8E9: dout <= 8'b01111111; // 2281 : 127 - 0x7f
      12'h8EA: dout <= 8'b01111111; // 2282 : 127 - 0x7f
      12'h8EB: dout <= 8'b01111111; // 2283 : 127 - 0x7f
      12'h8EC: dout <= 8'b01101110; // 2284 : 110 - 0x6e
      12'h8ED: dout <= 8'b01000110; // 2285 :  70 - 0x46
      12'h8EE: dout <= 8'b00000000; // 2286 :   0 - 0x0
      12'h8EF: dout <= 8'b00000000; // 2287 :   0 - 0x0
      12'h8F0: dout <= 8'b01100111; // 2288 : 103 - 0x67 -- Background 0x1e
      12'h8F1: dout <= 8'b01111111; // 2289 : 127 - 0x7f
      12'h8F2: dout <= 8'b01111111; // 2290 : 127 - 0x7f
      12'h8F3: dout <= 8'b01111111; // 2291 : 127 - 0x7f
      12'h8F4: dout <= 8'b01111011; // 2292 : 123 - 0x7b
      12'h8F5: dout <= 8'b00110001; // 2293 :  49 - 0x31
      12'h8F6: dout <= 8'b00000000; // 2294 :   0 - 0x0
      12'h8F7: dout <= 8'b00000000; // 2295 :   0 - 0x0
      12'h8F8: dout <= 8'b10011110; // 2296 : 158 - 0x9e -- Background 0x1f
      12'h8F9: dout <= 8'b11111110; // 2297 : 254 - 0xfe
      12'h8FA: dout <= 8'b11111110; // 2298 : 254 - 0xfe
      12'h8FB: dout <= 8'b11111110; // 2299 : 254 - 0xfe
      12'h8FC: dout <= 8'b01110110; // 2300 : 118 - 0x76
      12'h8FD: dout <= 8'b01100010; // 2301 :  98 - 0x62
      12'h8FE: dout <= 8'b00000000; // 2302 :   0 - 0x0
      12'h8FF: dout <= 8'b00000000; // 2303 :   0 - 0x0
      12'h900: dout <= 8'b10011110; // 2304 : 158 - 0x9e -- Background 0x20
      12'h901: dout <= 8'b11111110; // 2305 : 254 - 0xfe
      12'h902: dout <= 8'b11111110; // 2306 : 254 - 0xfe
      12'h903: dout <= 8'b11111110; // 2307 : 254 - 0xfe
      12'h904: dout <= 8'b11011110; // 2308 : 222 - 0xde
      12'h905: dout <= 8'b10001100; // 2309 : 140 - 0x8c
      12'h906: dout <= 8'b00000000; // 2310 :   0 - 0x0
      12'h907: dout <= 8'b00000000; // 2311 :   0 - 0x0
      12'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0 -- Background 0x21
      12'h909: dout <= 8'b00000011; // 2313 :   3 - 0x3
      12'h90A: dout <= 8'b00001111; // 2314 :  15 - 0xf
      12'h90B: dout <= 8'b00011111; // 2315 :  31 - 0x1f
      12'h90C: dout <= 8'b00111111; // 2316 :  63 - 0x3f
      12'h90D: dout <= 8'b00110011; // 2317 :  51 - 0x33
      12'h90E: dout <= 8'b00100001; // 2318 :  33 - 0x21
      12'h90F: dout <= 8'b01100001; // 2319 :  97 - 0x61
      12'h910: dout <= 8'b01100001; // 2320 :  97 - 0x61 -- Background 0x22
      12'h911: dout <= 8'b01110011; // 2321 : 115 - 0x73
      12'h912: dout <= 8'b01111111; // 2322 : 127 - 0x7f
      12'h913: dout <= 8'b01111111; // 2323 : 127 - 0x7f
      12'h914: dout <= 8'b01101110; // 2324 : 110 - 0x6e
      12'h915: dout <= 8'b01000110; // 2325 :  70 - 0x46
      12'h916: dout <= 8'b00000000; // 2326 :   0 - 0x0
      12'h917: dout <= 8'b00000000; // 2327 :   0 - 0x0
      12'h918: dout <= 8'b01100001; // 2328 :  97 - 0x61 -- Background 0x23
      12'h919: dout <= 8'b01110011; // 2329 : 115 - 0x73
      12'h91A: dout <= 8'b01111111; // 2330 : 127 - 0x7f
      12'h91B: dout <= 8'b01111111; // 2331 : 127 - 0x7f
      12'h91C: dout <= 8'b01110111; // 2332 : 119 - 0x77
      12'h91D: dout <= 8'b00100011; // 2333 :  35 - 0x23
      12'h91E: dout <= 8'b00000000; // 2334 :   0 - 0x0
      12'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout <= 8'b00000000; // 2336 :   0 - 0x0 -- Background 0x24
      12'h921: dout <= 8'b00000011; // 2337 :   3 - 0x3
      12'h922: dout <= 8'b00001111; // 2338 :  15 - 0xf
      12'h923: dout <= 8'b00011111; // 2339 :  31 - 0x1f
      12'h924: dout <= 8'b00111111; // 2340 :  63 - 0x3f
      12'h925: dout <= 8'b00111111; // 2341 :  63 - 0x3f
      12'h926: dout <= 8'b00111111; // 2342 :  63 - 0x3f
      12'h927: dout <= 8'b01111111; // 2343 : 127 - 0x7f
      12'h928: dout <= 8'b01111111; // 2344 : 127 - 0x7f -- Background 0x25
      12'h929: dout <= 8'b01111111; // 2345 : 127 - 0x7f
      12'h92A: dout <= 8'b01111111; // 2346 : 127 - 0x7f
      12'h92B: dout <= 8'b01111111; // 2347 : 127 - 0x7f
      12'h92C: dout <= 8'b01101110; // 2348 : 110 - 0x6e
      12'h92D: dout <= 8'b01000110; // 2349 :  70 - 0x46
      12'h92E: dout <= 8'b00000000; // 2350 :   0 - 0x0
      12'h92F: dout <= 8'b00000000; // 2351 :   0 - 0x0
      12'h930: dout <= 8'b01111111; // 2352 : 127 - 0x7f -- Background 0x26
      12'h931: dout <= 8'b01111111; // 2353 : 127 - 0x7f
      12'h932: dout <= 8'b01111111; // 2354 : 127 - 0x7f
      12'h933: dout <= 8'b01111111; // 2355 : 127 - 0x7f
      12'h934: dout <= 8'b01111011; // 2356 : 123 - 0x7b
      12'h935: dout <= 8'b00110001; // 2357 :  49 - 0x31
      12'h936: dout <= 8'b00000000; // 2358 :   0 - 0x0
      12'h937: dout <= 8'b00000000; // 2359 :   0 - 0x0
      12'h938: dout <= 8'b00000000; // 2360 :   0 - 0x0 -- Background 0x27
      12'h939: dout <= 8'b00000000; // 2361 :   0 - 0x0
      12'h93A: dout <= 8'b00000000; // 2362 :   0 - 0x0
      12'h93B: dout <= 8'b00000000; // 2363 :   0 - 0x0
      12'h93C: dout <= 8'b00000000; // 2364 :   0 - 0x0
      12'h93D: dout <= 8'b00000000; // 2365 :   0 - 0x0
      12'h93E: dout <= 8'b00000000; // 2366 :   0 - 0x0
      12'h93F: dout <= 8'b00000000; // 2367 :   0 - 0x0
      12'h940: dout <= 8'b00000000; // 2368 :   0 - 0x0 -- Background 0x28
      12'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout <= 8'b00000000; // 2370 :   0 - 0x0
      12'h943: dout <= 8'b00000000; // 2371 :   0 - 0x0
      12'h944: dout <= 8'b00000000; // 2372 :   0 - 0x0
      12'h945: dout <= 8'b00000000; // 2373 :   0 - 0x0
      12'h946: dout <= 8'b00000000; // 2374 :   0 - 0x0
      12'h947: dout <= 8'b00000000; // 2375 :   0 - 0x0
      12'h948: dout <= 8'b00000000; // 2376 :   0 - 0x0 -- Background 0x29
      12'h949: dout <= 8'b00000000; // 2377 :   0 - 0x0
      12'h94A: dout <= 8'b00000000; // 2378 :   0 - 0x0
      12'h94B: dout <= 8'b00000000; // 2379 :   0 - 0x0
      12'h94C: dout <= 8'b00000000; // 2380 :   0 - 0x0
      12'h94D: dout <= 8'b00000000; // 2381 :   0 - 0x0
      12'h94E: dout <= 8'b00000000; // 2382 :   0 - 0x0
      12'h94F: dout <= 8'b00000000; // 2383 :   0 - 0x0
      12'h950: dout <= 8'b00000000; // 2384 :   0 - 0x0 -- Background 0x2a
      12'h951: dout <= 8'b00000000; // 2385 :   0 - 0x0
      12'h952: dout <= 8'b00000000; // 2386 :   0 - 0x0
      12'h953: dout <= 8'b00000000; // 2387 :   0 - 0x0
      12'h954: dout <= 8'b00000000; // 2388 :   0 - 0x0
      12'h955: dout <= 8'b00000000; // 2389 :   0 - 0x0
      12'h956: dout <= 8'b00000000; // 2390 :   0 - 0x0
      12'h957: dout <= 8'b00000000; // 2391 :   0 - 0x0
      12'h958: dout <= 8'b00000000; // 2392 :   0 - 0x0 -- Background 0x2b
      12'h959: dout <= 8'b00000000; // 2393 :   0 - 0x0
      12'h95A: dout <= 8'b00000000; // 2394 :   0 - 0x0
      12'h95B: dout <= 8'b00000000; // 2395 :   0 - 0x0
      12'h95C: dout <= 8'b00000000; // 2396 :   0 - 0x0
      12'h95D: dout <= 8'b00000000; // 2397 :   0 - 0x0
      12'h95E: dout <= 8'b00000000; // 2398 :   0 - 0x0
      12'h95F: dout <= 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout <= 8'b00000000; // 2400 :   0 - 0x0 -- Background 0x2c
      12'h961: dout <= 8'b00000000; // 2401 :   0 - 0x0
      12'h962: dout <= 8'b00000000; // 2402 :   0 - 0x0
      12'h963: dout <= 8'b00000000; // 2403 :   0 - 0x0
      12'h964: dout <= 8'b00000000; // 2404 :   0 - 0x0
      12'h965: dout <= 8'b00000000; // 2405 :   0 - 0x0
      12'h966: dout <= 8'b00000000; // 2406 :   0 - 0x0
      12'h967: dout <= 8'b00000000; // 2407 :   0 - 0x0
      12'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0 -- Background 0x2d
      12'h969: dout <= 8'b00000000; // 2409 :   0 - 0x0
      12'h96A: dout <= 8'b00000000; // 2410 :   0 - 0x0
      12'h96B: dout <= 8'b00000000; // 2411 :   0 - 0x0
      12'h96C: dout <= 8'b00000000; // 2412 :   0 - 0x0
      12'h96D: dout <= 8'b00000000; // 2413 :   0 - 0x0
      12'h96E: dout <= 8'b00000000; // 2414 :   0 - 0x0
      12'h96F: dout <= 8'b00000000; // 2415 :   0 - 0x0
      12'h970: dout <= 8'b00000000; // 2416 :   0 - 0x0 -- Background 0x2e
      12'h971: dout <= 8'b00000000; // 2417 :   0 - 0x0
      12'h972: dout <= 8'b00000000; // 2418 :   0 - 0x0
      12'h973: dout <= 8'b00000000; // 2419 :   0 - 0x0
      12'h974: dout <= 8'b00000000; // 2420 :   0 - 0x0
      12'h975: dout <= 8'b00000000; // 2421 :   0 - 0x0
      12'h976: dout <= 8'b00000000; // 2422 :   0 - 0x0
      12'h977: dout <= 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout <= 8'b00000000; // 2424 :   0 - 0x0 -- Background 0x2f
      12'h979: dout <= 8'b00000000; // 2425 :   0 - 0x0
      12'h97A: dout <= 8'b00000000; // 2426 :   0 - 0x0
      12'h97B: dout <= 8'b00000000; // 2427 :   0 - 0x0
      12'h97C: dout <= 8'b00000000; // 2428 :   0 - 0x0
      12'h97D: dout <= 8'b00000000; // 2429 :   0 - 0x0
      12'h97E: dout <= 8'b00000000; // 2430 :   0 - 0x0
      12'h97F: dout <= 8'b00000000; // 2431 :   0 - 0x0
      12'h980: dout <= 8'b00000000; // 2432 :   0 - 0x0 -- Background 0x30
      12'h981: dout <= 8'b00000000; // 2433 :   0 - 0x0
      12'h982: dout <= 8'b00000000; // 2434 :   0 - 0x0
      12'h983: dout <= 8'b00000000; // 2435 :   0 - 0x0
      12'h984: dout <= 8'b00000000; // 2436 :   0 - 0x0
      12'h985: dout <= 8'b00000000; // 2437 :   0 - 0x0
      12'h986: dout <= 8'b00000000; // 2438 :   0 - 0x0
      12'h987: dout <= 8'b00000000; // 2439 :   0 - 0x0
      12'h988: dout <= 8'b00000000; // 2440 :   0 - 0x0 -- Background 0x31
      12'h989: dout <= 8'b00000000; // 2441 :   0 - 0x0
      12'h98A: dout <= 8'b00000000; // 2442 :   0 - 0x0
      12'h98B: dout <= 8'b00000000; // 2443 :   0 - 0x0
      12'h98C: dout <= 8'b00000000; // 2444 :   0 - 0x0
      12'h98D: dout <= 8'b00000000; // 2445 :   0 - 0x0
      12'h98E: dout <= 8'b00000000; // 2446 :   0 - 0x0
      12'h98F: dout <= 8'b00000000; // 2447 :   0 - 0x0
      12'h990: dout <= 8'b00000000; // 2448 :   0 - 0x0 -- Background 0x32
      12'h991: dout <= 8'b00000000; // 2449 :   0 - 0x0
      12'h992: dout <= 8'b00000000; // 2450 :   0 - 0x0
      12'h993: dout <= 8'b00000000; // 2451 :   0 - 0x0
      12'h994: dout <= 8'b00000000; // 2452 :   0 - 0x0
      12'h995: dout <= 8'b00000000; // 2453 :   0 - 0x0
      12'h996: dout <= 8'b00000000; // 2454 :   0 - 0x0
      12'h997: dout <= 8'b00000000; // 2455 :   0 - 0x0
      12'h998: dout <= 8'b00000000; // 2456 :   0 - 0x0 -- Background 0x33
      12'h999: dout <= 8'b00000000; // 2457 :   0 - 0x0
      12'h99A: dout <= 8'b00000000; // 2458 :   0 - 0x0
      12'h99B: dout <= 8'b00000000; // 2459 :   0 - 0x0
      12'h99C: dout <= 8'b00000000; // 2460 :   0 - 0x0
      12'h99D: dout <= 8'b00000000; // 2461 :   0 - 0x0
      12'h99E: dout <= 8'b00000000; // 2462 :   0 - 0x0
      12'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout <= 8'b00000000; // 2464 :   0 - 0x0 -- Background 0x34
      12'h9A1: dout <= 8'b00000000; // 2465 :   0 - 0x0
      12'h9A2: dout <= 8'b00000000; // 2466 :   0 - 0x0
      12'h9A3: dout <= 8'b00000000; // 2467 :   0 - 0x0
      12'h9A4: dout <= 8'b00000000; // 2468 :   0 - 0x0
      12'h9A5: dout <= 8'b00000000; // 2469 :   0 - 0x0
      12'h9A6: dout <= 8'b00000000; // 2470 :   0 - 0x0
      12'h9A7: dout <= 8'b00000000; // 2471 :   0 - 0x0
      12'h9A8: dout <= 8'b00000000; // 2472 :   0 - 0x0 -- Background 0x35
      12'h9A9: dout <= 8'b00000000; // 2473 :   0 - 0x0
      12'h9AA: dout <= 8'b00000000; // 2474 :   0 - 0x0
      12'h9AB: dout <= 8'b00000000; // 2475 :   0 - 0x0
      12'h9AC: dout <= 8'b00000000; // 2476 :   0 - 0x0
      12'h9AD: dout <= 8'b00000000; // 2477 :   0 - 0x0
      12'h9AE: dout <= 8'b00000000; // 2478 :   0 - 0x0
      12'h9AF: dout <= 8'b00000000; // 2479 :   0 - 0x0
      12'h9B0: dout <= 8'b00000000; // 2480 :   0 - 0x0 -- Background 0x36
      12'h9B1: dout <= 8'b00000000; // 2481 :   0 - 0x0
      12'h9B2: dout <= 8'b00000000; // 2482 :   0 - 0x0
      12'h9B3: dout <= 8'b00000000; // 2483 :   0 - 0x0
      12'h9B4: dout <= 8'b00000000; // 2484 :   0 - 0x0
      12'h9B5: dout <= 8'b00000000; // 2485 :   0 - 0x0
      12'h9B6: dout <= 8'b00000000; // 2486 :   0 - 0x0
      12'h9B7: dout <= 8'b00000000; // 2487 :   0 - 0x0
      12'h9B8: dout <= 8'b00000000; // 2488 :   0 - 0x0 -- Background 0x37
      12'h9B9: dout <= 8'b00000000; // 2489 :   0 - 0x0
      12'h9BA: dout <= 8'b00000000; // 2490 :   0 - 0x0
      12'h9BB: dout <= 8'b00000000; // 2491 :   0 - 0x0
      12'h9BC: dout <= 8'b00000000; // 2492 :   0 - 0x0
      12'h9BD: dout <= 8'b00000000; // 2493 :   0 - 0x0
      12'h9BE: dout <= 8'b00000000; // 2494 :   0 - 0x0
      12'h9BF: dout <= 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout <= 8'b00000000; // 2496 :   0 - 0x0 -- Background 0x38
      12'h9C1: dout <= 8'b00000000; // 2497 :   0 - 0x0
      12'h9C2: dout <= 8'b00000000; // 2498 :   0 - 0x0
      12'h9C3: dout <= 8'b00000000; // 2499 :   0 - 0x0
      12'h9C4: dout <= 8'b00000000; // 2500 :   0 - 0x0
      12'h9C5: dout <= 8'b00000000; // 2501 :   0 - 0x0
      12'h9C6: dout <= 8'b00000000; // 2502 :   0 - 0x0
      12'h9C7: dout <= 8'b00000000; // 2503 :   0 - 0x0
      12'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0 -- Background 0x39
      12'h9C9: dout <= 8'b00000000; // 2505 :   0 - 0x0
      12'h9CA: dout <= 8'b00000000; // 2506 :   0 - 0x0
      12'h9CB: dout <= 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout <= 8'b00000000; // 2508 :   0 - 0x0
      12'h9CD: dout <= 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout <= 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout <= 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout <= 8'b00000000; // 2512 :   0 - 0x0 -- Background 0x3a
      12'h9D1: dout <= 8'b00000000; // 2513 :   0 - 0x0
      12'h9D2: dout <= 8'b00000000; // 2514 :   0 - 0x0
      12'h9D3: dout <= 8'b00000000; // 2515 :   0 - 0x0
      12'h9D4: dout <= 8'b00000000; // 2516 :   0 - 0x0
      12'h9D5: dout <= 8'b00000000; // 2517 :   0 - 0x0
      12'h9D6: dout <= 8'b00000000; // 2518 :   0 - 0x0
      12'h9D7: dout <= 8'b00000000; // 2519 :   0 - 0x0
      12'h9D8: dout <= 8'b00000000; // 2520 :   0 - 0x0 -- Background 0x3b
      12'h9D9: dout <= 8'b00000000; // 2521 :   0 - 0x0
      12'h9DA: dout <= 8'b00000000; // 2522 :   0 - 0x0
      12'h9DB: dout <= 8'b00000000; // 2523 :   0 - 0x0
      12'h9DC: dout <= 8'b00000000; // 2524 :   0 - 0x0
      12'h9DD: dout <= 8'b00000000; // 2525 :   0 - 0x0
      12'h9DE: dout <= 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout <= 8'b00000000; // 2528 :   0 - 0x0 -- Background 0x3c
      12'h9E1: dout <= 8'b00000000; // 2529 :   0 - 0x0
      12'h9E2: dout <= 8'b00000000; // 2530 :   0 - 0x0
      12'h9E3: dout <= 8'b00000000; // 2531 :   0 - 0x0
      12'h9E4: dout <= 8'b00000000; // 2532 :   0 - 0x0
      12'h9E5: dout <= 8'b00000000; // 2533 :   0 - 0x0
      12'h9E6: dout <= 8'b00000000; // 2534 :   0 - 0x0
      12'h9E7: dout <= 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0 -- Background 0x3d
      12'h9E9: dout <= 8'b00000000; // 2537 :   0 - 0x0
      12'h9EA: dout <= 8'b00000000; // 2538 :   0 - 0x0
      12'h9EB: dout <= 8'b00000000; // 2539 :   0 - 0x0
      12'h9EC: dout <= 8'b00000000; // 2540 :   0 - 0x0
      12'h9ED: dout <= 8'b00000000; // 2541 :   0 - 0x0
      12'h9EE: dout <= 8'b00000000; // 2542 :   0 - 0x0
      12'h9EF: dout <= 8'b00000000; // 2543 :   0 - 0x0
      12'h9F0: dout <= 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x3e
      12'h9F1: dout <= 8'b00000000; // 2545 :   0 - 0x0
      12'h9F2: dout <= 8'b00000000; // 2546 :   0 - 0x0
      12'h9F3: dout <= 8'b00000000; // 2547 :   0 - 0x0
      12'h9F4: dout <= 8'b00000000; // 2548 :   0 - 0x0
      12'h9F5: dout <= 8'b00000000; // 2549 :   0 - 0x0
      12'h9F6: dout <= 8'b00000000; // 2550 :   0 - 0x0
      12'h9F7: dout <= 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- Background 0x3f
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout <= 8'b00000000; // 2560 :   0 - 0x0 -- Background 0x40
      12'hA01: dout <= 8'b00000000; // 2561 :   0 - 0x0
      12'hA02: dout <= 8'b00000000; // 2562 :   0 - 0x0
      12'hA03: dout <= 8'b00000000; // 2563 :   0 - 0x0
      12'hA04: dout <= 8'b00000000; // 2564 :   0 - 0x0
      12'hA05: dout <= 8'b00000000; // 2565 :   0 - 0x0
      12'hA06: dout <= 8'b00000000; // 2566 :   0 - 0x0
      12'hA07: dout <= 8'b00000000; // 2567 :   0 - 0x0
      12'hA08: dout <= 8'b00000000; // 2568 :   0 - 0x0 -- Background 0x41
      12'hA09: dout <= 8'b00000000; // 2569 :   0 - 0x0
      12'hA0A: dout <= 8'b00000000; // 2570 :   0 - 0x0
      12'hA0B: dout <= 8'b00000000; // 2571 :   0 - 0x0
      12'hA0C: dout <= 8'b00000000; // 2572 :   0 - 0x0
      12'hA0D: dout <= 8'b00000000; // 2573 :   0 - 0x0
      12'hA0E: dout <= 8'b00000000; // 2574 :   0 - 0x0
      12'hA0F: dout <= 8'b00000000; // 2575 :   0 - 0x0
      12'hA10: dout <= 8'b00000000; // 2576 :   0 - 0x0 -- Background 0x42
      12'hA11: dout <= 8'b00000000; // 2577 :   0 - 0x0
      12'hA12: dout <= 8'b00000000; // 2578 :   0 - 0x0
      12'hA13: dout <= 8'b00000000; // 2579 :   0 - 0x0
      12'hA14: dout <= 8'b00000000; // 2580 :   0 - 0x0
      12'hA15: dout <= 8'b00000000; // 2581 :   0 - 0x0
      12'hA16: dout <= 8'b00000000; // 2582 :   0 - 0x0
      12'hA17: dout <= 8'b00000000; // 2583 :   0 - 0x0
      12'hA18: dout <= 8'b00000000; // 2584 :   0 - 0x0 -- Background 0x43
      12'hA19: dout <= 8'b00000000; // 2585 :   0 - 0x0
      12'hA1A: dout <= 8'b00000000; // 2586 :   0 - 0x0
      12'hA1B: dout <= 8'b00000000; // 2587 :   0 - 0x0
      12'hA1C: dout <= 8'b00000000; // 2588 :   0 - 0x0
      12'hA1D: dout <= 8'b00000000; // 2589 :   0 - 0x0
      12'hA1E: dout <= 8'b00000000; // 2590 :   0 - 0x0
      12'hA1F: dout <= 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout <= 8'b00000000; // 2592 :   0 - 0x0 -- Background 0x44
      12'hA21: dout <= 8'b00000000; // 2593 :   0 - 0x0
      12'hA22: dout <= 8'b00000000; // 2594 :   0 - 0x0
      12'hA23: dout <= 8'b00000000; // 2595 :   0 - 0x0
      12'hA24: dout <= 8'b00000000; // 2596 :   0 - 0x0
      12'hA25: dout <= 8'b00000000; // 2597 :   0 - 0x0
      12'hA26: dout <= 8'b00000000; // 2598 :   0 - 0x0
      12'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0 -- Background 0x45
      12'hA29: dout <= 8'b00000000; // 2601 :   0 - 0x0
      12'hA2A: dout <= 8'b00000000; // 2602 :   0 - 0x0
      12'hA2B: dout <= 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout <= 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout <= 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout <= 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout <= 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout <= 8'b00000000; // 2608 :   0 - 0x0 -- Background 0x46
      12'hA31: dout <= 8'b00000000; // 2609 :   0 - 0x0
      12'hA32: dout <= 8'b00000000; // 2610 :   0 - 0x0
      12'hA33: dout <= 8'b00000000; // 2611 :   0 - 0x0
      12'hA34: dout <= 8'b00000000; // 2612 :   0 - 0x0
      12'hA35: dout <= 8'b00000000; // 2613 :   0 - 0x0
      12'hA36: dout <= 8'b00000000; // 2614 :   0 - 0x0
      12'hA37: dout <= 8'b00000000; // 2615 :   0 - 0x0
      12'hA38: dout <= 8'b00000000; // 2616 :   0 - 0x0 -- Background 0x47
      12'hA39: dout <= 8'b00000000; // 2617 :   0 - 0x0
      12'hA3A: dout <= 8'b00000000; // 2618 :   0 - 0x0
      12'hA3B: dout <= 8'b00000000; // 2619 :   0 - 0x0
      12'hA3C: dout <= 8'b00000000; // 2620 :   0 - 0x0
      12'hA3D: dout <= 8'b00000000; // 2621 :   0 - 0x0
      12'hA3E: dout <= 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout <= 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout <= 8'b00000000; // 2624 :   0 - 0x0 -- Background 0x48
      12'hA41: dout <= 8'b00000000; // 2625 :   0 - 0x0
      12'hA42: dout <= 8'b00000000; // 2626 :   0 - 0x0
      12'hA43: dout <= 8'b00000000; // 2627 :   0 - 0x0
      12'hA44: dout <= 8'b00000000; // 2628 :   0 - 0x0
      12'hA45: dout <= 8'b00000000; // 2629 :   0 - 0x0
      12'hA46: dout <= 8'b00000000; // 2630 :   0 - 0x0
      12'hA47: dout <= 8'b00000000; // 2631 :   0 - 0x0
      12'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0 -- Background 0x49
      12'hA49: dout <= 8'b00000000; // 2633 :   0 - 0x0
      12'hA4A: dout <= 8'b00000000; // 2634 :   0 - 0x0
      12'hA4B: dout <= 8'b00000000; // 2635 :   0 - 0x0
      12'hA4C: dout <= 8'b00000000; // 2636 :   0 - 0x0
      12'hA4D: dout <= 8'b00000000; // 2637 :   0 - 0x0
      12'hA4E: dout <= 8'b00000000; // 2638 :   0 - 0x0
      12'hA4F: dout <= 8'b00000000; // 2639 :   0 - 0x0
      12'hA50: dout <= 8'b00000000; // 2640 :   0 - 0x0 -- Background 0x4a
      12'hA51: dout <= 8'b00000000; // 2641 :   0 - 0x0
      12'hA52: dout <= 8'b00000000; // 2642 :   0 - 0x0
      12'hA53: dout <= 8'b00000000; // 2643 :   0 - 0x0
      12'hA54: dout <= 8'b00000000; // 2644 :   0 - 0x0
      12'hA55: dout <= 8'b00000000; // 2645 :   0 - 0x0
      12'hA56: dout <= 8'b00000000; // 2646 :   0 - 0x0
      12'hA57: dout <= 8'b00000000; // 2647 :   0 - 0x0
      12'hA58: dout <= 8'b00000000; // 2648 :   0 - 0x0 -- Background 0x4b
      12'hA59: dout <= 8'b00000000; // 2649 :   0 - 0x0
      12'hA5A: dout <= 8'b00000000; // 2650 :   0 - 0x0
      12'hA5B: dout <= 8'b00000000; // 2651 :   0 - 0x0
      12'hA5C: dout <= 8'b00000000; // 2652 :   0 - 0x0
      12'hA5D: dout <= 8'b00000000; // 2653 :   0 - 0x0
      12'hA5E: dout <= 8'b00000000; // 2654 :   0 - 0x0
      12'hA5F: dout <= 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout <= 8'b00000000; // 2656 :   0 - 0x0 -- Background 0x4c
      12'hA61: dout <= 8'b00000000; // 2657 :   0 - 0x0
      12'hA62: dout <= 8'b00000000; // 2658 :   0 - 0x0
      12'hA63: dout <= 8'b00000000; // 2659 :   0 - 0x0
      12'hA64: dout <= 8'b00000000; // 2660 :   0 - 0x0
      12'hA65: dout <= 8'b00000000; // 2661 :   0 - 0x0
      12'hA66: dout <= 8'b00000000; // 2662 :   0 - 0x0
      12'hA67: dout <= 8'b00000000; // 2663 :   0 - 0x0
      12'hA68: dout <= 8'b00000000; // 2664 :   0 - 0x0 -- Background 0x4d
      12'hA69: dout <= 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout <= 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout <= 8'b00000001; // 2667 :   1 - 0x1
      12'hA6C: dout <= 8'b00000011; // 2668 :   3 - 0x3
      12'hA6D: dout <= 8'b00000111; // 2669 :   7 - 0x7
      12'hA6E: dout <= 8'b00001111; // 2670 :  15 - 0xf
      12'hA6F: dout <= 8'b00011111; // 2671 :  31 - 0x1f
      12'hA70: dout <= 8'b00000000; // 2672 :   0 - 0x0 -- Background 0x4e
      12'hA71: dout <= 8'b00001111; // 2673 :  15 - 0xf
      12'hA72: dout <= 8'b01111111; // 2674 : 127 - 0x7f
      12'hA73: dout <= 8'b11111111; // 2675 : 255 - 0xff
      12'hA74: dout <= 8'b11111111; // 2676 : 255 - 0xff
      12'hA75: dout <= 8'b11111111; // 2677 : 255 - 0xff
      12'hA76: dout <= 8'b11111111; // 2678 : 255 - 0xff
      12'hA77: dout <= 8'b11111111; // 2679 : 255 - 0xff
      12'hA78: dout <= 8'b00011111; // 2680 :  31 - 0x1f -- Background 0x4f
      12'hA79: dout <= 8'b00111111; // 2681 :  63 - 0x3f
      12'hA7A: dout <= 8'b00111111; // 2682 :  63 - 0x3f
      12'hA7B: dout <= 8'b00111111; // 2683 :  63 - 0x3f
      12'hA7C: dout <= 8'b01111111; // 2684 : 127 - 0x7f
      12'hA7D: dout <= 8'b01111111; // 2685 : 127 - 0x7f
      12'hA7E: dout <= 8'b01111111; // 2686 : 127 - 0x7f
      12'hA7F: dout <= 8'b01111111; // 2687 : 127 - 0x7f
      12'hA80: dout <= 8'b11111111; // 2688 : 255 - 0xff -- Background 0x50
      12'hA81: dout <= 8'b11111111; // 2689 : 255 - 0xff
      12'hA82: dout <= 8'b11111111; // 2690 : 255 - 0xff
      12'hA83: dout <= 8'b11111111; // 2691 : 255 - 0xff
      12'hA84: dout <= 8'b11111111; // 2692 : 255 - 0xff
      12'hA85: dout <= 8'b11111111; // 2693 : 255 - 0xff
      12'hA86: dout <= 8'b11111111; // 2694 : 255 - 0xff
      12'hA87: dout <= 8'b11111111; // 2695 : 255 - 0xff
      12'hA88: dout <= 8'b11111111; // 2696 : 255 - 0xff -- Background 0x51
      12'hA89: dout <= 8'b11111111; // 2697 : 255 - 0xff
      12'hA8A: dout <= 8'b11111111; // 2698 : 255 - 0xff
      12'hA8B: dout <= 8'b11111111; // 2699 : 255 - 0xff
      12'hA8C: dout <= 8'b11111111; // 2700 : 255 - 0xff
      12'hA8D: dout <= 8'b11111111; // 2701 : 255 - 0xff
      12'hA8E: dout <= 8'b11111111; // 2702 : 255 - 0xff
      12'hA8F: dout <= 8'b11111110; // 2703 : 254 - 0xfe
      12'hA90: dout <= 8'b00000000; // 2704 :   0 - 0x0 -- Background 0x52
      12'hA91: dout <= 8'b00000000; // 2705 :   0 - 0x0
      12'hA92: dout <= 8'b00000000; // 2706 :   0 - 0x0
      12'hA93: dout <= 8'b10000000; // 2707 : 128 - 0x80
      12'hA94: dout <= 8'b11000000; // 2708 : 192 - 0xc0
      12'hA95: dout <= 8'b11100000; // 2709 : 224 - 0xe0
      12'hA96: dout <= 8'b11110000; // 2710 : 240 - 0xf0
      12'hA97: dout <= 8'b11110000; // 2711 : 240 - 0xf0
      12'hA98: dout <= 8'b11111111; // 2712 : 255 - 0xff -- Background 0x53
      12'hA99: dout <= 8'b11111111; // 2713 : 255 - 0xff
      12'hA9A: dout <= 8'b11111110; // 2714 : 254 - 0xfe
      12'hA9B: dout <= 8'b11111100; // 2715 : 252 - 0xfc
      12'hA9C: dout <= 8'b11110000; // 2716 : 240 - 0xf0
      12'hA9D: dout <= 8'b11100000; // 2717 : 224 - 0xe0
      12'hA9E: dout <= 8'b10000000; // 2718 : 128 - 0x80
      12'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout <= 8'b11000000; // 2720 : 192 - 0xc0 -- Background 0x54
      12'hAA1: dout <= 8'b10000000; // 2721 : 128 - 0x80
      12'hAA2: dout <= 8'b00000000; // 2722 :   0 - 0x0
      12'hAA3: dout <= 8'b00000000; // 2723 :   0 - 0x0
      12'hAA4: dout <= 8'b00000000; // 2724 :   0 - 0x0
      12'hAA5: dout <= 8'b00000000; // 2725 :   0 - 0x0
      12'hAA6: dout <= 8'b00000000; // 2726 :   0 - 0x0
      12'hAA7: dout <= 8'b00000000; // 2727 :   0 - 0x0
      12'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0 -- Background 0x55
      12'hAA9: dout <= 8'b11110000; // 2729 : 240 - 0xf0
      12'hAAA: dout <= 8'b11111110; // 2730 : 254 - 0xfe
      12'hAAB: dout <= 8'b11111110; // 2731 : 254 - 0xfe
      12'hAAC: dout <= 8'b11111110; // 2732 : 254 - 0xfe
      12'hAAD: dout <= 8'b11111100; // 2733 : 252 - 0xfc
      12'hAAE: dout <= 8'b11111000; // 2734 : 248 - 0xf8
      12'hAAF: dout <= 8'b11111000; // 2735 : 248 - 0xf8
      12'hAB0: dout <= 8'b11110000; // 2736 : 240 - 0xf0 -- Background 0x56
      12'hAB1: dout <= 8'b11100000; // 2737 : 224 - 0xe0
      12'hAB2: dout <= 8'b11100000; // 2738 : 224 - 0xe0
      12'hAB3: dout <= 8'b11000000; // 2739 : 192 - 0xc0
      12'hAB4: dout <= 8'b10000000; // 2740 : 128 - 0x80
      12'hAB5: dout <= 8'b10000000; // 2741 : 128 - 0x80
      12'hAB6: dout <= 8'b00000000; // 2742 :   0 - 0x0
      12'hAB7: dout <= 8'b00000000; // 2743 :   0 - 0x0
      12'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0 -- Background 0x57
      12'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout <= 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout <= 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout <= 8'b00000100; // 2751 :   4 - 0x4
      12'hAC0: dout <= 8'b00000110; // 2752 :   6 - 0x6 -- Background 0x58
      12'hAC1: dout <= 8'b00000110; // 2753 :   6 - 0x6
      12'hAC2: dout <= 8'b00000111; // 2754 :   7 - 0x7
      12'hAC3: dout <= 8'b00000111; // 2755 :   7 - 0x7
      12'hAC4: dout <= 8'b00000111; // 2756 :   7 - 0x7
      12'hAC5: dout <= 8'b00000111; // 2757 :   7 - 0x7
      12'hAC6: dout <= 8'b00000000; // 2758 :   0 - 0x0
      12'hAC7: dout <= 8'b00000000; // 2759 :   0 - 0x0
      12'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0 -- Background 0x59
      12'hAC9: dout <= 8'b00000000; // 2761 :   0 - 0x0
      12'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout <= 8'b00000000; // 2763 :   0 - 0x0
      12'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      12'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout <= 8'b00010000; // 2767 :  16 - 0x10
      12'hAD0: dout <= 8'b00011100; // 2768 :  28 - 0x1c -- Background 0x5a
      12'hAD1: dout <= 8'b00011110; // 2769 :  30 - 0x1e
      12'hAD2: dout <= 8'b00011111; // 2770 :  31 - 0x1f
      12'hAD3: dout <= 8'b00011111; // 2771 :  31 - 0x1f
      12'hAD4: dout <= 8'b00011111; // 2772 :  31 - 0x1f
      12'hAD5: dout <= 8'b00011111; // 2773 :  31 - 0x1f
      12'hAD6: dout <= 8'b00000000; // 2774 :   0 - 0x0
      12'hAD7: dout <= 8'b00000000; // 2775 :   0 - 0x0
      12'hAD8: dout <= 8'b00000000; // 2776 :   0 - 0x0 -- Background 0x5b
      12'hAD9: dout <= 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout <= 8'b00000000; // 2778 :   0 - 0x0
      12'hADB: dout <= 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout <= 8'b00000000; // 2780 :   0 - 0x0
      12'hADD: dout <= 8'b00000000; // 2781 :   0 - 0x0
      12'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      12'hADF: dout <= 8'b11000000; // 2783 : 192 - 0xc0
      12'hAE0: dout <= 8'b11110000; // 2784 : 240 - 0xf0 -- Background 0x5c
      12'hAE1: dout <= 8'b11111100; // 2785 : 252 - 0xfc
      12'hAE2: dout <= 8'b11111111; // 2786 : 255 - 0xff
      12'hAE3: dout <= 8'b11111111; // 2787 : 255 - 0xff
      12'hAE4: dout <= 8'b11111111; // 2788 : 255 - 0xff
      12'hAE5: dout <= 8'b11111111; // 2789 : 255 - 0xff
      12'hAE6: dout <= 8'b00000000; // 2790 :   0 - 0x0
      12'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0 -- Background 0x5d
      12'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout <= 8'b00000001; // 2794 :   1 - 0x1
      12'hAEB: dout <= 8'b00000011; // 2795 :   3 - 0x3
      12'hAEC: dout <= 8'b00001111; // 2796 :  15 - 0xf
      12'hAED: dout <= 8'b00001111; // 2797 :  15 - 0xf
      12'hAEE: dout <= 8'b00000000; // 2798 :   0 - 0x0
      12'hAEF: dout <= 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout <= 8'b11111100; // 2800 : 252 - 0xfc -- Background 0x5e
      12'hAF1: dout <= 8'b11111100; // 2801 : 252 - 0xfc
      12'hAF2: dout <= 8'b11111100; // 2802 : 252 - 0xfc
      12'hAF3: dout <= 8'b11111100; // 2803 : 252 - 0xfc
      12'hAF4: dout <= 8'b11111000; // 2804 : 248 - 0xf8
      12'hAF5: dout <= 8'b11111100; // 2805 : 252 - 0xfc
      12'hAF6: dout <= 8'b00111100; // 2806 :  60 - 0x3c
      12'hAF7: dout <= 8'b00000000; // 2807 :   0 - 0x0
      12'hAF8: dout <= 8'b00000100; // 2808 :   4 - 0x4 -- Background 0x5f
      12'hAF9: dout <= 8'b00001100; // 2809 :  12 - 0xc
      12'hAFA: dout <= 8'b00011100; // 2810 :  28 - 0x1c
      12'hAFB: dout <= 8'b00001100; // 2811 :  12 - 0xc
      12'hAFC: dout <= 8'b00011000; // 2812 :  24 - 0x18
      12'hAFD: dout <= 8'b00111100; // 2813 :  60 - 0x3c
      12'hAFE: dout <= 8'b00111100; // 2814 :  60 - 0x3c
      12'hAFF: dout <= 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout <= 8'b00000000; // 2816 :   0 - 0x0 -- Background 0x60
      12'hB01: dout <= 8'b00000011; // 2817 :   3 - 0x3
      12'hB02: dout <= 8'b00001111; // 2818 :  15 - 0xf
      12'hB03: dout <= 8'b00010011; // 2819 :  19 - 0x13
      12'hB04: dout <= 8'b00100001; // 2820 :  33 - 0x21
      12'hB05: dout <= 8'b00100001; // 2821 :  33 - 0x21
      12'hB06: dout <= 8'b00100001; // 2822 :  33 - 0x21
      12'hB07: dout <= 8'b01110011; // 2823 : 115 - 0x73
      12'hB08: dout <= 8'b00000000; // 2824 :   0 - 0x0 -- Background 0x61
      12'hB09: dout <= 8'b11000000; // 2825 : 192 - 0xc0
      12'hB0A: dout <= 8'b11110000; // 2826 : 240 - 0xf0
      12'hB0B: dout <= 8'b11001000; // 2827 : 200 - 0xc8
      12'hB0C: dout <= 8'b10000100; // 2828 : 132 - 0x84
      12'hB0D: dout <= 8'b10000100; // 2829 : 132 - 0x84
      12'hB0E: dout <= 8'b10000100; // 2830 : 132 - 0x84
      12'hB0F: dout <= 8'b11001110; // 2831 : 206 - 0xce
      12'hB10: dout <= 8'b10010100; // 2832 : 148 - 0x94 -- Background 0x62
      12'hB11: dout <= 8'b11101010; // 2833 : 234 - 0xea
      12'hB12: dout <= 8'b11011110; // 2834 : 222 - 0xde
      12'hB13: dout <= 8'b11101110; // 2835 : 238 - 0xee
      12'hB14: dout <= 8'b11011110; // 2836 : 222 - 0xde
      12'hB15: dout <= 8'b01100110; // 2837 : 102 - 0x66
      12'hB16: dout <= 8'b01000010; // 2838 :  66 - 0x42
      12'hB17: dout <= 8'b00000000; // 2839 :   0 - 0x0
      12'hB18: dout <= 8'b10010100; // 2840 : 148 - 0x94 -- Background 0x63
      12'hB19: dout <= 8'b11101010; // 2841 : 234 - 0xea
      12'hB1A: dout <= 8'b11011110; // 2842 : 222 - 0xde
      12'hB1B: dout <= 8'b11101110; // 2843 : 238 - 0xee
      12'hB1C: dout <= 8'b11011110; // 2844 : 222 - 0xde
      12'hB1D: dout <= 8'b11001110; // 2845 : 206 - 0xce
      12'hB1E: dout <= 8'b10001100; // 2846 : 140 - 0x8c
      12'hB1F: dout <= 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout <= 8'b00000000; // 2848 :   0 - 0x0 -- Background 0x64
      12'hB21: dout <= 8'b00000000; // 2849 :   0 - 0x0
      12'hB22: dout <= 8'b00000000; // 2850 :   0 - 0x0
      12'hB23: dout <= 8'b00000000; // 2851 :   0 - 0x0
      12'hB24: dout <= 8'b00000000; // 2852 :   0 - 0x0
      12'hB25: dout <= 8'b00000000; // 2853 :   0 - 0x0
      12'hB26: dout <= 8'b00000000; // 2854 :   0 - 0x0
      12'hB27: dout <= 8'b00000001; // 2855 :   1 - 0x1
      12'hB28: dout <= 8'b00000000; // 2856 :   0 - 0x0 -- Background 0x65
      12'hB29: dout <= 8'b00000000; // 2857 :   0 - 0x0
      12'hB2A: dout <= 8'b00000000; // 2858 :   0 - 0x0
      12'hB2B: dout <= 8'b00000000; // 2859 :   0 - 0x0
      12'hB2C: dout <= 8'b00000000; // 2860 :   0 - 0x0
      12'hB2D: dout <= 8'b00110110; // 2861 :  54 - 0x36
      12'hB2E: dout <= 8'b00110110; // 2862 :  54 - 0x36
      12'hB2F: dout <= 8'b10010000; // 2863 : 144 - 0x90
      12'hB30: dout <= 8'b00000001; // 2864 :   1 - 0x1 -- Background 0x66
      12'hB31: dout <= 8'b00000011; // 2865 :   3 - 0x3
      12'hB32: dout <= 8'b00000111; // 2866 :   7 - 0x7
      12'hB33: dout <= 8'b00000111; // 2867 :   7 - 0x7
      12'hB34: dout <= 8'b00011111; // 2868 :  31 - 0x1f
      12'hB35: dout <= 8'b00011111; // 2869 :  31 - 0x1f
      12'hB36: dout <= 8'b00011100; // 2870 :  28 - 0x1c
      12'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      12'hB38: dout <= 8'b11111000; // 2872 : 248 - 0xf8 -- Background 0x67
      12'hB39: dout <= 8'b11111000; // 2873 : 248 - 0xf8
      12'hB3A: dout <= 8'b11111000; // 2874 : 248 - 0xf8
      12'hB3B: dout <= 8'b11111000; // 2875 : 248 - 0xf8
      12'hB3C: dout <= 8'b11111110; // 2876 : 254 - 0xfe
      12'hB3D: dout <= 8'b11111110; // 2877 : 254 - 0xfe
      12'hB3E: dout <= 8'b00001110; // 2878 :  14 - 0xe
      12'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout <= 8'b00000111; // 2880 :   7 - 0x7 -- Background 0x68
      12'hB41: dout <= 8'b00001111; // 2881 :  15 - 0xf
      12'hB42: dout <= 8'b00011111; // 2882 :  31 - 0x1f
      12'hB43: dout <= 8'b00011111; // 2883 :  31 - 0x1f
      12'hB44: dout <= 8'b00111111; // 2884 :  63 - 0x3f
      12'hB45: dout <= 8'b00111111; // 2885 :  63 - 0x3f
      12'hB46: dout <= 8'b00111000; // 2886 :  56 - 0x38
      12'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout <= 8'b11111000; // 2888 : 248 - 0xf8 -- Background 0x69
      12'hB49: dout <= 8'b11110000; // 2889 : 240 - 0xf0
      12'hB4A: dout <= 8'b11110000; // 2890 : 240 - 0xf0
      12'hB4B: dout <= 8'b11100000; // 2891 : 224 - 0xe0
      12'hB4C: dout <= 8'b11111000; // 2892 : 248 - 0xf8
      12'hB4D: dout <= 8'b11111000; // 2893 : 248 - 0xf8
      12'hB4E: dout <= 8'b00111000; // 2894 :  56 - 0x38
      12'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout <= 8'b00000000; // 2896 :   0 - 0x0 -- Background 0x6a
      12'hB51: dout <= 8'b00011111; // 2897 :  31 - 0x1f
      12'hB52: dout <= 8'b01111111; // 2898 : 127 - 0x7f
      12'hB53: dout <= 8'b00111111; // 2899 :  63 - 0x3f
      12'hB54: dout <= 8'b00001111; // 2900 :  15 - 0xf
      12'hB55: dout <= 8'b00000111; // 2901 :   7 - 0x7
      12'hB56: dout <= 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout <= 8'b00000000; // 2904 :   0 - 0x0 -- Background 0x6b
      12'hB59: dout <= 8'b00000000; // 2905 :   0 - 0x0
      12'hB5A: dout <= 8'b11000000; // 2906 : 192 - 0xc0
      12'hB5B: dout <= 8'b11110000; // 2907 : 240 - 0xf0
      12'hB5C: dout <= 8'b11111000; // 2908 : 248 - 0xf8
      12'hB5D: dout <= 8'b11111000; // 2909 : 248 - 0xf8
      12'hB5E: dout <= 8'b11100000; // 2910 : 224 - 0xe0
      12'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout <= 8'b00000000; // 2912 :   0 - 0x0 -- Background 0x6c
      12'hB61: dout <= 8'b00000000; // 2913 :   0 - 0x0
      12'hB62: dout <= 8'b00000000; // 2914 :   0 - 0x0
      12'hB63: dout <= 8'b00000000; // 2915 :   0 - 0x0
      12'hB64: dout <= 8'b00000000; // 2916 :   0 - 0x0
      12'hB65: dout <= 8'b00000000; // 2917 :   0 - 0x0
      12'hB66: dout <= 8'b00000000; // 2918 :   0 - 0x0
      12'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout <= 8'b00000000; // 2920 :   0 - 0x0 -- Background 0x6d
      12'hB69: dout <= 8'b00000000; // 2921 :   0 - 0x0
      12'hB6A: dout <= 8'b00000000; // 2922 :   0 - 0x0
      12'hB6B: dout <= 8'b00000000; // 2923 :   0 - 0x0
      12'hB6C: dout <= 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout <= 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout <= 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout <= 8'b00000000; // 2928 :   0 - 0x0 -- Background 0x6e
      12'hB71: dout <= 8'b00000000; // 2929 :   0 - 0x0
      12'hB72: dout <= 8'b00000000; // 2930 :   0 - 0x0
      12'hB73: dout <= 8'b00000000; // 2931 :   0 - 0x0
      12'hB74: dout <= 8'b00000000; // 2932 :   0 - 0x0
      12'hB75: dout <= 8'b00000000; // 2933 :   0 - 0x0
      12'hB76: dout <= 8'b00000000; // 2934 :   0 - 0x0
      12'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout <= 8'b00000000; // 2936 :   0 - 0x0 -- Background 0x6f
      12'hB79: dout <= 8'b00000000; // 2937 :   0 - 0x0
      12'hB7A: dout <= 8'b00000000; // 2938 :   0 - 0x0
      12'hB7B: dout <= 8'b00000000; // 2939 :   0 - 0x0
      12'hB7C: dout <= 8'b00000000; // 2940 :   0 - 0x0
      12'hB7D: dout <= 8'b00000000; // 2941 :   0 - 0x0
      12'hB7E: dout <= 8'b00000000; // 2942 :   0 - 0x0
      12'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout <= 8'b11111111; // 2944 : 255 - 0xff -- Background 0x70
      12'hB81: dout <= 8'b11111111; // 2945 : 255 - 0xff
      12'hB82: dout <= 8'b11111111; // 2946 : 255 - 0xff
      12'hB83: dout <= 8'b11111111; // 2947 : 255 - 0xff
      12'hB84: dout <= 8'b11111111; // 2948 : 255 - 0xff
      12'hB85: dout <= 8'b11111111; // 2949 : 255 - 0xff
      12'hB86: dout <= 8'b11111111; // 2950 : 255 - 0xff
      12'hB87: dout <= 8'b11111111; // 2951 : 255 - 0xff
      12'hB88: dout <= 8'b11111111; // 2952 : 255 - 0xff -- Background 0x71
      12'hB89: dout <= 8'b11111111; // 2953 : 255 - 0xff
      12'hB8A: dout <= 8'b11111111; // 2954 : 255 - 0xff
      12'hB8B: dout <= 8'b11111111; // 2955 : 255 - 0xff
      12'hB8C: dout <= 8'b11111111; // 2956 : 255 - 0xff
      12'hB8D: dout <= 8'b11111111; // 2957 : 255 - 0xff
      12'hB8E: dout <= 8'b11111111; // 2958 : 255 - 0xff
      12'hB8F: dout <= 8'b11111111; // 2959 : 255 - 0xff
      12'hB90: dout <= 8'b11111111; // 2960 : 255 - 0xff -- Background 0x72
      12'hB91: dout <= 8'b11111111; // 2961 : 255 - 0xff
      12'hB92: dout <= 8'b11111111; // 2962 : 255 - 0xff
      12'hB93: dout <= 8'b11111111; // 2963 : 255 - 0xff
      12'hB94: dout <= 8'b11111111; // 2964 : 255 - 0xff
      12'hB95: dout <= 8'b11111111; // 2965 : 255 - 0xff
      12'hB96: dout <= 8'b11111111; // 2966 : 255 - 0xff
      12'hB97: dout <= 8'b11111111; // 2967 : 255 - 0xff
      12'hB98: dout <= 8'b11111111; // 2968 : 255 - 0xff -- Background 0x73
      12'hB99: dout <= 8'b11111111; // 2969 : 255 - 0xff
      12'hB9A: dout <= 8'b11111111; // 2970 : 255 - 0xff
      12'hB9B: dout <= 8'b11111111; // 2971 : 255 - 0xff
      12'hB9C: dout <= 8'b11111111; // 2972 : 255 - 0xff
      12'hB9D: dout <= 8'b11111111; // 2973 : 255 - 0xff
      12'hB9E: dout <= 8'b11111111; // 2974 : 255 - 0xff
      12'hB9F: dout <= 8'b11111111; // 2975 : 255 - 0xff
      12'hBA0: dout <= 8'b11111111; // 2976 : 255 - 0xff -- Background 0x74
      12'hBA1: dout <= 8'b11111111; // 2977 : 255 - 0xff
      12'hBA2: dout <= 8'b11111111; // 2978 : 255 - 0xff
      12'hBA3: dout <= 8'b11111111; // 2979 : 255 - 0xff
      12'hBA4: dout <= 8'b11111111; // 2980 : 255 - 0xff
      12'hBA5: dout <= 8'b11111111; // 2981 : 255 - 0xff
      12'hBA6: dout <= 8'b11111111; // 2982 : 255 - 0xff
      12'hBA7: dout <= 8'b11111111; // 2983 : 255 - 0xff
      12'hBA8: dout <= 8'b11111111; // 2984 : 255 - 0xff -- Background 0x75
      12'hBA9: dout <= 8'b11111111; // 2985 : 255 - 0xff
      12'hBAA: dout <= 8'b11111111; // 2986 : 255 - 0xff
      12'hBAB: dout <= 8'b11111111; // 2987 : 255 - 0xff
      12'hBAC: dout <= 8'b11111111; // 2988 : 255 - 0xff
      12'hBAD: dout <= 8'b11111111; // 2989 : 255 - 0xff
      12'hBAE: dout <= 8'b11111111; // 2990 : 255 - 0xff
      12'hBAF: dout <= 8'b11111111; // 2991 : 255 - 0xff
      12'hBB0: dout <= 8'b11111111; // 2992 : 255 - 0xff -- Background 0x76
      12'hBB1: dout <= 8'b11111111; // 2993 : 255 - 0xff
      12'hBB2: dout <= 8'b11111111; // 2994 : 255 - 0xff
      12'hBB3: dout <= 8'b11111111; // 2995 : 255 - 0xff
      12'hBB4: dout <= 8'b11111111; // 2996 : 255 - 0xff
      12'hBB5: dout <= 8'b11111111; // 2997 : 255 - 0xff
      12'hBB6: dout <= 8'b11111111; // 2998 : 255 - 0xff
      12'hBB7: dout <= 8'b11111111; // 2999 : 255 - 0xff
      12'hBB8: dout <= 8'b11111111; // 3000 : 255 - 0xff -- Background 0x77
      12'hBB9: dout <= 8'b11111111; // 3001 : 255 - 0xff
      12'hBBA: dout <= 8'b11111111; // 3002 : 255 - 0xff
      12'hBBB: dout <= 8'b11111111; // 3003 : 255 - 0xff
      12'hBBC: dout <= 8'b11111111; // 3004 : 255 - 0xff
      12'hBBD: dout <= 8'b11111111; // 3005 : 255 - 0xff
      12'hBBE: dout <= 8'b11111111; // 3006 : 255 - 0xff
      12'hBBF: dout <= 8'b11111111; // 3007 : 255 - 0xff
      12'hBC0: dout <= 8'b11111111; // 3008 : 255 - 0xff -- Background 0x78
      12'hBC1: dout <= 8'b11111111; // 3009 : 255 - 0xff
      12'hBC2: dout <= 8'b11111111; // 3010 : 255 - 0xff
      12'hBC3: dout <= 8'b11111111; // 3011 : 255 - 0xff
      12'hBC4: dout <= 8'b11111111; // 3012 : 255 - 0xff
      12'hBC5: dout <= 8'b11111111; // 3013 : 255 - 0xff
      12'hBC6: dout <= 8'b11111111; // 3014 : 255 - 0xff
      12'hBC7: dout <= 8'b11111111; // 3015 : 255 - 0xff
      12'hBC8: dout <= 8'b11111111; // 3016 : 255 - 0xff -- Background 0x79
      12'hBC9: dout <= 8'b11111111; // 3017 : 255 - 0xff
      12'hBCA: dout <= 8'b11111111; // 3018 : 255 - 0xff
      12'hBCB: dout <= 8'b11111111; // 3019 : 255 - 0xff
      12'hBCC: dout <= 8'b11111111; // 3020 : 255 - 0xff
      12'hBCD: dout <= 8'b11111111; // 3021 : 255 - 0xff
      12'hBCE: dout <= 8'b11111111; // 3022 : 255 - 0xff
      12'hBCF: dout <= 8'b11111111; // 3023 : 255 - 0xff
      12'hBD0: dout <= 8'b11111111; // 3024 : 255 - 0xff -- Background 0x7a
      12'hBD1: dout <= 8'b11111111; // 3025 : 255 - 0xff
      12'hBD2: dout <= 8'b11111111; // 3026 : 255 - 0xff
      12'hBD3: dout <= 8'b11111111; // 3027 : 255 - 0xff
      12'hBD4: dout <= 8'b11111111; // 3028 : 255 - 0xff
      12'hBD5: dout <= 8'b11111111; // 3029 : 255 - 0xff
      12'hBD6: dout <= 8'b11111111; // 3030 : 255 - 0xff
      12'hBD7: dout <= 8'b11111111; // 3031 : 255 - 0xff
      12'hBD8: dout <= 8'b11111111; // 3032 : 255 - 0xff -- Background 0x7b
      12'hBD9: dout <= 8'b11111111; // 3033 : 255 - 0xff
      12'hBDA: dout <= 8'b11111111; // 3034 : 255 - 0xff
      12'hBDB: dout <= 8'b11111111; // 3035 : 255 - 0xff
      12'hBDC: dout <= 8'b11111111; // 3036 : 255 - 0xff
      12'hBDD: dout <= 8'b11111111; // 3037 : 255 - 0xff
      12'hBDE: dout <= 8'b11111111; // 3038 : 255 - 0xff
      12'hBDF: dout <= 8'b11111111; // 3039 : 255 - 0xff
      12'hBE0: dout <= 8'b11111111; // 3040 : 255 - 0xff -- Background 0x7c
      12'hBE1: dout <= 8'b11111111; // 3041 : 255 - 0xff
      12'hBE2: dout <= 8'b11111111; // 3042 : 255 - 0xff
      12'hBE3: dout <= 8'b11111111; // 3043 : 255 - 0xff
      12'hBE4: dout <= 8'b11111111; // 3044 : 255 - 0xff
      12'hBE5: dout <= 8'b11111111; // 3045 : 255 - 0xff
      12'hBE6: dout <= 8'b11111111; // 3046 : 255 - 0xff
      12'hBE7: dout <= 8'b11111111; // 3047 : 255 - 0xff
      12'hBE8: dout <= 8'b11111111; // 3048 : 255 - 0xff -- Background 0x7d
      12'hBE9: dout <= 8'b11111111; // 3049 : 255 - 0xff
      12'hBEA: dout <= 8'b11111111; // 3050 : 255 - 0xff
      12'hBEB: dout <= 8'b11111111; // 3051 : 255 - 0xff
      12'hBEC: dout <= 8'b11111111; // 3052 : 255 - 0xff
      12'hBED: dout <= 8'b11111111; // 3053 : 255 - 0xff
      12'hBEE: dout <= 8'b11111111; // 3054 : 255 - 0xff
      12'hBEF: dout <= 8'b11111111; // 3055 : 255 - 0xff
      12'hBF0: dout <= 8'b11111111; // 3056 : 255 - 0xff -- Background 0x7e
      12'hBF1: dout <= 8'b11111111; // 3057 : 255 - 0xff
      12'hBF2: dout <= 8'b11111111; // 3058 : 255 - 0xff
      12'hBF3: dout <= 8'b11111111; // 3059 : 255 - 0xff
      12'hBF4: dout <= 8'b11111111; // 3060 : 255 - 0xff
      12'hBF5: dout <= 8'b11111111; // 3061 : 255 - 0xff
      12'hBF6: dout <= 8'b11111111; // 3062 : 255 - 0xff
      12'hBF7: dout <= 8'b11111111; // 3063 : 255 - 0xff
      12'hBF8: dout <= 8'b11111111; // 3064 : 255 - 0xff -- Background 0x7f
      12'hBF9: dout <= 8'b11111111; // 3065 : 255 - 0xff
      12'hBFA: dout <= 8'b11111111; // 3066 : 255 - 0xff
      12'hBFB: dout <= 8'b11111111; // 3067 : 255 - 0xff
      12'hBFC: dout <= 8'b11111111; // 3068 : 255 - 0xff
      12'hBFD: dout <= 8'b11111111; // 3069 : 255 - 0xff
      12'hBFE: dout <= 8'b11111111; // 3070 : 255 - 0xff
      12'hBFF: dout <= 8'b11111111; // 3071 : 255 - 0xff
      12'hC00: dout <= 8'b11111111; // 3072 : 255 - 0xff -- Background 0x80
      12'hC01: dout <= 8'b11111111; // 3073 : 255 - 0xff
      12'hC02: dout <= 8'b11111111; // 3074 : 255 - 0xff
      12'hC03: dout <= 8'b11111111; // 3075 : 255 - 0xff
      12'hC04: dout <= 8'b11111111; // 3076 : 255 - 0xff
      12'hC05: dout <= 8'b11111111; // 3077 : 255 - 0xff
      12'hC06: dout <= 8'b11111111; // 3078 : 255 - 0xff
      12'hC07: dout <= 8'b11111111; // 3079 : 255 - 0xff
      12'hC08: dout <= 8'b11111111; // 3080 : 255 - 0xff -- Background 0x81
      12'hC09: dout <= 8'b11111111; // 3081 : 255 - 0xff
      12'hC0A: dout <= 8'b11111111; // 3082 : 255 - 0xff
      12'hC0B: dout <= 8'b11111111; // 3083 : 255 - 0xff
      12'hC0C: dout <= 8'b11111111; // 3084 : 255 - 0xff
      12'hC0D: dout <= 8'b11111111; // 3085 : 255 - 0xff
      12'hC0E: dout <= 8'b11111111; // 3086 : 255 - 0xff
      12'hC0F: dout <= 8'b11111111; // 3087 : 255 - 0xff
      12'hC10: dout <= 8'b11111111; // 3088 : 255 - 0xff -- Background 0x82
      12'hC11: dout <= 8'b11111111; // 3089 : 255 - 0xff
      12'hC12: dout <= 8'b11111111; // 3090 : 255 - 0xff
      12'hC13: dout <= 8'b11111111; // 3091 : 255 - 0xff
      12'hC14: dout <= 8'b11111111; // 3092 : 255 - 0xff
      12'hC15: dout <= 8'b11111111; // 3093 : 255 - 0xff
      12'hC16: dout <= 8'b11111111; // 3094 : 255 - 0xff
      12'hC17: dout <= 8'b11111111; // 3095 : 255 - 0xff
      12'hC18: dout <= 8'b11111111; // 3096 : 255 - 0xff -- Background 0x83
      12'hC19: dout <= 8'b11111111; // 3097 : 255 - 0xff
      12'hC1A: dout <= 8'b11111111; // 3098 : 255 - 0xff
      12'hC1B: dout <= 8'b11111111; // 3099 : 255 - 0xff
      12'hC1C: dout <= 8'b11111111; // 3100 : 255 - 0xff
      12'hC1D: dout <= 8'b11111111; // 3101 : 255 - 0xff
      12'hC1E: dout <= 8'b11111111; // 3102 : 255 - 0xff
      12'hC1F: dout <= 8'b11111111; // 3103 : 255 - 0xff
      12'hC20: dout <= 8'b11111111; // 3104 : 255 - 0xff -- Background 0x84
      12'hC21: dout <= 8'b11111111; // 3105 : 255 - 0xff
      12'hC22: dout <= 8'b11111111; // 3106 : 255 - 0xff
      12'hC23: dout <= 8'b11111111; // 3107 : 255 - 0xff
      12'hC24: dout <= 8'b11111111; // 3108 : 255 - 0xff
      12'hC25: dout <= 8'b11111111; // 3109 : 255 - 0xff
      12'hC26: dout <= 8'b11111111; // 3110 : 255 - 0xff
      12'hC27: dout <= 8'b11111111; // 3111 : 255 - 0xff
      12'hC28: dout <= 8'b11111111; // 3112 : 255 - 0xff -- Background 0x85
      12'hC29: dout <= 8'b11111111; // 3113 : 255 - 0xff
      12'hC2A: dout <= 8'b11111111; // 3114 : 255 - 0xff
      12'hC2B: dout <= 8'b11111111; // 3115 : 255 - 0xff
      12'hC2C: dout <= 8'b11111111; // 3116 : 255 - 0xff
      12'hC2D: dout <= 8'b11111111; // 3117 : 255 - 0xff
      12'hC2E: dout <= 8'b11111111; // 3118 : 255 - 0xff
      12'hC2F: dout <= 8'b11111111; // 3119 : 255 - 0xff
      12'hC30: dout <= 8'b11111111; // 3120 : 255 - 0xff -- Background 0x86
      12'hC31: dout <= 8'b11111111; // 3121 : 255 - 0xff
      12'hC32: dout <= 8'b11111111; // 3122 : 255 - 0xff
      12'hC33: dout <= 8'b11111111; // 3123 : 255 - 0xff
      12'hC34: dout <= 8'b11111111; // 3124 : 255 - 0xff
      12'hC35: dout <= 8'b11111111; // 3125 : 255 - 0xff
      12'hC36: dout <= 8'b11111111; // 3126 : 255 - 0xff
      12'hC37: dout <= 8'b11111111; // 3127 : 255 - 0xff
      12'hC38: dout <= 8'b11111111; // 3128 : 255 - 0xff -- Background 0x87
      12'hC39: dout <= 8'b11111111; // 3129 : 255 - 0xff
      12'hC3A: dout <= 8'b11111111; // 3130 : 255 - 0xff
      12'hC3B: dout <= 8'b11111111; // 3131 : 255 - 0xff
      12'hC3C: dout <= 8'b11111111; // 3132 : 255 - 0xff
      12'hC3D: dout <= 8'b11111111; // 3133 : 255 - 0xff
      12'hC3E: dout <= 8'b11111111; // 3134 : 255 - 0xff
      12'hC3F: dout <= 8'b11111111; // 3135 : 255 - 0xff
      12'hC40: dout <= 8'b11111111; // 3136 : 255 - 0xff -- Background 0x88
      12'hC41: dout <= 8'b11111111; // 3137 : 255 - 0xff
      12'hC42: dout <= 8'b11111111; // 3138 : 255 - 0xff
      12'hC43: dout <= 8'b11111111; // 3139 : 255 - 0xff
      12'hC44: dout <= 8'b11111111; // 3140 : 255 - 0xff
      12'hC45: dout <= 8'b11111111; // 3141 : 255 - 0xff
      12'hC46: dout <= 8'b11111111; // 3142 : 255 - 0xff
      12'hC47: dout <= 8'b11111111; // 3143 : 255 - 0xff
      12'hC48: dout <= 8'b11111111; // 3144 : 255 - 0xff -- Background 0x89
      12'hC49: dout <= 8'b11111111; // 3145 : 255 - 0xff
      12'hC4A: dout <= 8'b11111111; // 3146 : 255 - 0xff
      12'hC4B: dout <= 8'b11111111; // 3147 : 255 - 0xff
      12'hC4C: dout <= 8'b11111111; // 3148 : 255 - 0xff
      12'hC4D: dout <= 8'b11111111; // 3149 : 255 - 0xff
      12'hC4E: dout <= 8'b11111111; // 3150 : 255 - 0xff
      12'hC4F: dout <= 8'b11111111; // 3151 : 255 - 0xff
      12'hC50: dout <= 8'b11111111; // 3152 : 255 - 0xff -- Background 0x8a
      12'hC51: dout <= 8'b11111111; // 3153 : 255 - 0xff
      12'hC52: dout <= 8'b11111111; // 3154 : 255 - 0xff
      12'hC53: dout <= 8'b11111111; // 3155 : 255 - 0xff
      12'hC54: dout <= 8'b11111111; // 3156 : 255 - 0xff
      12'hC55: dout <= 8'b11111111; // 3157 : 255 - 0xff
      12'hC56: dout <= 8'b11111111; // 3158 : 255 - 0xff
      12'hC57: dout <= 8'b11111111; // 3159 : 255 - 0xff
      12'hC58: dout <= 8'b11111111; // 3160 : 255 - 0xff -- Background 0x8b
      12'hC59: dout <= 8'b11111111; // 3161 : 255 - 0xff
      12'hC5A: dout <= 8'b11111111; // 3162 : 255 - 0xff
      12'hC5B: dout <= 8'b11111111; // 3163 : 255 - 0xff
      12'hC5C: dout <= 8'b11111111; // 3164 : 255 - 0xff
      12'hC5D: dout <= 8'b11111111; // 3165 : 255 - 0xff
      12'hC5E: dout <= 8'b11111111; // 3166 : 255 - 0xff
      12'hC5F: dout <= 8'b11111111; // 3167 : 255 - 0xff
      12'hC60: dout <= 8'b11111111; // 3168 : 255 - 0xff -- Background 0x8c
      12'hC61: dout <= 8'b11111111; // 3169 : 255 - 0xff
      12'hC62: dout <= 8'b11111111; // 3170 : 255 - 0xff
      12'hC63: dout <= 8'b11111111; // 3171 : 255 - 0xff
      12'hC64: dout <= 8'b11111111; // 3172 : 255 - 0xff
      12'hC65: dout <= 8'b11111111; // 3173 : 255 - 0xff
      12'hC66: dout <= 8'b11111111; // 3174 : 255 - 0xff
      12'hC67: dout <= 8'b11111111; // 3175 : 255 - 0xff
      12'hC68: dout <= 8'b11111111; // 3176 : 255 - 0xff -- Background 0x8d
      12'hC69: dout <= 8'b11111111; // 3177 : 255 - 0xff
      12'hC6A: dout <= 8'b11111111; // 3178 : 255 - 0xff
      12'hC6B: dout <= 8'b11111111; // 3179 : 255 - 0xff
      12'hC6C: dout <= 8'b11111111; // 3180 : 255 - 0xff
      12'hC6D: dout <= 8'b11111111; // 3181 : 255 - 0xff
      12'hC6E: dout <= 8'b11111111; // 3182 : 255 - 0xff
      12'hC6F: dout <= 8'b11111111; // 3183 : 255 - 0xff
      12'hC70: dout <= 8'b11111111; // 3184 : 255 - 0xff -- Background 0x8e
      12'hC71: dout <= 8'b11111111; // 3185 : 255 - 0xff
      12'hC72: dout <= 8'b11111111; // 3186 : 255 - 0xff
      12'hC73: dout <= 8'b11111111; // 3187 : 255 - 0xff
      12'hC74: dout <= 8'b11111111; // 3188 : 255 - 0xff
      12'hC75: dout <= 8'b11111111; // 3189 : 255 - 0xff
      12'hC76: dout <= 8'b11111111; // 3190 : 255 - 0xff
      12'hC77: dout <= 8'b11111111; // 3191 : 255 - 0xff
      12'hC78: dout <= 8'b11111111; // 3192 : 255 - 0xff -- Background 0x8f
      12'hC79: dout <= 8'b11111111; // 3193 : 255 - 0xff
      12'hC7A: dout <= 8'b11111111; // 3194 : 255 - 0xff
      12'hC7B: dout <= 8'b11111111; // 3195 : 255 - 0xff
      12'hC7C: dout <= 8'b11111111; // 3196 : 255 - 0xff
      12'hC7D: dout <= 8'b11111111; // 3197 : 255 - 0xff
      12'hC7E: dout <= 8'b11111111; // 3198 : 255 - 0xff
      12'hC7F: dout <= 8'b11111111; // 3199 : 255 - 0xff
      12'hC80: dout <= 8'b00000000; // 3200 :   0 - 0x0 -- Background 0x90
      12'hC81: dout <= 8'b00000000; // 3201 :   0 - 0x0
      12'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      12'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      12'hC84: dout <= 8'b00000000; // 3204 :   0 - 0x0
      12'hC85: dout <= 8'b00000001; // 3205 :   1 - 0x1
      12'hC86: dout <= 8'b00011110; // 3206 :  30 - 0x1e
      12'hC87: dout <= 8'b00111011; // 3207 :  59 - 0x3b
      12'hC88: dout <= 8'b00000000; // 3208 :   0 - 0x0 -- Background 0x91
      12'hC89: dout <= 8'b00000000; // 3209 :   0 - 0x0
      12'hC8A: dout <= 8'b00001100; // 3210 :  12 - 0xc
      12'hC8B: dout <= 8'b00111100; // 3211 :  60 - 0x3c
      12'hC8C: dout <= 8'b11010000; // 3212 : 208 - 0xd0
      12'hC8D: dout <= 8'b00010000; // 3213 :  16 - 0x10
      12'hC8E: dout <= 8'b00100000; // 3214 :  32 - 0x20
      12'hC8F: dout <= 8'b01000000; // 3215 :  64 - 0x40
      12'hC90: dout <= 8'b00111110; // 3216 :  62 - 0x3e -- Background 0x92
      12'hC91: dout <= 8'b00101101; // 3217 :  45 - 0x2d
      12'hC92: dout <= 8'b00110101; // 3218 :  53 - 0x35
      12'hC93: dout <= 8'b00011101; // 3219 :  29 - 0x1d
      12'hC94: dout <= 8'b00000001; // 3220 :   1 - 0x1
      12'hC95: dout <= 8'b00000000; // 3221 :   0 - 0x0
      12'hC96: dout <= 8'b00000000; // 3222 :   0 - 0x0
      12'hC97: dout <= 8'b00000000; // 3223 :   0 - 0x0
      12'hC98: dout <= 8'b10110000; // 3224 : 176 - 0xb0 -- Background 0x93
      12'hC99: dout <= 8'b10111000; // 3225 : 184 - 0xb8
      12'hC9A: dout <= 8'b11111000; // 3226 : 248 - 0xf8
      12'hC9B: dout <= 8'b01111000; // 3227 : 120 - 0x78
      12'hC9C: dout <= 8'b10011000; // 3228 : 152 - 0x98
      12'hC9D: dout <= 8'b11110000; // 3229 : 240 - 0xf0
      12'hC9E: dout <= 8'b00000000; // 3230 :   0 - 0x0
      12'hC9F: dout <= 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout <= 8'b00000000; // 3232 :   0 - 0x0 -- Background 0x94
      12'hCA1: dout <= 8'b00000000; // 3233 :   0 - 0x0
      12'hCA2: dout <= 8'b00000111; // 3234 :   7 - 0x7
      12'hCA3: dout <= 8'b00000011; // 3235 :   3 - 0x3
      12'hCA4: dout <= 8'b00001101; // 3236 :  13 - 0xd
      12'hCA5: dout <= 8'b00011110; // 3237 :  30 - 0x1e
      12'hCA6: dout <= 8'b00010111; // 3238 :  23 - 0x17
      12'hCA7: dout <= 8'b00011101; // 3239 :  29 - 0x1d
      12'hCA8: dout <= 8'b00000000; // 3240 :   0 - 0x0 -- Background 0x95
      12'hCA9: dout <= 8'b10000000; // 3241 : 128 - 0x80
      12'hCAA: dout <= 8'b01110000; // 3242 : 112 - 0x70
      12'hCAB: dout <= 8'b11100000; // 3243 : 224 - 0xe0
      12'hCAC: dout <= 8'b11011000; // 3244 : 216 - 0xd8
      12'hCAD: dout <= 8'b10111100; // 3245 : 188 - 0xbc
      12'hCAE: dout <= 8'b01110100; // 3246 : 116 - 0x74
      12'hCAF: dout <= 8'b11011100; // 3247 : 220 - 0xdc
      12'hCB0: dout <= 8'b00011111; // 3248 :  31 - 0x1f -- Background 0x96
      12'hCB1: dout <= 8'b00001011; // 3249 :  11 - 0xb
      12'hCB2: dout <= 8'b00001111; // 3250 :  15 - 0xf
      12'hCB3: dout <= 8'b00000101; // 3251 :   5 - 0x5
      12'hCB4: dout <= 8'b00000011; // 3252 :   3 - 0x3
      12'hCB5: dout <= 8'b00000001; // 3253 :   1 - 0x1
      12'hCB6: dout <= 8'b00000000; // 3254 :   0 - 0x0
      12'hCB7: dout <= 8'b00000000; // 3255 :   0 - 0x0
      12'hCB8: dout <= 8'b11111100; // 3256 : 252 - 0xfc -- Background 0x97
      12'hCB9: dout <= 8'b01101000; // 3257 : 104 - 0x68
      12'hCBA: dout <= 8'b11111000; // 3258 : 248 - 0xf8
      12'hCBB: dout <= 8'b10110000; // 3259 : 176 - 0xb0
      12'hCBC: dout <= 8'b11100000; // 3260 : 224 - 0xe0
      12'hCBD: dout <= 8'b10000000; // 3261 : 128 - 0x80
      12'hCBE: dout <= 8'b00000000; // 3262 :   0 - 0x0
      12'hCBF: dout <= 8'b00000000; // 3263 :   0 - 0x0
      12'hCC0: dout <= 8'b00000000; // 3264 :   0 - 0x0 -- Background 0x98
      12'hCC1: dout <= 8'b00000000; // 3265 :   0 - 0x0
      12'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      12'hCC3: dout <= 8'b00000001; // 3267 :   1 - 0x1
      12'hCC4: dout <= 8'b00000001; // 3268 :   1 - 0x1
      12'hCC5: dout <= 8'b00001011; // 3269 :  11 - 0xb
      12'hCC6: dout <= 8'b00011100; // 3270 :  28 - 0x1c
      12'hCC7: dout <= 8'b00111111; // 3271 :  63 - 0x3f
      12'hCC8: dout <= 8'b00000000; // 3272 :   0 - 0x0 -- Background 0x99
      12'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      12'hCCA: dout <= 8'b00110000; // 3274 :  48 - 0x30
      12'hCCB: dout <= 8'b01111000; // 3275 : 120 - 0x78
      12'hCCC: dout <= 8'b10000000; // 3276 : 128 - 0x80
      12'hCCD: dout <= 8'b11110000; // 3277 : 240 - 0xf0
      12'hCCE: dout <= 8'b11111000; // 3278 : 248 - 0xf8
      12'hCCF: dout <= 8'b11111100; // 3279 : 252 - 0xfc
      12'hCD0: dout <= 8'b00111111; // 3280 :  63 - 0x3f -- Background 0x9a
      12'hCD1: dout <= 8'b00111111; // 3281 :  63 - 0x3f
      12'hCD2: dout <= 8'b00111111; // 3282 :  63 - 0x3f
      12'hCD3: dout <= 8'b00011111; // 3283 :  31 - 0x1f
      12'hCD4: dout <= 8'b00011111; // 3284 :  31 - 0x1f
      12'hCD5: dout <= 8'b00000111; // 3285 :   7 - 0x7
      12'hCD6: dout <= 8'b00000000; // 3286 :   0 - 0x0
      12'hCD7: dout <= 8'b00000000; // 3287 :   0 - 0x0
      12'hCD8: dout <= 8'b11111100; // 3288 : 252 - 0xfc -- Background 0x9b
      12'hCD9: dout <= 8'b11101100; // 3289 : 236 - 0xec
      12'hCDA: dout <= 8'b11101100; // 3290 : 236 - 0xec
      12'hCDB: dout <= 8'b11011000; // 3291 : 216 - 0xd8
      12'hCDC: dout <= 8'b11111000; // 3292 : 248 - 0xf8
      12'hCDD: dout <= 8'b11100000; // 3293 : 224 - 0xe0
      12'hCDE: dout <= 8'b00000000; // 3294 :   0 - 0x0
      12'hCDF: dout <= 8'b00000000; // 3295 :   0 - 0x0
      12'hCE0: dout <= 8'b00000000; // 3296 :   0 - 0x0 -- Background 0x9c
      12'hCE1: dout <= 8'b00000000; // 3297 :   0 - 0x0
      12'hCE2: dout <= 8'b00000001; // 3298 :   1 - 0x1
      12'hCE3: dout <= 8'b00011101; // 3299 :  29 - 0x1d
      12'hCE4: dout <= 8'b00111110; // 3300 :  62 - 0x3e
      12'hCE5: dout <= 8'b00111111; // 3301 :  63 - 0x3f
      12'hCE6: dout <= 8'b00111111; // 3302 :  63 - 0x3f
      12'hCE7: dout <= 8'b00111111; // 3303 :  63 - 0x3f
      12'hCE8: dout <= 8'b00000000; // 3304 :   0 - 0x0 -- Background 0x9d
      12'hCE9: dout <= 8'b10000000; // 3305 : 128 - 0x80
      12'hCEA: dout <= 8'b00000000; // 3306 :   0 - 0x0
      12'hCEB: dout <= 8'b01110000; // 3307 : 112 - 0x70
      12'hCEC: dout <= 8'b11111000; // 3308 : 248 - 0xf8
      12'hCED: dout <= 8'b11111100; // 3309 : 252 - 0xfc
      12'hCEE: dout <= 8'b11111100; // 3310 : 252 - 0xfc
      12'hCEF: dout <= 8'b11111100; // 3311 : 252 - 0xfc
      12'hCF0: dout <= 8'b00111111; // 3312 :  63 - 0x3f -- Background 0x9e
      12'hCF1: dout <= 8'b00111111; // 3313 :  63 - 0x3f
      12'hCF2: dout <= 8'b00011111; // 3314 :  31 - 0x1f
      12'hCF3: dout <= 8'b00011111; // 3315 :  31 - 0x1f
      12'hCF4: dout <= 8'b00001111; // 3316 :  15 - 0xf
      12'hCF5: dout <= 8'b00000110; // 3317 :   6 - 0x6
      12'hCF6: dout <= 8'b00000000; // 3318 :   0 - 0x0
      12'hCF7: dout <= 8'b00000000; // 3319 :   0 - 0x0
      12'hCF8: dout <= 8'b11101100; // 3320 : 236 - 0xec -- Background 0x9f
      12'hCF9: dout <= 8'b11101100; // 3321 : 236 - 0xec
      12'hCFA: dout <= 8'b11011000; // 3322 : 216 - 0xd8
      12'hCFB: dout <= 8'b11111000; // 3323 : 248 - 0xf8
      12'hCFC: dout <= 8'b11110000; // 3324 : 240 - 0xf0
      12'hCFD: dout <= 8'b11100000; // 3325 : 224 - 0xe0
      12'hCFE: dout <= 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout <= 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout <= 8'b00000000; // 3328 :   0 - 0x0 -- Background 0xa0
      12'hD01: dout <= 8'b00000100; // 3329 :   4 - 0x4
      12'hD02: dout <= 8'b00000011; // 3330 :   3 - 0x3
      12'hD03: dout <= 8'b00000000; // 3331 :   0 - 0x0
      12'hD04: dout <= 8'b00000001; // 3332 :   1 - 0x1
      12'hD05: dout <= 8'b00000111; // 3333 :   7 - 0x7
      12'hD06: dout <= 8'b00001111; // 3334 :  15 - 0xf
      12'hD07: dout <= 8'b00001100; // 3335 :  12 - 0xc
      12'hD08: dout <= 8'b00000000; // 3336 :   0 - 0x0 -- Background 0xa1
      12'hD09: dout <= 8'b00000000; // 3337 :   0 - 0x0
      12'hD0A: dout <= 8'b11100000; // 3338 : 224 - 0xe0
      12'hD0B: dout <= 8'b10000000; // 3339 : 128 - 0x80
      12'hD0C: dout <= 8'b01000000; // 3340 :  64 - 0x40
      12'hD0D: dout <= 8'b11110000; // 3341 : 240 - 0xf0
      12'hD0E: dout <= 8'b10011000; // 3342 : 152 - 0x98
      12'hD0F: dout <= 8'b11111000; // 3343 : 248 - 0xf8
      12'hD10: dout <= 8'b00011111; // 3344 :  31 - 0x1f -- Background 0xa2
      12'hD11: dout <= 8'b00010011; // 3345 :  19 - 0x13
      12'hD12: dout <= 8'b00011111; // 3346 :  31 - 0x1f
      12'hD13: dout <= 8'b00001111; // 3347 :  15 - 0xf
      12'hD14: dout <= 8'b00001001; // 3348 :   9 - 0x9
      12'hD15: dout <= 8'b00000111; // 3349 :   7 - 0x7
      12'hD16: dout <= 8'b00000001; // 3350 :   1 - 0x1
      12'hD17: dout <= 8'b00000000; // 3351 :   0 - 0x0
      12'hD18: dout <= 8'b11100100; // 3352 : 228 - 0xe4 -- Background 0xa3
      12'hD19: dout <= 8'b00111100; // 3353 :  60 - 0x3c
      12'hD1A: dout <= 8'b11100100; // 3354 : 228 - 0xe4
      12'hD1B: dout <= 8'b00111000; // 3355 :  56 - 0x38
      12'hD1C: dout <= 8'b11111000; // 3356 : 248 - 0xf8
      12'hD1D: dout <= 8'b11110000; // 3357 : 240 - 0xf0
      12'hD1E: dout <= 8'b11000000; // 3358 : 192 - 0xc0
      12'hD1F: dout <= 8'b00000000; // 3359 :   0 - 0x0
      12'hD20: dout <= 8'b00000000; // 3360 :   0 - 0x0 -- Background 0xa4
      12'hD21: dout <= 8'b00000000; // 3361 :   0 - 0x0
      12'hD22: dout <= 8'b00000000; // 3362 :   0 - 0x0
      12'hD23: dout <= 8'b00000000; // 3363 :   0 - 0x0
      12'hD24: dout <= 8'b00010001; // 3364 :  17 - 0x11
      12'hD25: dout <= 8'b00010011; // 3365 :  19 - 0x13
      12'hD26: dout <= 8'b00011111; // 3366 :  31 - 0x1f
      12'hD27: dout <= 8'b00011111; // 3367 :  31 - 0x1f
      12'hD28: dout <= 8'b00000000; // 3368 :   0 - 0x0 -- Background 0xa5
      12'hD29: dout <= 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout <= 8'b00000000; // 3370 :   0 - 0x0
      12'hD2B: dout <= 8'b10000000; // 3371 : 128 - 0x80
      12'hD2C: dout <= 8'b11000100; // 3372 : 196 - 0xc4
      12'hD2D: dout <= 8'b11100100; // 3373 : 228 - 0xe4
      12'hD2E: dout <= 8'b11111100; // 3374 : 252 - 0xfc
      12'hD2F: dout <= 8'b11111100; // 3375 : 252 - 0xfc
      12'hD30: dout <= 8'b00011111; // 3376 :  31 - 0x1f -- Background 0xa6
      12'hD31: dout <= 8'b00001110; // 3377 :  14 - 0xe
      12'hD32: dout <= 8'b00000110; // 3378 :   6 - 0x6
      12'hD33: dout <= 8'b00000010; // 3379 :   2 - 0x2
      12'hD34: dout <= 8'b00000000; // 3380 :   0 - 0x0
      12'hD35: dout <= 8'b00000000; // 3381 :   0 - 0x0
      12'hD36: dout <= 8'b00000000; // 3382 :   0 - 0x0
      12'hD37: dout <= 8'b00000000; // 3383 :   0 - 0x0
      12'hD38: dout <= 8'b11111100; // 3384 : 252 - 0xfc -- Background 0xa7
      12'hD39: dout <= 8'b10111000; // 3385 : 184 - 0xb8
      12'hD3A: dout <= 8'b10110000; // 3386 : 176 - 0xb0
      12'hD3B: dout <= 8'b10100000; // 3387 : 160 - 0xa0
      12'hD3C: dout <= 8'b10000000; // 3388 : 128 - 0x80
      12'hD3D: dout <= 8'b00000000; // 3389 :   0 - 0x0
      12'hD3E: dout <= 8'b00000000; // 3390 :   0 - 0x0
      12'hD3F: dout <= 8'b00000000; // 3391 :   0 - 0x0
      12'hD40: dout <= 8'b00000000; // 3392 :   0 - 0x0 -- Background 0xa8
      12'hD41: dout <= 8'b00000000; // 3393 :   0 - 0x0
      12'hD42: dout <= 8'b00000000; // 3394 :   0 - 0x0
      12'hD43: dout <= 8'b00000001; // 3395 :   1 - 0x1
      12'hD44: dout <= 8'b00000011; // 3396 :   3 - 0x3
      12'hD45: dout <= 8'b00000110; // 3397 :   6 - 0x6
      12'hD46: dout <= 8'b00000110; // 3398 :   6 - 0x6
      12'hD47: dout <= 8'b00001111; // 3399 :  15 - 0xf
      12'hD48: dout <= 8'b00000000; // 3400 :   0 - 0x0 -- Background 0xa9
      12'hD49: dout <= 8'b00011000; // 3401 :  24 - 0x18
      12'hD4A: dout <= 8'b11110100; // 3402 : 244 - 0xf4
      12'hD4B: dout <= 8'b11111000; // 3403 : 248 - 0xf8
      12'hD4C: dout <= 8'b00111000; // 3404 :  56 - 0x38
      12'hD4D: dout <= 8'b01111100; // 3405 : 124 - 0x7c
      12'hD4E: dout <= 8'b11111100; // 3406 : 252 - 0xfc
      12'hD4F: dout <= 8'b11111100; // 3407 : 252 - 0xfc
      12'hD50: dout <= 8'b00001111; // 3408 :  15 - 0xf -- Background 0xaa
      12'hD51: dout <= 8'b00011111; // 3409 :  31 - 0x1f
      12'hD52: dout <= 8'b00110000; // 3410 :  48 - 0x30
      12'hD53: dout <= 8'b00111000; // 3411 :  56 - 0x38
      12'hD54: dout <= 8'b00011101; // 3412 :  29 - 0x1d
      12'hD55: dout <= 8'b00000011; // 3413 :   3 - 0x3
      12'hD56: dout <= 8'b00000011; // 3414 :   3 - 0x3
      12'hD57: dout <= 8'b00000000; // 3415 :   0 - 0x0
      12'hD58: dout <= 8'b11111100; // 3416 : 252 - 0xfc -- Background 0xab
      12'hD59: dout <= 8'b11111100; // 3417 : 252 - 0xfc
      12'hD5A: dout <= 8'b01111100; // 3418 : 124 - 0x7c
      12'hD5B: dout <= 8'b10001110; // 3419 : 142 - 0x8e
      12'hD5C: dout <= 8'b10000110; // 3420 : 134 - 0x86
      12'hD5D: dout <= 8'b10011100; // 3421 : 156 - 0x9c
      12'hD5E: dout <= 8'b01111000; // 3422 : 120 - 0x78
      12'hD5F: dout <= 8'b00000000; // 3423 :   0 - 0x0
      12'hD60: dout <= 8'b00000000; // 3424 :   0 - 0x0 -- Background 0xac
      12'hD61: dout <= 8'b00000001; // 3425 :   1 - 0x1
      12'hD62: dout <= 8'b00000110; // 3426 :   6 - 0x6
      12'hD63: dout <= 8'b00000111; // 3427 :   7 - 0x7
      12'hD64: dout <= 8'b00000111; // 3428 :   7 - 0x7
      12'hD65: dout <= 8'b00000111; // 3429 :   7 - 0x7
      12'hD66: dout <= 8'b00000001; // 3430 :   1 - 0x1
      12'hD67: dout <= 8'b00000011; // 3431 :   3 - 0x3
      12'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0 -- Background 0xad
      12'hD69: dout <= 8'b11000000; // 3433 : 192 - 0xc0
      12'hD6A: dout <= 8'b00110000; // 3434 :  48 - 0x30
      12'hD6B: dout <= 8'b11110000; // 3435 : 240 - 0xf0
      12'hD6C: dout <= 8'b11110000; // 3436 : 240 - 0xf0
      12'hD6D: dout <= 8'b11110000; // 3437 : 240 - 0xf0
      12'hD6E: dout <= 8'b01000000; // 3438 :  64 - 0x40
      12'hD6F: dout <= 8'b01000000; // 3439 :  64 - 0x40
      12'hD70: dout <= 8'b00000001; // 3440 :   1 - 0x1 -- Background 0xae
      12'hD71: dout <= 8'b00000000; // 3441 :   0 - 0x0
      12'hD72: dout <= 8'b00000001; // 3442 :   1 - 0x1
      12'hD73: dout <= 8'b00000011; // 3443 :   3 - 0x3
      12'hD74: dout <= 8'b00000001; // 3444 :   1 - 0x1
      12'hD75: dout <= 8'b00000000; // 3445 :   0 - 0x0
      12'hD76: dout <= 8'b00000000; // 3446 :   0 - 0x0
      12'hD77: dout <= 8'b00000000; // 3447 :   0 - 0x0
      12'hD78: dout <= 8'b01000000; // 3448 :  64 - 0x40 -- Background 0xaf
      12'hD79: dout <= 8'b01000000; // 3449 :  64 - 0x40
      12'hD7A: dout <= 8'b01000000; // 3450 :  64 - 0x40
      12'hD7B: dout <= 8'b01000000; // 3451 :  64 - 0x40
      12'hD7C: dout <= 8'b01000000; // 3452 :  64 - 0x40
      12'hD7D: dout <= 8'b10000000; // 3453 : 128 - 0x80
      12'hD7E: dout <= 8'b00000000; // 3454 :   0 - 0x0
      12'hD7F: dout <= 8'b00000000; // 3455 :   0 - 0x0
      12'hD80: dout <= 8'b01111110; // 3456 : 126 - 0x7e -- Background 0xb0
      12'hD81: dout <= 8'b01100011; // 3457 :  99 - 0x63
      12'hD82: dout <= 8'b01100011; // 3458 :  99 - 0x63
      12'hD83: dout <= 8'b01100011; // 3459 :  99 - 0x63
      12'hD84: dout <= 8'b01111110; // 3460 : 126 - 0x7e
      12'hD85: dout <= 8'b01100000; // 3461 :  96 - 0x60
      12'hD86: dout <= 8'b01100000; // 3462 :  96 - 0x60
      12'hD87: dout <= 8'b00000000; // 3463 :   0 - 0x0
      12'hD88: dout <= 8'b01100000; // 3464 :  96 - 0x60 -- Background 0xb1
      12'hD89: dout <= 8'b01100000; // 3465 :  96 - 0x60
      12'hD8A: dout <= 8'b01100000; // 3466 :  96 - 0x60
      12'hD8B: dout <= 8'b01100000; // 3467 :  96 - 0x60
      12'hD8C: dout <= 8'b01100000; // 3468 :  96 - 0x60
      12'hD8D: dout <= 8'b01100000; // 3469 :  96 - 0x60
      12'hD8E: dout <= 8'b01111111; // 3470 : 127 - 0x7f
      12'hD8F: dout <= 8'b00000000; // 3471 :   0 - 0x0
      12'hD90: dout <= 8'b00011100; // 3472 :  28 - 0x1c -- Background 0xb2
      12'hD91: dout <= 8'b00110110; // 3473 :  54 - 0x36
      12'hD92: dout <= 8'b01100011; // 3474 :  99 - 0x63
      12'hD93: dout <= 8'b01100011; // 3475 :  99 - 0x63
      12'hD94: dout <= 8'b01111111; // 3476 : 127 - 0x7f
      12'hD95: dout <= 8'b01100011; // 3477 :  99 - 0x63
      12'hD96: dout <= 8'b01100011; // 3478 :  99 - 0x63
      12'hD97: dout <= 8'b00000000; // 3479 :   0 - 0x0
      12'hD98: dout <= 8'b00110011; // 3480 :  51 - 0x33 -- Background 0xb3
      12'hD99: dout <= 8'b00110011; // 3481 :  51 - 0x33
      12'hD9A: dout <= 8'b00110011; // 3482 :  51 - 0x33
      12'hD9B: dout <= 8'b00011110; // 3483 :  30 - 0x1e
      12'hD9C: dout <= 8'b00001100; // 3484 :  12 - 0xc
      12'hD9D: dout <= 8'b00001100; // 3485 :  12 - 0xc
      12'hD9E: dout <= 8'b00001100; // 3486 :  12 - 0xc
      12'hD9F: dout <= 8'b00000000; // 3487 :   0 - 0x0
      12'hDA0: dout <= 8'b01111111; // 3488 : 127 - 0x7f -- Background 0xb4
      12'hDA1: dout <= 8'b01100000; // 3489 :  96 - 0x60
      12'hDA2: dout <= 8'b01100000; // 3490 :  96 - 0x60
      12'hDA3: dout <= 8'b01111110; // 3491 : 126 - 0x7e
      12'hDA4: dout <= 8'b01100000; // 3492 :  96 - 0x60
      12'hDA5: dout <= 8'b01100000; // 3493 :  96 - 0x60
      12'hDA6: dout <= 8'b01111111; // 3494 : 127 - 0x7f
      12'hDA7: dout <= 8'b00000000; // 3495 :   0 - 0x0
      12'hDA8: dout <= 8'b01111110; // 3496 : 126 - 0x7e -- Background 0xb5
      12'hDA9: dout <= 8'b01100011; // 3497 :  99 - 0x63
      12'hDAA: dout <= 8'b01100011; // 3498 :  99 - 0x63
      12'hDAB: dout <= 8'b01100111; // 3499 : 103 - 0x67
      12'hDAC: dout <= 8'b01111100; // 3500 : 124 - 0x7c
      12'hDAD: dout <= 8'b01101110; // 3501 : 110 - 0x6e
      12'hDAE: dout <= 8'b01100111; // 3502 : 103 - 0x67
      12'hDAF: dout <= 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout <= 8'b00111110; // 3504 :  62 - 0x3e -- Background 0xb6
      12'hDB1: dout <= 8'b01100011; // 3505 :  99 - 0x63
      12'hDB2: dout <= 8'b01100011; // 3506 :  99 - 0x63
      12'hDB3: dout <= 8'b01100011; // 3507 :  99 - 0x63
      12'hDB4: dout <= 8'b01100011; // 3508 :  99 - 0x63
      12'hDB5: dout <= 8'b01100011; // 3509 :  99 - 0x63
      12'hDB6: dout <= 8'b00111110; // 3510 :  62 - 0x3e
      12'hDB7: dout <= 8'b00000000; // 3511 :   0 - 0x0
      12'hDB8: dout <= 8'b01100011; // 3512 :  99 - 0x63 -- Background 0xb7
      12'hDB9: dout <= 8'b01110011; // 3513 : 115 - 0x73
      12'hDBA: dout <= 8'b01111011; // 3514 : 123 - 0x7b
      12'hDBB: dout <= 8'b01111111; // 3515 : 127 - 0x7f
      12'hDBC: dout <= 8'b01101111; // 3516 : 111 - 0x6f
      12'hDBD: dout <= 8'b01100111; // 3517 : 103 - 0x67
      12'hDBE: dout <= 8'b01100011; // 3518 :  99 - 0x63
      12'hDBF: dout <= 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout <= 8'b00111111; // 3520 :  63 - 0x3f -- Background 0xb8
      12'hDC1: dout <= 8'b00001100; // 3521 :  12 - 0xc
      12'hDC2: dout <= 8'b00001100; // 3522 :  12 - 0xc
      12'hDC3: dout <= 8'b00001100; // 3523 :  12 - 0xc
      12'hDC4: dout <= 8'b00001100; // 3524 :  12 - 0xc
      12'hDC5: dout <= 8'b00001100; // 3525 :  12 - 0xc
      12'hDC6: dout <= 8'b00001100; // 3526 :  12 - 0xc
      12'hDC7: dout <= 8'b00000000; // 3527 :   0 - 0x0
      12'hDC8: dout <= 8'b01100011; // 3528 :  99 - 0x63 -- Background 0xb9
      12'hDC9: dout <= 8'b01100011; // 3529 :  99 - 0x63
      12'hDCA: dout <= 8'b01101011; // 3530 : 107 - 0x6b
      12'hDCB: dout <= 8'b01111111; // 3531 : 127 - 0x7f
      12'hDCC: dout <= 8'b01111111; // 3532 : 127 - 0x7f
      12'hDCD: dout <= 8'b01110111; // 3533 : 119 - 0x77
      12'hDCE: dout <= 8'b01100011; // 3534 :  99 - 0x63
      12'hDCF: dout <= 8'b00000000; // 3535 :   0 - 0x0
      12'hDD0: dout <= 8'b01111100; // 3536 : 124 - 0x7c -- Background 0xba
      12'hDD1: dout <= 8'b01100110; // 3537 : 102 - 0x66
      12'hDD2: dout <= 8'b01100011; // 3538 :  99 - 0x63
      12'hDD3: dout <= 8'b01100011; // 3539 :  99 - 0x63
      12'hDD4: dout <= 8'b01100011; // 3540 :  99 - 0x63
      12'hDD5: dout <= 8'b01100110; // 3541 : 102 - 0x66
      12'hDD6: dout <= 8'b01111100; // 3542 : 124 - 0x7c
      12'hDD7: dout <= 8'b00000000; // 3543 :   0 - 0x0
      12'hDD8: dout <= 8'b00011100; // 3544 :  28 - 0x1c -- Background 0xbb
      12'hDD9: dout <= 8'b00011100; // 3545 :  28 - 0x1c
      12'hDDA: dout <= 8'b00011100; // 3546 :  28 - 0x1c
      12'hDDB: dout <= 8'b00011000; // 3547 :  24 - 0x18
      12'hDDC: dout <= 8'b00011000; // 3548 :  24 - 0x18
      12'hDDD: dout <= 8'b00000000; // 3549 :   0 - 0x0
      12'hDDE: dout <= 8'b00011000; // 3550 :  24 - 0x18
      12'hDDF: dout <= 8'b00000000; // 3551 :   0 - 0x0
      12'hDE0: dout <= 8'b00011111; // 3552 :  31 - 0x1f -- Background 0xbc
      12'hDE1: dout <= 8'b00110000; // 3553 :  48 - 0x30
      12'hDE2: dout <= 8'b01100000; // 3554 :  96 - 0x60
      12'hDE3: dout <= 8'b01100111; // 3555 : 103 - 0x67
      12'hDE4: dout <= 8'b01100011; // 3556 :  99 - 0x63
      12'hDE5: dout <= 8'b00110011; // 3557 :  51 - 0x33
      12'hDE6: dout <= 8'b00011111; // 3558 :  31 - 0x1f
      12'hDE7: dout <= 8'b00000000; // 3559 :   0 - 0x0
      12'hDE8: dout <= 8'b01100011; // 3560 :  99 - 0x63 -- Background 0xbd
      12'hDE9: dout <= 8'b01110111; // 3561 : 119 - 0x77
      12'hDEA: dout <= 8'b01111111; // 3562 : 127 - 0x7f
      12'hDEB: dout <= 8'b01111111; // 3563 : 127 - 0x7f
      12'hDEC: dout <= 8'b01101011; // 3564 : 107 - 0x6b
      12'hDED: dout <= 8'b01100011; // 3565 :  99 - 0x63
      12'hDEE: dout <= 8'b01100011; // 3566 :  99 - 0x63
      12'hDEF: dout <= 8'b00000000; // 3567 :   0 - 0x0
      12'hDF0: dout <= 8'b01100011; // 3568 :  99 - 0x63 -- Background 0xbe
      12'hDF1: dout <= 8'b01100011; // 3569 :  99 - 0x63
      12'hDF2: dout <= 8'b01100011; // 3570 :  99 - 0x63
      12'hDF3: dout <= 8'b01110111; // 3571 : 119 - 0x77
      12'hDF4: dout <= 8'b00111110; // 3572 :  62 - 0x3e
      12'hDF5: dout <= 8'b00011100; // 3573 :  28 - 0x1c
      12'hDF6: dout <= 8'b00001000; // 3574 :   8 - 0x8
      12'hDF7: dout <= 8'b00000000; // 3575 :   0 - 0x0
      12'hDF8: dout <= 8'b00000000; // 3576 :   0 - 0x0 -- Background 0xbf
      12'hDF9: dout <= 8'b00000000; // 3577 :   0 - 0x0
      12'hDFA: dout <= 8'b00000000; // 3578 :   0 - 0x0
      12'hDFB: dout <= 8'b00000000; // 3579 :   0 - 0x0
      12'hDFC: dout <= 8'b00000000; // 3580 :   0 - 0x0
      12'hDFD: dout <= 8'b00000000; // 3581 :   0 - 0x0
      12'hDFE: dout <= 8'b00000000; // 3582 :   0 - 0x0
      12'hDFF: dout <= 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout <= 8'b00011111; // 3584 :  31 - 0x1f -- Background 0xc0
      12'hE01: dout <= 8'b00110000; // 3585 :  48 - 0x30
      12'hE02: dout <= 8'b01100000; // 3586 :  96 - 0x60
      12'hE03: dout <= 8'b01100111; // 3587 : 103 - 0x67
      12'hE04: dout <= 8'b01100011; // 3588 :  99 - 0x63
      12'hE05: dout <= 8'b00110011; // 3589 :  51 - 0x33
      12'hE06: dout <= 8'b00011111; // 3590 :  31 - 0x1f
      12'hE07: dout <= 8'b00000000; // 3591 :   0 - 0x0
      12'hE08: dout <= 8'b00011100; // 3592 :  28 - 0x1c -- Background 0xc1
      12'hE09: dout <= 8'b00110110; // 3593 :  54 - 0x36
      12'hE0A: dout <= 8'b01100011; // 3594 :  99 - 0x63
      12'hE0B: dout <= 8'b01100011; // 3595 :  99 - 0x63
      12'hE0C: dout <= 8'b01111111; // 3596 : 127 - 0x7f
      12'hE0D: dout <= 8'b01100011; // 3597 :  99 - 0x63
      12'hE0E: dout <= 8'b01100011; // 3598 :  99 - 0x63
      12'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout <= 8'b01100011; // 3600 :  99 - 0x63 -- Background 0xc2
      12'hE11: dout <= 8'b01110111; // 3601 : 119 - 0x77
      12'hE12: dout <= 8'b01111111; // 3602 : 127 - 0x7f
      12'hE13: dout <= 8'b01111111; // 3603 : 127 - 0x7f
      12'hE14: dout <= 8'b01101011; // 3604 : 107 - 0x6b
      12'hE15: dout <= 8'b01100011; // 3605 :  99 - 0x63
      12'hE16: dout <= 8'b01100011; // 3606 :  99 - 0x63
      12'hE17: dout <= 8'b00000000; // 3607 :   0 - 0x0
      12'hE18: dout <= 8'b01111111; // 3608 : 127 - 0x7f -- Background 0xc3
      12'hE19: dout <= 8'b01100000; // 3609 :  96 - 0x60
      12'hE1A: dout <= 8'b01100000; // 3610 :  96 - 0x60
      12'hE1B: dout <= 8'b01111110; // 3611 : 126 - 0x7e
      12'hE1C: dout <= 8'b01100000; // 3612 :  96 - 0x60
      12'hE1D: dout <= 8'b01100000; // 3613 :  96 - 0x60
      12'hE1E: dout <= 8'b01111111; // 3614 : 127 - 0x7f
      12'hE1F: dout <= 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout <= 8'b00111110; // 3616 :  62 - 0x3e -- Background 0xc4
      12'hE21: dout <= 8'b01100011; // 3617 :  99 - 0x63
      12'hE22: dout <= 8'b01100011; // 3618 :  99 - 0x63
      12'hE23: dout <= 8'b01100011; // 3619 :  99 - 0x63
      12'hE24: dout <= 8'b01100011; // 3620 :  99 - 0x63
      12'hE25: dout <= 8'b01100011; // 3621 :  99 - 0x63
      12'hE26: dout <= 8'b00111110; // 3622 :  62 - 0x3e
      12'hE27: dout <= 8'b00000000; // 3623 :   0 - 0x0
      12'hE28: dout <= 8'b01100011; // 3624 :  99 - 0x63 -- Background 0xc5
      12'hE29: dout <= 8'b01100011; // 3625 :  99 - 0x63
      12'hE2A: dout <= 8'b01100011; // 3626 :  99 - 0x63
      12'hE2B: dout <= 8'b01110111; // 3627 : 119 - 0x77
      12'hE2C: dout <= 8'b00111110; // 3628 :  62 - 0x3e
      12'hE2D: dout <= 8'b00011100; // 3629 :  28 - 0x1c
      12'hE2E: dout <= 8'b00001000; // 3630 :   8 - 0x8
      12'hE2F: dout <= 8'b00000000; // 3631 :   0 - 0x0
      12'hE30: dout <= 8'b01111110; // 3632 : 126 - 0x7e -- Background 0xc6
      12'hE31: dout <= 8'b01100011; // 3633 :  99 - 0x63
      12'hE32: dout <= 8'b01100011; // 3634 :  99 - 0x63
      12'hE33: dout <= 8'b01100111; // 3635 : 103 - 0x67
      12'hE34: dout <= 8'b01111100; // 3636 : 124 - 0x7c
      12'hE35: dout <= 8'b01101110; // 3637 : 110 - 0x6e
      12'hE36: dout <= 8'b01100111; // 3638 : 103 - 0x67
      12'hE37: dout <= 8'b00000000; // 3639 :   0 - 0x0
      12'hE38: dout <= 8'b00110011; // 3640 :  51 - 0x33 -- Background 0xc7
      12'hE39: dout <= 8'b00110011; // 3641 :  51 - 0x33
      12'hE3A: dout <= 8'b00110011; // 3642 :  51 - 0x33
      12'hE3B: dout <= 8'b00011110; // 3643 :  30 - 0x1e
      12'hE3C: dout <= 8'b00001100; // 3644 :  12 - 0xc
      12'hE3D: dout <= 8'b00001100; // 3645 :  12 - 0xc
      12'hE3E: dout <= 8'b00001100; // 3646 :  12 - 0xc
      12'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout <= 8'b00000000; // 3648 :   0 - 0x0 -- Background 0xc8
      12'hE41: dout <= 8'b00000000; // 3649 :   0 - 0x0
      12'hE42: dout <= 8'b00000000; // 3650 :   0 - 0x0
      12'hE43: dout <= 8'b00000000; // 3651 :   0 - 0x0
      12'hE44: dout <= 8'b00000000; // 3652 :   0 - 0x0
      12'hE45: dout <= 8'b00000000; // 3653 :   0 - 0x0
      12'hE46: dout <= 8'b00000000; // 3654 :   0 - 0x0
      12'hE47: dout <= 8'b00000000; // 3655 :   0 - 0x0
      12'hE48: dout <= 8'b00000000; // 3656 :   0 - 0x0 -- Background 0xc9
      12'hE49: dout <= 8'b00000000; // 3657 :   0 - 0x0
      12'hE4A: dout <= 8'b00000000; // 3658 :   0 - 0x0
      12'hE4B: dout <= 8'b00000000; // 3659 :   0 - 0x0
      12'hE4C: dout <= 8'b00000000; // 3660 :   0 - 0x0
      12'hE4D: dout <= 8'b00000000; // 3661 :   0 - 0x0
      12'hE4E: dout <= 8'b00000000; // 3662 :   0 - 0x0
      12'hE4F: dout <= 8'b00000000; // 3663 :   0 - 0x0
      12'hE50: dout <= 8'b00000000; // 3664 :   0 - 0x0 -- Background 0xca
      12'hE51: dout <= 8'b00000000; // 3665 :   0 - 0x0
      12'hE52: dout <= 8'b00000000; // 3666 :   0 - 0x0
      12'hE53: dout <= 8'b00000000; // 3667 :   0 - 0x0
      12'hE54: dout <= 8'b00000000; // 3668 :   0 - 0x0
      12'hE55: dout <= 8'b00000000; // 3669 :   0 - 0x0
      12'hE56: dout <= 8'b00000000; // 3670 :   0 - 0x0
      12'hE57: dout <= 8'b00000000; // 3671 :   0 - 0x0
      12'hE58: dout <= 8'b00000000; // 3672 :   0 - 0x0 -- Background 0xcb
      12'hE59: dout <= 8'b00000000; // 3673 :   0 - 0x0
      12'hE5A: dout <= 8'b00000000; // 3674 :   0 - 0x0
      12'hE5B: dout <= 8'b00000000; // 3675 :   0 - 0x0
      12'hE5C: dout <= 8'b00000000; // 3676 :   0 - 0x0
      12'hE5D: dout <= 8'b00000000; // 3677 :   0 - 0x0
      12'hE5E: dout <= 8'b00000000; // 3678 :   0 - 0x0
      12'hE5F: dout <= 8'b00000000; // 3679 :   0 - 0x0
      12'hE60: dout <= 8'b00000000; // 3680 :   0 - 0x0 -- Background 0xcc
      12'hE61: dout <= 8'b00000000; // 3681 :   0 - 0x0
      12'hE62: dout <= 8'b00000000; // 3682 :   0 - 0x0
      12'hE63: dout <= 8'b00000000; // 3683 :   0 - 0x0
      12'hE64: dout <= 8'b00000000; // 3684 :   0 - 0x0
      12'hE65: dout <= 8'b00000000; // 3685 :   0 - 0x0
      12'hE66: dout <= 8'b00000000; // 3686 :   0 - 0x0
      12'hE67: dout <= 8'b00000000; // 3687 :   0 - 0x0
      12'hE68: dout <= 8'b00000000; // 3688 :   0 - 0x0 -- Background 0xcd
      12'hE69: dout <= 8'b00000000; // 3689 :   0 - 0x0
      12'hE6A: dout <= 8'b00000000; // 3690 :   0 - 0x0
      12'hE6B: dout <= 8'b00000000; // 3691 :   0 - 0x0
      12'hE6C: dout <= 8'b00000000; // 3692 :   0 - 0x0
      12'hE6D: dout <= 8'b00000000; // 3693 :   0 - 0x0
      12'hE6E: dout <= 8'b00000000; // 3694 :   0 - 0x0
      12'hE6F: dout <= 8'b00000000; // 3695 :   0 - 0x0
      12'hE70: dout <= 8'b00000000; // 3696 :   0 - 0x0 -- Background 0xce
      12'hE71: dout <= 8'b00000000; // 3697 :   0 - 0x0
      12'hE72: dout <= 8'b00000000; // 3698 :   0 - 0x0
      12'hE73: dout <= 8'b00000000; // 3699 :   0 - 0x0
      12'hE74: dout <= 8'b00000000; // 3700 :   0 - 0x0
      12'hE75: dout <= 8'b00000000; // 3701 :   0 - 0x0
      12'hE76: dout <= 8'b00000000; // 3702 :   0 - 0x0
      12'hE77: dout <= 8'b00000000; // 3703 :   0 - 0x0
      12'hE78: dout <= 8'b00000000; // 3704 :   0 - 0x0 -- Background 0xcf
      12'hE79: dout <= 8'b00000000; // 3705 :   0 - 0x0
      12'hE7A: dout <= 8'b00000000; // 3706 :   0 - 0x0
      12'hE7B: dout <= 8'b00000000; // 3707 :   0 - 0x0
      12'hE7C: dout <= 8'b00000000; // 3708 :   0 - 0x0
      12'hE7D: dout <= 8'b00000000; // 3709 :   0 - 0x0
      12'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout <= 8'b11111111; // 3712 : 255 - 0xff -- Background 0xd0
      12'hE81: dout <= 8'b11111111; // 3713 : 255 - 0xff
      12'hE82: dout <= 8'b11111111; // 3714 : 255 - 0xff
      12'hE83: dout <= 8'b11111111; // 3715 : 255 - 0xff
      12'hE84: dout <= 8'b11111111; // 3716 : 255 - 0xff
      12'hE85: dout <= 8'b11111111; // 3717 : 255 - 0xff
      12'hE86: dout <= 8'b11111111; // 3718 : 255 - 0xff
      12'hE87: dout <= 8'b11111111; // 3719 : 255 - 0xff
      12'hE88: dout <= 8'b11111111; // 3720 : 255 - 0xff -- Background 0xd1
      12'hE89: dout <= 8'b11111111; // 3721 : 255 - 0xff
      12'hE8A: dout <= 8'b11111111; // 3722 : 255 - 0xff
      12'hE8B: dout <= 8'b11111111; // 3723 : 255 - 0xff
      12'hE8C: dout <= 8'b11111111; // 3724 : 255 - 0xff
      12'hE8D: dout <= 8'b11111111; // 3725 : 255 - 0xff
      12'hE8E: dout <= 8'b11111111; // 3726 : 255 - 0xff
      12'hE8F: dout <= 8'b11111111; // 3727 : 255 - 0xff
      12'hE90: dout <= 8'b11111111; // 3728 : 255 - 0xff -- Background 0xd2
      12'hE91: dout <= 8'b11111111; // 3729 : 255 - 0xff
      12'hE92: dout <= 8'b11111111; // 3730 : 255 - 0xff
      12'hE93: dout <= 8'b11111111; // 3731 : 255 - 0xff
      12'hE94: dout <= 8'b11111111; // 3732 : 255 - 0xff
      12'hE95: dout <= 8'b11111111; // 3733 : 255 - 0xff
      12'hE96: dout <= 8'b11111111; // 3734 : 255 - 0xff
      12'hE97: dout <= 8'b11111111; // 3735 : 255 - 0xff
      12'hE98: dout <= 8'b11111111; // 3736 : 255 - 0xff -- Background 0xd3
      12'hE99: dout <= 8'b11111111; // 3737 : 255 - 0xff
      12'hE9A: dout <= 8'b11111111; // 3738 : 255 - 0xff
      12'hE9B: dout <= 8'b11111111; // 3739 : 255 - 0xff
      12'hE9C: dout <= 8'b11111111; // 3740 : 255 - 0xff
      12'hE9D: dout <= 8'b11111111; // 3741 : 255 - 0xff
      12'hE9E: dout <= 8'b11111111; // 3742 : 255 - 0xff
      12'hE9F: dout <= 8'b11111111; // 3743 : 255 - 0xff
      12'hEA0: dout <= 8'b11111111; // 3744 : 255 - 0xff -- Background 0xd4
      12'hEA1: dout <= 8'b11111111; // 3745 : 255 - 0xff
      12'hEA2: dout <= 8'b11111111; // 3746 : 255 - 0xff
      12'hEA3: dout <= 8'b11111111; // 3747 : 255 - 0xff
      12'hEA4: dout <= 8'b11111111; // 3748 : 255 - 0xff
      12'hEA5: dout <= 8'b11111111; // 3749 : 255 - 0xff
      12'hEA6: dout <= 8'b11111111; // 3750 : 255 - 0xff
      12'hEA7: dout <= 8'b11111111; // 3751 : 255 - 0xff
      12'hEA8: dout <= 8'b11111111; // 3752 : 255 - 0xff -- Background 0xd5
      12'hEA9: dout <= 8'b11111111; // 3753 : 255 - 0xff
      12'hEAA: dout <= 8'b11111111; // 3754 : 255 - 0xff
      12'hEAB: dout <= 8'b11111111; // 3755 : 255 - 0xff
      12'hEAC: dout <= 8'b11111111; // 3756 : 255 - 0xff
      12'hEAD: dout <= 8'b11111111; // 3757 : 255 - 0xff
      12'hEAE: dout <= 8'b11111111; // 3758 : 255 - 0xff
      12'hEAF: dout <= 8'b11111111; // 3759 : 255 - 0xff
      12'hEB0: dout <= 8'b11111111; // 3760 : 255 - 0xff -- Background 0xd6
      12'hEB1: dout <= 8'b11111111; // 3761 : 255 - 0xff
      12'hEB2: dout <= 8'b11111111; // 3762 : 255 - 0xff
      12'hEB3: dout <= 8'b11111111; // 3763 : 255 - 0xff
      12'hEB4: dout <= 8'b11111111; // 3764 : 255 - 0xff
      12'hEB5: dout <= 8'b11111111; // 3765 : 255 - 0xff
      12'hEB6: dout <= 8'b11111111; // 3766 : 255 - 0xff
      12'hEB7: dout <= 8'b11111111; // 3767 : 255 - 0xff
      12'hEB8: dout <= 8'b11111111; // 3768 : 255 - 0xff -- Background 0xd7
      12'hEB9: dout <= 8'b11111111; // 3769 : 255 - 0xff
      12'hEBA: dout <= 8'b11111111; // 3770 : 255 - 0xff
      12'hEBB: dout <= 8'b11111111; // 3771 : 255 - 0xff
      12'hEBC: dout <= 8'b11111111; // 3772 : 255 - 0xff
      12'hEBD: dout <= 8'b11111111; // 3773 : 255 - 0xff
      12'hEBE: dout <= 8'b11111111; // 3774 : 255 - 0xff
      12'hEBF: dout <= 8'b11111111; // 3775 : 255 - 0xff
      12'hEC0: dout <= 8'b11111111; // 3776 : 255 - 0xff -- Background 0xd8
      12'hEC1: dout <= 8'b11111111; // 3777 : 255 - 0xff
      12'hEC2: dout <= 8'b11111111; // 3778 : 255 - 0xff
      12'hEC3: dout <= 8'b11111111; // 3779 : 255 - 0xff
      12'hEC4: dout <= 8'b11111111; // 3780 : 255 - 0xff
      12'hEC5: dout <= 8'b11111111; // 3781 : 255 - 0xff
      12'hEC6: dout <= 8'b11111111; // 3782 : 255 - 0xff
      12'hEC7: dout <= 8'b11111111; // 3783 : 255 - 0xff
      12'hEC8: dout <= 8'b11111111; // 3784 : 255 - 0xff -- Background 0xd9
      12'hEC9: dout <= 8'b11111111; // 3785 : 255 - 0xff
      12'hECA: dout <= 8'b11111111; // 3786 : 255 - 0xff
      12'hECB: dout <= 8'b11111111; // 3787 : 255 - 0xff
      12'hECC: dout <= 8'b11111111; // 3788 : 255 - 0xff
      12'hECD: dout <= 8'b11111111; // 3789 : 255 - 0xff
      12'hECE: dout <= 8'b11111111; // 3790 : 255 - 0xff
      12'hECF: dout <= 8'b11111111; // 3791 : 255 - 0xff
      12'hED0: dout <= 8'b11111111; // 3792 : 255 - 0xff -- Background 0xda
      12'hED1: dout <= 8'b11111111; // 3793 : 255 - 0xff
      12'hED2: dout <= 8'b11111111; // 3794 : 255 - 0xff
      12'hED3: dout <= 8'b11111111; // 3795 : 255 - 0xff
      12'hED4: dout <= 8'b11111111; // 3796 : 255 - 0xff
      12'hED5: dout <= 8'b11111111; // 3797 : 255 - 0xff
      12'hED6: dout <= 8'b11111111; // 3798 : 255 - 0xff
      12'hED7: dout <= 8'b11111111; // 3799 : 255 - 0xff
      12'hED8: dout <= 8'b11111111; // 3800 : 255 - 0xff -- Background 0xdb
      12'hED9: dout <= 8'b11111111; // 3801 : 255 - 0xff
      12'hEDA: dout <= 8'b11111111; // 3802 : 255 - 0xff
      12'hEDB: dout <= 8'b11111111; // 3803 : 255 - 0xff
      12'hEDC: dout <= 8'b11111111; // 3804 : 255 - 0xff
      12'hEDD: dout <= 8'b11111111; // 3805 : 255 - 0xff
      12'hEDE: dout <= 8'b11111111; // 3806 : 255 - 0xff
      12'hEDF: dout <= 8'b11111111; // 3807 : 255 - 0xff
      12'hEE0: dout <= 8'b11111111; // 3808 : 255 - 0xff -- Background 0xdc
      12'hEE1: dout <= 8'b11111111; // 3809 : 255 - 0xff
      12'hEE2: dout <= 8'b11111111; // 3810 : 255 - 0xff
      12'hEE3: dout <= 8'b11111111; // 3811 : 255 - 0xff
      12'hEE4: dout <= 8'b11111111; // 3812 : 255 - 0xff
      12'hEE5: dout <= 8'b11111111; // 3813 : 255 - 0xff
      12'hEE6: dout <= 8'b11111111; // 3814 : 255 - 0xff
      12'hEE7: dout <= 8'b11111111; // 3815 : 255 - 0xff
      12'hEE8: dout <= 8'b11111111; // 3816 : 255 - 0xff -- Background 0xdd
      12'hEE9: dout <= 8'b11111111; // 3817 : 255 - 0xff
      12'hEEA: dout <= 8'b11111111; // 3818 : 255 - 0xff
      12'hEEB: dout <= 8'b11111111; // 3819 : 255 - 0xff
      12'hEEC: dout <= 8'b11111111; // 3820 : 255 - 0xff
      12'hEED: dout <= 8'b11111111; // 3821 : 255 - 0xff
      12'hEEE: dout <= 8'b11111111; // 3822 : 255 - 0xff
      12'hEEF: dout <= 8'b11111111; // 3823 : 255 - 0xff
      12'hEF0: dout <= 8'b11111111; // 3824 : 255 - 0xff -- Background 0xde
      12'hEF1: dout <= 8'b11111111; // 3825 : 255 - 0xff
      12'hEF2: dout <= 8'b11111111; // 3826 : 255 - 0xff
      12'hEF3: dout <= 8'b11111111; // 3827 : 255 - 0xff
      12'hEF4: dout <= 8'b11111111; // 3828 : 255 - 0xff
      12'hEF5: dout <= 8'b11111111; // 3829 : 255 - 0xff
      12'hEF6: dout <= 8'b11111111; // 3830 : 255 - 0xff
      12'hEF7: dout <= 8'b11111111; // 3831 : 255 - 0xff
      12'hEF8: dout <= 8'b11111111; // 3832 : 255 - 0xff -- Background 0xdf
      12'hEF9: dout <= 8'b11111111; // 3833 : 255 - 0xff
      12'hEFA: dout <= 8'b11111111; // 3834 : 255 - 0xff
      12'hEFB: dout <= 8'b11111111; // 3835 : 255 - 0xff
      12'hEFC: dout <= 8'b11111111; // 3836 : 255 - 0xff
      12'hEFD: dout <= 8'b11111111; // 3837 : 255 - 0xff
      12'hEFE: dout <= 8'b11111111; // 3838 : 255 - 0xff
      12'hEFF: dout <= 8'b11111111; // 3839 : 255 - 0xff
      12'hF00: dout <= 8'b11111111; // 3840 : 255 - 0xff -- Background 0xe0
      12'hF01: dout <= 8'b11111111; // 3841 : 255 - 0xff
      12'hF02: dout <= 8'b11111111; // 3842 : 255 - 0xff
      12'hF03: dout <= 8'b11111111; // 3843 : 255 - 0xff
      12'hF04: dout <= 8'b11111111; // 3844 : 255 - 0xff
      12'hF05: dout <= 8'b11111111; // 3845 : 255 - 0xff
      12'hF06: dout <= 8'b11111111; // 3846 : 255 - 0xff
      12'hF07: dout <= 8'b11111111; // 3847 : 255 - 0xff
      12'hF08: dout <= 8'b11111111; // 3848 : 255 - 0xff -- Background 0xe1
      12'hF09: dout <= 8'b11111111; // 3849 : 255 - 0xff
      12'hF0A: dout <= 8'b11111111; // 3850 : 255 - 0xff
      12'hF0B: dout <= 8'b11111111; // 3851 : 255 - 0xff
      12'hF0C: dout <= 8'b11111111; // 3852 : 255 - 0xff
      12'hF0D: dout <= 8'b11111111; // 3853 : 255 - 0xff
      12'hF0E: dout <= 8'b11111111; // 3854 : 255 - 0xff
      12'hF0F: dout <= 8'b11111111; // 3855 : 255 - 0xff
      12'hF10: dout <= 8'b11111111; // 3856 : 255 - 0xff -- Background 0xe2
      12'hF11: dout <= 8'b11111111; // 3857 : 255 - 0xff
      12'hF12: dout <= 8'b11111111; // 3858 : 255 - 0xff
      12'hF13: dout <= 8'b11111111; // 3859 : 255 - 0xff
      12'hF14: dout <= 8'b11111111; // 3860 : 255 - 0xff
      12'hF15: dout <= 8'b11111111; // 3861 : 255 - 0xff
      12'hF16: dout <= 8'b11111111; // 3862 : 255 - 0xff
      12'hF17: dout <= 8'b11111111; // 3863 : 255 - 0xff
      12'hF18: dout <= 8'b11111111; // 3864 : 255 - 0xff -- Background 0xe3
      12'hF19: dout <= 8'b11111111; // 3865 : 255 - 0xff
      12'hF1A: dout <= 8'b11111111; // 3866 : 255 - 0xff
      12'hF1B: dout <= 8'b11111111; // 3867 : 255 - 0xff
      12'hF1C: dout <= 8'b11111111; // 3868 : 255 - 0xff
      12'hF1D: dout <= 8'b11111111; // 3869 : 255 - 0xff
      12'hF1E: dout <= 8'b11111111; // 3870 : 255 - 0xff
      12'hF1F: dout <= 8'b11111111; // 3871 : 255 - 0xff
      12'hF20: dout <= 8'b11111111; // 3872 : 255 - 0xff -- Background 0xe4
      12'hF21: dout <= 8'b11111111; // 3873 : 255 - 0xff
      12'hF22: dout <= 8'b11111111; // 3874 : 255 - 0xff
      12'hF23: dout <= 8'b11111111; // 3875 : 255 - 0xff
      12'hF24: dout <= 8'b11111111; // 3876 : 255 - 0xff
      12'hF25: dout <= 8'b11111111; // 3877 : 255 - 0xff
      12'hF26: dout <= 8'b11111111; // 3878 : 255 - 0xff
      12'hF27: dout <= 8'b11111111; // 3879 : 255 - 0xff
      12'hF28: dout <= 8'b11111111; // 3880 : 255 - 0xff -- Background 0xe5
      12'hF29: dout <= 8'b11111111; // 3881 : 255 - 0xff
      12'hF2A: dout <= 8'b11111111; // 3882 : 255 - 0xff
      12'hF2B: dout <= 8'b11111111; // 3883 : 255 - 0xff
      12'hF2C: dout <= 8'b11111111; // 3884 : 255 - 0xff
      12'hF2D: dout <= 8'b11111111; // 3885 : 255 - 0xff
      12'hF2E: dout <= 8'b11111111; // 3886 : 255 - 0xff
      12'hF2F: dout <= 8'b11111111; // 3887 : 255 - 0xff
      12'hF30: dout <= 8'b11111111; // 3888 : 255 - 0xff -- Background 0xe6
      12'hF31: dout <= 8'b11111111; // 3889 : 255 - 0xff
      12'hF32: dout <= 8'b11111111; // 3890 : 255 - 0xff
      12'hF33: dout <= 8'b11111111; // 3891 : 255 - 0xff
      12'hF34: dout <= 8'b11111111; // 3892 : 255 - 0xff
      12'hF35: dout <= 8'b11111111; // 3893 : 255 - 0xff
      12'hF36: dout <= 8'b11111111; // 3894 : 255 - 0xff
      12'hF37: dout <= 8'b11111111; // 3895 : 255 - 0xff
      12'hF38: dout <= 8'b11111111; // 3896 : 255 - 0xff -- Background 0xe7
      12'hF39: dout <= 8'b11111111; // 3897 : 255 - 0xff
      12'hF3A: dout <= 8'b11111111; // 3898 : 255 - 0xff
      12'hF3B: dout <= 8'b11111111; // 3899 : 255 - 0xff
      12'hF3C: dout <= 8'b11111111; // 3900 : 255 - 0xff
      12'hF3D: dout <= 8'b11111111; // 3901 : 255 - 0xff
      12'hF3E: dout <= 8'b11111111; // 3902 : 255 - 0xff
      12'hF3F: dout <= 8'b11111111; // 3903 : 255 - 0xff
      12'hF40: dout <= 8'b11111111; // 3904 : 255 - 0xff -- Background 0xe8
      12'hF41: dout <= 8'b11111111; // 3905 : 255 - 0xff
      12'hF42: dout <= 8'b11111111; // 3906 : 255 - 0xff
      12'hF43: dout <= 8'b11111111; // 3907 : 255 - 0xff
      12'hF44: dout <= 8'b11111111; // 3908 : 255 - 0xff
      12'hF45: dout <= 8'b11111111; // 3909 : 255 - 0xff
      12'hF46: dout <= 8'b11111111; // 3910 : 255 - 0xff
      12'hF47: dout <= 8'b11111111; // 3911 : 255 - 0xff
      12'hF48: dout <= 8'b11111111; // 3912 : 255 - 0xff -- Background 0xe9
      12'hF49: dout <= 8'b11111111; // 3913 : 255 - 0xff
      12'hF4A: dout <= 8'b11111111; // 3914 : 255 - 0xff
      12'hF4B: dout <= 8'b11111111; // 3915 : 255 - 0xff
      12'hF4C: dout <= 8'b11111111; // 3916 : 255 - 0xff
      12'hF4D: dout <= 8'b11111111; // 3917 : 255 - 0xff
      12'hF4E: dout <= 8'b11111111; // 3918 : 255 - 0xff
      12'hF4F: dout <= 8'b11111111; // 3919 : 255 - 0xff
      12'hF50: dout <= 8'b11111111; // 3920 : 255 - 0xff -- Background 0xea
      12'hF51: dout <= 8'b11111111; // 3921 : 255 - 0xff
      12'hF52: dout <= 8'b11111111; // 3922 : 255 - 0xff
      12'hF53: dout <= 8'b11111111; // 3923 : 255 - 0xff
      12'hF54: dout <= 8'b11111111; // 3924 : 255 - 0xff
      12'hF55: dout <= 8'b11111111; // 3925 : 255 - 0xff
      12'hF56: dout <= 8'b11111111; // 3926 : 255 - 0xff
      12'hF57: dout <= 8'b11111111; // 3927 : 255 - 0xff
      12'hF58: dout <= 8'b11111111; // 3928 : 255 - 0xff -- Background 0xeb
      12'hF59: dout <= 8'b11111111; // 3929 : 255 - 0xff
      12'hF5A: dout <= 8'b11111111; // 3930 : 255 - 0xff
      12'hF5B: dout <= 8'b11111111; // 3931 : 255 - 0xff
      12'hF5C: dout <= 8'b11111111; // 3932 : 255 - 0xff
      12'hF5D: dout <= 8'b11111111; // 3933 : 255 - 0xff
      12'hF5E: dout <= 8'b11111111; // 3934 : 255 - 0xff
      12'hF5F: dout <= 8'b11111111; // 3935 : 255 - 0xff
      12'hF60: dout <= 8'b11111111; // 3936 : 255 - 0xff -- Background 0xec
      12'hF61: dout <= 8'b11111111; // 3937 : 255 - 0xff
      12'hF62: dout <= 8'b11111111; // 3938 : 255 - 0xff
      12'hF63: dout <= 8'b11111111; // 3939 : 255 - 0xff
      12'hF64: dout <= 8'b11111111; // 3940 : 255 - 0xff
      12'hF65: dout <= 8'b11111111; // 3941 : 255 - 0xff
      12'hF66: dout <= 8'b11111111; // 3942 : 255 - 0xff
      12'hF67: dout <= 8'b11111111; // 3943 : 255 - 0xff
      12'hF68: dout <= 8'b11111111; // 3944 : 255 - 0xff -- Background 0xed
      12'hF69: dout <= 8'b11111111; // 3945 : 255 - 0xff
      12'hF6A: dout <= 8'b11111111; // 3946 : 255 - 0xff
      12'hF6B: dout <= 8'b11111111; // 3947 : 255 - 0xff
      12'hF6C: dout <= 8'b11111111; // 3948 : 255 - 0xff
      12'hF6D: dout <= 8'b11111111; // 3949 : 255 - 0xff
      12'hF6E: dout <= 8'b11111111; // 3950 : 255 - 0xff
      12'hF6F: dout <= 8'b11111111; // 3951 : 255 - 0xff
      12'hF70: dout <= 8'b11111111; // 3952 : 255 - 0xff -- Background 0xee
      12'hF71: dout <= 8'b11111111; // 3953 : 255 - 0xff
      12'hF72: dout <= 8'b11111111; // 3954 : 255 - 0xff
      12'hF73: dout <= 8'b11111111; // 3955 : 255 - 0xff
      12'hF74: dout <= 8'b11111111; // 3956 : 255 - 0xff
      12'hF75: dout <= 8'b11111111; // 3957 : 255 - 0xff
      12'hF76: dout <= 8'b11111111; // 3958 : 255 - 0xff
      12'hF77: dout <= 8'b11111111; // 3959 : 255 - 0xff
      12'hF78: dout <= 8'b11111111; // 3960 : 255 - 0xff -- Background 0xef
      12'hF79: dout <= 8'b11111111; // 3961 : 255 - 0xff
      12'hF7A: dout <= 8'b11111111; // 3962 : 255 - 0xff
      12'hF7B: dout <= 8'b11111111; // 3963 : 255 - 0xff
      12'hF7C: dout <= 8'b11111111; // 3964 : 255 - 0xff
      12'hF7D: dout <= 8'b11111111; // 3965 : 255 - 0xff
      12'hF7E: dout <= 8'b11111111; // 3966 : 255 - 0xff
      12'hF7F: dout <= 8'b11111111; // 3967 : 255 - 0xff
      12'hF80: dout <= 8'b11111111; // 3968 : 255 - 0xff -- Background 0xf0
      12'hF81: dout <= 8'b11111111; // 3969 : 255 - 0xff
      12'hF82: dout <= 8'b11111111; // 3970 : 255 - 0xff
      12'hF83: dout <= 8'b11111111; // 3971 : 255 - 0xff
      12'hF84: dout <= 8'b11111111; // 3972 : 255 - 0xff
      12'hF85: dout <= 8'b11111111; // 3973 : 255 - 0xff
      12'hF86: dout <= 8'b11111111; // 3974 : 255 - 0xff
      12'hF87: dout <= 8'b11111111; // 3975 : 255 - 0xff
      12'hF88: dout <= 8'b11111111; // 3976 : 255 - 0xff -- Background 0xf1
      12'hF89: dout <= 8'b11111111; // 3977 : 255 - 0xff
      12'hF8A: dout <= 8'b11111111; // 3978 : 255 - 0xff
      12'hF8B: dout <= 8'b11111111; // 3979 : 255 - 0xff
      12'hF8C: dout <= 8'b11111111; // 3980 : 255 - 0xff
      12'hF8D: dout <= 8'b11111111; // 3981 : 255 - 0xff
      12'hF8E: dout <= 8'b11111111; // 3982 : 255 - 0xff
      12'hF8F: dout <= 8'b11111111; // 3983 : 255 - 0xff
      12'hF90: dout <= 8'b11111111; // 3984 : 255 - 0xff -- Background 0xf2
      12'hF91: dout <= 8'b11111111; // 3985 : 255 - 0xff
      12'hF92: dout <= 8'b11111111; // 3986 : 255 - 0xff
      12'hF93: dout <= 8'b11111111; // 3987 : 255 - 0xff
      12'hF94: dout <= 8'b11111111; // 3988 : 255 - 0xff
      12'hF95: dout <= 8'b11111111; // 3989 : 255 - 0xff
      12'hF96: dout <= 8'b11111111; // 3990 : 255 - 0xff
      12'hF97: dout <= 8'b11111111; // 3991 : 255 - 0xff
      12'hF98: dout <= 8'b11111111; // 3992 : 255 - 0xff -- Background 0xf3
      12'hF99: dout <= 8'b11111111; // 3993 : 255 - 0xff
      12'hF9A: dout <= 8'b11111111; // 3994 : 255 - 0xff
      12'hF9B: dout <= 8'b11111111; // 3995 : 255 - 0xff
      12'hF9C: dout <= 8'b11111111; // 3996 : 255 - 0xff
      12'hF9D: dout <= 8'b11111111; // 3997 : 255 - 0xff
      12'hF9E: dout <= 8'b11111111; // 3998 : 255 - 0xff
      12'hF9F: dout <= 8'b11111111; // 3999 : 255 - 0xff
      12'hFA0: dout <= 8'b11111111; // 4000 : 255 - 0xff -- Background 0xf4
      12'hFA1: dout <= 8'b11111111; // 4001 : 255 - 0xff
      12'hFA2: dout <= 8'b11111111; // 4002 : 255 - 0xff
      12'hFA3: dout <= 8'b11111111; // 4003 : 255 - 0xff
      12'hFA4: dout <= 8'b11111111; // 4004 : 255 - 0xff
      12'hFA5: dout <= 8'b11111111; // 4005 : 255 - 0xff
      12'hFA6: dout <= 8'b11111111; // 4006 : 255 - 0xff
      12'hFA7: dout <= 8'b11111111; // 4007 : 255 - 0xff
      12'hFA8: dout <= 8'b11111111; // 4008 : 255 - 0xff -- Background 0xf5
      12'hFA9: dout <= 8'b11111111; // 4009 : 255 - 0xff
      12'hFAA: dout <= 8'b11111111; // 4010 : 255 - 0xff
      12'hFAB: dout <= 8'b11111111; // 4011 : 255 - 0xff
      12'hFAC: dout <= 8'b11111111; // 4012 : 255 - 0xff
      12'hFAD: dout <= 8'b11111111; // 4013 : 255 - 0xff
      12'hFAE: dout <= 8'b11111111; // 4014 : 255 - 0xff
      12'hFAF: dout <= 8'b11111111; // 4015 : 255 - 0xff
      12'hFB0: dout <= 8'b11111111; // 4016 : 255 - 0xff -- Background 0xf6
      12'hFB1: dout <= 8'b11111111; // 4017 : 255 - 0xff
      12'hFB2: dout <= 8'b11111111; // 4018 : 255 - 0xff
      12'hFB3: dout <= 8'b11111111; // 4019 : 255 - 0xff
      12'hFB4: dout <= 8'b11111111; // 4020 : 255 - 0xff
      12'hFB5: dout <= 8'b11111111; // 4021 : 255 - 0xff
      12'hFB6: dout <= 8'b11111111; // 4022 : 255 - 0xff
      12'hFB7: dout <= 8'b11111111; // 4023 : 255 - 0xff
      12'hFB8: dout <= 8'b11111111; // 4024 : 255 - 0xff -- Background 0xf7
      12'hFB9: dout <= 8'b11111111; // 4025 : 255 - 0xff
      12'hFBA: dout <= 8'b11111111; // 4026 : 255 - 0xff
      12'hFBB: dout <= 8'b11111111; // 4027 : 255 - 0xff
      12'hFBC: dout <= 8'b11111111; // 4028 : 255 - 0xff
      12'hFBD: dout <= 8'b11111111; // 4029 : 255 - 0xff
      12'hFBE: dout <= 8'b11111111; // 4030 : 255 - 0xff
      12'hFBF: dout <= 8'b11111111; // 4031 : 255 - 0xff
      12'hFC0: dout <= 8'b11111111; // 4032 : 255 - 0xff -- Background 0xf8
      12'hFC1: dout <= 8'b11111111; // 4033 : 255 - 0xff
      12'hFC2: dout <= 8'b11111111; // 4034 : 255 - 0xff
      12'hFC3: dout <= 8'b11111111; // 4035 : 255 - 0xff
      12'hFC4: dout <= 8'b11111111; // 4036 : 255 - 0xff
      12'hFC5: dout <= 8'b11111111; // 4037 : 255 - 0xff
      12'hFC6: dout <= 8'b11111111; // 4038 : 255 - 0xff
      12'hFC7: dout <= 8'b11111111; // 4039 : 255 - 0xff
      12'hFC8: dout <= 8'b11111111; // 4040 : 255 - 0xff -- Background 0xf9
      12'hFC9: dout <= 8'b11111111; // 4041 : 255 - 0xff
      12'hFCA: dout <= 8'b11111111; // 4042 : 255 - 0xff
      12'hFCB: dout <= 8'b11111111; // 4043 : 255 - 0xff
      12'hFCC: dout <= 8'b11111111; // 4044 : 255 - 0xff
      12'hFCD: dout <= 8'b11111111; // 4045 : 255 - 0xff
      12'hFCE: dout <= 8'b11111111; // 4046 : 255 - 0xff
      12'hFCF: dout <= 8'b11111111; // 4047 : 255 - 0xff
      12'hFD0: dout <= 8'b11111111; // 4048 : 255 - 0xff -- Background 0xfa
      12'hFD1: dout <= 8'b11111111; // 4049 : 255 - 0xff
      12'hFD2: dout <= 8'b11111111; // 4050 : 255 - 0xff
      12'hFD3: dout <= 8'b11111111; // 4051 : 255 - 0xff
      12'hFD4: dout <= 8'b11111111; // 4052 : 255 - 0xff
      12'hFD5: dout <= 8'b11111111; // 4053 : 255 - 0xff
      12'hFD6: dout <= 8'b11111111; // 4054 : 255 - 0xff
      12'hFD7: dout <= 8'b11111111; // 4055 : 255 - 0xff
      12'hFD8: dout <= 8'b11111111; // 4056 : 255 - 0xff -- Background 0xfb
      12'hFD9: dout <= 8'b11111111; // 4057 : 255 - 0xff
      12'hFDA: dout <= 8'b11111111; // 4058 : 255 - 0xff
      12'hFDB: dout <= 8'b11111111; // 4059 : 255 - 0xff
      12'hFDC: dout <= 8'b11111111; // 4060 : 255 - 0xff
      12'hFDD: dout <= 8'b11111111; // 4061 : 255 - 0xff
      12'hFDE: dout <= 8'b11111111; // 4062 : 255 - 0xff
      12'hFDF: dout <= 8'b11111111; // 4063 : 255 - 0xff
      12'hFE0: dout <= 8'b11111111; // 4064 : 255 - 0xff -- Background 0xfc
      12'hFE1: dout <= 8'b11111111; // 4065 : 255 - 0xff
      12'hFE2: dout <= 8'b11111111; // 4066 : 255 - 0xff
      12'hFE3: dout <= 8'b11111111; // 4067 : 255 - 0xff
      12'hFE4: dout <= 8'b11111111; // 4068 : 255 - 0xff
      12'hFE5: dout <= 8'b11111111; // 4069 : 255 - 0xff
      12'hFE6: dout <= 8'b11111111; // 4070 : 255 - 0xff
      12'hFE7: dout <= 8'b11111111; // 4071 : 255 - 0xff
      12'hFE8: dout <= 8'b11111111; // 4072 : 255 - 0xff -- Background 0xfd
      12'hFE9: dout <= 8'b11111111; // 4073 : 255 - 0xff
      12'hFEA: dout <= 8'b11111111; // 4074 : 255 - 0xff
      12'hFEB: dout <= 8'b11111111; // 4075 : 255 - 0xff
      12'hFEC: dout <= 8'b11111111; // 4076 : 255 - 0xff
      12'hFED: dout <= 8'b11111111; // 4077 : 255 - 0xff
      12'hFEE: dout <= 8'b11111111; // 4078 : 255 - 0xff
      12'hFEF: dout <= 8'b11111111; // 4079 : 255 - 0xff
      12'hFF0: dout <= 8'b11111111; // 4080 : 255 - 0xff -- Background 0xfe
      12'hFF1: dout <= 8'b11111111; // 4081 : 255 - 0xff
      12'hFF2: dout <= 8'b11111111; // 4082 : 255 - 0xff
      12'hFF3: dout <= 8'b11111111; // 4083 : 255 - 0xff
      12'hFF4: dout <= 8'b11111111; // 4084 : 255 - 0xff
      12'hFF5: dout <= 8'b11111111; // 4085 : 255 - 0xff
      12'hFF6: dout <= 8'b11111111; // 4086 : 255 - 0xff
      12'hFF7: dout <= 8'b11111111; // 4087 : 255 - 0xff
      12'hFF8: dout <= 8'b11111111; // 4088 : 255 - 0xff -- Background 0xff
      12'hFF9: dout <= 8'b11111111; // 4089 : 255 - 0xff
      12'hFFA: dout <= 8'b11111111; // 4090 : 255 - 0xff
      12'hFFB: dout <= 8'b11111111; // 4091 : 255 - 0xff
      12'hFFC: dout <= 8'b11111111; // 4092 : 255 - 0xff
      12'hFFD: dout <= 8'b11111111; // 4093 : 255 - 0xff
      12'hFFE: dout <= 8'b11111111; // 4094 : 255 - 0xff
      12'hFFF: dout <= 8'b11111111; // 4095 : 255 - 0xff
    endcase
  end

endmodule
