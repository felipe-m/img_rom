//-   Background Pattern table COLOR PLANE 1
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: smario_traspas_patron.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_MARIO_TRASPAS_BG_PLN1
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table COLOR PLANE 1
      11'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Background 0x0
      11'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      11'h2: dout  = 8'b00000000; //    2 :   0 - 0x0
      11'h3: dout  = 8'b00000000; //    3 :   0 - 0x0
      11'h4: dout  = 8'b00000000; //    4 :   0 - 0x0
      11'h5: dout  = 8'b00000000; //    5 :   0 - 0x0
      11'h6: dout  = 8'b00000000; //    6 :   0 - 0x0
      11'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      11'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- Background 0x1
      11'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      11'hA: dout  = 8'b00000000; //   10 :   0 - 0x0
      11'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      11'hC: dout  = 8'b00000000; //   12 :   0 - 0x0
      11'hD: dout  = 8'b00000000; //   13 :   0 - 0x0
      11'hE: dout  = 8'b00000000; //   14 :   0 - 0x0
      11'hF: dout  = 8'b00000000; //   15 :   0 - 0x0
      11'h10: dout  = 8'b00000000; //   16 :   0 - 0x0 -- Background 0x2
      11'h11: dout  = 8'b00000000; //   17 :   0 - 0x0
      11'h12: dout  = 8'b00000000; //   18 :   0 - 0x0
      11'h13: dout  = 8'b00000000; //   19 :   0 - 0x0
      11'h14: dout  = 8'b00000000; //   20 :   0 - 0x0
      11'h15: dout  = 8'b00000000; //   21 :   0 - 0x0
      11'h16: dout  = 8'b00000000; //   22 :   0 - 0x0
      11'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      11'h18: dout  = 8'b00000000; //   24 :   0 - 0x0 -- Background 0x3
      11'h19: dout  = 8'b00000000; //   25 :   0 - 0x0
      11'h1A: dout  = 8'b00000000; //   26 :   0 - 0x0
      11'h1B: dout  = 8'b00000000; //   27 :   0 - 0x0
      11'h1C: dout  = 8'b00000000; //   28 :   0 - 0x0
      11'h1D: dout  = 8'b00000000; //   29 :   0 - 0x0
      11'h1E: dout  = 8'b00000000; //   30 :   0 - 0x0
      11'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      11'h20: dout  = 8'b00000000; //   32 :   0 - 0x0 -- Background 0x4
      11'h21: dout  = 8'b00000000; //   33 :   0 - 0x0
      11'h22: dout  = 8'b00000000; //   34 :   0 - 0x0
      11'h23: dout  = 8'b00000000; //   35 :   0 - 0x0
      11'h24: dout  = 8'b00000000; //   36 :   0 - 0x0
      11'h25: dout  = 8'b00000000; //   37 :   0 - 0x0
      11'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      11'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      11'h28: dout  = 8'b00000000; //   40 :   0 - 0x0 -- Background 0x5
      11'h29: dout  = 8'b00000000; //   41 :   0 - 0x0
      11'h2A: dout  = 8'b00000000; //   42 :   0 - 0x0
      11'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      11'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      11'h2D: dout  = 8'b00000000; //   45 :   0 - 0x0
      11'h2E: dout  = 8'b00000000; //   46 :   0 - 0x0
      11'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      11'h30: dout  = 8'b00000000; //   48 :   0 - 0x0 -- Background 0x6
      11'h31: dout  = 8'b00000000; //   49 :   0 - 0x0
      11'h32: dout  = 8'b00000000; //   50 :   0 - 0x0
      11'h33: dout  = 8'b00000000; //   51 :   0 - 0x0
      11'h34: dout  = 8'b00000000; //   52 :   0 - 0x0
      11'h35: dout  = 8'b00000000; //   53 :   0 - 0x0
      11'h36: dout  = 8'b00000000; //   54 :   0 - 0x0
      11'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      11'h38: dout  = 8'b00000000; //   56 :   0 - 0x0 -- Background 0x7
      11'h39: dout  = 8'b00000000; //   57 :   0 - 0x0
      11'h3A: dout  = 8'b00000000; //   58 :   0 - 0x0
      11'h3B: dout  = 8'b00000000; //   59 :   0 - 0x0
      11'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      11'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      11'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      11'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      11'h40: dout  = 8'b00000000; //   64 :   0 - 0x0 -- Background 0x8
      11'h41: dout  = 8'b00000000; //   65 :   0 - 0x0
      11'h42: dout  = 8'b00000000; //   66 :   0 - 0x0
      11'h43: dout  = 8'b00000000; //   67 :   0 - 0x0
      11'h44: dout  = 8'b00000000; //   68 :   0 - 0x0
      11'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      11'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      11'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      11'h48: dout  = 8'b00000000; //   72 :   0 - 0x0 -- Background 0x9
      11'h49: dout  = 8'b00000000; //   73 :   0 - 0x0
      11'h4A: dout  = 8'b00000000; //   74 :   0 - 0x0
      11'h4B: dout  = 8'b00000000; //   75 :   0 - 0x0
      11'h4C: dout  = 8'b00000000; //   76 :   0 - 0x0
      11'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      11'h4E: dout  = 8'b00000000; //   78 :   0 - 0x0
      11'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      11'h50: dout  = 8'b00000000; //   80 :   0 - 0x0 -- Background 0xa
      11'h51: dout  = 8'b00000000; //   81 :   0 - 0x0
      11'h52: dout  = 8'b00000000; //   82 :   0 - 0x0
      11'h53: dout  = 8'b00000000; //   83 :   0 - 0x0
      11'h54: dout  = 8'b00000000; //   84 :   0 - 0x0
      11'h55: dout  = 8'b00000000; //   85 :   0 - 0x0
      11'h56: dout  = 8'b00000000; //   86 :   0 - 0x0
      11'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      11'h58: dout  = 8'b00000000; //   88 :   0 - 0x0 -- Background 0xb
      11'h59: dout  = 8'b00000000; //   89 :   0 - 0x0
      11'h5A: dout  = 8'b00000000; //   90 :   0 - 0x0
      11'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      11'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      11'h5D: dout  = 8'b00000000; //   93 :   0 - 0x0
      11'h5E: dout  = 8'b00000000; //   94 :   0 - 0x0
      11'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      11'h60: dout  = 8'b00000000; //   96 :   0 - 0x0 -- Background 0xc
      11'h61: dout  = 8'b00000000; //   97 :   0 - 0x0
      11'h62: dout  = 8'b00000000; //   98 :   0 - 0x0
      11'h63: dout  = 8'b00000000; //   99 :   0 - 0x0
      11'h64: dout  = 8'b00000000; //  100 :   0 - 0x0
      11'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      11'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      11'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      11'h68: dout  = 8'b00000000; //  104 :   0 - 0x0 -- Background 0xd
      11'h69: dout  = 8'b00000000; //  105 :   0 - 0x0
      11'h6A: dout  = 8'b00000000; //  106 :   0 - 0x0
      11'h6B: dout  = 8'b00000000; //  107 :   0 - 0x0
      11'h6C: dout  = 8'b00000000; //  108 :   0 - 0x0
      11'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      11'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      11'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      11'h70: dout  = 8'b00000000; //  112 :   0 - 0x0 -- Background 0xe
      11'h71: dout  = 8'b00000000; //  113 :   0 - 0x0
      11'h72: dout  = 8'b00000000; //  114 :   0 - 0x0
      11'h73: dout  = 8'b00000000; //  115 :   0 - 0x0
      11'h74: dout  = 8'b00000000; //  116 :   0 - 0x0
      11'h75: dout  = 8'b00000000; //  117 :   0 - 0x0
      11'h76: dout  = 8'b00000000; //  118 :   0 - 0x0
      11'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      11'h78: dout  = 8'b00000000; //  120 :   0 - 0x0 -- Background 0xf
      11'h79: dout  = 8'b00000000; //  121 :   0 - 0x0
      11'h7A: dout  = 8'b00000000; //  122 :   0 - 0x0
      11'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      11'h7C: dout  = 8'b00000000; //  124 :   0 - 0x0
      11'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      11'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      11'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      11'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Background 0x10
      11'h81: dout  = 8'b00000000; //  129 :   0 - 0x0
      11'h82: dout  = 8'b00000000; //  130 :   0 - 0x0
      11'h83: dout  = 8'b00000000; //  131 :   0 - 0x0
      11'h84: dout  = 8'b00000000; //  132 :   0 - 0x0
      11'h85: dout  = 8'b00000000; //  133 :   0 - 0x0
      11'h86: dout  = 8'b00000000; //  134 :   0 - 0x0
      11'h87: dout  = 8'b00000000; //  135 :   0 - 0x0
      11'h88: dout  = 8'b00000000; //  136 :   0 - 0x0 -- Background 0x11
      11'h89: dout  = 8'b00000000; //  137 :   0 - 0x0
      11'h8A: dout  = 8'b00000000; //  138 :   0 - 0x0
      11'h8B: dout  = 8'b00000000; //  139 :   0 - 0x0
      11'h8C: dout  = 8'b00000000; //  140 :   0 - 0x0
      11'h8D: dout  = 8'b00000000; //  141 :   0 - 0x0
      11'h8E: dout  = 8'b00000000; //  142 :   0 - 0x0
      11'h8F: dout  = 8'b00000000; //  143 :   0 - 0x0
      11'h90: dout  = 8'b00000000; //  144 :   0 - 0x0 -- Background 0x12
      11'h91: dout  = 8'b00000000; //  145 :   0 - 0x0
      11'h92: dout  = 8'b00000000; //  146 :   0 - 0x0
      11'h93: dout  = 8'b00000000; //  147 :   0 - 0x0
      11'h94: dout  = 8'b00000000; //  148 :   0 - 0x0
      11'h95: dout  = 8'b00000000; //  149 :   0 - 0x0
      11'h96: dout  = 8'b00000000; //  150 :   0 - 0x0
      11'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      11'h98: dout  = 8'b00000000; //  152 :   0 - 0x0 -- Background 0x13
      11'h99: dout  = 8'b00000000; //  153 :   0 - 0x0
      11'h9A: dout  = 8'b00000000; //  154 :   0 - 0x0
      11'h9B: dout  = 8'b00000000; //  155 :   0 - 0x0
      11'h9C: dout  = 8'b00000000; //  156 :   0 - 0x0
      11'h9D: dout  = 8'b00000000; //  157 :   0 - 0x0
      11'h9E: dout  = 8'b00000000; //  158 :   0 - 0x0
      11'h9F: dout  = 8'b00000000; //  159 :   0 - 0x0
      11'hA0: dout  = 8'b00000000; //  160 :   0 - 0x0 -- Background 0x14
      11'hA1: dout  = 8'b00000000; //  161 :   0 - 0x0
      11'hA2: dout  = 8'b00000000; //  162 :   0 - 0x0
      11'hA3: dout  = 8'b00000000; //  163 :   0 - 0x0
      11'hA4: dout  = 8'b00000000; //  164 :   0 - 0x0
      11'hA5: dout  = 8'b00000000; //  165 :   0 - 0x0
      11'hA6: dout  = 8'b00000000; //  166 :   0 - 0x0
      11'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      11'hA8: dout  = 8'b00000000; //  168 :   0 - 0x0 -- Background 0x15
      11'hA9: dout  = 8'b00000000; //  169 :   0 - 0x0
      11'hAA: dout  = 8'b00000000; //  170 :   0 - 0x0
      11'hAB: dout  = 8'b00000000; //  171 :   0 - 0x0
      11'hAC: dout  = 8'b00000000; //  172 :   0 - 0x0
      11'hAD: dout  = 8'b00000000; //  173 :   0 - 0x0
      11'hAE: dout  = 8'b00000000; //  174 :   0 - 0x0
      11'hAF: dout  = 8'b00000000; //  175 :   0 - 0x0
      11'hB0: dout  = 8'b00000000; //  176 :   0 - 0x0 -- Background 0x16
      11'hB1: dout  = 8'b00000000; //  177 :   0 - 0x0
      11'hB2: dout  = 8'b00000000; //  178 :   0 - 0x0
      11'hB3: dout  = 8'b00000000; //  179 :   0 - 0x0
      11'hB4: dout  = 8'b00000000; //  180 :   0 - 0x0
      11'hB5: dout  = 8'b00000000; //  181 :   0 - 0x0
      11'hB6: dout  = 8'b00000000; //  182 :   0 - 0x0
      11'hB7: dout  = 8'b00000000; //  183 :   0 - 0x0
      11'hB8: dout  = 8'b00000000; //  184 :   0 - 0x0 -- Background 0x17
      11'hB9: dout  = 8'b00000000; //  185 :   0 - 0x0
      11'hBA: dout  = 8'b00000000; //  186 :   0 - 0x0
      11'hBB: dout  = 8'b00000000; //  187 :   0 - 0x0
      11'hBC: dout  = 8'b00000000; //  188 :   0 - 0x0
      11'hBD: dout  = 8'b00000000; //  189 :   0 - 0x0
      11'hBE: dout  = 8'b00000000; //  190 :   0 - 0x0
      11'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      11'hC0: dout  = 8'b00000000; //  192 :   0 - 0x0 -- Background 0x18
      11'hC1: dout  = 8'b00000000; //  193 :   0 - 0x0
      11'hC2: dout  = 8'b00000000; //  194 :   0 - 0x0
      11'hC3: dout  = 8'b00000000; //  195 :   0 - 0x0
      11'hC4: dout  = 8'b00000000; //  196 :   0 - 0x0
      11'hC5: dout  = 8'b00000000; //  197 :   0 - 0x0
      11'hC6: dout  = 8'b00000000; //  198 :   0 - 0x0
      11'hC7: dout  = 8'b00000000; //  199 :   0 - 0x0
      11'hC8: dout  = 8'b00000000; //  200 :   0 - 0x0 -- Background 0x19
      11'hC9: dout  = 8'b00000000; //  201 :   0 - 0x0
      11'hCA: dout  = 8'b00000000; //  202 :   0 - 0x0
      11'hCB: dout  = 8'b00000000; //  203 :   0 - 0x0
      11'hCC: dout  = 8'b00000000; //  204 :   0 - 0x0
      11'hCD: dout  = 8'b00000000; //  205 :   0 - 0x0
      11'hCE: dout  = 8'b00000000; //  206 :   0 - 0x0
      11'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      11'hD0: dout  = 8'b00000000; //  208 :   0 - 0x0 -- Background 0x1a
      11'hD1: dout  = 8'b00000000; //  209 :   0 - 0x0
      11'hD2: dout  = 8'b00000000; //  210 :   0 - 0x0
      11'hD3: dout  = 8'b00000000; //  211 :   0 - 0x0
      11'hD4: dout  = 8'b00000000; //  212 :   0 - 0x0
      11'hD5: dout  = 8'b00000000; //  213 :   0 - 0x0
      11'hD6: dout  = 8'b00000000; //  214 :   0 - 0x0
      11'hD7: dout  = 8'b00000000; //  215 :   0 - 0x0
      11'hD8: dout  = 8'b00000000; //  216 :   0 - 0x0 -- Background 0x1b
      11'hD9: dout  = 8'b00000000; //  217 :   0 - 0x0
      11'hDA: dout  = 8'b00000000; //  218 :   0 - 0x0
      11'hDB: dout  = 8'b00000000; //  219 :   0 - 0x0
      11'hDC: dout  = 8'b00000000; //  220 :   0 - 0x0
      11'hDD: dout  = 8'b00000000; //  221 :   0 - 0x0
      11'hDE: dout  = 8'b00000000; //  222 :   0 - 0x0
      11'hDF: dout  = 8'b00000000; //  223 :   0 - 0x0
      11'hE0: dout  = 8'b00000000; //  224 :   0 - 0x0 -- Background 0x1c
      11'hE1: dout  = 8'b00000000; //  225 :   0 - 0x0
      11'hE2: dout  = 8'b00000000; //  226 :   0 - 0x0
      11'hE3: dout  = 8'b00000000; //  227 :   0 - 0x0
      11'hE4: dout  = 8'b00000000; //  228 :   0 - 0x0
      11'hE5: dout  = 8'b00000000; //  229 :   0 - 0x0
      11'hE6: dout  = 8'b00000000; //  230 :   0 - 0x0
      11'hE7: dout  = 8'b00000000; //  231 :   0 - 0x0
      11'hE8: dout  = 8'b00000000; //  232 :   0 - 0x0 -- Background 0x1d
      11'hE9: dout  = 8'b00000000; //  233 :   0 - 0x0
      11'hEA: dout  = 8'b00000000; //  234 :   0 - 0x0
      11'hEB: dout  = 8'b00000000; //  235 :   0 - 0x0
      11'hEC: dout  = 8'b00000000; //  236 :   0 - 0x0
      11'hED: dout  = 8'b00000000; //  237 :   0 - 0x0
      11'hEE: dout  = 8'b00000000; //  238 :   0 - 0x0
      11'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      11'hF0: dout  = 8'b00000000; //  240 :   0 - 0x0 -- Background 0x1e
      11'hF1: dout  = 8'b00000000; //  241 :   0 - 0x0
      11'hF2: dout  = 8'b00000000; //  242 :   0 - 0x0
      11'hF3: dout  = 8'b00000000; //  243 :   0 - 0x0
      11'hF4: dout  = 8'b00000000; //  244 :   0 - 0x0
      11'hF5: dout  = 8'b00000000; //  245 :   0 - 0x0
      11'hF6: dout  = 8'b00000000; //  246 :   0 - 0x0
      11'hF7: dout  = 8'b00000000; //  247 :   0 - 0x0
      11'hF8: dout  = 8'b00000000; //  248 :   0 - 0x0 -- Background 0x1f
      11'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      11'hFA: dout  = 8'b00000000; //  250 :   0 - 0x0
      11'hFB: dout  = 8'b00000000; //  251 :   0 - 0x0
      11'hFC: dout  = 8'b00000000; //  252 :   0 - 0x0
      11'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      11'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      11'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Background 0x20
      11'h101: dout  = 8'b00000000; //  257 :   0 - 0x0
      11'h102: dout  = 8'b00000000; //  258 :   0 - 0x0
      11'h103: dout  = 8'b00000000; //  259 :   0 - 0x0
      11'h104: dout  = 8'b00000000; //  260 :   0 - 0x0
      11'h105: dout  = 8'b00000000; //  261 :   0 - 0x0
      11'h106: dout  = 8'b00000000; //  262 :   0 - 0x0
      11'h107: dout  = 8'b00000000; //  263 :   0 - 0x0
      11'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- Background 0x21
      11'h109: dout  = 8'b00000000; //  265 :   0 - 0x0
      11'h10A: dout  = 8'b00000000; //  266 :   0 - 0x0
      11'h10B: dout  = 8'b00000000; //  267 :   0 - 0x0
      11'h10C: dout  = 8'b00000000; //  268 :   0 - 0x0
      11'h10D: dout  = 8'b00000000; //  269 :   0 - 0x0
      11'h10E: dout  = 8'b00000000; //  270 :   0 - 0x0
      11'h10F: dout  = 8'b00000000; //  271 :   0 - 0x0
      11'h110: dout  = 8'b00000000; //  272 :   0 - 0x0 -- Background 0x22
      11'h111: dout  = 8'b00000000; //  273 :   0 - 0x0
      11'h112: dout  = 8'b00000000; //  274 :   0 - 0x0
      11'h113: dout  = 8'b00000000; //  275 :   0 - 0x0
      11'h114: dout  = 8'b00000000; //  276 :   0 - 0x0
      11'h115: dout  = 8'b00000000; //  277 :   0 - 0x0
      11'h116: dout  = 8'b00000000; //  278 :   0 - 0x0
      11'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      11'h118: dout  = 8'b00000000; //  280 :   0 - 0x0 -- Background 0x23
      11'h119: dout  = 8'b00000000; //  281 :   0 - 0x0
      11'h11A: dout  = 8'b00000000; //  282 :   0 - 0x0
      11'h11B: dout  = 8'b00000000; //  283 :   0 - 0x0
      11'h11C: dout  = 8'b00000000; //  284 :   0 - 0x0
      11'h11D: dout  = 8'b00000000; //  285 :   0 - 0x0
      11'h11E: dout  = 8'b00000000; //  286 :   0 - 0x0
      11'h11F: dout  = 8'b00000000; //  287 :   0 - 0x0
      11'h120: dout  = 8'b00000000; //  288 :   0 - 0x0 -- Background 0x24
      11'h121: dout  = 8'b00000000; //  289 :   0 - 0x0
      11'h122: dout  = 8'b00000000; //  290 :   0 - 0x0
      11'h123: dout  = 8'b00000000; //  291 :   0 - 0x0
      11'h124: dout  = 8'b00000000; //  292 :   0 - 0x0
      11'h125: dout  = 8'b00000000; //  293 :   0 - 0x0
      11'h126: dout  = 8'b00000000; //  294 :   0 - 0x0
      11'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      11'h128: dout  = 8'b00000000; //  296 :   0 - 0x0 -- Background 0x25
      11'h129: dout  = 8'b00000000; //  297 :   0 - 0x0
      11'h12A: dout  = 8'b00000000; //  298 :   0 - 0x0
      11'h12B: dout  = 8'b00000000; //  299 :   0 - 0x0
      11'h12C: dout  = 8'b00000000; //  300 :   0 - 0x0
      11'h12D: dout  = 8'b00000000; //  301 :   0 - 0x0
      11'h12E: dout  = 8'b00000000; //  302 :   0 - 0x0
      11'h12F: dout  = 8'b00000000; //  303 :   0 - 0x0
      11'h130: dout  = 8'b11111111; //  304 : 255 - 0xff -- Background 0x26
      11'h131: dout  = 8'b11111111; //  305 : 255 - 0xff
      11'h132: dout  = 8'b11111111; //  306 : 255 - 0xff
      11'h133: dout  = 8'b11111111; //  307 : 255 - 0xff
      11'h134: dout  = 8'b11111111; //  308 : 255 - 0xff
      11'h135: dout  = 8'b11111111; //  309 : 255 - 0xff
      11'h136: dout  = 8'b11111111; //  310 : 255 - 0xff
      11'h137: dout  = 8'b11111111; //  311 : 255 - 0xff
      11'h138: dout  = 8'b11111111; //  312 : 255 - 0xff -- Background 0x27
      11'h139: dout  = 8'b11111111; //  313 : 255 - 0xff
      11'h13A: dout  = 8'b11111111; //  314 : 255 - 0xff
      11'h13B: dout  = 8'b11111111; //  315 : 255 - 0xff
      11'h13C: dout  = 8'b11111111; //  316 : 255 - 0xff
      11'h13D: dout  = 8'b11111111; //  317 : 255 - 0xff
      11'h13E: dout  = 8'b11111111; //  318 : 255 - 0xff
      11'h13F: dout  = 8'b11111111; //  319 : 255 - 0xff
      11'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Background 0x28
      11'h141: dout  = 8'b00000000; //  321 :   0 - 0x0
      11'h142: dout  = 8'b00000000; //  322 :   0 - 0x0
      11'h143: dout  = 8'b00000000; //  323 :   0 - 0x0
      11'h144: dout  = 8'b00000000; //  324 :   0 - 0x0
      11'h145: dout  = 8'b00000000; //  325 :   0 - 0x0
      11'h146: dout  = 8'b00000000; //  326 :   0 - 0x0
      11'h147: dout  = 8'b00000000; //  327 :   0 - 0x0
      11'h148: dout  = 8'b00000000; //  328 :   0 - 0x0 -- Background 0x29
      11'h149: dout  = 8'b00000000; //  329 :   0 - 0x0
      11'h14A: dout  = 8'b00000000; //  330 :   0 - 0x0
      11'h14B: dout  = 8'b00000000; //  331 :   0 - 0x0
      11'h14C: dout  = 8'b00000000; //  332 :   0 - 0x0
      11'h14D: dout  = 8'b00000000; //  333 :   0 - 0x0
      11'h14E: dout  = 8'b00000000; //  334 :   0 - 0x0
      11'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      11'h150: dout  = 8'b01111111; //  336 : 127 - 0x7f -- Background 0x2a
      11'h151: dout  = 8'b01111111; //  337 : 127 - 0x7f
      11'h152: dout  = 8'b01111111; //  338 : 127 - 0x7f
      11'h153: dout  = 8'b01111111; //  339 : 127 - 0x7f
      11'h154: dout  = 8'b01111111; //  340 : 127 - 0x7f
      11'h155: dout  = 8'b01111111; //  341 : 127 - 0x7f
      11'h156: dout  = 8'b01111111; //  342 : 127 - 0x7f
      11'h157: dout  = 8'b01111111; //  343 : 127 - 0x7f
      11'h158: dout  = 8'b00000000; //  344 :   0 - 0x0 -- Background 0x2b
      11'h159: dout  = 8'b00000000; //  345 :   0 - 0x0
      11'h15A: dout  = 8'b00000000; //  346 :   0 - 0x0
      11'h15B: dout  = 8'b00000000; //  347 :   0 - 0x0
      11'h15C: dout  = 8'b00000000; //  348 :   0 - 0x0
      11'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      11'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      11'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      11'h160: dout  = 8'b11111111; //  352 : 255 - 0xff -- Background 0x2c
      11'h161: dout  = 8'b10000000; //  353 : 128 - 0x80
      11'h162: dout  = 8'b10000000; //  354 : 128 - 0x80
      11'h163: dout  = 8'b10000000; //  355 : 128 - 0x80
      11'h164: dout  = 8'b10000000; //  356 : 128 - 0x80
      11'h165: dout  = 8'b00000000; //  357 :   0 - 0x0
      11'h166: dout  = 8'b00011100; //  358 :  28 - 0x1c
      11'h167: dout  = 8'b00111110; //  359 :  62 - 0x3e
      11'h168: dout  = 8'b01111111; //  360 : 127 - 0x7f -- Background 0x2d
      11'h169: dout  = 8'b01111111; //  361 : 127 - 0x7f
      11'h16A: dout  = 8'b01111111; //  362 : 127 - 0x7f
      11'h16B: dout  = 8'b00111110; //  363 :  62 - 0x3e
      11'h16C: dout  = 8'b00011100; //  364 :  28 - 0x1c
      11'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      11'h16E: dout  = 8'b00000000; //  366 :   0 - 0x0
      11'h16F: dout  = 8'b11111111; //  367 : 255 - 0xff
      11'h170: dout  = 8'b00001000; //  368 :   8 - 0x8 -- Background 0x2e
      11'h171: dout  = 8'b00000100; //  369 :   4 - 0x4
      11'h172: dout  = 8'b00000100; //  370 :   4 - 0x4
      11'h173: dout  = 8'b00000100; //  371 :   4 - 0x4
      11'h174: dout  = 8'b00000100; //  372 :   4 - 0x4
      11'h175: dout  = 8'b00000100; //  373 :   4 - 0x4
      11'h176: dout  = 8'b00001000; //  374 :   8 - 0x8
      11'h177: dout  = 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout  = 8'b00000011; //  376 :   3 - 0x3 -- Background 0x2f
      11'h179: dout  = 8'b00000101; //  377 :   5 - 0x5
      11'h17A: dout  = 8'b00001011; //  378 :  11 - 0xb
      11'h17B: dout  = 8'b00001011; //  379 :  11 - 0xb
      11'h17C: dout  = 8'b00001111; //  380 :  15 - 0xf
      11'h17D: dout  = 8'b00001111; //  381 :  15 - 0xf
      11'h17E: dout  = 8'b00000111; //  382 :   7 - 0x7
      11'h17F: dout  = 8'b00000011; //  383 :   3 - 0x3
      11'h180: dout  = 8'b00000001; //  384 :   1 - 0x1 -- Background 0x30
      11'h181: dout  = 8'b00000011; //  385 :   3 - 0x3
      11'h182: dout  = 8'b00000111; //  386 :   7 - 0x7
      11'h183: dout  = 8'b00001111; //  387 :  15 - 0xf
      11'h184: dout  = 8'b00011111; //  388 :  31 - 0x1f
      11'h185: dout  = 8'b00111111; //  389 :  63 - 0x3f
      11'h186: dout  = 8'b01111111; //  390 : 127 - 0x7f
      11'h187: dout  = 8'b11111111; //  391 : 255 - 0xff
      11'h188: dout  = 8'b00000000; //  392 :   0 - 0x0 -- Background 0x31
      11'h189: dout  = 8'b00000000; //  393 :   0 - 0x0
      11'h18A: dout  = 8'b00000000; //  394 :   0 - 0x0
      11'h18B: dout  = 8'b00000000; //  395 :   0 - 0x0
      11'h18C: dout  = 8'b00000000; //  396 :   0 - 0x0
      11'h18D: dout  = 8'b00000111; //  397 :   7 - 0x7
      11'h18E: dout  = 8'b00111111; //  398 :  63 - 0x3f
      11'h18F: dout  = 8'b11111111; //  399 : 255 - 0xff
      11'h190: dout  = 8'b00000000; //  400 :   0 - 0x0 -- Background 0x32
      11'h191: dout  = 8'b00000000; //  401 :   0 - 0x0
      11'h192: dout  = 8'b00000000; //  402 :   0 - 0x0
      11'h193: dout  = 8'b00000000; //  403 :   0 - 0x0
      11'h194: dout  = 8'b00000000; //  404 :   0 - 0x0
      11'h195: dout  = 8'b11100000; //  405 : 224 - 0xe0
      11'h196: dout  = 8'b11111100; //  406 : 252 - 0xfc
      11'h197: dout  = 8'b11111111; //  407 : 255 - 0xff
      11'h198: dout  = 8'b10000000; //  408 : 128 - 0x80 -- Background 0x33
      11'h199: dout  = 8'b11000000; //  409 : 192 - 0xc0
      11'h19A: dout  = 8'b11100000; //  410 : 224 - 0xe0
      11'h19B: dout  = 8'b11110000; //  411 : 240 - 0xf0
      11'h19C: dout  = 8'b11111000; //  412 : 248 - 0xf8
      11'h19D: dout  = 8'b11111100; //  413 : 252 - 0xfc
      11'h19E: dout  = 8'b11111110; //  414 : 254 - 0xfe
      11'h19F: dout  = 8'b11111111; //  415 : 255 - 0xff
      11'h1A0: dout  = 8'b11111111; //  416 : 255 - 0xff -- Background 0x34
      11'h1A1: dout  = 8'b11111111; //  417 : 255 - 0xff
      11'h1A2: dout  = 8'b11111111; //  418 : 255 - 0xff
      11'h1A3: dout  = 8'b11111111; //  419 : 255 - 0xff
      11'h1A4: dout  = 8'b11111111; //  420 : 255 - 0xff
      11'h1A5: dout  = 8'b11111111; //  421 : 255 - 0xff
      11'h1A6: dout  = 8'b11111111; //  422 : 255 - 0xff
      11'h1A7: dout  = 8'b11111111; //  423 : 255 - 0xff
      11'h1A8: dout  = 8'b00000111; //  424 :   7 - 0x7 -- Background 0x35
      11'h1A9: dout  = 8'b00001000; //  425 :   8 - 0x8
      11'h1AA: dout  = 8'b00010000; //  426 :  16 - 0x10
      11'h1AB: dout  = 8'b00000000; //  427 :   0 - 0x0
      11'h1AC: dout  = 8'b01100000; //  428 :  96 - 0x60
      11'h1AD: dout  = 8'b10000000; //  429 : 128 - 0x80
      11'h1AE: dout  = 8'b10000000; //  430 : 128 - 0x80
      11'h1AF: dout  = 8'b01000000; //  431 :  64 - 0x40
      11'h1B0: dout  = 8'b00000011; //  432 :   3 - 0x3 -- Background 0x36
      11'h1B1: dout  = 8'b00000100; //  433 :   4 - 0x4
      11'h1B2: dout  = 8'b00011000; //  434 :  24 - 0x18
      11'h1B3: dout  = 8'b00100000; //  435 :  32 - 0x20
      11'h1B4: dout  = 8'b00100000; //  436 :  32 - 0x20
      11'h1B5: dout  = 8'b00100000; //  437 :  32 - 0x20
      11'h1B6: dout  = 8'b01000110; //  438 :  70 - 0x46
      11'h1B7: dout  = 8'b10001000; //  439 : 136 - 0x88
      11'h1B8: dout  = 8'b11000000; //  440 : 192 - 0xc0 -- Background 0x37
      11'h1B9: dout  = 8'b00100000; //  441 :  32 - 0x20
      11'h1BA: dout  = 8'b00010000; //  442 :  16 - 0x10
      11'h1BB: dout  = 8'b00010100; //  443 :  20 - 0x14
      11'h1BC: dout  = 8'b00001010; //  444 :  10 - 0xa
      11'h1BD: dout  = 8'b01000001; //  445 :  65 - 0x41
      11'h1BE: dout  = 8'b00100001; //  446 :  33 - 0x21
      11'h1BF: dout  = 8'b00000001; //  447 :   1 - 0x1
      11'h1C0: dout  = 8'b10010000; //  448 : 144 - 0x90 -- Background 0x38
      11'h1C1: dout  = 8'b10101000; //  449 : 168 - 0xa8
      11'h1C2: dout  = 8'b01001000; //  450 :  72 - 0x48
      11'h1C3: dout  = 8'b00001010; //  451 :  10 - 0xa
      11'h1C4: dout  = 8'b00000101; //  452 :   5 - 0x5
      11'h1C5: dout  = 8'b00000001; //  453 :   1 - 0x1
      11'h1C6: dout  = 8'b00000001; //  454 :   1 - 0x1
      11'h1C7: dout  = 8'b00000010; //  455 :   2 - 0x2
      11'h1C8: dout  = 8'b00100100; //  456 :  36 - 0x24 -- Background 0x39
      11'h1C9: dout  = 8'b00010010; //  457 :  18 - 0x12
      11'h1CA: dout  = 8'b00001001; //  458 :   9 - 0x9
      11'h1CB: dout  = 8'b00001000; //  459 :   8 - 0x8
      11'h1CC: dout  = 8'b00000111; //  460 :   7 - 0x7
      11'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Background 0x3a
      11'h1D1: dout  = 8'b01000000; //  465 :  64 - 0x40
      11'h1D2: dout  = 8'b11100011; //  466 : 227 - 0xe3
      11'h1D3: dout  = 8'b00111111; //  467 :  63 - 0x3f
      11'h1D4: dout  = 8'b00001100; //  468 :  12 - 0xc
      11'h1D5: dout  = 8'b10000001; //  469 : 129 - 0x81
      11'h1D6: dout  = 8'b01100010; //  470 :  98 - 0x62
      11'h1D7: dout  = 8'b00011100; //  471 :  28 - 0x1c
      11'h1D8: dout  = 8'b01000000; //  472 :  64 - 0x40 -- Background 0x3b
      11'h1D9: dout  = 8'b10000000; //  473 : 128 - 0x80
      11'h1DA: dout  = 8'b11000010; //  474 : 194 - 0xc2
      11'h1DB: dout  = 8'b01111100; //  475 : 124 - 0x7c
      11'h1DC: dout  = 8'b00111000; //  476 :  56 - 0x38
      11'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      11'h1DE: dout  = 8'b11000011; //  478 : 195 - 0xc3
      11'h1DF: dout  = 8'b00111100; //  479 :  60 - 0x3c
      11'h1E0: dout  = 8'b00000100; //  480 :   4 - 0x4 -- Background 0x3c
      11'h1E1: dout  = 8'b00000010; //  481 :   2 - 0x2
      11'h1E2: dout  = 8'b00000001; //  482 :   1 - 0x1
      11'h1E3: dout  = 8'b00000000; //  483 :   0 - 0x0
      11'h1E4: dout  = 8'b00000110; //  484 :   6 - 0x6
      11'h1E5: dout  = 8'b10011000; //  485 : 152 - 0x98
      11'h1E6: dout  = 8'b01100000; //  486 :  96 - 0x60
      11'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout  = 8'b11000000; //  488 : 192 - 0xc0 -- Background 0x3d
      11'h1E9: dout  = 8'b11100000; //  489 : 224 - 0xe0
      11'h1EA: dout  = 8'b11110000; //  490 : 240 - 0xf0
      11'h1EB: dout  = 8'b11110000; //  491 : 240 - 0xf0
      11'h1EC: dout  = 8'b11110000; //  492 : 240 - 0xf0
      11'h1ED: dout  = 8'b11110000; //  493 : 240 - 0xf0
      11'h1EE: dout  = 8'b11100000; //  494 : 224 - 0xe0
      11'h1EF: dout  = 8'b11000000; //  495 : 192 - 0xc0
      11'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Background 0x3e
      11'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      11'h1F2: dout  = 8'b00000000; //  498 :   0 - 0x0
      11'h1F3: dout  = 8'b00000000; //  499 :   0 - 0x0
      11'h1F4: dout  = 8'b00000000; //  500 :   0 - 0x0
      11'h1F5: dout  = 8'b00000000; //  501 :   0 - 0x0
      11'h1F6: dout  = 8'b00011100; //  502 :  28 - 0x1c
      11'h1F7: dout  = 8'b00111110; //  503 :  62 - 0x3e
      11'h1F8: dout  = 8'b01111111; //  504 : 127 - 0x7f -- Background 0x3f
      11'h1F9: dout  = 8'b01111111; //  505 : 127 - 0x7f
      11'h1FA: dout  = 8'b01111111; //  506 : 127 - 0x7f
      11'h1FB: dout  = 8'b00111110; //  507 :  62 - 0x3e
      11'h1FC: dout  = 8'b00011100; //  508 :  28 - 0x1c
      11'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      11'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      11'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      11'h200: dout  = 8'b11111111; //  512 : 255 - 0xff -- Background 0x40
      11'h201: dout  = 8'b11111111; //  513 : 255 - 0xff
      11'h202: dout  = 8'b11111111; //  514 : 255 - 0xff
      11'h203: dout  = 8'b11111111; //  515 : 255 - 0xff
      11'h204: dout  = 8'b11111111; //  516 : 255 - 0xff
      11'h205: dout  = 8'b11111111; //  517 : 255 - 0xff
      11'h206: dout  = 8'b11111111; //  518 : 255 - 0xff
      11'h207: dout  = 8'b11111111; //  519 : 255 - 0xff
      11'h208: dout  = 8'b00000000; //  520 :   0 - 0x0 -- Background 0x41
      11'h209: dout  = 8'b00001000; //  521 :   8 - 0x8
      11'h20A: dout  = 8'b00011000; //  522 :  24 - 0x18
      11'h20B: dout  = 8'b00111000; //  523 :  56 - 0x38
      11'h20C: dout  = 8'b11111100; //  524 : 252 - 0xfc
      11'h20D: dout  = 8'b10111111; //  525 : 191 - 0xbf
      11'h20E: dout  = 8'b01011110; //  526 :  94 - 0x5e
      11'h20F: dout  = 8'b11011001; //  527 : 217 - 0xd9
      11'h210: dout  = 8'b10000001; //  528 : 129 - 0x81 -- Background 0x42
      11'h211: dout  = 8'b10000001; //  529 : 129 - 0x81
      11'h212: dout  = 8'b10000001; //  530 : 129 - 0x81
      11'h213: dout  = 8'b10000001; //  531 : 129 - 0x81
      11'h214: dout  = 8'b10000001; //  532 : 129 - 0x81
      11'h215: dout  = 8'b10000001; //  533 : 129 - 0x81
      11'h216: dout  = 8'b10000001; //  534 : 129 - 0x81
      11'h217: dout  = 8'b10000001; //  535 : 129 - 0x81
      11'h218: dout  = 8'b00000001; //  536 :   1 - 0x1 -- Background 0x43
      11'h219: dout  = 8'b00000001; //  537 :   1 - 0x1
      11'h21A: dout  = 8'b00000001; //  538 :   1 - 0x1
      11'h21B: dout  = 8'b00000001; //  539 :   1 - 0x1
      11'h21C: dout  = 8'b00000001; //  540 :   1 - 0x1
      11'h21D: dout  = 8'b00000001; //  541 :   1 - 0x1
      11'h21E: dout  = 8'b00000001; //  542 :   1 - 0x1
      11'h21F: dout  = 8'b00000001; //  543 :   1 - 0x1
      11'h220: dout  = 8'b00000000; //  544 :   0 - 0x0 -- Background 0x44
      11'h221: dout  = 8'b01111111; //  545 : 127 - 0x7f
      11'h222: dout  = 8'b01111111; //  546 : 127 - 0x7f
      11'h223: dout  = 8'b01100111; //  547 : 103 - 0x67
      11'h224: dout  = 8'b01100111; //  548 : 103 - 0x67
      11'h225: dout  = 8'b01111111; //  549 : 127 - 0x7f
      11'h226: dout  = 8'b01111111; //  550 : 127 - 0x7f
      11'h227: dout  = 8'b01111111; //  551 : 127 - 0x7f
      11'h228: dout  = 8'b00000000; //  552 :   0 - 0x0 -- Background 0x45
      11'h229: dout  = 8'b11111111; //  553 : 255 - 0xff
      11'h22A: dout  = 8'b11111111; //  554 : 255 - 0xff
      11'h22B: dout  = 8'b11111111; //  555 : 255 - 0xff
      11'h22C: dout  = 8'b11111111; //  556 : 255 - 0xff
      11'h22D: dout  = 8'b11111111; //  557 : 255 - 0xff
      11'h22E: dout  = 8'b11111111; //  558 : 255 - 0xff
      11'h22F: dout  = 8'b11111111; //  559 : 255 - 0xff
      11'h230: dout  = 8'b01111111; //  560 : 127 - 0x7f -- Background 0x46
      11'h231: dout  = 8'b01111111; //  561 : 127 - 0x7f
      11'h232: dout  = 8'b01111111; //  562 : 127 - 0x7f
      11'h233: dout  = 8'b01111111; //  563 : 127 - 0x7f
      11'h234: dout  = 8'b01111111; //  564 : 127 - 0x7f
      11'h235: dout  = 8'b01111111; //  565 : 127 - 0x7f
      11'h236: dout  = 8'b01111111; //  566 : 127 - 0x7f
      11'h237: dout  = 8'b01111111; //  567 : 127 - 0x7f
      11'h238: dout  = 8'b11111111; //  568 : 255 - 0xff -- Background 0x47
      11'h239: dout  = 8'b11111111; //  569 : 255 - 0xff
      11'h23A: dout  = 8'b11111111; //  570 : 255 - 0xff
      11'h23B: dout  = 8'b11111111; //  571 : 255 - 0xff
      11'h23C: dout  = 8'b11111111; //  572 : 255 - 0xff
      11'h23D: dout  = 8'b11111111; //  573 : 255 - 0xff
      11'h23E: dout  = 8'b11111111; //  574 : 255 - 0xff
      11'h23F: dout  = 8'b11111111; //  575 : 255 - 0xff
      11'h240: dout  = 8'b00000000; //  576 :   0 - 0x0 -- Background 0x48
      11'h241: dout  = 8'b11111111; //  577 : 255 - 0xff
      11'h242: dout  = 8'b11111111; //  578 : 255 - 0xff
      11'h243: dout  = 8'b11111111; //  579 : 255 - 0xff
      11'h244: dout  = 8'b11111111; //  580 : 255 - 0xff
      11'h245: dout  = 8'b11111111; //  581 : 255 - 0xff
      11'h246: dout  = 8'b11111111; //  582 : 255 - 0xff
      11'h247: dout  = 8'b11111111; //  583 : 255 - 0xff
      11'h248: dout  = 8'b00000000; //  584 :   0 - 0x0 -- Background 0x49
      11'h249: dout  = 8'b11111111; //  585 : 255 - 0xff
      11'h24A: dout  = 8'b11111111; //  586 : 255 - 0xff
      11'h24B: dout  = 8'b11100111; //  587 : 231 - 0xe7
      11'h24C: dout  = 8'b11100111; //  588 : 231 - 0xe7
      11'h24D: dout  = 8'b11111111; //  589 : 255 - 0xff
      11'h24E: dout  = 8'b11111111; //  590 : 255 - 0xff
      11'h24F: dout  = 8'b11111111; //  591 : 255 - 0xff
      11'h250: dout  = 8'b11111111; //  592 : 255 - 0xff -- Background 0x4a
      11'h251: dout  = 8'b11111111; //  593 : 255 - 0xff
      11'h252: dout  = 8'b11111111; //  594 : 255 - 0xff
      11'h253: dout  = 8'b11111111; //  595 : 255 - 0xff
      11'h254: dout  = 8'b11111111; //  596 : 255 - 0xff
      11'h255: dout  = 8'b11111111; //  597 : 255 - 0xff
      11'h256: dout  = 8'b11111111; //  598 : 255 - 0xff
      11'h257: dout  = 8'b11111111; //  599 : 255 - 0xff
      11'h258: dout  = 8'b00111111; //  600 :  63 - 0x3f -- Background 0x4b
      11'h259: dout  = 8'b01100000; //  601 :  96 - 0x60
      11'h25A: dout  = 8'b01000000; //  602 :  64 - 0x40
      11'h25B: dout  = 8'b11000000; //  603 : 192 - 0xc0
      11'h25C: dout  = 8'b10000000; //  604 : 128 - 0x80
      11'h25D: dout  = 8'b10000000; //  605 : 128 - 0x80
      11'h25E: dout  = 8'b10000000; //  606 : 128 - 0x80
      11'h25F: dout  = 8'b10000000; //  607 : 128 - 0x80
      11'h260: dout  = 8'b10000000; //  608 : 128 - 0x80 -- Background 0x4c
      11'h261: dout  = 8'b10000000; //  609 : 128 - 0x80
      11'h262: dout  = 8'b10000000; //  610 : 128 - 0x80
      11'h263: dout  = 8'b10000000; //  611 : 128 - 0x80
      11'h264: dout  = 8'b10000000; //  612 : 128 - 0x80
      11'h265: dout  = 8'b10000001; //  613 : 129 - 0x81
      11'h266: dout  = 8'b01000010; //  614 :  66 - 0x42
      11'h267: dout  = 8'b00111100; //  615 :  60 - 0x3c
      11'h268: dout  = 8'b11111111; //  616 : 255 - 0xff -- Background 0x4d
      11'h269: dout  = 8'b00000000; //  617 :   0 - 0x0
      11'h26A: dout  = 8'b00000000; //  618 :   0 - 0x0
      11'h26B: dout  = 8'b00000000; //  619 :   0 - 0x0
      11'h26C: dout  = 8'b00000000; //  620 :   0 - 0x0
      11'h26D: dout  = 8'b00000000; //  621 :   0 - 0x0
      11'h26E: dout  = 8'b00000000; //  622 :   0 - 0x0
      11'h26F: dout  = 8'b00000000; //  623 :   0 - 0x0
      11'h270: dout  = 8'b00000000; //  624 :   0 - 0x0 -- Background 0x4e
      11'h271: dout  = 8'b00000000; //  625 :   0 - 0x0
      11'h272: dout  = 8'b00000000; //  626 :   0 - 0x0
      11'h273: dout  = 8'b00000000; //  627 :   0 - 0x0
      11'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      11'h275: dout  = 8'b00000001; //  629 :   1 - 0x1
      11'h276: dout  = 8'b10000010; //  630 : 130 - 0x82
      11'h277: dout  = 8'b01111100; //  631 : 124 - 0x7c
      11'h278: dout  = 8'b00000000; //  632 :   0 - 0x0 -- Background 0x4f
      11'h279: dout  = 8'b00000000; //  633 :   0 - 0x0
      11'h27A: dout  = 8'b00000000; //  634 :   0 - 0x0
      11'h27B: dout  = 8'b00000000; //  635 :   0 - 0x0
      11'h27C: dout  = 8'b00000000; //  636 :   0 - 0x0
      11'h27D: dout  = 8'b00000001; //  637 :   1 - 0x1
      11'h27E: dout  = 8'b10000011; //  638 : 131 - 0x83
      11'h27F: dout  = 8'b11111111; //  639 : 255 - 0xff
      11'h280: dout  = 8'b11111000; //  640 : 248 - 0xf8 -- Background 0x50
      11'h281: dout  = 8'b00000100; //  641 :   4 - 0x4
      11'h282: dout  = 8'b00000010; //  642 :   2 - 0x2
      11'h283: dout  = 8'b00000010; //  643 :   2 - 0x2
      11'h284: dout  = 8'b00000001; //  644 :   1 - 0x1
      11'h285: dout  = 8'b00000001; //  645 :   1 - 0x1
      11'h286: dout  = 8'b00000001; //  646 :   1 - 0x1
      11'h287: dout  = 8'b00000001; //  647 :   1 - 0x1
      11'h288: dout  = 8'b00000001; //  648 :   1 - 0x1 -- Background 0x51
      11'h289: dout  = 8'b00000001; //  649 :   1 - 0x1
      11'h28A: dout  = 8'b00000001; //  650 :   1 - 0x1
      11'h28B: dout  = 8'b00000001; //  651 :   1 - 0x1
      11'h28C: dout  = 8'b00000001; //  652 :   1 - 0x1
      11'h28D: dout  = 8'b10000001; //  653 : 129 - 0x81
      11'h28E: dout  = 8'b01000010; //  654 :  66 - 0x42
      11'h28F: dout  = 8'b00111100; //  655 :  60 - 0x3c
      11'h290: dout  = 8'b11111111; //  656 : 255 - 0xff -- Background 0x52
      11'h291: dout  = 8'b11111111; //  657 : 255 - 0xff
      11'h292: dout  = 8'b11111111; //  658 : 255 - 0xff
      11'h293: dout  = 8'b11111111; //  659 : 255 - 0xff
      11'h294: dout  = 8'b11111111; //  660 : 255 - 0xff
      11'h295: dout  = 8'b11111111; //  661 : 255 - 0xff
      11'h296: dout  = 8'b11111111; //  662 : 255 - 0xff
      11'h297: dout  = 8'b11111111; //  663 : 255 - 0xff
      11'h298: dout  = 8'b01111111; //  664 : 127 - 0x7f -- Background 0x53
      11'h299: dout  = 8'b10000000; //  665 : 128 - 0x80
      11'h29A: dout  = 8'b10100000; //  666 : 160 - 0xa0
      11'h29B: dout  = 8'b10000111; //  667 : 135 - 0x87
      11'h29C: dout  = 8'b10001111; //  668 : 143 - 0x8f
      11'h29D: dout  = 8'b10001110; //  669 : 142 - 0x8e
      11'h29E: dout  = 8'b10001110; //  670 : 142 - 0x8e
      11'h29F: dout  = 8'b10000110; //  671 : 134 - 0x86
      11'h2A0: dout  = 8'b11111110; //  672 : 254 - 0xfe -- Background 0x54
      11'h2A1: dout  = 8'b00000001; //  673 :   1 - 0x1
      11'h2A2: dout  = 8'b00000101; //  674 :   5 - 0x5
      11'h2A3: dout  = 8'b11000001; //  675 : 193 - 0xc1
      11'h2A4: dout  = 8'b11100001; //  676 : 225 - 0xe1
      11'h2A5: dout  = 8'b01110001; //  677 : 113 - 0x71
      11'h2A6: dout  = 8'b01110001; //  678 : 113 - 0x71
      11'h2A7: dout  = 8'b11110001; //  679 : 241 - 0xf1
      11'h2A8: dout  = 8'b10000001; //  680 : 129 - 0x81 -- Background 0x55
      11'h2A9: dout  = 8'b10000001; //  681 : 129 - 0x81
      11'h2AA: dout  = 8'b10000000; //  682 : 128 - 0x80
      11'h2AB: dout  = 8'b10000001; //  683 : 129 - 0x81
      11'h2AC: dout  = 8'b10000001; //  684 : 129 - 0x81
      11'h2AD: dout  = 8'b10100000; //  685 : 160 - 0xa0
      11'h2AE: dout  = 8'b10000000; //  686 : 128 - 0x80
      11'h2AF: dout  = 8'b11111111; //  687 : 255 - 0xff
      11'h2B0: dout  = 8'b11110001; //  688 : 241 - 0xf1 -- Background 0x56
      11'h2B1: dout  = 8'b11000001; //  689 : 193 - 0xc1
      11'h2B2: dout  = 8'b11000001; //  690 : 193 - 0xc1
      11'h2B3: dout  = 8'b10000001; //  691 : 129 - 0x81
      11'h2B4: dout  = 8'b11000001; //  692 : 193 - 0xc1
      11'h2B5: dout  = 8'b11000101; //  693 : 197 - 0xc5
      11'h2B6: dout  = 8'b00000001; //  694 :   1 - 0x1
      11'h2B7: dout  = 8'b11111111; //  695 : 255 - 0xff
      11'h2B8: dout  = 8'b01111111; //  696 : 127 - 0x7f -- Background 0x57
      11'h2B9: dout  = 8'b11111111; //  697 : 255 - 0xff
      11'h2BA: dout  = 8'b11111111; //  698 : 255 - 0xff
      11'h2BB: dout  = 8'b11111111; //  699 : 255 - 0xff
      11'h2BC: dout  = 8'b11111111; //  700 : 255 - 0xff
      11'h2BD: dout  = 8'b11111111; //  701 : 255 - 0xff
      11'h2BE: dout  = 8'b11111111; //  702 : 255 - 0xff
      11'h2BF: dout  = 8'b11111111; //  703 : 255 - 0xff
      11'h2C0: dout  = 8'b11111110; //  704 : 254 - 0xfe -- Background 0x58
      11'h2C1: dout  = 8'b11111111; //  705 : 255 - 0xff
      11'h2C2: dout  = 8'b11111111; //  706 : 255 - 0xff
      11'h2C3: dout  = 8'b11111111; //  707 : 255 - 0xff
      11'h2C4: dout  = 8'b11111111; //  708 : 255 - 0xff
      11'h2C5: dout  = 8'b11111111; //  709 : 255 - 0xff
      11'h2C6: dout  = 8'b11111111; //  710 : 255 - 0xff
      11'h2C7: dout  = 8'b11111111; //  711 : 255 - 0xff
      11'h2C8: dout  = 8'b11111111; //  712 : 255 - 0xff -- Background 0x59
      11'h2C9: dout  = 8'b11111111; //  713 : 255 - 0xff
      11'h2CA: dout  = 8'b11111111; //  714 : 255 - 0xff
      11'h2CB: dout  = 8'b11111111; //  715 : 255 - 0xff
      11'h2CC: dout  = 8'b11111111; //  716 : 255 - 0xff
      11'h2CD: dout  = 8'b11111111; //  717 : 255 - 0xff
      11'h2CE: dout  = 8'b11111111; //  718 : 255 - 0xff
      11'h2CF: dout  = 8'b01111111; //  719 : 127 - 0x7f
      11'h2D0: dout  = 8'b11111111; //  720 : 255 - 0xff -- Background 0x5a
      11'h2D1: dout  = 8'b11111111; //  721 : 255 - 0xff
      11'h2D2: dout  = 8'b11111111; //  722 : 255 - 0xff
      11'h2D3: dout  = 8'b11111111; //  723 : 255 - 0xff
      11'h2D4: dout  = 8'b11111111; //  724 : 255 - 0xff
      11'h2D5: dout  = 8'b11111111; //  725 : 255 - 0xff
      11'h2D6: dout  = 8'b11111111; //  726 : 255 - 0xff
      11'h2D7: dout  = 8'b11111110; //  727 : 254 - 0xfe
      11'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- Background 0x5b
      11'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      11'h2DA: dout  = 8'b00000000; //  730 :   0 - 0x0
      11'h2DB: dout  = 8'b00000000; //  731 :   0 - 0x0
      11'h2DC: dout  = 8'b00000000; //  732 :   0 - 0x0
      11'h2DD: dout  = 8'b00000000; //  733 :   0 - 0x0
      11'h2DE: dout  = 8'b00111000; //  734 :  56 - 0x38
      11'h2DF: dout  = 8'b01111100; //  735 : 124 - 0x7c
      11'h2E0: dout  = 8'b11111110; //  736 : 254 - 0xfe -- Background 0x5c
      11'h2E1: dout  = 8'b11111110; //  737 : 254 - 0xfe
      11'h2E2: dout  = 8'b11111110; //  738 : 254 - 0xfe
      11'h2E3: dout  = 8'b01111100; //  739 : 124 - 0x7c
      11'h2E4: dout  = 8'b00111000; //  740 :  56 - 0x38
      11'h2E5: dout  = 8'b00000000; //  741 :   0 - 0x0
      11'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      11'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      11'h2E8: dout  = 8'b00100000; //  744 :  32 - 0x20 -- Background 0x5d
      11'h2E9: dout  = 8'b11100111; //  745 : 231 - 0xe7
      11'h2EA: dout  = 8'b11100111; //  746 : 231 - 0xe7
      11'h2EB: dout  = 8'b11100111; //  747 : 231 - 0xe7
      11'h2EC: dout  = 8'b11100111; //  748 : 231 - 0xe7
      11'h2ED: dout  = 8'b11100111; //  749 : 231 - 0xe7
      11'h2EE: dout  = 8'b11101111; //  750 : 239 - 0xef
      11'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      11'h2F0: dout  = 8'b00000010; //  752 :   2 - 0x2 -- Background 0x5e
      11'h2F1: dout  = 8'b01111110; //  753 : 126 - 0x7e
      11'h2F2: dout  = 8'b01111110; //  754 : 126 - 0x7e
      11'h2F3: dout  = 8'b01111110; //  755 : 126 - 0x7e
      11'h2F4: dout  = 8'b01111110; //  756 : 126 - 0x7e
      11'h2F5: dout  = 8'b01111110; //  757 : 126 - 0x7e
      11'h2F6: dout  = 8'b11111110; //  758 : 254 - 0xfe
      11'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      11'h2F8: dout  = 8'b01111111; //  760 : 127 - 0x7f -- Background 0x5f
      11'h2F9: dout  = 8'b01111111; //  761 : 127 - 0x7f
      11'h2FA: dout  = 8'b01111111; //  762 : 127 - 0x7f
      11'h2FB: dout  = 8'b01100111; //  763 : 103 - 0x67
      11'h2FC: dout  = 8'b01100111; //  764 : 103 - 0x67
      11'h2FD: dout  = 8'b01111111; //  765 : 127 - 0x7f
      11'h2FE: dout  = 8'b01111111; //  766 : 127 - 0x7f
      11'h2FF: dout  = 8'b01111111; //  767 : 127 - 0x7f
      11'h300: dout  = 8'b11111111; //  768 : 255 - 0xff -- Background 0x60
      11'h301: dout  = 8'b10000000; //  769 : 128 - 0x80
      11'h302: dout  = 8'b11111100; //  770 : 252 - 0xfc
      11'h303: dout  = 8'b10001100; //  771 : 140 - 0x8c
      11'h304: dout  = 8'b10001100; //  772 : 140 - 0x8c
      11'h305: dout  = 8'b10001100; //  773 : 140 - 0x8c
      11'h306: dout  = 8'b10001100; //  774 : 140 - 0x8c
      11'h307: dout  = 8'b10001100; //  775 : 140 - 0x8c
      11'h308: dout  = 8'b11111111; //  776 : 255 - 0xff -- Background 0x61
      11'h309: dout  = 8'b00000000; //  777 :   0 - 0x0
      11'h30A: dout  = 8'b00001111; //  778 :  15 - 0xf
      11'h30B: dout  = 8'b00001001; //  779 :   9 - 0x9
      11'h30C: dout  = 8'b00001001; //  780 :   9 - 0x9
      11'h30D: dout  = 8'b00001001; //  781 :   9 - 0x9
      11'h30E: dout  = 8'b00001001; //  782 :   9 - 0x9
      11'h30F: dout  = 8'b00001001; //  783 :   9 - 0x9
      11'h310: dout  = 8'b11111111; //  784 : 255 - 0xff -- Background 0x62
      11'h311: dout  = 8'b00000000; //  785 :   0 - 0x0
      11'h312: dout  = 8'b11111111; //  786 : 255 - 0xff
      11'h313: dout  = 8'b11111111; //  787 : 255 - 0xff
      11'h314: dout  = 8'b11111111; //  788 : 255 - 0xff
      11'h315: dout  = 8'b11111111; //  789 : 255 - 0xff
      11'h316: dout  = 8'b11111111; //  790 : 255 - 0xff
      11'h317: dout  = 8'b11111111; //  791 : 255 - 0xff
      11'h318: dout  = 8'b11111111; //  792 : 255 - 0xff -- Background 0x63
      11'h319: dout  = 8'b00000001; //  793 :   1 - 0x1
      11'h31A: dout  = 8'b11111111; //  794 : 255 - 0xff
      11'h31B: dout  = 8'b10101001; //  795 : 169 - 0xa9
      11'h31C: dout  = 8'b11010001; //  796 : 209 - 0xd1
      11'h31D: dout  = 8'b10101001; //  797 : 169 - 0xa9
      11'h31E: dout  = 8'b11010001; //  798 : 209 - 0xd1
      11'h31F: dout  = 8'b10101001; //  799 : 169 - 0xa9
      11'h320: dout  = 8'b10001100; //  800 : 140 - 0x8c -- Background 0x64
      11'h321: dout  = 8'b10001100; //  801 : 140 - 0x8c
      11'h322: dout  = 8'b10001100; //  802 : 140 - 0x8c
      11'h323: dout  = 8'b10001100; //  803 : 140 - 0x8c
      11'h324: dout  = 8'b10001100; //  804 : 140 - 0x8c
      11'h325: dout  = 8'b10001100; //  805 : 140 - 0x8c
      11'h326: dout  = 8'b11111111; //  806 : 255 - 0xff
      11'h327: dout  = 8'b00111111; //  807 :  63 - 0x3f
      11'h328: dout  = 8'b00001001; //  808 :   9 - 0x9 -- Background 0x65
      11'h329: dout  = 8'b00001001; //  809 :   9 - 0x9
      11'h32A: dout  = 8'b00001001; //  810 :   9 - 0x9
      11'h32B: dout  = 8'b00001001; //  811 :   9 - 0x9
      11'h32C: dout  = 8'b00001001; //  812 :   9 - 0x9
      11'h32D: dout  = 8'b00001001; //  813 :   9 - 0x9
      11'h32E: dout  = 8'b11111111; //  814 : 255 - 0xff
      11'h32F: dout  = 8'b11111111; //  815 : 255 - 0xff
      11'h330: dout  = 8'b11111111; //  816 : 255 - 0xff -- Background 0x66
      11'h331: dout  = 8'b11111111; //  817 : 255 - 0xff
      11'h332: dout  = 8'b11111111; //  818 : 255 - 0xff
      11'h333: dout  = 8'b11111111; //  819 : 255 - 0xff
      11'h334: dout  = 8'b11111111; //  820 : 255 - 0xff
      11'h335: dout  = 8'b11111111; //  821 : 255 - 0xff
      11'h336: dout  = 8'b11111111; //  822 : 255 - 0xff
      11'h337: dout  = 8'b11111111; //  823 : 255 - 0xff
      11'h338: dout  = 8'b11010001; //  824 : 209 - 0xd1 -- Background 0x67
      11'h339: dout  = 8'b10101001; //  825 : 169 - 0xa9
      11'h33A: dout  = 8'b11010001; //  826 : 209 - 0xd1
      11'h33B: dout  = 8'b10101001; //  827 : 169 - 0xa9
      11'h33C: dout  = 8'b11010001; //  828 : 209 - 0xd1
      11'h33D: dout  = 8'b10101001; //  829 : 169 - 0xa9
      11'h33E: dout  = 8'b11111111; //  830 : 255 - 0xff
      11'h33F: dout  = 8'b11111100; //  831 : 252 - 0xfc
      11'h340: dout  = 8'b00100011; //  832 :  35 - 0x23 -- Background 0x68
      11'h341: dout  = 8'b00100011; //  833 :  35 - 0x23
      11'h342: dout  = 8'b00100011; //  834 :  35 - 0x23
      11'h343: dout  = 8'b00100011; //  835 :  35 - 0x23
      11'h344: dout  = 8'b00100011; //  836 :  35 - 0x23
      11'h345: dout  = 8'b00100011; //  837 :  35 - 0x23
      11'h346: dout  = 8'b00100011; //  838 :  35 - 0x23
      11'h347: dout  = 8'b00100011; //  839 :  35 - 0x23
      11'h348: dout  = 8'b00000100; //  840 :   4 - 0x4 -- Background 0x69
      11'h349: dout  = 8'b00000100; //  841 :   4 - 0x4
      11'h34A: dout  = 8'b00000100; //  842 :   4 - 0x4
      11'h34B: dout  = 8'b00000100; //  843 :   4 - 0x4
      11'h34C: dout  = 8'b00000100; //  844 :   4 - 0x4
      11'h34D: dout  = 8'b00000100; //  845 :   4 - 0x4
      11'h34E: dout  = 8'b00000100; //  846 :   4 - 0x4
      11'h34F: dout  = 8'b00000100; //  847 :   4 - 0x4
      11'h350: dout  = 8'b01000100; //  848 :  68 - 0x44 -- Background 0x6a
      11'h351: dout  = 8'b10100100; //  849 : 164 - 0xa4
      11'h352: dout  = 8'b01000100; //  850 :  68 - 0x44
      11'h353: dout  = 8'b10100100; //  851 : 164 - 0xa4
      11'h354: dout  = 8'b01000100; //  852 :  68 - 0x44
      11'h355: dout  = 8'b10100100; //  853 : 164 - 0xa4
      11'h356: dout  = 8'b01000100; //  854 :  68 - 0x44
      11'h357: dout  = 8'b10100100; //  855 : 164 - 0xa4
      11'h358: dout  = 8'b00011111; //  856 :  31 - 0x1f -- Background 0x6b
      11'h359: dout  = 8'b00111111; //  857 :  63 - 0x3f
      11'h35A: dout  = 8'b01111111; //  858 : 127 - 0x7f
      11'h35B: dout  = 8'b01111111; //  859 : 127 - 0x7f
      11'h35C: dout  = 8'b11111111; //  860 : 255 - 0xff
      11'h35D: dout  = 8'b11111111; //  861 : 255 - 0xff
      11'h35E: dout  = 8'b11111111; //  862 : 255 - 0xff
      11'h35F: dout  = 8'b11111110; //  863 : 254 - 0xfe
      11'h360: dout  = 8'b11111111; //  864 : 255 - 0xff -- Background 0x6c
      11'h361: dout  = 8'b01111111; //  865 : 127 - 0x7f
      11'h362: dout  = 8'b01111111; //  866 : 127 - 0x7f
      11'h363: dout  = 8'b00111111; //  867 :  63 - 0x3f
      11'h364: dout  = 8'b00000000; //  868 :   0 - 0x0
      11'h365: dout  = 8'b00000000; //  869 :   0 - 0x0
      11'h366: dout  = 8'b00000001; //  870 :   1 - 0x1
      11'h367: dout  = 8'b00000001; //  871 :   1 - 0x1
      11'h368: dout  = 8'b11111111; //  872 : 255 - 0xff -- Background 0x6d
      11'h369: dout  = 8'b10000000; //  873 : 128 - 0x80
      11'h36A: dout  = 8'b10000000; //  874 : 128 - 0x80
      11'h36B: dout  = 8'b00000000; //  875 :   0 - 0x0
      11'h36C: dout  = 8'b00000000; //  876 :   0 - 0x0
      11'h36D: dout  = 8'b11111000; //  877 : 248 - 0xf8
      11'h36E: dout  = 8'b11111100; //  878 : 252 - 0xfc
      11'h36F: dout  = 8'b11111100; //  879 : 252 - 0xfc
      11'h370: dout  = 8'b11111111; //  880 : 255 - 0xff -- Background 0x6e
      11'h371: dout  = 8'b11111111; //  881 : 255 - 0xff
      11'h372: dout  = 8'b11111111; //  882 : 255 - 0xff
      11'h373: dout  = 8'b11111111; //  883 : 255 - 0xff
      11'h374: dout  = 8'b11111111; //  884 : 255 - 0xff
      11'h375: dout  = 8'b01111110; //  885 : 126 - 0x7e
      11'h376: dout  = 8'b00111100; //  886 :  60 - 0x3c
      11'h377: dout  = 8'b00000000; //  887 :   0 - 0x0
      11'h378: dout  = 8'b11111000; //  888 : 248 - 0xf8 -- Background 0x6f
      11'h379: dout  = 8'b00000100; //  889 :   4 - 0x4
      11'h37A: dout  = 8'b00000010; //  890 :   2 - 0x2
      11'h37B: dout  = 8'b00000010; //  891 :   2 - 0x2
      11'h37C: dout  = 8'b00011101; //  892 :  29 - 0x1d
      11'h37D: dout  = 8'b00111111; //  893 :  63 - 0x3f
      11'h37E: dout  = 8'b01111111; //  894 : 127 - 0x7f
      11'h37F: dout  = 8'b01111111; //  895 : 127 - 0x7f
      11'h380: dout  = 8'b11111100; //  896 : 252 - 0xfc -- Background 0x70
      11'h381: dout  = 8'b10000000; //  897 : 128 - 0x80
      11'h382: dout  = 8'b10000000; //  898 : 128 - 0x80
      11'h383: dout  = 8'b10000000; //  899 : 128 - 0x80
      11'h384: dout  = 8'b10000000; //  900 : 128 - 0x80
      11'h385: dout  = 8'b10000000; //  901 : 128 - 0x80
      11'h386: dout  = 8'b01100000; //  902 :  96 - 0x60
      11'h387: dout  = 8'b00011111; //  903 :  31 - 0x1f
      11'h388: dout  = 8'b00000011; //  904 :   3 - 0x3 -- Background 0x71
      11'h389: dout  = 8'b00000011; //  905 :   3 - 0x3
      11'h38A: dout  = 8'b00000011; //  906 :   3 - 0x3
      11'h38B: dout  = 8'b00000011; //  907 :   3 - 0x3
      11'h38C: dout  = 8'b00000001; //  908 :   1 - 0x1
      11'h38D: dout  = 8'b00000001; //  909 :   1 - 0x1
      11'h38E: dout  = 8'b00000000; //  910 :   0 - 0x0
      11'h38F: dout  = 8'b11111111; //  911 : 255 - 0xff
      11'h390: dout  = 8'b11111110; //  912 : 254 - 0xfe -- Background 0x72
      11'h391: dout  = 8'b11111110; //  913 : 254 - 0xfe
      11'h392: dout  = 8'b11111110; //  914 : 254 - 0xfe
      11'h393: dout  = 8'b11111110; //  915 : 254 - 0xfe
      11'h394: dout  = 8'b11111100; //  916 : 252 - 0xfc
      11'h395: dout  = 8'b11111100; //  917 : 252 - 0xfc
      11'h396: dout  = 8'b11111000; //  918 : 248 - 0xf8
      11'h397: dout  = 8'b11111111; //  919 : 255 - 0xff
      11'h398: dout  = 8'b00000000; //  920 :   0 - 0x0 -- Background 0x73
      11'h399: dout  = 8'b00000000; //  921 :   0 - 0x0
      11'h39A: dout  = 8'b00000000; //  922 :   0 - 0x0
      11'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      11'h39C: dout  = 8'b00000000; //  924 :   0 - 0x0
      11'h39D: dout  = 8'b00000000; //  925 :   0 - 0x0
      11'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      11'h39F: dout  = 8'b11111111; //  927 : 255 - 0xff
      11'h3A0: dout  = 8'b01111111; //  928 : 127 - 0x7f -- Background 0x74
      11'h3A1: dout  = 8'b00111111; //  929 :  63 - 0x3f
      11'h3A2: dout  = 8'b00011101; //  930 :  29 - 0x1d
      11'h3A3: dout  = 8'b00000001; //  931 :   1 - 0x1
      11'h3A4: dout  = 8'b00000001; //  932 :   1 - 0x1
      11'h3A5: dout  = 8'b00000001; //  933 :   1 - 0x1
      11'h3A6: dout  = 8'b00000011; //  934 :   3 - 0x3
      11'h3A7: dout  = 8'b11111110; //  935 : 254 - 0xfe
      11'h3A8: dout  = 8'b10000000; //  936 : 128 - 0x80 -- Background 0x75
      11'h3A9: dout  = 8'b10000000; //  937 : 128 - 0x80
      11'h3AA: dout  = 8'b10000000; //  938 : 128 - 0x80
      11'h3AB: dout  = 8'b10000000; //  939 : 128 - 0x80
      11'h3AC: dout  = 8'b10000000; //  940 : 128 - 0x80
      11'h3AD: dout  = 8'b10000100; //  941 : 132 - 0x84
      11'h3AE: dout  = 8'b11001010; //  942 : 202 - 0xca
      11'h3AF: dout  = 8'b10110001; //  943 : 177 - 0xb1
      11'h3B0: dout  = 8'b00000001; //  944 :   1 - 0x1 -- Background 0x76
      11'h3B1: dout  = 8'b00000001; //  945 :   1 - 0x1
      11'h3B2: dout  = 8'b00000001; //  946 :   1 - 0x1
      11'h3B3: dout  = 8'b00000001; //  947 :   1 - 0x1
      11'h3B4: dout  = 8'b00000001; //  948 :   1 - 0x1
      11'h3B5: dout  = 8'b00100001; //  949 :  33 - 0x21
      11'h3B6: dout  = 8'b01010011; //  950 :  83 - 0x53
      11'h3B7: dout  = 8'b10001101; //  951 : 141 - 0x8d
      11'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0 -- Background 0x77
      11'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      11'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      11'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      11'h3BC: dout  = 8'b01110111; //  956 : 119 - 0x77
      11'h3BD: dout  = 8'b11111111; //  957 : 255 - 0xff
      11'h3BE: dout  = 8'b11111111; //  958 : 255 - 0xff
      11'h3BF: dout  = 8'b11111111; //  959 : 255 - 0xff
      11'h3C0: dout  = 8'b11111111; //  960 : 255 - 0xff -- Background 0x78
      11'h3C1: dout  = 8'b11111111; //  961 : 255 - 0xff
      11'h3C2: dout  = 8'b11111111; //  962 : 255 - 0xff
      11'h3C3: dout  = 8'b11111111; //  963 : 255 - 0xff
      11'h3C4: dout  = 8'b11111111; //  964 : 255 - 0xff
      11'h3C5: dout  = 8'b11111111; //  965 : 255 - 0xff
      11'h3C6: dout  = 8'b11111111; //  966 : 255 - 0xff
      11'h3C7: dout  = 8'b11111111; //  967 : 255 - 0xff
      11'h3C8: dout  = 8'b11111111; //  968 : 255 - 0xff -- Background 0x79
      11'h3C9: dout  = 8'b11111111; //  969 : 255 - 0xff
      11'h3CA: dout  = 8'b11111111; //  970 : 255 - 0xff
      11'h3CB: dout  = 8'b01110111; //  971 : 119 - 0x77
      11'h3CC: dout  = 8'b01110111; //  972 : 119 - 0x77
      11'h3CD: dout  = 8'b01110111; //  973 : 119 - 0x77
      11'h3CE: dout  = 8'b01110111; //  974 : 119 - 0x77
      11'h3CF: dout  = 8'b01110111; //  975 : 119 - 0x77
      11'h3D0: dout  = 8'b11111111; //  976 : 255 - 0xff -- Background 0x7a
      11'h3D1: dout  = 8'b11111111; //  977 : 255 - 0xff
      11'h3D2: dout  = 8'b11111111; //  978 : 255 - 0xff
      11'h3D3: dout  = 8'b11100111; //  979 : 231 - 0xe7
      11'h3D4: dout  = 8'b11100111; //  980 : 231 - 0xe7
      11'h3D5: dout  = 8'b11111111; //  981 : 255 - 0xff
      11'h3D6: dout  = 8'b11111111; //  982 : 255 - 0xff
      11'h3D7: dout  = 8'b11111110; //  983 : 254 - 0xfe
      11'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0 -- Background 0x7b
      11'h3D9: dout  = 8'b00100001; //  985 :  33 - 0x21
      11'h3DA: dout  = 8'b00100001; //  986 :  33 - 0x21
      11'h3DB: dout  = 8'b01000001; //  987 :  65 - 0x41
      11'h3DC: dout  = 8'b01000001; //  988 :  65 - 0x41
      11'h3DD: dout  = 8'b01000001; //  989 :  65 - 0x41
      11'h3DE: dout  = 8'b01000001; //  990 :  65 - 0x41
      11'h3DF: dout  = 8'b01000001; //  991 :  65 - 0x41
      11'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Background 0x7c
      11'h3E1: dout  = 8'b10000000; //  993 : 128 - 0x80
      11'h3E2: dout  = 8'b10000000; //  994 : 128 - 0x80
      11'h3E3: dout  = 8'b10000000; //  995 : 128 - 0x80
      11'h3E4: dout  = 8'b10000000; //  996 : 128 - 0x80
      11'h3E5: dout  = 8'b10000000; //  997 : 128 - 0x80
      11'h3E6: dout  = 8'b10000000; //  998 : 128 - 0x80
      11'h3E7: dout  = 8'b10000000; //  999 : 128 - 0x80
      11'h3E8: dout  = 8'b00100001; // 1000 :  33 - 0x21 -- Background 0x7d
      11'h3E9: dout  = 8'b00100001; // 1001 :  33 - 0x21
      11'h3EA: dout  = 8'b00000001; // 1002 :   1 - 0x1
      11'h3EB: dout  = 8'b00000001; // 1003 :   1 - 0x1
      11'h3EC: dout  = 8'b00000001; // 1004 :   1 - 0x1
      11'h3ED: dout  = 8'b00000001; // 1005 :   1 - 0x1
      11'h3EE: dout  = 8'b00000001; // 1006 :   1 - 0x1
      11'h3EF: dout  = 8'b00000001; // 1007 :   1 - 0x1
      11'h3F0: dout  = 8'b10000000; // 1008 : 128 - 0x80 -- Background 0x7e
      11'h3F1: dout  = 8'b10000000; // 1009 : 128 - 0x80
      11'h3F2: dout  = 8'b10000000; // 1010 : 128 - 0x80
      11'h3F3: dout  = 8'b10000000; // 1011 : 128 - 0x80
      11'h3F4: dout  = 8'b10000000; // 1012 : 128 - 0x80
      11'h3F5: dout  = 8'b10000000; // 1013 : 128 - 0x80
      11'h3F6: dout  = 8'b10000000; // 1014 : 128 - 0x80
      11'h3F7: dout  = 8'b10000000; // 1015 : 128 - 0x80
      11'h3F8: dout  = 8'b00000001; // 1016 :   1 - 0x1 -- Background 0x7f
      11'h3F9: dout  = 8'b00000001; // 1017 :   1 - 0x1
      11'h3FA: dout  = 8'b00000110; // 1018 :   6 - 0x6
      11'h3FB: dout  = 8'b00001000; // 1019 :   8 - 0x8
      11'h3FC: dout  = 8'b00011000; // 1020 :  24 - 0x18
      11'h3FD: dout  = 8'b00100000; // 1021 :  32 - 0x20
      11'h3FE: dout  = 8'b00100000; // 1022 :  32 - 0x20
      11'h3FF: dout  = 8'b11000000; // 1023 : 192 - 0xc0
      11'h400: dout  = 8'b00000100; // 1024 :   4 - 0x4 -- Background 0x80
      11'h401: dout  = 8'b00000100; // 1025 :   4 - 0x4
      11'h402: dout  = 8'b11000100; // 1026 : 196 - 0xc4
      11'h403: dout  = 8'b11110100; // 1027 : 244 - 0xf4
      11'h404: dout  = 8'b11110100; // 1028 : 244 - 0xf4
      11'h405: dout  = 8'b00000100; // 1029 :   4 - 0x4
      11'h406: dout  = 8'b00000100; // 1030 :   4 - 0x4
      11'h407: dout  = 8'b00000101; // 1031 :   5 - 0x5
      11'h408: dout  = 8'b01110000; // 1032 : 112 - 0x70 -- Background 0x81
      11'h409: dout  = 8'b11110000; // 1033 : 240 - 0xf0
      11'h40A: dout  = 8'b11110000; // 1034 : 240 - 0xf0
      11'h40B: dout  = 8'b11111111; // 1035 : 255 - 0xff
      11'h40C: dout  = 8'b11111111; // 1036 : 255 - 0xff
      11'h40D: dout  = 8'b11110000; // 1037 : 240 - 0xf0
      11'h40E: dout  = 8'b11110000; // 1038 : 240 - 0xf0
      11'h40F: dout  = 8'b01110000; // 1039 : 112 - 0x70
      11'h410: dout  = 8'b11000000; // 1040 : 192 - 0xc0 -- Background 0x82
      11'h411: dout  = 8'b10000111; // 1041 : 135 - 0x87
      11'h412: dout  = 8'b00011000; // 1042 :  24 - 0x18
      11'h413: dout  = 8'b10110000; // 1043 : 176 - 0xb0
      11'h414: dout  = 8'b11100111; // 1044 : 231 - 0xe7
      11'h415: dout  = 8'b11100111; // 1045 : 231 - 0xe7
      11'h416: dout  = 8'b11101111; // 1046 : 239 - 0xef
      11'h417: dout  = 8'b11101111; // 1047 : 239 - 0xef
      11'h418: dout  = 8'b01101111; // 1048 : 111 - 0x6f -- Background 0x83
      11'h419: dout  = 8'b01000011; // 1049 :  67 - 0x43
      11'h41A: dout  = 8'b01011101; // 1050 :  93 - 0x5d
      11'h41B: dout  = 8'b00111111; // 1051 :  63 - 0x3f
      11'h41C: dout  = 8'b00111111; // 1052 :  63 - 0x3f
      11'h41D: dout  = 8'b01111111; // 1053 : 127 - 0x7f
      11'h41E: dout  = 8'b01111111; // 1054 : 127 - 0x7f
      11'h41F: dout  = 8'b11111111; // 1055 : 255 - 0xff
      11'h420: dout  = 8'b00000011; // 1056 :   3 - 0x3 -- Background 0x84
      11'h421: dout  = 8'b11111111; // 1057 : 255 - 0xff
      11'h422: dout  = 8'b11110001; // 1058 : 241 - 0xf1
      11'h423: dout  = 8'b01101110; // 1059 : 110 - 0x6e
      11'h424: dout  = 8'b11001111; // 1060 : 207 - 0xcf
      11'h425: dout  = 8'b11011111; // 1061 : 223 - 0xdf
      11'h426: dout  = 8'b11111111; // 1062 : 255 - 0xff
      11'h427: dout  = 8'b11111111; // 1063 : 255 - 0xff
      11'h428: dout  = 8'b11111101; // 1064 : 253 - 0xfd -- Background 0x85
      11'h429: dout  = 8'b11111011; // 1065 : 251 - 0xfb
      11'h42A: dout  = 8'b11111011; // 1066 : 251 - 0xfb
      11'h42B: dout  = 8'b11110111; // 1067 : 247 - 0xf7
      11'h42C: dout  = 8'b11110111; // 1068 : 247 - 0xf7
      11'h42D: dout  = 8'b00001111; // 1069 :  15 - 0xf
      11'h42E: dout  = 8'b01111111; // 1070 : 127 - 0x7f
      11'h42F: dout  = 8'b11111111; // 1071 : 255 - 0xff
      11'h430: dout  = 8'b11111111; // 1072 : 255 - 0xff -- Background 0x86
      11'h431: dout  = 8'b10000000; // 1073 : 128 - 0x80
      11'h432: dout  = 8'b10000000; // 1074 : 128 - 0x80
      11'h433: dout  = 8'b10000000; // 1075 : 128 - 0x80
      11'h434: dout  = 8'b10000000; // 1076 : 128 - 0x80
      11'h435: dout  = 8'b11111111; // 1077 : 255 - 0xff
      11'h436: dout  = 8'b11111111; // 1078 : 255 - 0xff
      11'h437: dout  = 8'b10000000; // 1079 : 128 - 0x80
      11'h438: dout  = 8'b11111110; // 1080 : 254 - 0xfe -- Background 0x87
      11'h439: dout  = 8'b00000011; // 1081 :   3 - 0x3
      11'h43A: dout  = 8'b00000011; // 1082 :   3 - 0x3
      11'h43B: dout  = 8'b00000011; // 1083 :   3 - 0x3
      11'h43C: dout  = 8'b00000011; // 1084 :   3 - 0x3
      11'h43D: dout  = 8'b11111111; // 1085 : 255 - 0xff
      11'h43E: dout  = 8'b11111111; // 1086 : 255 - 0xff
      11'h43F: dout  = 8'b00000011; // 1087 :   3 - 0x3
      11'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Background 0x88
      11'h441: dout  = 8'b11111111; // 1089 : 255 - 0xff
      11'h442: dout  = 8'b00000000; // 1090 :   0 - 0x0
      11'h443: dout  = 8'b00000000; // 1091 :   0 - 0x0
      11'h444: dout  = 8'b00000000; // 1092 :   0 - 0x0
      11'h445: dout  = 8'b00000000; // 1093 :   0 - 0x0
      11'h446: dout  = 8'b11111111; // 1094 : 255 - 0xff
      11'h447: dout  = 8'b11111111; // 1095 : 255 - 0xff
      11'h448: dout  = 8'b00100011; // 1096 :  35 - 0x23 -- Background 0x89
      11'h449: dout  = 8'b11110011; // 1097 : 243 - 0xf3
      11'h44A: dout  = 8'b00001011; // 1098 :  11 - 0xb
      11'h44B: dout  = 8'b00001011; // 1099 :  11 - 0xb
      11'h44C: dout  = 8'b00001011; // 1100 :  11 - 0xb
      11'h44D: dout  = 8'b00000111; // 1101 :   7 - 0x7
      11'h44E: dout  = 8'b11111111; // 1102 : 255 - 0xff
      11'h44F: dout  = 8'b11111111; // 1103 : 255 - 0xff
      11'h450: dout  = 8'b10000000; // 1104 : 128 - 0x80 -- Background 0x8a
      11'h451: dout  = 8'b10000000; // 1105 : 128 - 0x80
      11'h452: dout  = 8'b10000000; // 1106 : 128 - 0x80
      11'h453: dout  = 8'b10000000; // 1107 : 128 - 0x80
      11'h454: dout  = 8'b11111111; // 1108 : 255 - 0xff
      11'h455: dout  = 8'b10000000; // 1109 : 128 - 0x80
      11'h456: dout  = 8'b10000000; // 1110 : 128 - 0x80
      11'h457: dout  = 8'b10000000; // 1111 : 128 - 0x80
      11'h458: dout  = 8'b00000011; // 1112 :   3 - 0x3 -- Background 0x8b
      11'h459: dout  = 8'b00000011; // 1113 :   3 - 0x3
      11'h45A: dout  = 8'b00000011; // 1114 :   3 - 0x3
      11'h45B: dout  = 8'b00000011; // 1115 :   3 - 0x3
      11'h45C: dout  = 8'b11111111; // 1116 : 255 - 0xff
      11'h45D: dout  = 8'b00000011; // 1117 :   3 - 0x3
      11'h45E: dout  = 8'b00000011; // 1118 :   3 - 0x3
      11'h45F: dout  = 8'b00000011; // 1119 :   3 - 0x3
      11'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Background 0x8c
      11'h461: dout  = 8'b00000000; // 1121 :   0 - 0x0
      11'h462: dout  = 8'b00000000; // 1122 :   0 - 0x0
      11'h463: dout  = 8'b00000000; // 1123 :   0 - 0x0
      11'h464: dout  = 8'b00000000; // 1124 :   0 - 0x0
      11'h465: dout  = 8'b11111111; // 1125 : 255 - 0xff
      11'h466: dout  = 8'b00000000; // 1126 :   0 - 0x0
      11'h467: dout  = 8'b00000000; // 1127 :   0 - 0x0
      11'h468: dout  = 8'b00000111; // 1128 :   7 - 0x7 -- Background 0x8d
      11'h469: dout  = 8'b00000111; // 1129 :   7 - 0x7
      11'h46A: dout  = 8'b00000011; // 1130 :   3 - 0x3
      11'h46B: dout  = 8'b00000011; // 1131 :   3 - 0x3
      11'h46C: dout  = 8'b00000011; // 1132 :   3 - 0x3
      11'h46D: dout  = 8'b11111111; // 1133 : 255 - 0xff
      11'h46E: dout  = 8'b00000011; // 1134 :   3 - 0x3
      11'h46F: dout  = 8'b00000011; // 1135 :   3 - 0x3
      11'h470: dout  = 8'b10000000; // 1136 : 128 - 0x80 -- Background 0x8e
      11'h471: dout  = 8'b11111111; // 1137 : 255 - 0xff
      11'h472: dout  = 8'b11111111; // 1138 : 255 - 0xff
      11'h473: dout  = 8'b11111111; // 1139 : 255 - 0xff
      11'h474: dout  = 8'b11111111; // 1140 : 255 - 0xff
      11'h475: dout  = 8'b11111111; // 1141 : 255 - 0xff
      11'h476: dout  = 8'b11111111; // 1142 : 255 - 0xff
      11'h477: dout  = 8'b11111111; // 1143 : 255 - 0xff
      11'h478: dout  = 8'b00000011; // 1144 :   3 - 0x3 -- Background 0x8f
      11'h479: dout  = 8'b11111111; // 1145 : 255 - 0xff
      11'h47A: dout  = 8'b11111111; // 1146 : 255 - 0xff
      11'h47B: dout  = 8'b11111111; // 1147 : 255 - 0xff
      11'h47C: dout  = 8'b11111111; // 1148 : 255 - 0xff
      11'h47D: dout  = 8'b11111111; // 1149 : 255 - 0xff
      11'h47E: dout  = 8'b11111111; // 1150 : 255 - 0xff
      11'h47F: dout  = 8'b11111111; // 1151 : 255 - 0xff
      11'h480: dout  = 8'b11111111; // 1152 : 255 - 0xff -- Background 0x90
      11'h481: dout  = 8'b11111111; // 1153 : 255 - 0xff
      11'h482: dout  = 8'b11111111; // 1154 : 255 - 0xff
      11'h483: dout  = 8'b11111111; // 1155 : 255 - 0xff
      11'h484: dout  = 8'b11111111; // 1156 : 255 - 0xff
      11'h485: dout  = 8'b11111111; // 1157 : 255 - 0xff
      11'h486: dout  = 8'b11111111; // 1158 : 255 - 0xff
      11'h487: dout  = 8'b11111111; // 1159 : 255 - 0xff
      11'h488: dout  = 8'b11111111; // 1160 : 255 - 0xff -- Background 0x91
      11'h489: dout  = 8'b11111111; // 1161 : 255 - 0xff
      11'h48A: dout  = 8'b11010101; // 1162 : 213 - 0xd5
      11'h48B: dout  = 8'b10101010; // 1163 : 170 - 0xaa
      11'h48C: dout  = 8'b11010101; // 1164 : 213 - 0xd5
      11'h48D: dout  = 8'b10000000; // 1165 : 128 - 0x80
      11'h48E: dout  = 8'b10000000; // 1166 : 128 - 0x80
      11'h48F: dout  = 8'b11111111; // 1167 : 255 - 0xff
      11'h490: dout  = 8'b11111111; // 1168 : 255 - 0xff -- Background 0x92
      11'h491: dout  = 8'b11111111; // 1169 : 255 - 0xff
      11'h492: dout  = 8'b01010111; // 1170 :  87 - 0x57
      11'h493: dout  = 8'b10101011; // 1171 : 171 - 0xab
      11'h494: dout  = 8'b01010111; // 1172 :  87 - 0x57
      11'h495: dout  = 8'b00000011; // 1173 :   3 - 0x3
      11'h496: dout  = 8'b00000011; // 1174 :   3 - 0x3
      11'h497: dout  = 8'b11111110; // 1175 : 254 - 0xfe
      11'h498: dout  = 8'b11111111; // 1176 : 255 - 0xff -- Background 0x93
      11'h499: dout  = 8'b10101010; // 1177 : 170 - 0xaa
      11'h49A: dout  = 8'b01010101; // 1178 :  85 - 0x55
      11'h49B: dout  = 8'b10101010; // 1179 : 170 - 0xaa
      11'h49C: dout  = 8'b00000000; // 1180 :   0 - 0x0
      11'h49D: dout  = 8'b00000000; // 1181 :   0 - 0x0
      11'h49E: dout  = 8'b11111111; // 1182 : 255 - 0xff
      11'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      11'h4A0: dout  = 8'b11111111; // 1184 : 255 - 0xff -- Background 0x94
      11'h4A1: dout  = 8'b10101111; // 1185 : 175 - 0xaf
      11'h4A2: dout  = 8'b01010111; // 1186 :  87 - 0x57
      11'h4A3: dout  = 8'b10101011; // 1187 : 171 - 0xab
      11'h4A4: dout  = 8'b00001011; // 1188 :  11 - 0xb
      11'h4A5: dout  = 8'b00001011; // 1189 :  11 - 0xb
      11'h4A6: dout  = 8'b11110011; // 1190 : 243 - 0xf3
      11'h4A7: dout  = 8'b00100011; // 1191 :  35 - 0x23
      11'h4A8: dout  = 8'b11111111; // 1192 : 255 - 0xff -- Background 0x95
      11'h4A9: dout  = 8'b11111111; // 1193 : 255 - 0xff
      11'h4AA: dout  = 8'b11111111; // 1194 : 255 - 0xff
      11'h4AB: dout  = 8'b11111111; // 1195 : 255 - 0xff
      11'h4AC: dout  = 8'b11111111; // 1196 : 255 - 0xff
      11'h4AD: dout  = 8'b11111111; // 1197 : 255 - 0xff
      11'h4AE: dout  = 8'b11111111; // 1198 : 255 - 0xff
      11'h4AF: dout  = 8'b11111111; // 1199 : 255 - 0xff
      11'h4B0: dout  = 8'b11111111; // 1200 : 255 - 0xff -- Background 0x96
      11'h4B1: dout  = 8'b11111111; // 1201 : 255 - 0xff
      11'h4B2: dout  = 8'b11111111; // 1202 : 255 - 0xff
      11'h4B3: dout  = 8'b11111111; // 1203 : 255 - 0xff
      11'h4B4: dout  = 8'b11111111; // 1204 : 255 - 0xff
      11'h4B5: dout  = 8'b11111111; // 1205 : 255 - 0xff
      11'h4B6: dout  = 8'b11111111; // 1206 : 255 - 0xff
      11'h4B7: dout  = 8'b11111111; // 1207 : 255 - 0xff
      11'h4B8: dout  = 8'b11111111; // 1208 : 255 - 0xff -- Background 0x97
      11'h4B9: dout  = 8'b11111111; // 1209 : 255 - 0xff
      11'h4BA: dout  = 8'b11111111; // 1210 : 255 - 0xff
      11'h4BB: dout  = 8'b11111111; // 1211 : 255 - 0xff
      11'h4BC: dout  = 8'b11111111; // 1212 : 255 - 0xff
      11'h4BD: dout  = 8'b11111111; // 1213 : 255 - 0xff
      11'h4BE: dout  = 8'b11111111; // 1214 : 255 - 0xff
      11'h4BF: dout  = 8'b11111111; // 1215 : 255 - 0xff
      11'h4C0: dout  = 8'b11111111; // 1216 : 255 - 0xff -- Background 0x98
      11'h4C1: dout  = 8'b11111111; // 1217 : 255 - 0xff
      11'h4C2: dout  = 8'b11111111; // 1218 : 255 - 0xff
      11'h4C3: dout  = 8'b11111111; // 1219 : 255 - 0xff
      11'h4C4: dout  = 8'b11111111; // 1220 : 255 - 0xff
      11'h4C5: dout  = 8'b11111111; // 1221 : 255 - 0xff
      11'h4C6: dout  = 8'b11111111; // 1222 : 255 - 0xff
      11'h4C7: dout  = 8'b11111111; // 1223 : 255 - 0xff
      11'h4C8: dout  = 8'b00000000; // 1224 :   0 - 0x0 -- Background 0x99
      11'h4C9: dout  = 8'b00000000; // 1225 :   0 - 0x0
      11'h4CA: dout  = 8'b00000000; // 1226 :   0 - 0x0
      11'h4CB: dout  = 8'b00000000; // 1227 :   0 - 0x0
      11'h4CC: dout  = 8'b00000000; // 1228 :   0 - 0x0
      11'h4CD: dout  = 8'b00000000; // 1229 :   0 - 0x0
      11'h4CE: dout  = 8'b00000000; // 1230 :   0 - 0x0
      11'h4CF: dout  = 8'b00000000; // 1231 :   0 - 0x0
      11'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Background 0x9a
      11'h4D1: dout  = 8'b00000000; // 1233 :   0 - 0x0
      11'h4D2: dout  = 8'b00000000; // 1234 :   0 - 0x0
      11'h4D3: dout  = 8'b00000000; // 1235 :   0 - 0x0
      11'h4D4: dout  = 8'b00000000; // 1236 :   0 - 0x0
      11'h4D5: dout  = 8'b00000000; // 1237 :   0 - 0x0
      11'h4D6: dout  = 8'b00000000; // 1238 :   0 - 0x0
      11'h4D7: dout  = 8'b00000000; // 1239 :   0 - 0x0
      11'h4D8: dout  = 8'b11111111; // 1240 : 255 - 0xff -- Background 0x9b
      11'h4D9: dout  = 8'b11111111; // 1241 : 255 - 0xff
      11'h4DA: dout  = 8'b11111111; // 1242 : 255 - 0xff
      11'h4DB: dout  = 8'b11111111; // 1243 : 255 - 0xff
      11'h4DC: dout  = 8'b11111111; // 1244 : 255 - 0xff
      11'h4DD: dout  = 8'b11111111; // 1245 : 255 - 0xff
      11'h4DE: dout  = 8'b11111111; // 1246 : 255 - 0xff
      11'h4DF: dout  = 8'b11111111; // 1247 : 255 - 0xff
      11'h4E0: dout  = 8'b11111111; // 1248 : 255 - 0xff -- Background 0x9c
      11'h4E1: dout  = 8'b11111111; // 1249 : 255 - 0xff
      11'h4E2: dout  = 8'b11111111; // 1250 : 255 - 0xff
      11'h4E3: dout  = 8'b11111111; // 1251 : 255 - 0xff
      11'h4E4: dout  = 8'b11111111; // 1252 : 255 - 0xff
      11'h4E5: dout  = 8'b11111111; // 1253 : 255 - 0xff
      11'h4E6: dout  = 8'b11111111; // 1254 : 255 - 0xff
      11'h4E7: dout  = 8'b11111111; // 1255 : 255 - 0xff
      11'h4E8: dout  = 8'b00000000; // 1256 :   0 - 0x0 -- Background 0x9d
      11'h4E9: dout  = 8'b11100000; // 1257 : 224 - 0xe0
      11'h4EA: dout  = 8'b11100000; // 1258 : 224 - 0xe0
      11'h4EB: dout  = 8'b11100000; // 1259 : 224 - 0xe0
      11'h4EC: dout  = 8'b11100000; // 1260 : 224 - 0xe0
      11'h4ED: dout  = 8'b11100000; // 1261 : 224 - 0xe0
      11'h4EE: dout  = 8'b11100000; // 1262 : 224 - 0xe0
      11'h4EF: dout  = 8'b11100000; // 1263 : 224 - 0xe0
      11'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Background 0x9e
      11'h4F1: dout  = 8'b00001111; // 1265 :  15 - 0xf
      11'h4F2: dout  = 8'b00001111; // 1266 :  15 - 0xf
      11'h4F3: dout  = 8'b00001111; // 1267 :  15 - 0xf
      11'h4F4: dout  = 8'b00001111; // 1268 :  15 - 0xf
      11'h4F5: dout  = 8'b00001111; // 1269 :  15 - 0xf
      11'h4F6: dout  = 8'b00001111; // 1270 :  15 - 0xf
      11'h4F7: dout  = 8'b00001111; // 1271 :  15 - 0xf
      11'h4F8: dout  = 8'b01001000; // 1272 :  72 - 0x48 -- Background 0x9f
      11'h4F9: dout  = 8'b01001000; // 1273 :  72 - 0x48
      11'h4FA: dout  = 8'b01101100; // 1274 : 108 - 0x6c
      11'h4FB: dout  = 8'b00000000; // 1275 :   0 - 0x0
      11'h4FC: dout  = 8'b00000000; // 1276 :   0 - 0x0
      11'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      11'h4FE: dout  = 8'b11111110; // 1278 : 254 - 0xfe
      11'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout  = 8'b00000101; // 1280 :   5 - 0x5 -- Background 0xa0
      11'h501: dout  = 8'b00000101; // 1281 :   5 - 0x5
      11'h502: dout  = 8'b11000101; // 1282 : 197 - 0xc5
      11'h503: dout  = 8'b11110101; // 1283 : 245 - 0xf5
      11'h504: dout  = 8'b11110100; // 1284 : 244 - 0xf4
      11'h505: dout  = 8'b00000100; // 1285 :   4 - 0x4
      11'h506: dout  = 8'b00000100; // 1286 :   4 - 0x4
      11'h507: dout  = 8'b00000100; // 1287 :   4 - 0x4
      11'h508: dout  = 8'b01110000; // 1288 : 112 - 0x70 -- Background 0xa1
      11'h509: dout  = 8'b01110000; // 1289 : 112 - 0x70
      11'h50A: dout  = 8'b01110000; // 1290 : 112 - 0x70
      11'h50B: dout  = 8'b01111111; // 1291 : 127 - 0x7f
      11'h50C: dout  = 8'b01111111; // 1292 : 127 - 0x7f
      11'h50D: dout  = 8'b01110000; // 1293 : 112 - 0x70
      11'h50E: dout  = 8'b01110000; // 1294 : 112 - 0x70
      11'h50F: dout  = 8'b01110000; // 1295 : 112 - 0x70
      11'h510: dout  = 8'b00000000; // 1296 :   0 - 0x0 -- Background 0xa2
      11'h511: dout  = 8'b00000000; // 1297 :   0 - 0x0
      11'h512: dout  = 8'b00000000; // 1298 :   0 - 0x0
      11'h513: dout  = 8'b00000000; // 1299 :   0 - 0x0
      11'h514: dout  = 8'b00000000; // 1300 :   0 - 0x0
      11'h515: dout  = 8'b00000000; // 1301 :   0 - 0x0
      11'h516: dout  = 8'b00000000; // 1302 :   0 - 0x0
      11'h517: dout  = 8'b00000000; // 1303 :   0 - 0x0
      11'h518: dout  = 8'b00000000; // 1304 :   0 - 0x0 -- Background 0xa3
      11'h519: dout  = 8'b00000000; // 1305 :   0 - 0x0
      11'h51A: dout  = 8'b00000000; // 1306 :   0 - 0x0
      11'h51B: dout  = 8'b00000000; // 1307 :   0 - 0x0
      11'h51C: dout  = 8'b00000000; // 1308 :   0 - 0x0
      11'h51D: dout  = 8'b00000000; // 1309 :   0 - 0x0
      11'h51E: dout  = 8'b00000000; // 1310 :   0 - 0x0
      11'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      11'h520: dout  = 8'b11111111; // 1312 : 255 - 0xff -- Background 0xa4
      11'h521: dout  = 8'b11111111; // 1313 : 255 - 0xff
      11'h522: dout  = 8'b11111111; // 1314 : 255 - 0xff
      11'h523: dout  = 8'b11111111; // 1315 : 255 - 0xff
      11'h524: dout  = 8'b11111111; // 1316 : 255 - 0xff
      11'h525: dout  = 8'b11111110; // 1317 : 254 - 0xfe
      11'h526: dout  = 8'b10111110; // 1318 : 190 - 0xbe
      11'h527: dout  = 8'b11001110; // 1319 : 206 - 0xce
      11'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- Background 0xa5
      11'h529: dout  = 8'b00000000; // 1321 :   0 - 0x0
      11'h52A: dout  = 8'b00000000; // 1322 :   0 - 0x0
      11'h52B: dout  = 8'b00000000; // 1323 :   0 - 0x0
      11'h52C: dout  = 8'b00000011; // 1324 :   3 - 0x3
      11'h52D: dout  = 8'b00000100; // 1325 :   4 - 0x4
      11'h52E: dout  = 8'b00000100; // 1326 :   4 - 0x4
      11'h52F: dout  = 8'b00000100; // 1327 :   4 - 0x4
      11'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Background 0xa6
      11'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      11'h532: dout  = 8'b01100000; // 1330 :  96 - 0x60
      11'h533: dout  = 8'b00110000; // 1331 :  48 - 0x30
      11'h534: dout  = 8'b00110000; // 1332 :  48 - 0x30
      11'h535: dout  = 8'b10011000; // 1333 : 152 - 0x98
      11'h536: dout  = 8'b10011000; // 1334 : 152 - 0x98
      11'h537: dout  = 8'b10011000; // 1335 : 152 - 0x98
      11'h538: dout  = 8'b00000100; // 1336 :   4 - 0x4 -- Background 0xa7
      11'h539: dout  = 8'b00000100; // 1337 :   4 - 0x4
      11'h53A: dout  = 8'b00000100; // 1338 :   4 - 0x4
      11'h53B: dout  = 8'b00000100; // 1339 :   4 - 0x4
      11'h53C: dout  = 8'b00000100; // 1340 :   4 - 0x4
      11'h53D: dout  = 8'b00000011; // 1341 :   3 - 0x3
      11'h53E: dout  = 8'b00000000; // 1342 :   0 - 0x0
      11'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      11'h540: dout  = 8'b10011000; // 1344 : 152 - 0x98 -- Background 0xa8
      11'h541: dout  = 8'b10011000; // 1345 : 152 - 0x98
      11'h542: dout  = 8'b10011000; // 1346 : 152 - 0x98
      11'h543: dout  = 8'b10011000; // 1347 : 152 - 0x98
      11'h544: dout  = 8'b10011000; // 1348 : 152 - 0x98
      11'h545: dout  = 8'b00110000; // 1349 :  48 - 0x30
      11'h546: dout  = 8'b00110000; // 1350 :  48 - 0x30
      11'h547: dout  = 8'b01100000; // 1351 :  96 - 0x60
      11'h548: dout  = 8'b00001111; // 1352 :  15 - 0xf -- Background 0xa9
      11'h549: dout  = 8'b11101111; // 1353 : 239 - 0xef
      11'h54A: dout  = 8'b11101111; // 1354 : 239 - 0xef
      11'h54B: dout  = 8'b11101111; // 1355 : 239 - 0xef
      11'h54C: dout  = 8'b11101111; // 1356 : 239 - 0xef
      11'h54D: dout  = 8'b11101111; // 1357 : 239 - 0xef
      11'h54E: dout  = 8'b11101111; // 1358 : 239 - 0xef
      11'h54F: dout  = 8'b11100000; // 1359 : 224 - 0xe0
      11'h550: dout  = 8'b11100000; // 1360 : 224 - 0xe0 -- Background 0xaa
      11'h551: dout  = 8'b11101111; // 1361 : 239 - 0xef
      11'h552: dout  = 8'b11101111; // 1362 : 239 - 0xef
      11'h553: dout  = 8'b11101111; // 1363 : 239 - 0xef
      11'h554: dout  = 8'b11101111; // 1364 : 239 - 0xef
      11'h555: dout  = 8'b11101111; // 1365 : 239 - 0xef
      11'h556: dout  = 8'b11101111; // 1366 : 239 - 0xef
      11'h557: dout  = 8'b00001111; // 1367 :  15 - 0xf
      11'h558: dout  = 8'b10000000; // 1368 : 128 - 0x80 -- Background 0xab
      11'h559: dout  = 8'b01000000; // 1369 :  64 - 0x40
      11'h55A: dout  = 8'b00100000; // 1370 :  32 - 0x20
      11'h55B: dout  = 8'b00010000; // 1371 :  16 - 0x10
      11'h55C: dout  = 8'b00001111; // 1372 :  15 - 0xf
      11'h55D: dout  = 8'b00001111; // 1373 :  15 - 0xf
      11'h55E: dout  = 8'b00001111; // 1374 :  15 - 0xf
      11'h55F: dout  = 8'b00001111; // 1375 :  15 - 0xf
      11'h560: dout  = 8'b00001111; // 1376 :  15 - 0xf -- Background 0xac
      11'h561: dout  = 8'b00001111; // 1377 :  15 - 0xf
      11'h562: dout  = 8'b00001111; // 1378 :  15 - 0xf
      11'h563: dout  = 8'b00001111; // 1379 :  15 - 0xf
      11'h564: dout  = 8'b00011111; // 1380 :  31 - 0x1f
      11'h565: dout  = 8'b00111111; // 1381 :  63 - 0x3f
      11'h566: dout  = 8'b01111111; // 1382 : 127 - 0x7f
      11'h567: dout  = 8'b11111111; // 1383 : 255 - 0xff
      11'h568: dout  = 8'b00000001; // 1384 :   1 - 0x1 -- Background 0xad
      11'h569: dout  = 8'b00000011; // 1385 :   3 - 0x3
      11'h56A: dout  = 8'b00000111; // 1386 :   7 - 0x7
      11'h56B: dout  = 8'b00001111; // 1387 :  15 - 0xf
      11'h56C: dout  = 8'b11111111; // 1388 : 255 - 0xff
      11'h56D: dout  = 8'b11111111; // 1389 : 255 - 0xff
      11'h56E: dout  = 8'b11111111; // 1390 : 255 - 0xff
      11'h56F: dout  = 8'b11111111; // 1391 : 255 - 0xff
      11'h570: dout  = 8'b11111111; // 1392 : 255 - 0xff -- Background 0xae
      11'h571: dout  = 8'b11111111; // 1393 : 255 - 0xff
      11'h572: dout  = 8'b11111111; // 1394 : 255 - 0xff
      11'h573: dout  = 8'b11111111; // 1395 : 255 - 0xff
      11'h574: dout  = 8'b11111111; // 1396 : 255 - 0xff
      11'h575: dout  = 8'b11111111; // 1397 : 255 - 0xff
      11'h576: dout  = 8'b11111111; // 1398 : 255 - 0xff
      11'h577: dout  = 8'b11111111; // 1399 : 255 - 0xff
      11'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Background 0xaf
      11'h579: dout  = 8'b00000000; // 1401 :   0 - 0x0
      11'h57A: dout  = 8'b00000000; // 1402 :   0 - 0x0
      11'h57B: dout  = 8'b00000000; // 1403 :   0 - 0x0
      11'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      11'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      11'h57E: dout  = 8'b00000000; // 1406 :   0 - 0x0
      11'h57F: dout  = 8'b00000000; // 1407 :   0 - 0x0
      11'h580: dout  = 8'b00011111; // 1408 :  31 - 0x1f -- Background 0xb0
      11'h581: dout  = 8'b00100000; // 1409 :  32 - 0x20
      11'h582: dout  = 8'b01000000; // 1410 :  64 - 0x40
      11'h583: dout  = 8'b01000000; // 1411 :  64 - 0x40
      11'h584: dout  = 8'b01000000; // 1412 :  64 - 0x40
      11'h585: dout  = 8'b10000000; // 1413 : 128 - 0x80
      11'h586: dout  = 8'b10000010; // 1414 : 130 - 0x82
      11'h587: dout  = 8'b10000010; // 1415 : 130 - 0x82
      11'h588: dout  = 8'b10000010; // 1416 : 130 - 0x82 -- Background 0xb1
      11'h589: dout  = 8'b10000000; // 1417 : 128 - 0x80
      11'h58A: dout  = 8'b10100000; // 1418 : 160 - 0xa0
      11'h58B: dout  = 8'b01000100; // 1419 :  68 - 0x44
      11'h58C: dout  = 8'b01000011; // 1420 :  67 - 0x43
      11'h58D: dout  = 8'b01000000; // 1421 :  64 - 0x40
      11'h58E: dout  = 8'b00100001; // 1422 :  33 - 0x21
      11'h58F: dout  = 8'b00011110; // 1423 :  30 - 0x1e
      11'h590: dout  = 8'b11111000; // 1424 : 248 - 0xf8 -- Background 0xb2
      11'h591: dout  = 8'b00000100; // 1425 :   4 - 0x4
      11'h592: dout  = 8'b00000010; // 1426 :   2 - 0x2
      11'h593: dout  = 8'b00000010; // 1427 :   2 - 0x2
      11'h594: dout  = 8'b00000010; // 1428 :   2 - 0x2
      11'h595: dout  = 8'b00000001; // 1429 :   1 - 0x1
      11'h596: dout  = 8'b01000001; // 1430 :  65 - 0x41
      11'h597: dout  = 8'b01000001; // 1431 :  65 - 0x41
      11'h598: dout  = 8'b01000001; // 1432 :  65 - 0x41 -- Background 0xb3
      11'h599: dout  = 8'b00000001; // 1433 :   1 - 0x1
      11'h59A: dout  = 8'b00000101; // 1434 :   5 - 0x5
      11'h59B: dout  = 8'b00100010; // 1435 :  34 - 0x22
      11'h59C: dout  = 8'b11000010; // 1436 : 194 - 0xc2
      11'h59D: dout  = 8'b00000010; // 1437 :   2 - 0x2
      11'h59E: dout  = 8'b10000100; // 1438 : 132 - 0x84
      11'h59F: dout  = 8'b01111000; // 1439 : 120 - 0x78
      11'h5A0: dout  = 8'b10000000; // 1440 : 128 - 0x80 -- Background 0xb4
      11'h5A1: dout  = 8'b01111111; // 1441 : 127 - 0x7f
      11'h5A2: dout  = 8'b01111111; // 1442 : 127 - 0x7f
      11'h5A3: dout  = 8'b01111111; // 1443 : 127 - 0x7f
      11'h5A4: dout  = 8'b01111111; // 1444 : 127 - 0x7f
      11'h5A5: dout  = 8'b01111111; // 1445 : 127 - 0x7f
      11'h5A6: dout  = 8'b01111111; // 1446 : 127 - 0x7f
      11'h5A7: dout  = 8'b01111111; // 1447 : 127 - 0x7f
      11'h5A8: dout  = 8'b01100001; // 1448 :  97 - 0x61 -- Background 0xb5
      11'h5A9: dout  = 8'b11011111; // 1449 : 223 - 0xdf
      11'h5AA: dout  = 8'b11011111; // 1450 : 223 - 0xdf
      11'h5AB: dout  = 8'b11011111; // 1451 : 223 - 0xdf
      11'h5AC: dout  = 8'b11011111; // 1452 : 223 - 0xdf
      11'h5AD: dout  = 8'b11111111; // 1453 : 255 - 0xff
      11'h5AE: dout  = 8'b11000001; // 1454 : 193 - 0xc1
      11'h5AF: dout  = 8'b11011111; // 1455 : 223 - 0xdf
      11'h5B0: dout  = 8'b01111111; // 1456 : 127 - 0x7f -- Background 0xb6
      11'h5B1: dout  = 8'b01111111; // 1457 : 127 - 0x7f
      11'h5B2: dout  = 8'b11111111; // 1458 : 255 - 0xff
      11'h5B3: dout  = 8'b00111111; // 1459 :  63 - 0x3f
      11'h5B4: dout  = 8'b01001111; // 1460 :  79 - 0x4f
      11'h5B5: dout  = 8'b01110001; // 1461 : 113 - 0x71
      11'h5B6: dout  = 8'b01111111; // 1462 : 127 - 0x7f
      11'h5B7: dout  = 8'b11111111; // 1463 : 255 - 0xff
      11'h5B8: dout  = 8'b11011111; // 1464 : 223 - 0xdf -- Background 0xb7
      11'h5B9: dout  = 8'b11011111; // 1465 : 223 - 0xdf
      11'h5BA: dout  = 8'b10111111; // 1466 : 191 - 0xbf
      11'h5BB: dout  = 8'b10111111; // 1467 : 191 - 0xbf
      11'h5BC: dout  = 8'b01111111; // 1468 : 127 - 0x7f
      11'h5BD: dout  = 8'b01111111; // 1469 : 127 - 0x7f
      11'h5BE: dout  = 8'b01111111; // 1470 : 127 - 0x7f
      11'h5BF: dout  = 8'b01111111; // 1471 : 127 - 0x7f
      11'h5C0: dout  = 8'b00000000; // 1472 :   0 - 0x0 -- Background 0xb8
      11'h5C1: dout  = 8'b00000000; // 1473 :   0 - 0x0
      11'h5C2: dout  = 8'b00000011; // 1474 :   3 - 0x3
      11'h5C3: dout  = 8'b00001100; // 1475 :  12 - 0xc
      11'h5C4: dout  = 8'b00010000; // 1476 :  16 - 0x10
      11'h5C5: dout  = 8'b00100000; // 1477 :  32 - 0x20
      11'h5C6: dout  = 8'b01000000; // 1478 :  64 - 0x40
      11'h5C7: dout  = 8'b01000000; // 1479 :  64 - 0x40
      11'h5C8: dout  = 8'b00000000; // 1480 :   0 - 0x0 -- Background 0xb9
      11'h5C9: dout  = 8'b00000000; // 1481 :   0 - 0x0
      11'h5CA: dout  = 8'b11000000; // 1482 : 192 - 0xc0
      11'h5CB: dout  = 8'b00110000; // 1483 :  48 - 0x30
      11'h5CC: dout  = 8'b00001000; // 1484 :   8 - 0x8
      11'h5CD: dout  = 8'b00000100; // 1485 :   4 - 0x4
      11'h5CE: dout  = 8'b00000010; // 1486 :   2 - 0x2
      11'h5CF: dout  = 8'b00000010; // 1487 :   2 - 0x2
      11'h5D0: dout  = 8'b10000000; // 1488 : 128 - 0x80 -- Background 0xba
      11'h5D1: dout  = 8'b10000000; // 1489 : 128 - 0x80
      11'h5D2: dout  = 8'b10000000; // 1490 : 128 - 0x80
      11'h5D3: dout  = 8'b10000000; // 1491 : 128 - 0x80
      11'h5D4: dout  = 8'b10000000; // 1492 : 128 - 0x80
      11'h5D5: dout  = 8'b10000000; // 1493 : 128 - 0x80
      11'h5D6: dout  = 8'b10000000; // 1494 : 128 - 0x80
      11'h5D7: dout  = 8'b10000000; // 1495 : 128 - 0x80
      11'h5D8: dout  = 8'b00000001; // 1496 :   1 - 0x1 -- Background 0xbb
      11'h5D9: dout  = 8'b00000001; // 1497 :   1 - 0x1
      11'h5DA: dout  = 8'b00000001; // 1498 :   1 - 0x1
      11'h5DB: dout  = 8'b00000001; // 1499 :   1 - 0x1
      11'h5DC: dout  = 8'b00000001; // 1500 :   1 - 0x1
      11'h5DD: dout  = 8'b00000001; // 1501 :   1 - 0x1
      11'h5DE: dout  = 8'b00000001; // 1502 :   1 - 0x1
      11'h5DF: dout  = 8'b00000001; // 1503 :   1 - 0x1
      11'h5E0: dout  = 8'b01000000; // 1504 :  64 - 0x40 -- Background 0xbc
      11'h5E1: dout  = 8'b01000000; // 1505 :  64 - 0x40
      11'h5E2: dout  = 8'b01000000; // 1506 :  64 - 0x40
      11'h5E3: dout  = 8'b00100000; // 1507 :  32 - 0x20
      11'h5E4: dout  = 8'b00110000; // 1508 :  48 - 0x30
      11'h5E5: dout  = 8'b00011100; // 1509 :  28 - 0x1c
      11'h5E6: dout  = 8'b00001111; // 1510 :  15 - 0xf
      11'h5E7: dout  = 8'b00000111; // 1511 :   7 - 0x7
      11'h5E8: dout  = 8'b00000010; // 1512 :   2 - 0x2 -- Background 0xbd
      11'h5E9: dout  = 8'b00000010; // 1513 :   2 - 0x2
      11'h5EA: dout  = 8'b00000010; // 1514 :   2 - 0x2
      11'h5EB: dout  = 8'b00000100; // 1515 :   4 - 0x4
      11'h5EC: dout  = 8'b00001100; // 1516 :  12 - 0xc
      11'h5ED: dout  = 8'b00111000; // 1517 :  56 - 0x38
      11'h5EE: dout  = 8'b11110000; // 1518 : 240 - 0xf0
      11'h5EF: dout  = 8'b11110000; // 1519 : 240 - 0xf0
      11'h5F0: dout  = 8'b00001000; // 1520 :   8 - 0x8 -- Background 0xbe
      11'h5F1: dout  = 8'b00001000; // 1521 :   8 - 0x8
      11'h5F2: dout  = 8'b00001000; // 1522 :   8 - 0x8
      11'h5F3: dout  = 8'b00001000; // 1523 :   8 - 0x8
      11'h5F4: dout  = 8'b00001000; // 1524 :   8 - 0x8
      11'h5F5: dout  = 8'b00001100; // 1525 :  12 - 0xc
      11'h5F6: dout  = 8'b00000101; // 1526 :   5 - 0x5
      11'h5F7: dout  = 8'b00001010; // 1527 :  10 - 0xa
      11'h5F8: dout  = 8'b00010000; // 1528 :  16 - 0x10 -- Background 0xbf
      11'h5F9: dout  = 8'b01010000; // 1529 :  80 - 0x50
      11'h5FA: dout  = 8'b01010000; // 1530 :  80 - 0x50
      11'h5FB: dout  = 8'b01010000; // 1531 :  80 - 0x50
      11'h5FC: dout  = 8'b01010000; // 1532 :  80 - 0x50
      11'h5FD: dout  = 8'b00110000; // 1533 :  48 - 0x30
      11'h5FE: dout  = 8'b10100000; // 1534 : 160 - 0xa0
      11'h5FF: dout  = 8'b01010000; // 1535 :  80 - 0x50
      11'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Background 0xc0
      11'h601: dout  = 8'b01000001; // 1537 :  65 - 0x41
      11'h602: dout  = 8'b00100010; // 1538 :  34 - 0x22
      11'h603: dout  = 8'b00100010; // 1539 :  34 - 0x22
      11'h604: dout  = 8'b00011100; // 1540 :  28 - 0x1c
      11'h605: dout  = 8'b00000000; // 1541 :   0 - 0x0
      11'h606: dout  = 8'b00000000; // 1542 :   0 - 0x0
      11'h607: dout  = 8'b00000000; // 1543 :   0 - 0x0
      11'h608: dout  = 8'b11100011; // 1544 : 227 - 0xe3 -- Background 0xc1
      11'h609: dout  = 8'b00010100; // 1545 :  20 - 0x14
      11'h60A: dout  = 8'b00111110; // 1546 :  62 - 0x3e
      11'h60B: dout  = 8'b00111110; // 1547 :  62 - 0x3e
      11'h60C: dout  = 8'b00111110; // 1548 :  62 - 0x3e
      11'h60D: dout  = 8'b00111110; // 1549 :  62 - 0x3e
      11'h60E: dout  = 8'b00010100; // 1550 :  20 - 0x14
      11'h60F: dout  = 8'b11100011; // 1551 : 227 - 0xe3
      11'h610: dout  = 8'b11111111; // 1552 : 255 - 0xff -- Background 0xc2
      11'h611: dout  = 8'b11111111; // 1553 : 255 - 0xff
      11'h612: dout  = 8'b11111000; // 1554 : 248 - 0xf8
      11'h613: dout  = 8'b11110000; // 1555 : 240 - 0xf0
      11'h614: dout  = 8'b11110000; // 1556 : 240 - 0xf0
      11'h615: dout  = 8'b11100000; // 1557 : 224 - 0xe0
      11'h616: dout  = 8'b11100000; // 1558 : 224 - 0xe0
      11'h617: dout  = 8'b11100000; // 1559 : 224 - 0xe0
      11'h618: dout  = 8'b11111111; // 1560 : 255 - 0xff -- Background 0xc3
      11'h619: dout  = 8'b11111111; // 1561 : 255 - 0xff
      11'h61A: dout  = 8'b01111111; // 1562 : 127 - 0x7f
      11'h61B: dout  = 8'b00111111; // 1563 :  63 - 0x3f
      11'h61C: dout  = 8'b00111111; // 1564 :  63 - 0x3f
      11'h61D: dout  = 8'b10011111; // 1565 : 159 - 0x9f
      11'h61E: dout  = 8'b10011111; // 1566 : 159 - 0x9f
      11'h61F: dout  = 8'b10011111; // 1567 : 159 - 0x9f
      11'h620: dout  = 8'b11100000; // 1568 : 224 - 0xe0 -- Background 0xc4
      11'h621: dout  = 8'b11100000; // 1569 : 224 - 0xe0
      11'h622: dout  = 8'b11100000; // 1570 : 224 - 0xe0
      11'h623: dout  = 8'b11100000; // 1571 : 224 - 0xe0
      11'h624: dout  = 8'b11100000; // 1572 : 224 - 0xe0
      11'h625: dout  = 8'b11110011; // 1573 : 243 - 0xf3
      11'h626: dout  = 8'b11110000; // 1574 : 240 - 0xf0
      11'h627: dout  = 8'b11111000; // 1575 : 248 - 0xf8
      11'h628: dout  = 8'b10011111; // 1576 : 159 - 0x9f -- Background 0xc5
      11'h629: dout  = 8'b10011111; // 1577 : 159 - 0x9f
      11'h62A: dout  = 8'b10011111; // 1578 : 159 - 0x9f
      11'h62B: dout  = 8'b10011111; // 1579 : 159 - 0x9f
      11'h62C: dout  = 8'b10011111; // 1580 : 159 - 0x9f
      11'h62D: dout  = 8'b00111111; // 1581 :  63 - 0x3f
      11'h62E: dout  = 8'b00111111; // 1582 :  63 - 0x3f
      11'h62F: dout  = 8'b01111111; // 1583 : 127 - 0x7f
      11'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Background 0xc6
      11'h631: dout  = 8'b01110000; // 1585 : 112 - 0x70
      11'h632: dout  = 8'b00011111; // 1586 :  31 - 0x1f
      11'h633: dout  = 8'b00010000; // 1587 :  16 - 0x10
      11'h634: dout  = 8'b01110000; // 1588 : 112 - 0x70
      11'h635: dout  = 8'b01111111; // 1589 : 127 - 0x7f
      11'h636: dout  = 8'b01111111; // 1590 : 127 - 0x7f
      11'h637: dout  = 8'b01111111; // 1591 : 127 - 0x7f
      11'h638: dout  = 8'b00000000; // 1592 :   0 - 0x0 -- Background 0xc7
      11'h639: dout  = 8'b00000011; // 1593 :   3 - 0x3
      11'h63A: dout  = 8'b11111000; // 1594 : 248 - 0xf8
      11'h63B: dout  = 8'b00000000; // 1595 :   0 - 0x0
      11'h63C: dout  = 8'b00000011; // 1596 :   3 - 0x3
      11'h63D: dout  = 8'b11111011; // 1597 : 251 - 0xfb
      11'h63E: dout  = 8'b11111011; // 1598 : 251 - 0xfb
      11'h63F: dout  = 8'b11111011; // 1599 : 251 - 0xfb
      11'h640: dout  = 8'b01111100; // 1600 : 124 - 0x7c -- Background 0xc8
      11'h641: dout  = 8'b01111011; // 1601 : 123 - 0x7b
      11'h642: dout  = 8'b01110110; // 1602 : 118 - 0x76
      11'h643: dout  = 8'b01110101; // 1603 : 117 - 0x75
      11'h644: dout  = 8'b01110101; // 1604 : 117 - 0x75
      11'h645: dout  = 8'b01110111; // 1605 : 119 - 0x77
      11'h646: dout  = 8'b00010111; // 1606 :  23 - 0x17
      11'h647: dout  = 8'b01100111; // 1607 : 103 - 0x67
      11'h648: dout  = 8'b00111011; // 1608 :  59 - 0x3b -- Background 0xc9
      11'h649: dout  = 8'b11111011; // 1609 : 251 - 0xfb
      11'h64A: dout  = 8'b01111011; // 1610 : 123 - 0x7b
      11'h64B: dout  = 8'b11111011; // 1611 : 251 - 0xfb
      11'h64C: dout  = 8'b11111011; // 1612 : 251 - 0xfb
      11'h64D: dout  = 8'b11110011; // 1613 : 243 - 0xf3
      11'h64E: dout  = 8'b11111000; // 1614 : 248 - 0xf8
      11'h64F: dout  = 8'b11110011; // 1615 : 243 - 0xf3
      11'h650: dout  = 8'b00001111; // 1616 :  15 - 0xf -- Background 0xca
      11'h651: dout  = 8'b00001111; // 1617 :  15 - 0xf
      11'h652: dout  = 8'b00011111; // 1618 :  31 - 0x1f
      11'h653: dout  = 8'b00011111; // 1619 :  31 - 0x1f
      11'h654: dout  = 8'b00111111; // 1620 :  63 - 0x3f
      11'h655: dout  = 8'b00111100; // 1621 :  60 - 0x3c
      11'h656: dout  = 8'b01111000; // 1622 : 120 - 0x78
      11'h657: dout  = 8'b01111010; // 1623 : 122 - 0x7a
      11'h658: dout  = 8'b11111000; // 1624 : 248 - 0xf8 -- Background 0xcb
      11'h659: dout  = 8'b11111000; // 1625 : 248 - 0xf8
      11'h65A: dout  = 8'b11111100; // 1626 : 252 - 0xfc
      11'h65B: dout  = 8'b11111100; // 1627 : 252 - 0xfc
      11'h65C: dout  = 8'b11111110; // 1628 : 254 - 0xfe
      11'h65D: dout  = 8'b00111110; // 1629 :  62 - 0x3e
      11'h65E: dout  = 8'b00011110; // 1630 :  30 - 0x1e
      11'h65F: dout  = 8'b01011111; // 1631 :  95 - 0x5f
      11'h660: dout  = 8'b01110110; // 1632 : 118 - 0x76 -- Background 0xcc
      11'h661: dout  = 8'b01110110; // 1633 : 118 - 0x76
      11'h662: dout  = 8'b01110110; // 1634 : 118 - 0x76
      11'h663: dout  = 8'b01110000; // 1635 : 112 - 0x70
      11'h664: dout  = 8'b01111101; // 1636 : 125 - 0x7d
      11'h665: dout  = 8'b01111100; // 1637 : 124 - 0x7c
      11'h666: dout  = 8'b01111111; // 1638 : 127 - 0x7f
      11'h667: dout  = 8'b01111111; // 1639 : 127 - 0x7f
      11'h668: dout  = 8'b01101111; // 1640 : 111 - 0x6f -- Background 0xcd
      11'h669: dout  = 8'b01101111; // 1641 : 111 - 0x6f
      11'h66A: dout  = 8'b01101111; // 1642 : 111 - 0x6f
      11'h66B: dout  = 8'b00001111; // 1643 :  15 - 0xf
      11'h66C: dout  = 8'b10111111; // 1644 : 191 - 0xbf
      11'h66D: dout  = 8'b00111111; // 1645 :  63 - 0x3f
      11'h66E: dout  = 8'b11111111; // 1646 : 255 - 0xff
      11'h66F: dout  = 8'b11111111; // 1647 : 255 - 0xff
      11'h670: dout  = 8'b00111100; // 1648 :  60 - 0x3c -- Background 0xce
      11'h671: dout  = 8'b01111110; // 1649 : 126 - 0x7e
      11'h672: dout  = 8'b01111110; // 1650 : 126 - 0x7e
      11'h673: dout  = 8'b11111111; // 1651 : 255 - 0xff
      11'h674: dout  = 8'b11111111; // 1652 : 255 - 0xff
      11'h675: dout  = 8'b11111111; // 1653 : 255 - 0xff
      11'h676: dout  = 8'b01000010; // 1654 :  66 - 0x42
      11'h677: dout  = 8'b00000000; // 1655 :   0 - 0x0
      11'h678: dout  = 8'b00000000; // 1656 :   0 - 0x0 -- Background 0xcf
      11'h679: dout  = 8'b00000000; // 1657 :   0 - 0x0
      11'h67A: dout  = 8'b00000000; // 1658 :   0 - 0x0
      11'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      11'h67C: dout  = 8'b00000000; // 1660 :   0 - 0x0
      11'h67D: dout  = 8'b00000000; // 1661 :   0 - 0x0
      11'h67E: dout  = 8'b00000000; // 1662 :   0 - 0x0
      11'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      11'h680: dout  = 8'b11110000; // 1664 : 240 - 0xf0 -- Background 0xd0
      11'h681: dout  = 8'b11100000; // 1665 : 224 - 0xe0
      11'h682: dout  = 8'b11100000; // 1666 : 224 - 0xe0
      11'h683: dout  = 8'b11000000; // 1667 : 192 - 0xc0
      11'h684: dout  = 8'b11000000; // 1668 : 192 - 0xc0
      11'h685: dout  = 8'b10000000; // 1669 : 128 - 0x80
      11'h686: dout  = 8'b10000000; // 1670 : 128 - 0x80
      11'h687: dout  = 8'b10000000; // 1671 : 128 - 0x80
      11'h688: dout  = 8'b00001111; // 1672 :  15 - 0xf -- Background 0xd1
      11'h689: dout  = 8'b00000111; // 1673 :   7 - 0x7
      11'h68A: dout  = 8'b00000111; // 1674 :   7 - 0x7
      11'h68B: dout  = 8'b00000011; // 1675 :   3 - 0x3
      11'h68C: dout  = 8'b00000011; // 1676 :   3 - 0x3
      11'h68D: dout  = 8'b00000001; // 1677 :   1 - 0x1
      11'h68E: dout  = 8'b00000001; // 1678 :   1 - 0x1
      11'h68F: dout  = 8'b00000001; // 1679 :   1 - 0x1
      11'h690: dout  = 8'b10000000; // 1680 : 128 - 0x80 -- Background 0xd2
      11'h691: dout  = 8'b10000000; // 1681 : 128 - 0x80
      11'h692: dout  = 8'b11000000; // 1682 : 192 - 0xc0
      11'h693: dout  = 8'b11000000; // 1683 : 192 - 0xc0
      11'h694: dout  = 8'b11100000; // 1684 : 224 - 0xe0
      11'h695: dout  = 8'b11111000; // 1685 : 248 - 0xf8
      11'h696: dout  = 8'b11111110; // 1686 : 254 - 0xfe
      11'h697: dout  = 8'b11111111; // 1687 : 255 - 0xff
      11'h698: dout  = 8'b11111111; // 1688 : 255 - 0xff -- Background 0xd3
      11'h699: dout  = 8'b01111111; // 1689 : 127 - 0x7f
      11'h69A: dout  = 8'b00011111; // 1690 :  31 - 0x1f
      11'h69B: dout  = 8'b00000111; // 1691 :   7 - 0x7
      11'h69C: dout  = 8'b00000011; // 1692 :   3 - 0x3
      11'h69D: dout  = 8'b00000011; // 1693 :   3 - 0x3
      11'h69E: dout  = 8'b00000001; // 1694 :   1 - 0x1
      11'h69F: dout  = 8'b10000001; // 1695 : 129 - 0x81
      11'h6A0: dout  = 8'b10000000; // 1696 : 128 - 0x80 -- Background 0xd4
      11'h6A1: dout  = 8'b10000000; // 1697 : 128 - 0x80
      11'h6A2: dout  = 8'b10000000; // 1698 : 128 - 0x80
      11'h6A3: dout  = 8'b11000000; // 1699 : 192 - 0xc0
      11'h6A4: dout  = 8'b11000000; // 1700 : 192 - 0xc0
      11'h6A5: dout  = 8'b11100000; // 1701 : 224 - 0xe0
      11'h6A6: dout  = 8'b11100000; // 1702 : 224 - 0xe0
      11'h6A7: dout  = 8'b11110000; // 1703 : 240 - 0xf0
      11'h6A8: dout  = 8'b00000001; // 1704 :   1 - 0x1 -- Background 0xd5
      11'h6A9: dout  = 8'b00000001; // 1705 :   1 - 0x1
      11'h6AA: dout  = 8'b00000001; // 1706 :   1 - 0x1
      11'h6AB: dout  = 8'b00000011; // 1707 :   3 - 0x3
      11'h6AC: dout  = 8'b00000011; // 1708 :   3 - 0x3
      11'h6AD: dout  = 8'b00000111; // 1709 :   7 - 0x7
      11'h6AE: dout  = 8'b00000111; // 1710 :   7 - 0x7
      11'h6AF: dout  = 8'b00001111; // 1711 :  15 - 0xf
      11'h6B0: dout  = 8'b11111111; // 1712 : 255 - 0xff -- Background 0xd6
      11'h6B1: dout  = 8'b11111111; // 1713 : 255 - 0xff
      11'h6B2: dout  = 8'b11111111; // 1714 : 255 - 0xff
      11'h6B3: dout  = 8'b11111111; // 1715 : 255 - 0xff
      11'h6B4: dout  = 8'b11111111; // 1716 : 255 - 0xff
      11'h6B5: dout  = 8'b11111111; // 1717 : 255 - 0xff
      11'h6B6: dout  = 8'b11111111; // 1718 : 255 - 0xff
      11'h6B7: dout  = 8'b11111111; // 1719 : 255 - 0xff
      11'h6B8: dout  = 8'b11111111; // 1720 : 255 - 0xff -- Background 0xd7
      11'h6B9: dout  = 8'b11111111; // 1721 : 255 - 0xff
      11'h6BA: dout  = 8'b11111111; // 1722 : 255 - 0xff
      11'h6BB: dout  = 8'b11111111; // 1723 : 255 - 0xff
      11'h6BC: dout  = 8'b11111111; // 1724 : 255 - 0xff
      11'h6BD: dout  = 8'b11111111; // 1725 : 255 - 0xff
      11'h6BE: dout  = 8'b11111111; // 1726 : 255 - 0xff
      11'h6BF: dout  = 8'b11111111; // 1727 : 255 - 0xff
      11'h6C0: dout  = 8'b10000001; // 1728 : 129 - 0x81 -- Background 0xd8
      11'h6C1: dout  = 8'b10000001; // 1729 : 129 - 0x81
      11'h6C2: dout  = 8'b10000001; // 1730 : 129 - 0x81
      11'h6C3: dout  = 8'b10000001; // 1731 : 129 - 0x81
      11'h6C4: dout  = 8'b10000001; // 1732 : 129 - 0x81
      11'h6C5: dout  = 8'b10000001; // 1733 : 129 - 0x81
      11'h6C6: dout  = 8'b10000001; // 1734 : 129 - 0x81
      11'h6C7: dout  = 8'b10000001; // 1735 : 129 - 0x81
      11'h6C8: dout  = 8'b00000001; // 1736 :   1 - 0x1 -- Background 0xd9
      11'h6C9: dout  = 8'b00000001; // 1737 :   1 - 0x1
      11'h6CA: dout  = 8'b00000001; // 1738 :   1 - 0x1
      11'h6CB: dout  = 8'b00000011; // 1739 :   3 - 0x3
      11'h6CC: dout  = 8'b00000011; // 1740 :   3 - 0x3
      11'h6CD: dout  = 8'b00000111; // 1741 :   7 - 0x7
      11'h6CE: dout  = 8'b00000111; // 1742 :   7 - 0x7
      11'h6CF: dout  = 8'b00001111; // 1743 :  15 - 0xf
      11'h6D0: dout  = 8'b00000001; // 1744 :   1 - 0x1 -- Background 0xda
      11'h6D1: dout  = 8'b00000001; // 1745 :   1 - 0x1
      11'h6D2: dout  = 8'b00000001; // 1746 :   1 - 0x1
      11'h6D3: dout  = 8'b00000001; // 1747 :   1 - 0x1
      11'h6D4: dout  = 8'b00000001; // 1748 :   1 - 0x1
      11'h6D5: dout  = 8'b00000001; // 1749 :   1 - 0x1
      11'h6D6: dout  = 8'b00000001; // 1750 :   1 - 0x1
      11'h6D7: dout  = 8'b00000001; // 1751 :   1 - 0x1
      11'h6D8: dout  = 8'b10000001; // 1752 : 129 - 0x81 -- Background 0xdb
      11'h6D9: dout  = 8'b10000001; // 1753 : 129 - 0x81
      11'h6DA: dout  = 8'b10000001; // 1754 : 129 - 0x81
      11'h6DB: dout  = 8'b10000001; // 1755 : 129 - 0x81
      11'h6DC: dout  = 8'b10000001; // 1756 : 129 - 0x81
      11'h6DD: dout  = 8'b10000001; // 1757 : 129 - 0x81
      11'h6DE: dout  = 8'b10000001; // 1758 : 129 - 0x81
      11'h6DF: dout  = 8'b10000001; // 1759 : 129 - 0x81
      11'h6E0: dout  = 8'b11111111; // 1760 : 255 - 0xff -- Background 0xdc
      11'h6E1: dout  = 8'b00000011; // 1761 :   3 - 0x3
      11'h6E2: dout  = 8'b00000011; // 1762 :   3 - 0x3
      11'h6E3: dout  = 8'b00000011; // 1763 :   3 - 0x3
      11'h6E4: dout  = 8'b00000011; // 1764 :   3 - 0x3
      11'h6E5: dout  = 8'b00000011; // 1765 :   3 - 0x3
      11'h6E6: dout  = 8'b00000011; // 1766 :   3 - 0x3
      11'h6E7: dout  = 8'b11111111; // 1767 : 255 - 0xff
      11'h6E8: dout  = 8'b11111111; // 1768 : 255 - 0xff -- Background 0xdd
      11'h6E9: dout  = 8'b11111111; // 1769 : 255 - 0xff
      11'h6EA: dout  = 8'b11111111; // 1770 : 255 - 0xff
      11'h6EB: dout  = 8'b11111111; // 1771 : 255 - 0xff
      11'h6EC: dout  = 8'b11111111; // 1772 : 255 - 0xff
      11'h6ED: dout  = 8'b11111111; // 1773 : 255 - 0xff
      11'h6EE: dout  = 8'b11111111; // 1774 : 255 - 0xff
      11'h6EF: dout  = 8'b11111111; // 1775 : 255 - 0xff
      11'h6F0: dout  = 8'b10000000; // 1776 : 128 - 0x80 -- Background 0xde
      11'h6F1: dout  = 8'b10000000; // 1777 : 128 - 0x80
      11'h6F2: dout  = 8'b10000000; // 1778 : 128 - 0x80
      11'h6F3: dout  = 8'b10000000; // 1779 : 128 - 0x80
      11'h6F4: dout  = 8'b10000000; // 1780 : 128 - 0x80
      11'h6F5: dout  = 8'b10000000; // 1781 : 128 - 0x80
      11'h6F6: dout  = 8'b10000000; // 1782 : 128 - 0x80
      11'h6F7: dout  = 8'b10000000; // 1783 : 128 - 0x80
      11'h6F8: dout  = 8'b00000001; // 1784 :   1 - 0x1 -- Background 0xdf
      11'h6F9: dout  = 8'b00000001; // 1785 :   1 - 0x1
      11'h6FA: dout  = 8'b00000001; // 1786 :   1 - 0x1
      11'h6FB: dout  = 8'b00000011; // 1787 :   3 - 0x3
      11'h6FC: dout  = 8'b00000111; // 1788 :   7 - 0x7
      11'h6FD: dout  = 8'b00000011; // 1789 :   3 - 0x3
      11'h6FE: dout  = 8'b00000001; // 1790 :   1 - 0x1
      11'h6FF: dout  = 8'b00000001; // 1791 :   1 - 0x1
      11'h700: dout  = 8'b10000001; // 1792 : 129 - 0x81 -- Background 0xe0
      11'h701: dout  = 8'b10000001; // 1793 : 129 - 0x81
      11'h702: dout  = 8'b10000001; // 1794 : 129 - 0x81
      11'h703: dout  = 8'b10000001; // 1795 : 129 - 0x81
      11'h704: dout  = 8'b10000001; // 1796 : 129 - 0x81
      11'h705: dout  = 8'b10000001; // 1797 : 129 - 0x81
      11'h706: dout  = 8'b10000001; // 1798 : 129 - 0x81
      11'h707: dout  = 8'b10000001; // 1799 : 129 - 0x81
      11'h708: dout  = 8'b11111111; // 1800 : 255 - 0xff -- Background 0xe1
      11'h709: dout  = 8'b11111111; // 1801 : 255 - 0xff
      11'h70A: dout  = 8'b11111111; // 1802 : 255 - 0xff
      11'h70B: dout  = 8'b11111111; // 1803 : 255 - 0xff
      11'h70C: dout  = 8'b11111111; // 1804 : 255 - 0xff
      11'h70D: dout  = 8'b11111111; // 1805 : 255 - 0xff
      11'h70E: dout  = 8'b11111111; // 1806 : 255 - 0xff
      11'h70F: dout  = 8'b11111111; // 1807 : 255 - 0xff
      11'h710: dout  = 8'b11111111; // 1808 : 255 - 0xff -- Background 0xe2
      11'h711: dout  = 8'b11111111; // 1809 : 255 - 0xff
      11'h712: dout  = 8'b11111111; // 1810 : 255 - 0xff
      11'h713: dout  = 8'b11111111; // 1811 : 255 - 0xff
      11'h714: dout  = 8'b11111111; // 1812 : 255 - 0xff
      11'h715: dout  = 8'b11111111; // 1813 : 255 - 0xff
      11'h716: dout  = 8'b11111111; // 1814 : 255 - 0xff
      11'h717: dout  = 8'b11111111; // 1815 : 255 - 0xff
      11'h718: dout  = 8'b10000001; // 1816 : 129 - 0x81 -- Background 0xe3
      11'h719: dout  = 8'b10000001; // 1817 : 129 - 0x81
      11'h71A: dout  = 8'b10000001; // 1818 : 129 - 0x81
      11'h71B: dout  = 8'b10000001; // 1819 : 129 - 0x81
      11'h71C: dout  = 8'b10000001; // 1820 : 129 - 0x81
      11'h71D: dout  = 8'b10000001; // 1821 : 129 - 0x81
      11'h71E: dout  = 8'b10000001; // 1822 : 129 - 0x81
      11'h71F: dout  = 8'b10000001; // 1823 : 129 - 0x81
      11'h720: dout  = 8'b10000000; // 1824 : 128 - 0x80 -- Background 0xe4
      11'h721: dout  = 8'b10000000; // 1825 : 128 - 0x80
      11'h722: dout  = 8'b11000000; // 1826 : 192 - 0xc0
      11'h723: dout  = 8'b11000000; // 1827 : 192 - 0xc0
      11'h724: dout  = 8'b11100000; // 1828 : 224 - 0xe0
      11'h725: dout  = 8'b11111000; // 1829 : 248 - 0xf8
      11'h726: dout  = 8'b11111110; // 1830 : 254 - 0xfe
      11'h727: dout  = 8'b11111111; // 1831 : 255 - 0xff
      11'h728: dout  = 8'b11111111; // 1832 : 255 - 0xff -- Background 0xe5
      11'h729: dout  = 8'b01111111; // 1833 : 127 - 0x7f
      11'h72A: dout  = 8'b00011111; // 1834 :  31 - 0x1f
      11'h72B: dout  = 8'b00000111; // 1835 :   7 - 0x7
      11'h72C: dout  = 8'b00000011; // 1836 :   3 - 0x3
      11'h72D: dout  = 8'b00000011; // 1837 :   3 - 0x3
      11'h72E: dout  = 8'b00000001; // 1838 :   1 - 0x1
      11'h72F: dout  = 8'b10000001; // 1839 : 129 - 0x81
      11'h730: dout  = 8'b10000001; // 1840 : 129 - 0x81 -- Background 0xe6
      11'h731: dout  = 8'b10000001; // 1841 : 129 - 0x81
      11'h732: dout  = 8'b10000001; // 1842 : 129 - 0x81
      11'h733: dout  = 8'b10000001; // 1843 : 129 - 0x81
      11'h734: dout  = 8'b10000001; // 1844 : 129 - 0x81
      11'h735: dout  = 8'b10000001; // 1845 : 129 - 0x81
      11'h736: dout  = 8'b10000001; // 1846 : 129 - 0x81
      11'h737: dout  = 8'b10000001; // 1847 : 129 - 0x81
      11'h738: dout  = 8'b10000001; // 1848 : 129 - 0x81 -- Background 0xe7
      11'h739: dout  = 8'b10000001; // 1849 : 129 - 0x81
      11'h73A: dout  = 8'b10000001; // 1850 : 129 - 0x81
      11'h73B: dout  = 8'b10000001; // 1851 : 129 - 0x81
      11'h73C: dout  = 8'b10000001; // 1852 : 129 - 0x81
      11'h73D: dout  = 8'b10000001; // 1853 : 129 - 0x81
      11'h73E: dout  = 8'b10000001; // 1854 : 129 - 0x81
      11'h73F: dout  = 8'b10000001; // 1855 : 129 - 0x81
      11'h740: dout  = 8'b01111110; // 1856 : 126 - 0x7e -- Background 0xe8
      11'h741: dout  = 8'b00111100; // 1857 :  60 - 0x3c
      11'h742: dout  = 8'b00111100; // 1858 :  60 - 0x3c
      11'h743: dout  = 8'b00011000; // 1859 :  24 - 0x18
      11'h744: dout  = 8'b00011000; // 1860 :  24 - 0x18
      11'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      11'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      11'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      11'h748: dout  = 8'b11110010; // 1864 : 242 - 0xf2 -- Background 0xe9
      11'h749: dout  = 8'b11111110; // 1865 : 254 - 0xfe
      11'h74A: dout  = 8'b11111110; // 1866 : 254 - 0xfe
      11'h74B: dout  = 8'b11111111; // 1867 : 255 - 0xff
      11'h74C: dout  = 8'b11111111; // 1868 : 255 - 0xff
      11'h74D: dout  = 8'b11101111; // 1869 : 239 - 0xef
      11'h74E: dout  = 8'b11110111; // 1870 : 247 - 0xf7
      11'h74F: dout  = 8'b11111000; // 1871 : 248 - 0xf8
      11'h750: dout  = 8'b10111111; // 1872 : 191 - 0xbf -- Background 0xea
      11'h751: dout  = 8'b10111110; // 1873 : 190 - 0xbe
      11'h752: dout  = 8'b10111101; // 1874 : 189 - 0xbd
      11'h753: dout  = 8'b01111011; // 1875 : 123 - 0x7b
      11'h754: dout  = 8'b01111011; // 1876 : 123 - 0x7b
      11'h755: dout  = 8'b00000111; // 1877 :   7 - 0x7
      11'h756: dout  = 8'b11110011; // 1878 : 243 - 0xf3
      11'h757: dout  = 8'b11111101; // 1879 : 253 - 0xfd
      11'h758: dout  = 8'b11111111; // 1880 : 255 - 0xff -- Background 0xeb
      11'h759: dout  = 8'b11111111; // 1881 : 255 - 0xff
      11'h75A: dout  = 8'b11111111; // 1882 : 255 - 0xff
      11'h75B: dout  = 8'b01100111; // 1883 : 103 - 0x67
      11'h75C: dout  = 8'b01011001; // 1884 :  89 - 0x59
      11'h75D: dout  = 8'b10011110; // 1885 : 158 - 0x9e
      11'h75E: dout  = 8'b10111111; // 1886 : 191 - 0xbf
      11'h75F: dout  = 8'b10111111; // 1887 : 191 - 0xbf
      11'h760: dout  = 8'b00100000; // 1888 :  32 - 0x20 -- Background 0xec
      11'h761: dout  = 8'b11100110; // 1889 : 230 - 0xe6
      11'h762: dout  = 8'b01010100; // 1890 :  84 - 0x54
      11'h763: dout  = 8'b00100110; // 1891 :  38 - 0x26
      11'h764: dout  = 8'b00100001; // 1892 :  33 - 0x21
      11'h765: dout  = 8'b00000110; // 1893 :   6 - 0x6
      11'h766: dout  = 8'b01010100; // 1894 :  84 - 0x54
      11'h767: dout  = 8'b00100110; // 1895 :  38 - 0x26
      11'h768: dout  = 8'b00100000; // 1896 :  32 - 0x20 -- Background 0xed
      11'h769: dout  = 8'b10011010; // 1897 : 154 - 0x9a
      11'h76A: dout  = 8'b00000001; // 1898 :   1 - 0x1
      11'h76B: dout  = 8'b01001001; // 1899 :  73 - 0x49
      11'h76C: dout  = 8'b00100000; // 1900 :  32 - 0x20
      11'h76D: dout  = 8'b10100101; // 1901 : 165 - 0xa5
      11'h76E: dout  = 8'b11001001; // 1902 : 201 - 0xc9
      11'h76F: dout  = 8'b01000110; // 1903 :  70 - 0x46
      11'h770: dout  = 8'b11010001; // 1904 : 209 - 0xd1 -- Background 0xee
      11'h771: dout  = 8'b11011000; // 1905 : 216 - 0xd8
      11'h772: dout  = 8'b11011000; // 1906 : 216 - 0xd8
      11'h773: dout  = 8'b11011110; // 1907 : 222 - 0xde
      11'h774: dout  = 8'b11010001; // 1908 : 209 - 0xd1
      11'h775: dout  = 8'b11010000; // 1909 : 208 - 0xd0
      11'h776: dout  = 8'b11011010; // 1910 : 218 - 0xda
      11'h777: dout  = 8'b11011110; // 1911 : 222 - 0xde
      11'h778: dout  = 8'b11011011; // 1912 : 219 - 0xdb -- Background 0xef
      11'h779: dout  = 8'b11011001; // 1913 : 217 - 0xd9
      11'h77A: dout  = 8'b11011011; // 1914 : 219 - 0xdb
      11'h77B: dout  = 8'b11011100; // 1915 : 220 - 0xdc
      11'h77C: dout  = 8'b11011011; // 1916 : 219 - 0xdb
      11'h77D: dout  = 8'b11011111; // 1917 : 223 - 0xdf
      11'h77E: dout  = 8'b00100000; // 1918 :  32 - 0x20
      11'h77F: dout  = 8'b11100110; // 1919 : 230 - 0xe6
      11'h780: dout  = 8'b11011010; // 1920 : 218 - 0xda -- Background 0xf0
      11'h781: dout  = 8'b11011011; // 1921 : 219 - 0xdb
      11'h782: dout  = 8'b11100000; // 1922 : 224 - 0xe0
      11'h783: dout  = 8'b00100001; // 1923 :  33 - 0x21
      11'h784: dout  = 8'b00000110; // 1924 :   6 - 0x6
      11'h785: dout  = 8'b00001010; // 1925 :  10 - 0xa
      11'h786: dout  = 8'b11010110; // 1926 : 214 - 0xd6
      11'h787: dout  = 8'b11010111; // 1927 : 215 - 0xd7
      11'h788: dout  = 8'b00100001; // 1928 :  33 - 0x21 -- Background 0xf1
      11'h789: dout  = 8'b00100110; // 1929 :  38 - 0x26
      11'h78A: dout  = 8'b00010100; // 1930 :  20 - 0x14
      11'h78B: dout  = 8'b11010000; // 1931 : 208 - 0xd0
      11'h78C: dout  = 8'b11101000; // 1932 : 232 - 0xe8
      11'h78D: dout  = 8'b11010001; // 1933 : 209 - 0xd1
      11'h78E: dout  = 8'b11010000; // 1934 : 208 - 0xd0
      11'h78F: dout  = 8'b11010001; // 1935 : 209 - 0xd1
      11'h790: dout  = 8'b11011110; // 1936 : 222 - 0xde -- Background 0xf2
      11'h791: dout  = 8'b11010001; // 1937 : 209 - 0xd1
      11'h792: dout  = 8'b11010000; // 1938 : 208 - 0xd0
      11'h793: dout  = 8'b11010001; // 1939 : 209 - 0xd1
      11'h794: dout  = 8'b11010000; // 1940 : 208 - 0xd0
      11'h795: dout  = 8'b11010001; // 1941 : 209 - 0xd1
      11'h796: dout  = 8'b00100110; // 1942 :  38 - 0x26
      11'h797: dout  = 8'b00100001; // 1943 :  33 - 0x21
      11'h798: dout  = 8'b01000010; // 1944 :  66 - 0x42 -- Background 0xf3
      11'h799: dout  = 8'b11011011; // 1945 : 219 - 0xdb
      11'h79A: dout  = 8'b11011011; // 1946 : 219 - 0xdb
      11'h79B: dout  = 8'b01000010; // 1947 :  66 - 0x42
      11'h79C: dout  = 8'b00100110; // 1948 :  38 - 0x26
      11'h79D: dout  = 8'b11011011; // 1949 : 219 - 0xdb
      11'h79E: dout  = 8'b01000010; // 1950 :  66 - 0x42
      11'h79F: dout  = 8'b11011011; // 1951 : 219 - 0xdb
      11'h7A0: dout  = 8'b01000110; // 1952 :  70 - 0x46 -- Background 0xf4
      11'h7A1: dout  = 8'b11011011; // 1953 : 219 - 0xdb
      11'h7A2: dout  = 8'b00100001; // 1954 :  33 - 0x21
      11'h7A3: dout  = 8'b01101100; // 1955 : 108 - 0x6c
      11'h7A4: dout  = 8'b00001110; // 1956 :  14 - 0xe
      11'h7A5: dout  = 8'b11011111; // 1957 : 223 - 0xdf
      11'h7A6: dout  = 8'b11011011; // 1958 : 219 - 0xdb
      11'h7A7: dout  = 8'b11011011; // 1959 : 219 - 0xdb
      11'h7A8: dout  = 8'b11100100; // 1960 : 228 - 0xe4 -- Background 0xf5
      11'h7A9: dout  = 8'b11100101; // 1961 : 229 - 0xe5
      11'h7AA: dout  = 8'b00100110; // 1962 :  38 - 0x26
      11'h7AB: dout  = 8'b00100001; // 1963 :  33 - 0x21
      11'h7AC: dout  = 8'b10000110; // 1964 : 134 - 0x86
      11'h7AD: dout  = 8'b00010100; // 1965 :  20 - 0x14
      11'h7AE: dout  = 8'b11011011; // 1966 : 219 - 0xdb
      11'h7AF: dout  = 8'b11011011; // 1967 : 219 - 0xdb
      11'h7B0: dout  = 8'b00100110; // 1968 :  38 - 0x26 -- Background 0xf6
      11'h7B1: dout  = 8'b11011011; // 1969 : 219 - 0xdb
      11'h7B2: dout  = 8'b11100011; // 1970 : 227 - 0xe3
      11'h7B3: dout  = 8'b11011011; // 1971 : 219 - 0xdb
      11'h7B4: dout  = 8'b11100000; // 1972 : 224 - 0xe0
      11'h7B5: dout  = 8'b11011011; // 1973 : 219 - 0xdb
      11'h7B6: dout  = 8'b11011011; // 1974 : 219 - 0xdb
      11'h7B7: dout  = 8'b11100110; // 1975 : 230 - 0xe6
      11'h7B8: dout  = 8'b11011011; // 1976 : 219 - 0xdb -- Background 0xf7
      11'h7B9: dout  = 8'b01000010; // 1977 :  66 - 0x42
      11'h7BA: dout  = 8'b11011011; // 1978 : 219 - 0xdb
      11'h7BB: dout  = 8'b11011011; // 1979 : 219 - 0xdb
      11'h7BC: dout  = 8'b11011011; // 1980 : 219 - 0xdb
      11'h7BD: dout  = 8'b11010100; // 1981 : 212 - 0xd4
      11'h7BE: dout  = 8'b11011001; // 1982 : 217 - 0xd9
      11'h7BF: dout  = 8'b00100110; // 1983 :  38 - 0x26
      11'h7C0: dout  = 8'b11100111; // 1984 : 231 - 0xe7 -- Background 0xf8
      11'h7C1: dout  = 8'b00100001; // 1985 :  33 - 0x21
      11'h7C2: dout  = 8'b11000101; // 1986 : 197 - 0xc5
      11'h7C3: dout  = 8'b00010110; // 1987 :  22 - 0x16
      11'h7C4: dout  = 8'b01011111; // 1988 :  95 - 0x5f
      11'h7C5: dout  = 8'b10010101; // 1989 : 149 - 0x95
      11'h7C6: dout  = 8'b10010101; // 1990 : 149 - 0x95
      11'h7C7: dout  = 8'b10010101; // 1991 : 149 - 0x95
      11'h7C8: dout  = 8'b10010101; // 1992 : 149 - 0x95 -- Background 0xf9
      11'h7C9: dout  = 8'b10010110; // 1993 : 150 - 0x96
      11'h7CA: dout  = 8'b10010101; // 1994 : 149 - 0x95
      11'h7CB: dout  = 8'b10010101; // 1995 : 149 - 0x95
      11'h7CC: dout  = 8'b10010111; // 1996 : 151 - 0x97
      11'h7CD: dout  = 8'b10011000; // 1997 : 152 - 0x98
      11'h7CE: dout  = 8'b10010111; // 1998 : 151 - 0x97
      11'h7CF: dout  = 8'b10011000; // 1999 : 152 - 0x98
      11'h7D0: dout  = 8'b00001000; // 2000 :   8 - 0x8 -- Background 0xfa
      11'h7D1: dout  = 8'b00000101; // 2001 :   5 - 0x5
      11'h7D2: dout  = 8'b00100100; // 2002 :  36 - 0x24
      11'h7D3: dout  = 8'b00010111; // 2003 :  23 - 0x17
      11'h7D4: dout  = 8'b00010010; // 2004 :  18 - 0x12
      11'h7D5: dout  = 8'b00010111; // 2005 :  23 - 0x17
      11'h7D6: dout  = 8'b00011101; // 2006 :  29 - 0x1d
      11'h7D7: dout  = 8'b00001110; // 2007 :  14 - 0xe
      11'h7D8: dout  = 8'b00011001; // 2008 :  25 - 0x19 -- Background 0xfb
      11'h7D9: dout  = 8'b00010101; // 2009 :  21 - 0x15
      11'h7DA: dout  = 8'b00001010; // 2010 :  10 - 0xa
      11'h7DB: dout  = 8'b00100010; // 2011 :  34 - 0x22
      11'h7DC: dout  = 8'b00001110; // 2012 :  14 - 0xe
      11'h7DD: dout  = 8'b00011011; // 2013 :  27 - 0x1b
      11'h7DE: dout  = 8'b00100100; // 2014 :  36 - 0x24
      11'h7DF: dout  = 8'b00010000; // 2015 :  16 - 0x10
      11'h7E0: dout  = 8'b00011001; // 2016 :  25 - 0x19 -- Background 0xfc
      11'h7E1: dout  = 8'b00010101; // 2017 :  21 - 0x15
      11'h7E2: dout  = 8'b00001010; // 2018 :  10 - 0xa
      11'h7E3: dout  = 8'b00100010; // 2019 :  34 - 0x22
      11'h7E4: dout  = 8'b00001110; // 2020 :  14 - 0xe
      11'h7E5: dout  = 8'b00011011; // 2021 :  27 - 0x1b
      11'h7E6: dout  = 8'b00100100; // 2022 :  36 - 0x24
      11'h7E7: dout  = 8'b00010000; // 2023 :  16 - 0x10
      11'h7E8: dout  = 8'b00011001; // 2024 :  25 - 0x19 -- Background 0xfd
      11'h7E9: dout  = 8'b00101000; // 2025 :  40 - 0x28
      11'h7EA: dout  = 8'b00100010; // 2026 :  34 - 0x22
      11'h7EB: dout  = 8'b11110110; // 2027 : 246 - 0xf6
      11'h7EC: dout  = 8'b00000001; // 2028 :   1 - 0x1
      11'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      11'h7EE: dout  = 8'b00100011; // 2030 :  35 - 0x23
      11'h7EF: dout  = 8'b11001001; // 2031 : 201 - 0xc9
      11'h7F0: dout  = 8'b10101010; // 2032 : 170 - 0xaa -- Background 0xfe
      11'h7F1: dout  = 8'b00100011; // 2033 :  35 - 0x23
      11'h7F2: dout  = 8'b11101010; // 2034 : 234 - 0xea
      11'h7F3: dout  = 8'b00000100; // 2035 :   4 - 0x4
      11'h7F4: dout  = 8'b10011001; // 2036 : 153 - 0x99
      11'h7F5: dout  = 8'b10101010; // 2037 : 170 - 0xaa
      11'h7F6: dout  = 8'b10101010; // 2038 : 170 - 0xaa
      11'h7F7: dout  = 8'b10101010; // 2039 : 170 - 0xaa
      11'h7F8: dout  = 8'b11111111; // 2040 : 255 - 0xff -- Background 0xff
      11'h7F9: dout  = 8'b11111111; // 2041 : 255 - 0xff
      11'h7FA: dout  = 8'b11111111; // 2042 : 255 - 0xff
      11'h7FB: dout  = 8'b11111111; // 2043 : 255 - 0xff
      11'h7FC: dout  = 8'b11111111; // 2044 : 255 - 0xff
      11'h7FD: dout  = 8'b11111111; // 2045 : 255 - 0xff
      11'h7FE: dout  = 8'b11111111; // 2046 : 255 - 0xff
      11'h7FF: dout  = 8'b11111111; // 2047 : 255 - 0xff
    endcase
  end

endmodule
