--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: sprilo_endscr.bin --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_SPRILO_ENDSCREEN is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_SPRILO_ENDSCREEN;

architecture BEHAVIORAL of ROM_NTABLE_SPRILO_ENDSCREEN is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "11111010", --    0 -  0x0  :  250 - 0xfa -- line 0x0
    "11111010", --    1 -  0x1  :  250 - 0xfa
    "11111010", --    2 -  0x2  :  250 - 0xfa
    "11101010", --    3 -  0x3  :  234 - 0xea
    "11111010", --    4 -  0x4  :  250 - 0xfa
    "11111010", --    5 -  0x5  :  250 - 0xfa
    "11111010", --    6 -  0x6  :  250 - 0xfa
    "11111010", --    7 -  0x7  :  250 - 0xfa
    "11111010", --    8 -  0x8  :  250 - 0xfa
    "11111010", --    9 -  0x9  :  250 - 0xfa
    "11111010", --   10 -  0xa  :  250 - 0xfa
    "11111010", --   11 -  0xb  :  250 - 0xfa
    "11111010", --   12 -  0xc  :  250 - 0xfa
    "11111010", --   13 -  0xd  :  250 - 0xfa
    "11101010", --   14 -  0xe  :  234 - 0xea
    "11111010", --   15 -  0xf  :  250 - 0xfa
    "11111010", --   16 - 0x10  :  250 - 0xfa
    "11111010", --   17 - 0x11  :  250 - 0xfa
    "11111010", --   18 - 0x12  :  250 - 0xfa
    "11111010", --   19 - 0x13  :  250 - 0xfa
    "11111010", --   20 - 0x14  :  250 - 0xfa
    "11111010", --   21 - 0x15  :  250 - 0xfa
    "11111010", --   22 - 0x16  :  250 - 0xfa
    "11111010", --   23 - 0x17  :  250 - 0xfa
    "11111010", --   24 - 0x18  :  250 - 0xfa
    "11111010", --   25 - 0x19  :  250 - 0xfa
    "11111010", --   26 - 0x1a  :  250 - 0xfa
    "11111010", --   27 - 0x1b  :  250 - 0xfa
    "11111010", --   28 - 0x1c  :  250 - 0xfa
    "11111010", --   29 - 0x1d  :  250 - 0xfa
    "11111010", --   30 - 0x1e  :  250 - 0xfa
    "11111010", --   31 - 0x1f  :  250 - 0xfa
    "11111010", --   32 - 0x20  :  250 - 0xfa -- line 0x1
    "11111010", --   33 - 0x21  :  250 - 0xfa
    "11111010", --   34 - 0x22  :  250 - 0xfa
    "11111010", --   35 - 0x23  :  250 - 0xfa
    "11111010", --   36 - 0x24  :  250 - 0xfa
    "11111010", --   37 - 0x25  :  250 - 0xfa
    "11111010", --   38 - 0x26  :  250 - 0xfa
    "11111001", --   39 - 0x27  :  249 - 0xf9
    "11111001", --   40 - 0x28  :  249 - 0xf9
    "11111010", --   41 - 0x29  :  250 - 0xfa
    "11111010", --   42 - 0x2a  :  250 - 0xfa
    "11111010", --   43 - 0x2b  :  250 - 0xfa
    "11111010", --   44 - 0x2c  :  250 - 0xfa
    "11111010", --   45 - 0x2d  :  250 - 0xfa
    "11111010", --   46 - 0x2e  :  250 - 0xfa
    "11111010", --   47 - 0x2f  :  250 - 0xfa
    "11111010", --   48 - 0x30  :  250 - 0xfa
    "11111010", --   49 - 0x31  :  250 - 0xfa
    "11101001", --   50 - 0x32  :  233 - 0xe9
    "11111010", --   51 - 0x33  :  250 - 0xfa
    "11111010", --   52 - 0x34  :  250 - 0xfa
    "11111010", --   53 - 0x35  :  250 - 0xfa
    "11111010", --   54 - 0x36  :  250 - 0xfa
    "11111010", --   55 - 0x37  :  250 - 0xfa
    "11111010", --   56 - 0x38  :  250 - 0xfa
    "11111010", --   57 - 0x39  :  250 - 0xfa
    "11111001", --   58 - 0x3a  :  249 - 0xf9
    "11111010", --   59 - 0x3b  :  250 - 0xfa
    "11111010", --   60 - 0x3c  :  250 - 0xfa
    "11111010", --   61 - 0x3d  :  250 - 0xfa
    "11111010", --   62 - 0x3e  :  250 - 0xfa
    "11111010", --   63 - 0x3f  :  250 - 0xfa
    "11111010", --   64 - 0x40  :  250 - 0xfa -- line 0x2
    "11111001", --   65 - 0x41  :  249 - 0xf9
    "11111010", --   66 - 0x42  :  250 - 0xfa
    "11111010", --   67 - 0x43  :  250 - 0xfa
    "11111010", --   68 - 0x44  :  250 - 0xfa
    "11111010", --   69 - 0x45  :  250 - 0xfa
    "11111010", --   70 - 0x46  :  250 - 0xfa
    "11111010", --   71 - 0x47  :  250 - 0xfa
    "11111010", --   72 - 0x48  :  250 - 0xfa
    "11111010", --   73 - 0x49  :  250 - 0xfa
    "11111010", --   74 - 0x4a  :  250 - 0xfa
    "11111010", --   75 - 0x4b  :  250 - 0xfa
    "11111010", --   76 - 0x4c  :  250 - 0xfa
    "11111010", --   77 - 0x4d  :  250 - 0xfa
    "11111010", --   78 - 0x4e  :  250 - 0xfa
    "11101001", --   79 - 0x4f  :  233 - 0xe9
    "11111010", --   80 - 0x50  :  250 - 0xfa
    "11111010", --   81 - 0x51  :  250 - 0xfa
    "11111010", --   82 - 0x52  :  250 - 0xfa
    "11111010", --   83 - 0x53  :  250 - 0xfa
    "11111010", --   84 - 0x54  :  250 - 0xfa
    "11111010", --   85 - 0x55  :  250 - 0xfa
    "11111010", --   86 - 0x56  :  250 - 0xfa
    "11111010", --   87 - 0x57  :  250 - 0xfa
    "11111010", --   88 - 0x58  :  250 - 0xfa
    "11111010", --   89 - 0x59  :  250 - 0xfa
    "11111010", --   90 - 0x5a  :  250 - 0xfa
    "11111010", --   91 - 0x5b  :  250 - 0xfa
    "11111010", --   92 - 0x5c  :  250 - 0xfa
    "11111010", --   93 - 0x5d  :  250 - 0xfa
    "11111010", --   94 - 0x5e  :  250 - 0xfa
    "11111010", --   95 - 0x5f  :  250 - 0xfa
    "11111010", --   96 - 0x60  :  250 - 0xfa -- line 0x3
    "11111010", --   97 - 0x61  :  250 - 0xfa
    "11111010", --   98 - 0x62  :  250 - 0xfa
    "11111010", --   99 - 0x63  :  250 - 0xfa
    "11111010", --  100 - 0x64  :  250 - 0xfa
    "11111010", --  101 - 0x65  :  250 - 0xfa
    "11111010", --  102 - 0x66  :  250 - 0xfa
    "11101001", --  103 - 0x67  :  233 - 0xe9
    "11111010", --  104 - 0x68  :  250 - 0xfa
    "11111010", --  105 - 0x69  :  250 - 0xfa
    "11111010", --  106 - 0x6a  :  250 - 0xfa
    "11111010", --  107 - 0x6b  :  250 - 0xfa
    "11111010", --  108 - 0x6c  :  250 - 0xfa
    "11111010", --  109 - 0x6d  :  250 - 0xfa
    "11111010", --  110 - 0x6e  :  250 - 0xfa
    "11111010", --  111 - 0x6f  :  250 - 0xfa
    "11111010", --  112 - 0x70  :  250 - 0xfa
    "11111010", --  113 - 0x71  :  250 - 0xfa
    "11111010", --  114 - 0x72  :  250 - 0xfa
    "11111010", --  115 - 0x73  :  250 - 0xfa
    "11111010", --  116 - 0x74  :  250 - 0xfa
    "11111010", --  117 - 0x75  :  250 - 0xfa
    "11101010", --  118 - 0x76  :  234 - 0xea
    "11111010", --  119 - 0x77  :  250 - 0xfa
    "11111010", --  120 - 0x78  :  250 - 0xfa
    "11111010", --  121 - 0x79  :  250 - 0xfa
    "11111010", --  122 - 0x7a  :  250 - 0xfa
    "11111010", --  123 - 0x7b  :  250 - 0xfa
    "11111010", --  124 - 0x7c  :  250 - 0xfa
    "11111010", --  125 - 0x7d  :  250 - 0xfa
    "11111010", --  126 - 0x7e  :  250 - 0xfa
    "11111010", --  127 - 0x7f  :  250 - 0xfa
    "11111010", --  128 - 0x80  :  250 - 0xfa -- line 0x4
    "11111010", --  129 - 0x81  :  250 - 0xfa
    "11111010", --  130 - 0x82  :  250 - 0xfa
    "11111010", --  131 - 0x83  :  250 - 0xfa
    "11111010", --  132 - 0x84  :  250 - 0xfa
    "11111010", --  133 - 0x85  :  250 - 0xfa
    "11111010", --  134 - 0x86  :  250 - 0xfa
    "11111010", --  135 - 0x87  :  250 - 0xfa
    "11111010", --  136 - 0x88  :  250 - 0xfa
    "11111010", --  137 - 0x89  :  250 - 0xfa
    "11111010", --  138 - 0x8a  :  250 - 0xfa
    "11111010", --  139 - 0x8b  :  250 - 0xfa
    "11111010", --  140 - 0x8c  :  250 - 0xfa
    "11111010", --  141 - 0x8d  :  250 - 0xfa
    "11111010", --  142 - 0x8e  :  250 - 0xfa
    "11111010", --  143 - 0x8f  :  250 - 0xfa
    "11111010", --  144 - 0x90  :  250 - 0xfa
    "11111010", --  145 - 0x91  :  250 - 0xfa
    "11111010", --  146 - 0x92  :  250 - 0xfa
    "11111010", --  147 - 0x93  :  250 - 0xfa
    "11111010", --  148 - 0x94  :  250 - 0xfa
    "11111010", --  149 - 0x95  :  250 - 0xfa
    "11111010", --  150 - 0x96  :  250 - 0xfa
    "11111010", --  151 - 0x97  :  250 - 0xfa
    "11111010", --  152 - 0x98  :  250 - 0xfa
    "11111010", --  153 - 0x99  :  250 - 0xfa
    "11111010", --  154 - 0x9a  :  250 - 0xfa
    "11111010", --  155 - 0x9b  :  250 - 0xfa
    "11111001", --  156 - 0x9c  :  249 - 0xf9
    "11111010", --  157 - 0x9d  :  250 - 0xfa
    "11111010", --  158 - 0x9e  :  250 - 0xfa
    "11111010", --  159 - 0x9f  :  250 - 0xfa
    "11111010", --  160 - 0xa0  :  250 - 0xfa -- line 0x5
    "11111010", --  161 - 0xa1  :  250 - 0xfa
    "11111010", --  162 - 0xa2  :  250 - 0xfa
    "11111010", --  163 - 0xa3  :  250 - 0xfa
    "11111010", --  164 - 0xa4  :  250 - 0xfa
    "11111010", --  165 - 0xa5  :  250 - 0xfa
    "11111010", --  166 - 0xa6  :  250 - 0xfa
    "11111010", --  167 - 0xa7  :  250 - 0xfa
    "11111010", --  168 - 0xa8  :  250 - 0xfa
    "11111010", --  169 - 0xa9  :  250 - 0xfa
    "11111010", --  170 - 0xaa  :  250 - 0xfa
    "11101010", --  171 - 0xab  :  234 - 0xea
    "11111010", --  172 - 0xac  :  250 - 0xfa
    "11111010", --  173 - 0xad  :  250 - 0xfa
    "11111010", --  174 - 0xae  :  250 - 0xfa
    "11111010", --  175 - 0xaf  :  250 - 0xfa
    "11111010", --  176 - 0xb0  :  250 - 0xfa
    "11111010", --  177 - 0xb1  :  250 - 0xfa
    "11111010", --  178 - 0xb2  :  250 - 0xfa
    "11111001", --  179 - 0xb3  :  249 - 0xf9
    "11111010", --  180 - 0xb4  :  250 - 0xfa
    "11111010", --  181 - 0xb5  :  250 - 0xfa
    "11111010", --  182 - 0xb6  :  250 - 0xfa
    "11111010", --  183 - 0xb7  :  250 - 0xfa
    "11111010", --  184 - 0xb8  :  250 - 0xfa
    "11111010", --  185 - 0xb9  :  250 - 0xfa
    "11111010", --  186 - 0xba  :  250 - 0xfa
    "11111010", --  187 - 0xbb  :  250 - 0xfa
    "11111010", --  188 - 0xbc  :  250 - 0xfa
    "11111010", --  189 - 0xbd  :  250 - 0xfa
    "11111010", --  190 - 0xbe  :  250 - 0xfa
    "11111010", --  191 - 0xbf  :  250 - 0xfa
    "11111010", --  192 - 0xc0  :  250 - 0xfa -- line 0x6
    "11111010", --  193 - 0xc1  :  250 - 0xfa
    "11111010", --  194 - 0xc2  :  250 - 0xfa
    "11111010", --  195 - 0xc3  :  250 - 0xfa
    "11101010", --  196 - 0xc4  :  234 - 0xea
    "11111010", --  197 - 0xc5  :  250 - 0xfa
    "11111010", --  198 - 0xc6  :  250 - 0xfa
    "11111010", --  199 - 0xc7  :  250 - 0xfa
    "11111010", --  200 - 0xc8  :  250 - 0xfa
    "11111010", --  201 - 0xc9  :  250 - 0xfa
    "11111010", --  202 - 0xca  :  250 - 0xfa
    "11111010", --  203 - 0xcb  :  250 - 0xfa
    "11111010", --  204 - 0xcc  :  250 - 0xfa
    "11111010", --  205 - 0xcd  :  250 - 0xfa
    "11111010", --  206 - 0xce  :  250 - 0xfa
    "11111010", --  207 - 0xcf  :  250 - 0xfa
    "11111010", --  208 - 0xd0  :  250 - 0xfa
    "11111010", --  209 - 0xd1  :  250 - 0xfa
    "11111010", --  210 - 0xd2  :  250 - 0xfa
    "11111010", --  211 - 0xd3  :  250 - 0xfa
    "11111010", --  212 - 0xd4  :  250 - 0xfa
    "11101010", --  213 - 0xd5  :  234 - 0xea
    "11111010", --  214 - 0xd6  :  250 - 0xfa
    "11111010", --  215 - 0xd7  :  250 - 0xfa
    "11111010", --  216 - 0xd8  :  250 - 0xfa
    "11111010", --  217 - 0xd9  :  250 - 0xfa
    "11111010", --  218 - 0xda  :  250 - 0xfa
    "11111010", --  219 - 0xdb  :  250 - 0xfa
    "11111010", --  220 - 0xdc  :  250 - 0xfa
    "11111010", --  221 - 0xdd  :  250 - 0xfa
    "11111010", --  222 - 0xde  :  250 - 0xfa
    "11111010", --  223 - 0xdf  :  250 - 0xfa
    "11111010", --  224 - 0xe0  :  250 - 0xfa -- line 0x7
    "11111010", --  225 - 0xe1  :  250 - 0xfa
    "11111010", --  226 - 0xe2  :  250 - 0xfa
    "11111010", --  227 - 0xe3  :  250 - 0xfa
    "11111010", --  228 - 0xe4  :  250 - 0xfa
    "11111010", --  229 - 0xe5  :  250 - 0xfa
    "11111010", --  230 - 0xe6  :  250 - 0xfa
    "11111010", --  231 - 0xe7  :  250 - 0xfa
    "11111010", --  232 - 0xe8  :  250 - 0xfa
    "11111001", --  233 - 0xe9  :  249 - 0xf9
    "11111010", --  234 - 0xea  :  250 - 0xfa
    "11111010", --  235 - 0xeb  :  250 - 0xfa
    "11111010", --  236 - 0xec  :  250 - 0xfa
    "11111010", --  237 - 0xed  :  250 - 0xfa
    "11111010", --  238 - 0xee  :  250 - 0xfa
    "11111010", --  239 - 0xef  :  250 - 0xfa
    "11111010", --  240 - 0xf0  :  250 - 0xfa
    "11111001", --  241 - 0xf1  :  249 - 0xf9
    "11111010", --  242 - 0xf2  :  250 - 0xfa
    "11111010", --  243 - 0xf3  :  250 - 0xfa
    "11111010", --  244 - 0xf4  :  250 - 0xfa
    "11111010", --  245 - 0xf5  :  250 - 0xfa
    "11101001", --  246 - 0xf6  :  233 - 0xe9
    "11111010", --  247 - 0xf7  :  250 - 0xfa
    "11111010", --  248 - 0xf8  :  250 - 0xfa
    "11111010", --  249 - 0xf9  :  250 - 0xfa
    "11111010", --  250 - 0xfa  :  250 - 0xfa
    "11111010", --  251 - 0xfb  :  250 - 0xfa
    "11111010", --  252 - 0xfc  :  250 - 0xfa
    "11111010", --  253 - 0xfd  :  250 - 0xfa
    "11111010", --  254 - 0xfe  :  250 - 0xfa
    "11101010", --  255 - 0xff  :  234 - 0xea
    "11111010", --  256 - 0x100  :  250 - 0xfa -- line 0x8
    "11111010", --  257 - 0x101  :  250 - 0xfa
    "11111010", --  258 - 0x102  :  250 - 0xfa
    "11111010", --  259 - 0x103  :  250 - 0xfa
    "11111010", --  260 - 0x104  :  250 - 0xfa
    "11111001", --  261 - 0x105  :  249 - 0xf9
    "11111010", --  262 - 0x106  :  250 - 0xfa
    "11111010", --  263 - 0x107  :  250 - 0xfa
    "11111001", --  264 - 0x108  :  249 - 0xf9
    "11111001", --  265 - 0x109  :  249 - 0xf9
    "00101001", --  266 - 0x10a  :   41 - 0x29
    "00011111", --  267 - 0x10b  :   31 - 0x1f
    "00100101", --  268 - 0x10c  :   37 - 0x25
    "11111010", --  269 - 0x10d  :  250 - 0xfa
    "00010011", --  270 - 0x10e  :   19 - 0x13
    "00011111", --  271 - 0x10f  :   31 - 0x1f
    "00011101", --  272 - 0x110  :   29 - 0x1d
    "00100000", --  273 - 0x111  :   32 - 0x20
    "00011100", --  274 - 0x112  :   28 - 0x1c
    "00010101", --  275 - 0x113  :   21 - 0x15
    "00100100", --  276 - 0x114  :   36 - 0x24
    "00010101", --  277 - 0x115  :   21 - 0x15
    "00010100", --  278 - 0x116  :   20 - 0x14
    "11111010", --  279 - 0x117  :  250 - 0xfa
    "11111010", --  280 - 0x118  :  250 - 0xfa
    "11111010", --  281 - 0x119  :  250 - 0xfa
    "11111010", --  282 - 0x11a  :  250 - 0xfa
    "11111010", --  283 - 0x11b  :  250 - 0xfa
    "11111010", --  284 - 0x11c  :  250 - 0xfa
    "11111010", --  285 - 0x11d  :  250 - 0xfa
    "11111010", --  286 - 0x11e  :  250 - 0xfa
    "11111010", --  287 - 0x11f  :  250 - 0xfa
    "11111010", --  288 - 0x120  :  250 - 0xfa -- line 0x9
    "11111010", --  289 - 0x121  :  250 - 0xfa
    "11101001", --  290 - 0x122  :  233 - 0xe9
    "11111010", --  291 - 0x123  :  250 - 0xfa
    "11111010", --  292 - 0x124  :  250 - 0xfa
    "11111010", --  293 - 0x125  :  250 - 0xfa
    "11111010", --  294 - 0x126  :  250 - 0xfa
    "11111010", --  295 - 0x127  :  250 - 0xfa
    "11111010", --  296 - 0x128  :  250 - 0xfa
    "11111010", --  297 - 0x129  :  250 - 0xfa
    "11111010", --  298 - 0x12a  :  250 - 0xfa
    "11111010", --  299 - 0x12b  :  250 - 0xfa
    "11111010", --  300 - 0x12c  :  250 - 0xfa
    "11111010", --  301 - 0x12d  :  250 - 0xfa
    "11111010", --  302 - 0x12e  :  250 - 0xfa
    "11101001", --  303 - 0x12f  :  233 - 0xe9
    "11111010", --  304 - 0x130  :  250 - 0xfa
    "11111010", --  305 - 0x131  :  250 - 0xfa
    "11111010", --  306 - 0x132  :  250 - 0xfa
    "11111010", --  307 - 0x133  :  250 - 0xfa
    "11111010", --  308 - 0x134  :  250 - 0xfa
    "11111010", --  309 - 0x135  :  250 - 0xfa
    "11111010", --  310 - 0x136  :  250 - 0xfa
    "11101010", --  311 - 0x137  :  234 - 0xea
    "11111010", --  312 - 0x138  :  250 - 0xfa
    "11111010", --  313 - 0x139  :  250 - 0xfa
    "11111010", --  314 - 0x13a  :  250 - 0xfa
    "11111010", --  315 - 0x13b  :  250 - 0xfa
    "11111010", --  316 - 0x13c  :  250 - 0xfa
    "11111010", --  317 - 0x13d  :  250 - 0xfa
    "11111010", --  318 - 0x13e  :  250 - 0xfa
    "11111010", --  319 - 0x13f  :  250 - 0xfa
    "11111010", --  320 - 0x140  :  250 - 0xfa -- line 0xa
    "11111010", --  321 - 0x141  :  250 - 0xfa
    "11111010", --  322 - 0x142  :  250 - 0xfa
    "11111010", --  323 - 0x143  :  250 - 0xfa
    "11111010", --  324 - 0x144  :  250 - 0xfa
    "11111010", --  325 - 0x145  :  250 - 0xfa
    "11111010", --  326 - 0x146  :  250 - 0xfa
    "11111010", --  327 - 0x147  :  250 - 0xfa
    "11111010", --  328 - 0x148  :  250 - 0xfa
    "11111010", --  329 - 0x149  :  250 - 0xfa
    "00001111", --  330 - 0x14a  :   15 - 0xf
    "11111010", --  331 - 0x14b  :  250 - 0xfa
    "11111010", --  332 - 0x14c  :  250 - 0xfa
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00011000", --  334 - 0x14e  :   24 - 0x18
    "11111010", --  335 - 0x14f  :  250 - 0xfa
    "00011100", --  336 - 0x150  :   28 - 0x1c
    "00010001", --  337 - 0x151  :   17 - 0x11
    "00100000", --  338 - 0x152  :   32 - 0x20
    "00100011", --  339 - 0x153  :   35 - 0x23
    "11111010", --  340 - 0x154  :  250 - 0xfa
    "11101001", --  341 - 0x155  :  233 - 0xe9
    "00001111", --  342 - 0x156  :   15 - 0xf
    "11111010", --  343 - 0x157  :  250 - 0xfa
    "11111010", --  344 - 0x158  :  250 - 0xfa
    "11111010", --  345 - 0x159  :  250 - 0xfa
    "11111010", --  346 - 0x15a  :  250 - 0xfa
    "11111010", --  347 - 0x15b  :  250 - 0xfa
    "11111010", --  348 - 0x15c  :  250 - 0xfa
    "11101010", --  349 - 0x15d  :  234 - 0xea
    "11111010", --  350 - 0x15e  :  250 - 0xfa
    "11111010", --  351 - 0x15f  :  250 - 0xfa
    "11111010", --  352 - 0x160  :  250 - 0xfa -- line 0xb
    "11111010", --  353 - 0x161  :  250 - 0xfa
    "11111010", --  354 - 0x162  :  250 - 0xfa
    "11111010", --  355 - 0x163  :  250 - 0xfa
    "11111010", --  356 - 0x164  :  250 - 0xfa
    "11111010", --  357 - 0x165  :  250 - 0xfa
    "11111010", --  358 - 0x166  :  250 - 0xfa
    "11111010", --  359 - 0x167  :  250 - 0xfa
    "11111010", --  360 - 0x168  :  250 - 0xfa
    "11111010", --  361 - 0x169  :  250 - 0xfa
    "11111010", --  362 - 0x16a  :  250 - 0xfa
    "11111010", --  363 - 0x16b  :  250 - 0xfa
    "11101010", --  364 - 0x16c  :  234 - 0xea
    "11111010", --  365 - 0x16d  :  250 - 0xfa
    "11111010", --  366 - 0x16e  :  250 - 0xfa
    "11111010", --  367 - 0x16f  :  250 - 0xfa
    "11111010", --  368 - 0x170  :  250 - 0xfa
    "11111010", --  369 - 0x171  :  250 - 0xfa
    "11111010", --  370 - 0x172  :  250 - 0xfa
    "11111010", --  371 - 0x173  :  250 - 0xfa
    "11111010", --  372 - 0x174  :  250 - 0xfa
    "11111010", --  373 - 0x175  :  250 - 0xfa
    "11111010", --  374 - 0x176  :  250 - 0xfa
    "11101010", --  375 - 0x177  :  234 - 0xea
    "11111010", --  376 - 0x178  :  250 - 0xfa
    "11111010", --  377 - 0x179  :  250 - 0xfa
    "11111010", --  378 - 0x17a  :  250 - 0xfa
    "11111010", --  379 - 0x17b  :  250 - 0xfa
    "11111010", --  380 - 0x17c  :  250 - 0xfa
    "11111010", --  381 - 0x17d  :  250 - 0xfa
    "11111010", --  382 - 0x17e  :  250 - 0xfa
    "11111010", --  383 - 0x17f  :  250 - 0xfa
    "11111010", --  384 - 0x180  :  250 - 0xfa -- line 0xc
    "11111010", --  385 - 0x181  :  250 - 0xfa
    "11111010", --  386 - 0x182  :  250 - 0xfa
    "11111010", --  387 - 0x183  :  250 - 0xfa
    "11111010", --  388 - 0x184  :  250 - 0xfa
    "11111010", --  389 - 0x185  :  250 - 0xfa
    "11111010", --  390 - 0x186  :  250 - 0xfa
    "11111010", --  391 - 0x187  :  250 - 0xfa
    "11111010", --  392 - 0x188  :  250 - 0xfa
    "11111010", --  393 - 0x189  :  250 - 0xfa
    "11111010", --  394 - 0x18a  :  250 - 0xfa
    "11111010", --  395 - 0x18b  :  250 - 0xfa
    "11111010", --  396 - 0x18c  :  250 - 0xfa
    "11111010", --  397 - 0x18d  :  250 - 0xfa
    "11111010", --  398 - 0x18e  :  250 - 0xfa
    "00011001", --  399 - 0x18f  :   25 - 0x19
    "00011110", --  400 - 0x190  :   30 - 0x1e
    "11101001", --  401 - 0x191  :  233 - 0xe9
    "11111001", --  402 - 0x192  :  249 - 0xf9
    "11111010", --  403 - 0x193  :  250 - 0xfa
    "11111010", --  404 - 0x194  :  250 - 0xfa
    "11111010", --  405 - 0x195  :  250 - 0xfa
    "11111010", --  406 - 0x196  :  250 - 0xfa
    "11111010", --  407 - 0x197  :  250 - 0xfa
    "11111010", --  408 - 0x198  :  250 - 0xfa
    "11111010", --  409 - 0x199  :  250 - 0xfa
    "11111010", --  410 - 0x19a  :  250 - 0xfa
    "11111010", --  411 - 0x19b  :  250 - 0xfa
    "11111010", --  412 - 0x19c  :  250 - 0xfa
    "11111010", --  413 - 0x19d  :  250 - 0xfa
    "11111010", --  414 - 0x19e  :  250 - 0xfa
    "11111010", --  415 - 0x19f  :  250 - 0xfa
    "11111010", --  416 - 0x1a0  :  250 - 0xfa -- line 0xd
    "11111010", --  417 - 0x1a1  :  250 - 0xfa
    "11111010", --  418 - 0x1a2  :  250 - 0xfa
    "11111010", --  419 - 0x1a3  :  250 - 0xfa
    "11101010", --  420 - 0x1a4  :  234 - 0xea
    "11111010", --  421 - 0x1a5  :  250 - 0xfa
    "11111010", --  422 - 0x1a6  :  250 - 0xfa
    "11111010", --  423 - 0x1a7  :  250 - 0xfa
    "11111001", --  424 - 0x1a8  :  249 - 0xf9
    "11111010", --  425 - 0x1a9  :  250 - 0xfa
    "11111010", --  426 - 0x1aa  :  250 - 0xfa
    "11111010", --  427 - 0x1ab  :  250 - 0xfa
    "11111010", --  428 - 0x1ac  :  250 - 0xfa
    "11111010", --  429 - 0x1ad  :  250 - 0xfa
    "11111010", --  430 - 0x1ae  :  250 - 0xfa
    "11111010", --  431 - 0x1af  :  250 - 0xfa
    "11111010", --  432 - 0x1b0  :  250 - 0xfa
    "11111010", --  433 - 0x1b1  :  250 - 0xfa
    "11111010", --  434 - 0x1b2  :  250 - 0xfa
    "11111010", --  435 - 0x1b3  :  250 - 0xfa
    "11111010", --  436 - 0x1b4  :  250 - 0xfa
    "11111010", --  437 - 0x1b5  :  250 - 0xfa
    "11111010", --  438 - 0x1b6  :  250 - 0xfa
    "11111010", --  439 - 0x1b7  :  250 - 0xfa
    "11111010", --  440 - 0x1b8  :  250 - 0xfa
    "11111010", --  441 - 0x1b9  :  250 - 0xfa
    "11111010", --  442 - 0x1ba  :  250 - 0xfa
    "11111010", --  443 - 0x1bb  :  250 - 0xfa
    "11111010", --  444 - 0x1bc  :  250 - 0xfa
    "11111010", --  445 - 0x1bd  :  250 - 0xfa
    "11111010", --  446 - 0x1be  :  250 - 0xfa
    "11111010", --  447 - 0x1bf  :  250 - 0xfa
    "11111010", --  448 - 0x1c0  :  250 - 0xfa -- line 0xe
    "11111010", --  449 - 0x1c1  :  250 - 0xfa
    "11111010", --  450 - 0x1c2  :  250 - 0xfa
    "11111010", --  451 - 0x1c3  :  250 - 0xfa
    "11111010", --  452 - 0x1c4  :  250 - 0xfa
    "11111010", --  453 - 0x1c5  :  250 - 0xfa
    "11111010", --  454 - 0x1c6  :  250 - 0xfa
    "11111010", --  455 - 0x1c7  :  250 - 0xfa
    "11111010", --  456 - 0x1c8  :  250 - 0xfa
    "11111010", --  457 - 0x1c9  :  250 - 0xfa
    "00001101", --  458 - 0x1ca  :   13 - 0xd
    "11111010", --  459 - 0x1cb  :  250 - 0xfa
    "00010010", --  460 - 0x1cc  :   18 - 0x12
    "00010001", --  461 - 0x1cd  :   17 - 0x11
    "00010010", --  462 - 0x1ce  :   18 - 0x12
    "11111010", --  463 - 0x1cf  :  250 - 0xfa
    "00100011", --  464 - 0x1d0  :   35 - 0x23
    "00010101", --  465 - 0x1d1  :   21 - 0x15
    "00010011", --  466 - 0x1d2  :   19 - 0x13
    "00100011", --  467 - 0x1d3  :   35 - 0x23
    "00001011", --  468 - 0x1d4  :   11 - 0xb
    "11111010", --  469 - 0x1d5  :  250 - 0xfa
    "00001101", --  470 - 0x1d6  :   13 - 0xd
    "11111010", --  471 - 0x1d7  :  250 - 0xfa
    "11111010", --  472 - 0x1d8  :  250 - 0xfa
    "11111010", --  473 - 0x1d9  :  250 - 0xfa
    "11111010", --  474 - 0x1da  :  250 - 0xfa
    "11111010", --  475 - 0x1db  :  250 - 0xfa
    "11111010", --  476 - 0x1dc  :  250 - 0xfa
    "11111010", --  477 - 0x1dd  :  250 - 0xfa
    "11111010", --  478 - 0x1de  :  250 - 0xfa
    "11111010", --  479 - 0x1df  :  250 - 0xfa
    "11111010", --  480 - 0x1e0  :  250 - 0xfa -- line 0xf
    "11111001", --  481 - 0x1e1  :  249 - 0xf9
    "11111010", --  482 - 0x1e2  :  250 - 0xfa
    "11111010", --  483 - 0x1e3  :  250 - 0xfa
    "11111010", --  484 - 0x1e4  :  250 - 0xfa
    "11111010", --  485 - 0x1e5  :  250 - 0xfa
    "11111010", --  486 - 0x1e6  :  250 - 0xfa
    "11111010", --  487 - 0x1e7  :  250 - 0xfa
    "11111010", --  488 - 0x1e8  :  250 - 0xfa
    "11111010", --  489 - 0x1e9  :  250 - 0xfa
    "11111010", --  490 - 0x1ea  :  250 - 0xfa
    "11111010", --  491 - 0x1eb  :  250 - 0xfa
    "11111010", --  492 - 0x1ec  :  250 - 0xfa
    "11111010", --  493 - 0x1ed  :  250 - 0xfa
    "11111010", --  494 - 0x1ee  :  250 - 0xfa
    "11111010", --  495 - 0x1ef  :  250 - 0xfa
    "11111010", --  496 - 0x1f0  :  250 - 0xfa
    "11111010", --  497 - 0x1f1  :  250 - 0xfa
    "11111010", --  498 - 0x1f2  :  250 - 0xfa
    "11111010", --  499 - 0x1f3  :  250 - 0xfa
    "11111010", --  500 - 0x1f4  :  250 - 0xfa
    "11111010", --  501 - 0x1f5  :  250 - 0xfa
    "11111010", --  502 - 0x1f6  :  250 - 0xfa
    "11101001", --  503 - 0x1f7  :  233 - 0xe9
    "11111010", --  504 - 0x1f8  :  250 - 0xfa
    "11101001", --  505 - 0x1f9  :  233 - 0xe9
    "11111010", --  506 - 0x1fa  :  250 - 0xfa
    "11111010", --  507 - 0x1fb  :  250 - 0xfa
    "11111010", --  508 - 0x1fc  :  250 - 0xfa
    "11111010", --  509 - 0x1fd  :  250 - 0xfa
    "11111010", --  510 - 0x1fe  :  250 - 0xfa
    "11111010", --  511 - 0x1ff  :  250 - 0xfa
    "11111010", --  512 - 0x200  :  250 - 0xfa -- line 0x10
    "11111010", --  513 - 0x201  :  250 - 0xfa
    "11111010", --  514 - 0x202  :  250 - 0xfa
    "11111010", --  515 - 0x203  :  250 - 0xfa
    "11111010", --  516 - 0x204  :  250 - 0xfa
    "11111010", --  517 - 0x205  :  250 - 0xfa
    "11111010", --  518 - 0x206  :  250 - 0xfa
    "11111010", --  519 - 0x207  :  250 - 0xfa
    "11111010", --  520 - 0x208  :  250 - 0xfa
    "11111001", --  521 - 0x209  :  249 - 0xf9
    "11111010", --  522 - 0x20a  :  250 - 0xfa
    "11111010", --  523 - 0x20b  :  250 - 0xfa
    "11111010", --  524 - 0x20c  :  250 - 0xfa
    "11111010", --  525 - 0x20d  :  250 - 0xfa
    "11111010", --  526 - 0x20e  :  250 - 0xfa
    "11111010", --  527 - 0x20f  :  250 - 0xfa
    "11111010", --  528 - 0x210  :  250 - 0xfa
    "11111010", --  529 - 0x211  :  250 - 0xfa
    "11111010", --  530 - 0x212  :  250 - 0xfa
    "11111010", --  531 - 0x213  :  250 - 0xfa
    "11101001", --  532 - 0x214  :  233 - 0xe9
    "11111010", --  533 - 0x215  :  250 - 0xfa
    "11111010", --  534 - 0x216  :  250 - 0xfa
    "11111010", --  535 - 0x217  :  250 - 0xfa
    "11111010", --  536 - 0x218  :  250 - 0xfa
    "11111010", --  537 - 0x219  :  250 - 0xfa
    "11111010", --  538 - 0x21a  :  250 - 0xfa
    "11111010", --  539 - 0x21b  :  250 - 0xfa
    "11111010", --  540 - 0x21c  :  250 - 0xfa
    "11101010", --  541 - 0x21d  :  234 - 0xea
    "11111010", --  542 - 0x21e  :  250 - 0xfa
    "11111010", --  543 - 0x21f  :  250 - 0xfa
    "11111010", --  544 - 0x220  :  250 - 0xfa -- line 0x11
    "11111010", --  545 - 0x221  :  250 - 0xfa
    "11111010", --  546 - 0x222  :  250 - 0xfa
    "11111010", --  547 - 0x223  :  250 - 0xfa
    "11111010", --  548 - 0x224  :  250 - 0xfa
    "11111010", --  549 - 0x225  :  250 - 0xfa
    "11111010", --  550 - 0x226  :  250 - 0xfa
    "11111010", --  551 - 0x227  :  250 - 0xfa
    "11111010", --  552 - 0x228  :  250 - 0xfa
    "11111010", --  553 - 0x229  :  250 - 0xfa
    "11111010", --  554 - 0x22a  :  250 - 0xfa
    "11111010", --  555 - 0x22b  :  250 - 0xfa
    "11101010", --  556 - 0x22c  :  234 - 0xea
    "11111010", --  557 - 0x22d  :  250 - 0xfa
    "11111010", --  558 - 0x22e  :  250 - 0xfa
    "11111010", --  559 - 0x22f  :  250 - 0xfa
    "11111010", --  560 - 0x230  :  250 - 0xfa
    "11111010", --  561 - 0x231  :  250 - 0xfa
    "11111010", --  562 - 0x232  :  250 - 0xfa
    "11111010", --  563 - 0x233  :  250 - 0xfa
    "11101010", --  564 - 0x234  :  234 - 0xea
    "11111010", --  565 - 0x235  :  250 - 0xfa
    "11111010", --  566 - 0x236  :  250 - 0xfa
    "11111010", --  567 - 0x237  :  250 - 0xfa
    "11111010", --  568 - 0x238  :  250 - 0xfa
    "11111010", --  569 - 0x239  :  250 - 0xfa
    "11111010", --  570 - 0x23a  :  250 - 0xfa
    "11111001", --  571 - 0x23b  :  249 - 0xf9
    "11111010", --  572 - 0x23c  :  250 - 0xfa
    "11111010", --  573 - 0x23d  :  250 - 0xfa
    "11111010", --  574 - 0x23e  :  250 - 0xfa
    "11111010", --  575 - 0x23f  :  250 - 0xfa
    "11111010", --  576 - 0x240  :  250 - 0xfa -- line 0x12
    "11111010", --  577 - 0x241  :  250 - 0xfa
    "11111010", --  578 - 0x242  :  250 - 0xfa
    "11111010", --  579 - 0x243  :  250 - 0xfa
    "11111001", --  580 - 0x244  :  249 - 0xf9
    "11111010", --  581 - 0x245  :  250 - 0xfa
    "11111010", --  582 - 0x246  :  250 - 0xfa
    "11111010", --  583 - 0x247  :  250 - 0xfa
    "11111010", --  584 - 0x248  :  250 - 0xfa
    "11111010", --  585 - 0x249  :  250 - 0xfa
    "11111010", --  586 - 0x24a  :  250 - 0xfa
    "11111010", --  587 - 0x24b  :  250 - 0xfa
    "11111010", --  588 - 0x24c  :  250 - 0xfa
    "11111010", --  589 - 0x24d  :  250 - 0xfa
    "11111010", --  590 - 0x24e  :  250 - 0xfa
    "11111010", --  591 - 0x24f  :  250 - 0xfa
    "11111010", --  592 - 0x250  :  250 - 0xfa
    "11111010", --  593 - 0x251  :  250 - 0xfa
    "11111010", --  594 - 0x252  :  250 - 0xfa
    "11111001", --  595 - 0x253  :  249 - 0xf9
    "11111010", --  596 - 0x254  :  250 - 0xfa
    "11111010", --  597 - 0x255  :  250 - 0xfa
    "11111010", --  598 - 0x256  :  250 - 0xfa
    "11111010", --  599 - 0x257  :  250 - 0xfa
    "11111010", --  600 - 0x258  :  250 - 0xfa
    "11111010", --  601 - 0x259  :  250 - 0xfa
    "11111010", --  602 - 0x25a  :  250 - 0xfa
    "11111010", --  603 - 0x25b  :  250 - 0xfa
    "11111010", --  604 - 0x25c  :  250 - 0xfa
    "11111010", --  605 - 0x25d  :  250 - 0xfa
    "11111010", --  606 - 0x25e  :  250 - 0xfa
    "11111010", --  607 - 0x25f  :  250 - 0xfa
    "11111010", --  608 - 0x260  :  250 - 0xfa -- line 0x13
    "11111010", --  609 - 0x261  :  250 - 0xfa
    "11111010", --  610 - 0x262  :  250 - 0xfa
    "11111010", --  611 - 0x263  :  250 - 0xfa
    "11111010", --  612 - 0x264  :  250 - 0xfa
    "11111010", --  613 - 0x265  :  250 - 0xfa
    "11111010", --  614 - 0x266  :  250 - 0xfa
    "11111010", --  615 - 0x267  :  250 - 0xfa
    "11101001", --  616 - 0x268  :  233 - 0xe9
    "11111010", --  617 - 0x269  :  250 - 0xfa
    "11111010", --  618 - 0x26a  :  250 - 0xfa
    "11111010", --  619 - 0x26b  :  250 - 0xfa
    "11111010", --  620 - 0x26c  :  250 - 0xfa
    "11111010", --  621 - 0x26d  :  250 - 0xfa
    "11101001", --  622 - 0x26e  :  233 - 0xe9
    "11111010", --  623 - 0x26f  :  250 - 0xfa
    "11111010", --  624 - 0x270  :  250 - 0xfa
    "11111010", --  625 - 0x271  :  250 - 0xfa
    "11111010", --  626 - 0x272  :  250 - 0xfa
    "11111010", --  627 - 0x273  :  250 - 0xfa
    "11111010", --  628 - 0x274  :  250 - 0xfa
    "11111010", --  629 - 0x275  :  250 - 0xfa
    "11111010", --  630 - 0x276  :  250 - 0xfa
    "11101010", --  631 - 0x277  :  234 - 0xea
    "11101001", --  632 - 0x278  :  233 - 0xe9
    "11111010", --  633 - 0x279  :  250 - 0xfa
    "11111010", --  634 - 0x27a  :  250 - 0xfa
    "11111010", --  635 - 0x27b  :  250 - 0xfa
    "11111001", --  636 - 0x27c  :  249 - 0xf9
    "11111010", --  637 - 0x27d  :  250 - 0xfa
    "11111010", --  638 - 0x27e  :  250 - 0xfa
    "11111010", --  639 - 0x27f  :  250 - 0xfa
    "11111010", --  640 - 0x280  :  250 - 0xfa -- line 0x14
    "11111010", --  641 - 0x281  :  250 - 0xfa
    "11111010", --  642 - 0x282  :  250 - 0xfa
    "11111010", --  643 - 0x283  :  250 - 0xfa
    "11111010", --  644 - 0x284  :  250 - 0xfa
    "11111010", --  645 - 0x285  :  250 - 0xfa
    "11111010", --  646 - 0x286  :  250 - 0xfa
    "11111010", --  647 - 0x287  :  250 - 0xfa
    "11111010", --  648 - 0x288  :  250 - 0xfa
    "00100000", --  649 - 0x289  :   32 - 0x20
    "00100010", --  650 - 0x28a  :   34 - 0x22
    "00010101", --  651 - 0x28b  :   21 - 0x15
    "00100011", --  652 - 0x28c  :   35 - 0x23
    "00100011", --  653 - 0x28d  :   35 - 0x23
    "11111010", --  654 - 0x28e  :  250 - 0xfa
    "00100011", --  655 - 0x28f  :   35 - 0x23
    "00100100", --  656 - 0x290  :   36 - 0x24
    "00010001", --  657 - 0x291  :   17 - 0x11
    "00100010", --  658 - 0x292  :   34 - 0x22
    "00100100", --  659 - 0x293  :   36 - 0x24
    "11111010", --  660 - 0x294  :  250 - 0xfa
    "00100100", --  661 - 0x295  :   36 - 0x24
    "00011111", --  662 - 0x296  :   31 - 0x1f
    "11111010", --  663 - 0x297  :  250 - 0xfa
    "11111010", --  664 - 0x298  :  250 - 0xfa
    "11111010", --  665 - 0x299  :  250 - 0xfa
    "11111010", --  666 - 0x29a  :  250 - 0xfa
    "11111010", --  667 - 0x29b  :  250 - 0xfa
    "11111010", --  668 - 0x29c  :  250 - 0xfa
    "11111010", --  669 - 0x29d  :  250 - 0xfa
    "11111010", --  670 - 0x29e  :  250 - 0xfa
    "11111010", --  671 - 0x29f  :  250 - 0xfa
    "11111010", --  672 - 0x2a0  :  250 - 0xfa -- line 0x15
    "11111010", --  673 - 0x2a1  :  250 - 0xfa
    "11101010", --  674 - 0x2a2  :  234 - 0xea
    "11111010", --  675 - 0x2a3  :  250 - 0xfa
    "11111010", --  676 - 0x2a4  :  250 - 0xfa
    "11111010", --  677 - 0x2a5  :  250 - 0xfa
    "11111010", --  678 - 0x2a6  :  250 - 0xfa
    "11111010", --  679 - 0x2a7  :  250 - 0xfa
    "11111010", --  680 - 0x2a8  :  250 - 0xfa
    "11111010", --  681 - 0x2a9  :  250 - 0xfa
    "11111010", --  682 - 0x2aa  :  250 - 0xfa
    "11111010", --  683 - 0x2ab  :  250 - 0xfa
    "11111010", --  684 - 0x2ac  :  250 - 0xfa
    "11111010", --  685 - 0x2ad  :  250 - 0xfa
    "11111010", --  686 - 0x2ae  :  250 - 0xfa
    "11111010", --  687 - 0x2af  :  250 - 0xfa
    "11111010", --  688 - 0x2b0  :  250 - 0xfa
    "11111010", --  689 - 0x2b1  :  250 - 0xfa
    "11111010", --  690 - 0x2b2  :  250 - 0xfa
    "11111010", --  691 - 0x2b3  :  250 - 0xfa
    "11111010", --  692 - 0x2b4  :  250 - 0xfa
    "11111010", --  693 - 0x2b5  :  250 - 0xfa
    "11111010", --  694 - 0x2b6  :  250 - 0xfa
    "11111010", --  695 - 0x2b7  :  250 - 0xfa
    "11111010", --  696 - 0x2b8  :  250 - 0xfa
    "11111010", --  697 - 0x2b9  :  250 - 0xfa
    "11111010", --  698 - 0x2ba  :  250 - 0xfa
    "11111010", --  699 - 0x2bb  :  250 - 0xfa
    "11111010", --  700 - 0x2bc  :  250 - 0xfa
    "11111010", --  701 - 0x2bd  :  250 - 0xfa
    "11111010", --  702 - 0x2be  :  250 - 0xfa
    "11111010", --  703 - 0x2bf  :  250 - 0xfa
    "11111010", --  704 - 0x2c0  :  250 - 0xfa -- line 0x16
    "11111010", --  705 - 0x2c1  :  250 - 0xfa
    "11111010", --  706 - 0x2c2  :  250 - 0xfa
    "11111010", --  707 - 0x2c3  :  250 - 0xfa
    "11111010", --  708 - 0x2c4  :  250 - 0xfa
    "11111010", --  709 - 0x2c5  :  250 - 0xfa
    "11111010", --  710 - 0x2c6  :  250 - 0xfa
    "11111010", --  711 - 0x2c7  :  250 - 0xfa
    "11111010", --  712 - 0x2c8  :  250 - 0xfa
    "00010111", --  713 - 0x2c9  :   23 - 0x17
    "00011111", --  714 - 0x2ca  :   31 - 0x1f
    "11111010", --  715 - 0x2cb  :  250 - 0xfa
    "00010010", --  716 - 0x2cc  :   18 - 0x12
    "00010001", --  717 - 0x2cd  :   17 - 0x11
    "00010011", --  718 - 0x2ce  :   19 - 0x13
    "00011011", --  719 - 0x2cf  :   27 - 0x1b
    "11111010", --  720 - 0x2d0  :  250 - 0xfa
    "00100100", --  721 - 0x2d1  :   36 - 0x24
    "00011111", --  722 - 0x2d2  :   31 - 0x1f
    "11111010", --  723 - 0x2d3  :  250 - 0xfa
    "00011101", --  724 - 0x2d4  :   29 - 0x1d
    "00010101", --  725 - 0x2d5  :   21 - 0x15
    "00011110", --  726 - 0x2d6  :   30 - 0x1e
    "00100101", --  727 - 0x2d7  :   37 - 0x25
    "11111010", --  728 - 0x2d8  :  250 - 0xfa
    "11111010", --  729 - 0x2d9  :  250 - 0xfa
    "11111010", --  730 - 0x2da  :  250 - 0xfa
    "11111010", --  731 - 0x2db  :  250 - 0xfa
    "11111010", --  732 - 0x2dc  :  250 - 0xfa
    "11111010", --  733 - 0x2dd  :  250 - 0xfa
    "11111010", --  734 - 0x2de  :  250 - 0xfa
    "11111010", --  735 - 0x2df  :  250 - 0xfa
    "11111010", --  736 - 0x2e0  :  250 - 0xfa -- line 0x17
    "11111010", --  737 - 0x2e1  :  250 - 0xfa
    "11111010", --  738 - 0x2e2  :  250 - 0xfa
    "11111010", --  739 - 0x2e3  :  250 - 0xfa
    "11111010", --  740 - 0x2e4  :  250 - 0xfa
    "11111010", --  741 - 0x2e5  :  250 - 0xfa
    "11111010", --  742 - 0x2e6  :  250 - 0xfa
    "11111001", --  743 - 0x2e7  :  249 - 0xf9
    "11111010", --  744 - 0x2e8  :  250 - 0xfa
    "11111001", --  745 - 0x2e9  :  249 - 0xf9
    "11111010", --  746 - 0x2ea  :  250 - 0xfa
    "11111010", --  747 - 0x2eb  :  250 - 0xfa
    "11111010", --  748 - 0x2ec  :  250 - 0xfa
    "11111010", --  749 - 0x2ed  :  250 - 0xfa
    "11111010", --  750 - 0x2ee  :  250 - 0xfa
    "11111010", --  751 - 0x2ef  :  250 - 0xfa
    "11111010", --  752 - 0x2f0  :  250 - 0xfa
    "11111010", --  753 - 0x2f1  :  250 - 0xfa
    "11111010", --  754 - 0x2f2  :  250 - 0xfa
    "11111010", --  755 - 0x2f3  :  250 - 0xfa
    "11111010", --  756 - 0x2f4  :  250 - 0xfa
    "11111010", --  757 - 0x2f5  :  250 - 0xfa
    "11111010", --  758 - 0x2f6  :  250 - 0xfa
    "11111010", --  759 - 0x2f7  :  250 - 0xfa
    "11111010", --  760 - 0x2f8  :  250 - 0xfa
    "11111010", --  761 - 0x2f9  :  250 - 0xfa
    "11111010", --  762 - 0x2fa  :  250 - 0xfa
    "11111010", --  763 - 0x2fb  :  250 - 0xfa
    "11111010", --  764 - 0x2fc  :  250 - 0xfa
    "11111010", --  765 - 0x2fd  :  250 - 0xfa
    "11101010", --  766 - 0x2fe  :  234 - 0xea
    "11111010", --  767 - 0x2ff  :  250 - 0xfa
    "11111010", --  768 - 0x300  :  250 - 0xfa -- line 0x18
    "11111010", --  769 - 0x301  :  250 - 0xfa
    "11111010", --  770 - 0x302  :  250 - 0xfa
    "11111010", --  771 - 0x303  :  250 - 0xfa
    "11111010", --  772 - 0x304  :  250 - 0xfa
    "11111010", --  773 - 0x305  :  250 - 0xfa
    "11111010", --  774 - 0x306  :  250 - 0xfa
    "11111010", --  775 - 0x307  :  250 - 0xfa
    "11111010", --  776 - 0x308  :  250 - 0xfa
    "11111010", --  777 - 0x309  :  250 - 0xfa
    "11111010", --  778 - 0x30a  :  250 - 0xfa
    "11111010", --  779 - 0x30b  :  250 - 0xfa
    "11111010", --  780 - 0x30c  :  250 - 0xfa
    "11111010", --  781 - 0x30d  :  250 - 0xfa
    "11111010", --  782 - 0x30e  :  250 - 0xfa
    "11111010", --  783 - 0x30f  :  250 - 0xfa
    "11111001", --  784 - 0x310  :  249 - 0xf9
    "11111010", --  785 - 0x311  :  250 - 0xfa
    "11111010", --  786 - 0x312  :  250 - 0xfa
    "11111010", --  787 - 0x313  :  250 - 0xfa
    "11111010", --  788 - 0x314  :  250 - 0xfa
    "11111010", --  789 - 0x315  :  250 - 0xfa
    "11101001", --  790 - 0x316  :  233 - 0xe9
    "11111001", --  791 - 0x317  :  249 - 0xf9
    "11111010", --  792 - 0x318  :  250 - 0xfa
    "11111010", --  793 - 0x319  :  250 - 0xfa
    "11111001", --  794 - 0x31a  :  249 - 0xf9
    "11111010", --  795 - 0x31b  :  250 - 0xfa
    "11111010", --  796 - 0x31c  :  250 - 0xfa
    "11111010", --  797 - 0x31d  :  250 - 0xfa
    "11111010", --  798 - 0x31e  :  250 - 0xfa
    "11101001", --  799 - 0x31f  :  233 - 0xe9
    "11111010", --  800 - 0x320  :  250 - 0xfa -- line 0x19
    "11111010", --  801 - 0x321  :  250 - 0xfa
    "11111010", --  802 - 0x322  :  250 - 0xfa
    "11111010", --  803 - 0x323  :  250 - 0xfa
    "11111010", --  804 - 0x324  :  250 - 0xfa
    "11111010", --  805 - 0x325  :  250 - 0xfa
    "11111010", --  806 - 0x326  :  250 - 0xfa
    "11111010", --  807 - 0x327  :  250 - 0xfa
    "11111010", --  808 - 0x328  :  250 - 0xfa
    "11111010", --  809 - 0x329  :  250 - 0xfa
    "11111010", --  810 - 0x32a  :  250 - 0xfa
    "11111010", --  811 - 0x32b  :  250 - 0xfa
    "11111010", --  812 - 0x32c  :  250 - 0xfa
    "11111010", --  813 - 0x32d  :  250 - 0xfa
    "11111010", --  814 - 0x32e  :  250 - 0xfa
    "11111010", --  815 - 0x32f  :  250 - 0xfa
    "11111010", --  816 - 0x330  :  250 - 0xfa
    "11111010", --  817 - 0x331  :  250 - 0xfa
    "11111010", --  818 - 0x332  :  250 - 0xfa
    "11111010", --  819 - 0x333  :  250 - 0xfa
    "11111010", --  820 - 0x334  :  250 - 0xfa
    "11111010", --  821 - 0x335  :  250 - 0xfa
    "11111010", --  822 - 0x336  :  250 - 0xfa
    "11111010", --  823 - 0x337  :  250 - 0xfa
    "11111010", --  824 - 0x338  :  250 - 0xfa
    "11111010", --  825 - 0x339  :  250 - 0xfa
    "11111010", --  826 - 0x33a  :  250 - 0xfa
    "11111010", --  827 - 0x33b  :  250 - 0xfa
    "11111010", --  828 - 0x33c  :  250 - 0xfa
    "11111010", --  829 - 0x33d  :  250 - 0xfa
    "11111010", --  830 - 0x33e  :  250 - 0xfa
    "11111010", --  831 - 0x33f  :  250 - 0xfa
    "11111010", --  832 - 0x340  :  250 - 0xfa -- line 0x1a
    "11111010", --  833 - 0x341  :  250 - 0xfa
    "11111010", --  834 - 0x342  :  250 - 0xfa
    "11111010", --  835 - 0x343  :  250 - 0xfa
    "11111010", --  836 - 0x344  :  250 - 0xfa
    "11111010", --  837 - 0x345  :  250 - 0xfa
    "11111010", --  838 - 0x346  :  250 - 0xfa
    "11111010", --  839 - 0x347  :  250 - 0xfa
    "11111010", --  840 - 0x348  :  250 - 0xfa
    "11111010", --  841 - 0x349  :  250 - 0xfa
    "11111010", --  842 - 0x34a  :  250 - 0xfa
    "11101010", --  843 - 0x34b  :  234 - 0xea
    "11111010", --  844 - 0x34c  :  250 - 0xfa
    "11111010", --  845 - 0x34d  :  250 - 0xfa
    "11111010", --  846 - 0x34e  :  250 - 0xfa
    "11111010", --  847 - 0x34f  :  250 - 0xfa
    "11111010", --  848 - 0x350  :  250 - 0xfa
    "11111010", --  849 - 0x351  :  250 - 0xfa
    "11111010", --  850 - 0x352  :  250 - 0xfa
    "11111010", --  851 - 0x353  :  250 - 0xfa
    "11111010", --  852 - 0x354  :  250 - 0xfa
    "11111010", --  853 - 0x355  :  250 - 0xfa
    "11111010", --  854 - 0x356  :  250 - 0xfa
    "11111010", --  855 - 0x357  :  250 - 0xfa
    "11111010", --  856 - 0x358  :  250 - 0xfa
    "11111010", --  857 - 0x359  :  250 - 0xfa
    "11111010", --  858 - 0x35a  :  250 - 0xfa
    "11111010", --  859 - 0x35b  :  250 - 0xfa
    "11111010", --  860 - 0x35c  :  250 - 0xfa
    "11111010", --  861 - 0x35d  :  250 - 0xfa
    "11111010", --  862 - 0x35e  :  250 - 0xfa
    "11111010", --  863 - 0x35f  :  250 - 0xfa
    "11111010", --  864 - 0x360  :  250 - 0xfa -- line 0x1b
    "11111010", --  865 - 0x361  :  250 - 0xfa
    "11111010", --  866 - 0x362  :  250 - 0xfa
    "11111010", --  867 - 0x363  :  250 - 0xfa
    "11111010", --  868 - 0x364  :  250 - 0xfa
    "11111010", --  869 - 0x365  :  250 - 0xfa
    "11111010", --  870 - 0x366  :  250 - 0xfa
    "11111010", --  871 - 0x367  :  250 - 0xfa
    "11111010", --  872 - 0x368  :  250 - 0xfa
    "11111010", --  873 - 0x369  :  250 - 0xfa
    "11111010", --  874 - 0x36a  :  250 - 0xfa
    "11111010", --  875 - 0x36b  :  250 - 0xfa
    "11111010", --  876 - 0x36c  :  250 - 0xfa
    "11111010", --  877 - 0x36d  :  250 - 0xfa
    "11101001", --  878 - 0x36e  :  233 - 0xe9
    "11111010", --  879 - 0x36f  :  250 - 0xfa
    "11111010", --  880 - 0x370  :  250 - 0xfa
    "11111010", --  881 - 0x371  :  250 - 0xfa
    "11111010", --  882 - 0x372  :  250 - 0xfa
    "11111010", --  883 - 0x373  :  250 - 0xfa
    "11111010", --  884 - 0x374  :  250 - 0xfa
    "11111010", --  885 - 0x375  :  250 - 0xfa
    "11111010", --  886 - 0x376  :  250 - 0xfa
    "11111010", --  887 - 0x377  :  250 - 0xfa
    "11111010", --  888 - 0x378  :  250 - 0xfa
    "11111010", --  889 - 0x379  :  250 - 0xfa
    "11101010", --  890 - 0x37a  :  234 - 0xea
    "11111010", --  891 - 0x37b  :  250 - 0xfa
    "11111010", --  892 - 0x37c  :  250 - 0xfa
    "11111010", --  893 - 0x37d  :  250 - 0xfa
    "11111010", --  894 - 0x37e  :  250 - 0xfa
    "11111010", --  895 - 0x37f  :  250 - 0xfa
    "11111010", --  896 - 0x380  :  250 - 0xfa -- line 0x1c
    "11111010", --  897 - 0x381  :  250 - 0xfa
    "11111001", --  898 - 0x382  :  249 - 0xf9
    "11111010", --  899 - 0x383  :  250 - 0xfa
    "11111010", --  900 - 0x384  :  250 - 0xfa
    "11101010", --  901 - 0x385  :  234 - 0xea
    "11111010", --  902 - 0x386  :  250 - 0xfa
    "11111010", --  903 - 0x387  :  250 - 0xfa
    "11111010", --  904 - 0x388  :  250 - 0xfa
    "11101001", --  905 - 0x389  :  233 - 0xe9
    "11111010", --  906 - 0x38a  :  250 - 0xfa
    "11111010", --  907 - 0x38b  :  250 - 0xfa
    "11111010", --  908 - 0x38c  :  250 - 0xfa
    "11111010", --  909 - 0x38d  :  250 - 0xfa
    "11111010", --  910 - 0x38e  :  250 - 0xfa
    "11111010", --  911 - 0x38f  :  250 - 0xfa
    "11111010", --  912 - 0x390  :  250 - 0xfa
    "11111010", --  913 - 0x391  :  250 - 0xfa
    "11111001", --  914 - 0x392  :  249 - 0xf9
    "11111010", --  915 - 0x393  :  250 - 0xfa
    "11111010", --  916 - 0x394  :  250 - 0xfa
    "11111010", --  917 - 0x395  :  250 - 0xfa
    "11111010", --  918 - 0x396  :  250 - 0xfa
    "11111010", --  919 - 0x397  :  250 - 0xfa
    "11111010", --  920 - 0x398  :  250 - 0xfa
    "11111001", --  921 - 0x399  :  249 - 0xf9
    "11111010", --  922 - 0x39a  :  250 - 0xfa
    "11111010", --  923 - 0x39b  :  250 - 0xfa
    "11111010", --  924 - 0x39c  :  250 - 0xfa
    "11111010", --  925 - 0x39d  :  250 - 0xfa
    "11111001", --  926 - 0x39e  :  249 - 0xf9
    "11111010", --  927 - 0x39f  :  250 - 0xfa
    "11111010", --  928 - 0x3a0  :  250 - 0xfa -- line 0x1d
    "11111001", --  929 - 0x3a1  :  249 - 0xf9
    "11111010", --  930 - 0x3a2  :  250 - 0xfa
    "11111010", --  931 - 0x3a3  :  250 - 0xfa
    "11111010", --  932 - 0x3a4  :  250 - 0xfa
    "11111010", --  933 - 0x3a5  :  250 - 0xfa
    "11111010", --  934 - 0x3a6  :  250 - 0xfa
    "11111010", --  935 - 0x3a7  :  250 - 0xfa
    "11111010", --  936 - 0x3a8  :  250 - 0xfa
    "11111010", --  937 - 0x3a9  :  250 - 0xfa
    "11111010", --  938 - 0x3aa  :  250 - 0xfa
    "11111010", --  939 - 0x3ab  :  250 - 0xfa
    "11111010", --  940 - 0x3ac  :  250 - 0xfa
    "11111010", --  941 - 0x3ad  :  250 - 0xfa
    "11111010", --  942 - 0x3ae  :  250 - 0xfa
    "11111010", --  943 - 0x3af  :  250 - 0xfa
    "11111010", --  944 - 0x3b0  :  250 - 0xfa
    "11111010", --  945 - 0x3b1  :  250 - 0xfa
    "11111010", --  946 - 0x3b2  :  250 - 0xfa
    "11111010", --  947 - 0x3b3  :  250 - 0xfa
    "11111010", --  948 - 0x3b4  :  250 - 0xfa
    "11111010", --  949 - 0x3b5  :  250 - 0xfa
    "11111010", --  950 - 0x3b6  :  250 - 0xfa
    "11111010", --  951 - 0x3b7  :  250 - 0xfa
    "11111010", --  952 - 0x3b8  :  250 - 0xfa
    "11111010", --  953 - 0x3b9  :  250 - 0xfa
    "11111010", --  954 - 0x3ba  :  250 - 0xfa
    "11111010", --  955 - 0x3bb  :  250 - 0xfa
    "11111010", --  956 - 0x3bc  :  250 - 0xfa
    "11111010", --  957 - 0x3bd  :  250 - 0xfa
    "11111010", --  958 - 0x3be  :  250 - 0xfa
    "11111010", --  959 - 0x3bf  :  250 - 0xfa
        ---- Attribute Table 0----
    "01010101", --  960 - 0x3c0  :   85 - 0x55
    "01010101", --  961 - 0x3c1  :   85 - 0x55
    "01010101", --  962 - 0x3c2  :   85 - 0x55
    "01010101", --  963 - 0x3c3  :   85 - 0x55
    "01010101", --  964 - 0x3c4  :   85 - 0x55
    "01010101", --  965 - 0x3c5  :   85 - 0x55
    "01010101", --  966 - 0x3c6  :   85 - 0x55
    "01010101", --  967 - 0x3c7  :   85 - 0x55
    "01010101", --  968 - 0x3c8  :   85 - 0x55
    "01010101", --  969 - 0x3c9  :   85 - 0x55
    "01010101", --  970 - 0x3ca  :   85 - 0x55
    "01010101", --  971 - 0x3cb  :   85 - 0x55
    "01010101", --  972 - 0x3cc  :   85 - 0x55
    "01010101", --  973 - 0x3cd  :   85 - 0x55
    "01010101", --  974 - 0x3ce  :   85 - 0x55
    "01010101", --  975 - 0x3cf  :   85 - 0x55
    "01010101", --  976 - 0x3d0  :   85 - 0x55
    "01010101", --  977 - 0x3d1  :   85 - 0x55
    "01010101", --  978 - 0x3d2  :   85 - 0x55
    "01010101", --  979 - 0x3d3  :   85 - 0x55
    "01010101", --  980 - 0x3d4  :   85 - 0x55
    "01010101", --  981 - 0x3d5  :   85 - 0x55
    "01010101", --  982 - 0x3d6  :   85 - 0x55
    "01010101", --  983 - 0x3d7  :   85 - 0x55
    "01010101", --  984 - 0x3d8  :   85 - 0x55
    "01010101", --  985 - 0x3d9  :   85 - 0x55
    "01010101", --  986 - 0x3da  :   85 - 0x55
    "01010101", --  987 - 0x3db  :   85 - 0x55
    "01010101", --  988 - 0x3dc  :   85 - 0x55
    "01010101", --  989 - 0x3dd  :   85 - 0x55
    "01010101", --  990 - 0x3de  :   85 - 0x55
    "01010101", --  991 - 0x3df  :   85 - 0x55
    "01010101", --  992 - 0x3e0  :   85 - 0x55
    "01010101", --  993 - 0x3e1  :   85 - 0x55
    "01010101", --  994 - 0x3e2  :   85 - 0x55
    "01010101", --  995 - 0x3e3  :   85 - 0x55
    "01010101", --  996 - 0x3e4  :   85 - 0x55
    "01010101", --  997 - 0x3e5  :   85 - 0x55
    "01010101", --  998 - 0x3e6  :   85 - 0x55
    "01010101", --  999 - 0x3e7  :   85 - 0x55
    "01010101", -- 1000 - 0x3e8  :   85 - 0x55
    "01010101", -- 1001 - 0x3e9  :   85 - 0x55
    "01010101", -- 1002 - 0x3ea  :   85 - 0x55
    "01010101", -- 1003 - 0x3eb  :   85 - 0x55
    "01010101", -- 1004 - 0x3ec  :   85 - 0x55
    "01010101", -- 1005 - 0x3ed  :   85 - 0x55
    "01010101", -- 1006 - 0x3ee  :   85 - 0x55
    "01010101", -- 1007 - 0x3ef  :   85 - 0x55
    "01010101", -- 1008 - 0x3f0  :   85 - 0x55
    "01010101", -- 1009 - 0x3f1  :   85 - 0x55
    "01010101", -- 1010 - 0x3f2  :   85 - 0x55
    "01010101", -- 1011 - 0x3f3  :   85 - 0x55
    "01010101", -- 1012 - 0x3f4  :   85 - 0x55
    "01010101", -- 1013 - 0x3f5  :   85 - 0x55
    "01010101", -- 1014 - 0x3f6  :   85 - 0x55
    "01010101", -- 1015 - 0x3f7  :   85 - 0x55
    "00000101", -- 1016 - 0x3f8  :    5 - 0x5
    "00000101", -- 1017 - 0x3f9  :    5 - 0x5
    "00000101", -- 1018 - 0x3fa  :    5 - 0x5
    "00000101", -- 1019 - 0x3fb  :    5 - 0x5
    "00000101", -- 1020 - 0x3fc  :    5 - 0x5
    "00000101", -- 1021 - 0x3fd  :    5 - 0x5
    "00000101", -- 1022 - 0x3fe  :    5 - 0x5
    "00000101"  -- 1023 - 0x3ff  :    5 - 0x5
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
