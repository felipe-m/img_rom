//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_NOVA_color0
  (
     //input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout  = 8'b00001111; //    1 :  15 - 0xf
      12'h2: dout  = 8'b00000100; //    2 :   4 - 0x4
      12'h3: dout  = 8'b00000011; //    3 :   3 - 0x3
      12'h4: dout  = 8'b00000011; //    4 :   3 - 0x3
      12'h5: dout  = 8'b00000011; //    5 :   3 - 0x3
      12'h6: dout  = 8'b00000100; //    6 :   4 - 0x4
      12'h7: dout  = 8'b00111010; //    7 :  58 - 0x3a
      12'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      12'h9: dout  = 8'b00111000; //    9 :  56 - 0x38
      12'hA: dout  = 8'b11000110; //   10 : 198 - 0xc6
      12'hB: dout  = 8'b11001011; //   11 : 203 - 0xcb
      12'hC: dout  = 8'b11011100; //   12 : 220 - 0xdc
      12'hD: dout  = 8'b00111010; //   13 :  58 - 0x3a
      12'hE: dout  = 8'b10011010; //   14 : 154 - 0x9a
      12'hF: dout  = 8'b10000001; //   15 : 129 - 0x81
      12'h10: dout  = 8'b01000101; //   16 :  69 - 0x45 -- Sprite 0x2
      12'h11: dout  = 8'b10000111; //   17 : 135 - 0x87
      12'h12: dout  = 8'b10000011; //   18 : 131 - 0x83
      12'h13: dout  = 8'b10000001; //   19 : 129 - 0x81
      12'h14: dout  = 8'b10000001; //   20 : 129 - 0x81
      12'h15: dout  = 8'b10000001; //   21 : 129 - 0x81
      12'h16: dout  = 8'b01000001; //   22 :  65 - 0x41
      12'h17: dout  = 8'b00100001; //   23 :  33 - 0x21
      12'h18: dout  = 8'b01111111; //   24 : 127 - 0x7f -- Sprite 0x3
      12'h19: dout  = 8'b01111110; //   25 : 126 - 0x7e
      12'h1A: dout  = 8'b11111100; //   26 : 252 - 0xfc
      12'h1B: dout  = 8'b00111000; //   27 :  56 - 0x38
      12'h1C: dout  = 8'b00011000; //   28 :  24 - 0x18
      12'h1D: dout  = 8'b10001100; //   29 : 140 - 0x8c
      12'h1E: dout  = 8'b11000100; //   30 : 196 - 0xc4
      12'h1F: dout  = 8'b11111100; //   31 : 252 - 0xfc
      12'h20: dout  = 8'b00100011; //   32 :  35 - 0x23 -- Sprite 0x4
      12'h21: dout  = 8'b00100011; //   33 :  35 - 0x23
      12'h22: dout  = 8'b00100001; //   34 :  33 - 0x21
      12'h23: dout  = 8'b00100000; //   35 :  32 - 0x20
      12'h24: dout  = 8'b00010011; //   36 :  19 - 0x13
      12'h25: dout  = 8'b00001100; //   37 :  12 - 0xc
      12'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      12'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout  = 8'b11111100; //   40 : 252 - 0xfc -- Sprite 0x5
      12'h29: dout  = 8'b11111100; //   41 : 252 - 0xfc
      12'h2A: dout  = 8'b11111100; //   42 : 252 - 0xfc
      12'h2B: dout  = 8'b11111100; //   43 : 252 - 0xfc
      12'h2C: dout  = 8'b10010000; //   44 : 144 - 0x90
      12'h2D: dout  = 8'b10010000; //   45 : 144 - 0x90
      12'h2E: dout  = 8'b10001000; //   46 : 136 - 0x88
      12'h2F: dout  = 8'b11111000; //   47 : 248 - 0xf8
      12'h30: dout  = 8'b00100011; //   48 :  35 - 0x23 -- Sprite 0x6
      12'h31: dout  = 8'b00100011; //   49 :  35 - 0x23
      12'h32: dout  = 8'b00100001; //   50 :  33 - 0x21
      12'h33: dout  = 8'b00100000; //   51 :  32 - 0x20
      12'h34: dout  = 8'b00010011; //   52 :  19 - 0x13
      12'h35: dout  = 8'b00001101; //   53 :  13 - 0xd
      12'h36: dout  = 8'b00000010; //   54 :   2 - 0x2
      12'h37: dout  = 8'b00000001; //   55 :   1 - 0x1
      12'h38: dout  = 8'b11111100; //   56 : 252 - 0xfc -- Sprite 0x7
      12'h39: dout  = 8'b11111100; //   57 : 252 - 0xfc
      12'h3A: dout  = 8'b11111100; //   58 : 252 - 0xfc
      12'h3B: dout  = 8'b11111100; //   59 : 252 - 0xfc
      12'h3C: dout  = 8'b10100100; //   60 : 164 - 0xa4
      12'h3D: dout  = 8'b00100100; //   61 :  36 - 0x24
      12'h3E: dout  = 8'b01010010; //   62 :  82 - 0x52
      12'h3F: dout  = 8'b11101110; //   63 : 238 - 0xee
      12'h40: dout  = 8'b00100011; //   64 :  35 - 0x23 -- Sprite 0x8
      12'h41: dout  = 8'b00100011; //   65 :  35 - 0x23
      12'h42: dout  = 8'b00100001; //   66 :  33 - 0x21
      12'h43: dout  = 8'b00100000; //   67 :  32 - 0x20
      12'h44: dout  = 8'b00010011; //   68 :  19 - 0x13
      12'h45: dout  = 8'b00001101; //   69 :  13 - 0xd
      12'h46: dout  = 8'b00000001; //   70 :   1 - 0x1
      12'h47: dout  = 8'b00000001; //   71 :   1 - 0x1
      12'h48: dout  = 8'b11111110; //   72 : 254 - 0xfe -- Sprite 0x9
      12'h49: dout  = 8'b11111110; //   73 : 254 - 0xfe
      12'h4A: dout  = 8'b11111110; //   74 : 254 - 0xfe
      12'h4B: dout  = 8'b11111111; //   75 : 255 - 0xff
      12'h4C: dout  = 8'b10010001; //   76 : 145 - 0x91
      12'h4D: dout  = 8'b00101111; //   77 :  47 - 0x2f
      12'h4E: dout  = 8'b01000000; //   78 :  64 - 0x40
      12'h4F: dout  = 8'b11100000; //   79 : 224 - 0xe0
      12'h50: dout  = 8'b00100011; //   80 :  35 - 0x23 -- Sprite 0xa
      12'h51: dout  = 8'b00100011; //   81 :  35 - 0x23
      12'h52: dout  = 8'b00100001; //   82 :  33 - 0x21
      12'h53: dout  = 8'b00100000; //   83 :  32 - 0x20
      12'h54: dout  = 8'b00010011; //   84 :  19 - 0x13
      12'h55: dout  = 8'b00001110; //   85 :  14 - 0xe
      12'h56: dout  = 8'b00000001; //   86 :   1 - 0x1
      12'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      12'h58: dout  = 8'b11111110; //   88 : 254 - 0xfe -- Sprite 0xb
      12'h59: dout  = 8'b11111110; //   89 : 254 - 0xfe
      12'h5A: dout  = 8'b11111110; //   90 : 254 - 0xfe
      12'h5B: dout  = 8'b11111100; //   91 : 252 - 0xfc
      12'h5C: dout  = 8'b00100100; //   92 :  36 - 0x24
      12'h5D: dout  = 8'b00100010; //   93 :  34 - 0x22
      12'h5E: dout  = 8'b11010010; //   94 : 210 - 0xd2
      12'h5F: dout  = 8'b00001111; //   95 :  15 - 0xf
      12'h60: dout  = 8'b01111111; //   96 : 127 - 0x7f -- Sprite 0xc
      12'h61: dout  = 8'b01111110; //   97 : 126 - 0x7e
      12'h62: dout  = 8'b11111100; //   98 : 252 - 0xfc
      12'h63: dout  = 8'b00000010; //   99 :   2 - 0x2
      12'h64: dout  = 8'b00000100; //  100 :   4 - 0x4
      12'h65: dout  = 8'b11111100; //  101 : 252 - 0xfc
      12'h66: dout  = 8'b11111100; //  102 : 252 - 0xfc
      12'h67: dout  = 8'b11111110; //  103 : 254 - 0xfe
      12'h68: dout  = 8'b01000101; //  104 :  69 - 0x45 -- Sprite 0xd
      12'h69: dout  = 8'b10000111; //  105 : 135 - 0x87
      12'h6A: dout  = 8'b10000011; //  106 : 131 - 0x83
      12'h6B: dout  = 8'b10000010; //  107 : 130 - 0x82
      12'h6C: dout  = 8'b10000010; //  108 : 130 - 0x82
      12'h6D: dout  = 8'b10000100; //  109 : 132 - 0x84
      12'h6E: dout  = 8'b01000100; //  110 :  68 - 0x44
      12'h6F: dout  = 8'b00100100; //  111 :  36 - 0x24
      12'h70: dout  = 8'b01111111; //  112 : 127 - 0x7f -- Sprite 0xe
      12'h71: dout  = 8'b01111110; //  113 : 126 - 0x7e
      12'h72: dout  = 8'b11111100; //  114 : 252 - 0xfc
      12'h73: dout  = 8'b11111000; //  115 : 248 - 0xf8
      12'h74: dout  = 8'b01111000; //  116 : 120 - 0x78
      12'h75: dout  = 8'b01111100; //  117 : 124 - 0x7c
      12'h76: dout  = 8'b11111100; //  118 : 252 - 0xfc
      12'h77: dout  = 8'b11111110; //  119 : 254 - 0xfe
      12'h78: dout  = 8'b00000000; //  120 :   0 - 0x0 -- Sprite 0xf
      12'h79: dout  = 8'b00001111; //  121 :  15 - 0xf
      12'h7A: dout  = 8'b00000100; //  122 :   4 - 0x4
      12'h7B: dout  = 8'b00000011; //  123 :   3 - 0x3
      12'h7C: dout  = 8'b00000011; //  124 :   3 - 0x3
      12'h7D: dout  = 8'b00000011; //  125 :   3 - 0x3
      12'h7E: dout  = 8'b00000100; //  126 :   4 - 0x4
      12'h7F: dout  = 8'b00000010; //  127 :   2 - 0x2
      12'h80: dout  = 8'b00000111; //  128 :   7 - 0x7 -- Sprite 0x10
      12'h81: dout  = 8'b00001100; //  129 :  12 - 0xc
      12'h82: dout  = 8'b00010000; //  130 :  16 - 0x10
      12'h83: dout  = 8'b00010000; //  131 :  16 - 0x10
      12'h84: dout  = 8'b00010000; //  132 :  16 - 0x10
      12'h85: dout  = 8'b00100000; //  133 :  32 - 0x20
      12'h86: dout  = 8'b00100000; //  134 :  32 - 0x20
      12'h87: dout  = 8'b00100001; //  135 :  33 - 0x21
      12'h88: dout  = 8'b11111111; //  136 : 255 - 0xff -- Sprite 0x11
      12'h89: dout  = 8'b01111110; //  137 : 126 - 0x7e
      12'h8A: dout  = 8'b01111100; //  138 : 124 - 0x7c
      12'h8B: dout  = 8'b01111000; //  139 : 120 - 0x78
      12'h8C: dout  = 8'b01011000; //  140 :  88 - 0x58
      12'h8D: dout  = 8'b10001100; //  141 : 140 - 0x8c
      12'h8E: dout  = 8'b11000100; //  142 : 196 - 0xc4
      12'h8F: dout  = 8'b11111100; //  143 : 252 - 0xfc
      12'h90: dout  = 8'b00100011; //  144 :  35 - 0x23 -- Sprite 0x12
      12'h91: dout  = 8'b00100011; //  145 :  35 - 0x23
      12'h92: dout  = 8'b00100001; //  146 :  33 - 0x21
      12'h93: dout  = 8'b00100000; //  147 :  32 - 0x20
      12'h94: dout  = 8'b00010011; //  148 :  19 - 0x13
      12'h95: dout  = 8'b00001100; //  149 :  12 - 0xc
      12'h96: dout  = 8'b00000000; //  150 :   0 - 0x0
      12'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      12'h98: dout  = 8'b00000001; //  152 :   1 - 0x1 -- Sprite 0x13
      12'h99: dout  = 8'b00000001; //  153 :   1 - 0x1
      12'h9A: dout  = 8'b00000011; //  154 :   3 - 0x3
      12'h9B: dout  = 8'b00000100; //  155 :   4 - 0x4
      12'h9C: dout  = 8'b00001000; //  156 :   8 - 0x8
      12'h9D: dout  = 8'b00010000; //  157 :  16 - 0x10
      12'h9E: dout  = 8'b00010000; //  158 :  16 - 0x10
      12'h9F: dout  = 8'b00100000; //  159 :  32 - 0x20
      12'hA0: dout  = 8'b01111111; //  160 : 127 - 0x7f -- Sprite 0x14
      12'hA1: dout  = 8'b11111110; //  161 : 254 - 0xfe
      12'hA2: dout  = 8'b00000110; //  162 :   6 - 0x6
      12'hA3: dout  = 8'b00000001; //  163 :   1 - 0x1
      12'hA4: dout  = 8'b00000001; //  164 :   1 - 0x1
      12'hA5: dout  = 8'b00000001; //  165 :   1 - 0x1
      12'hA6: dout  = 8'b00000111; //  166 :   7 - 0x7
      12'hA7: dout  = 8'b11111110; //  167 : 254 - 0xfe
      12'hA8: dout  = 8'b00000101; //  168 :   5 - 0x5 -- Sprite 0x15
      12'hA9: dout  = 8'b00000101; //  169 :   5 - 0x5
      12'hAA: dout  = 8'b00000111; //  170 :   7 - 0x7
      12'hAB: dout  = 8'b00000100; //  171 :   4 - 0x4
      12'hAC: dout  = 8'b00000100; //  172 :   4 - 0x4
      12'hAD: dout  = 8'b00001111; //  173 :  15 - 0xf
      12'hAE: dout  = 8'b00110000; //  174 :  48 - 0x30
      12'hAF: dout  = 8'b01000000; //  175 :  64 - 0x40
      12'hB0: dout  = 8'b11111100; //  176 : 252 - 0xfc -- Sprite 0x16
      12'hB1: dout  = 8'b11111000; //  177 : 248 - 0xf8
      12'hB2: dout  = 8'b11110000; //  178 : 240 - 0xf0
      12'hB3: dout  = 8'b11100000; //  179 : 224 - 0xe0
      12'hB4: dout  = 8'b01100000; //  180 :  96 - 0x60
      12'hB5: dout  = 8'b11110000; //  181 : 240 - 0xf0
      12'hB6: dout  = 8'b00011100; //  182 :  28 - 0x1c
      12'hB7: dout  = 8'b00000010; //  183 :   2 - 0x2
      12'hB8: dout  = 8'b10000000; //  184 : 128 - 0x80 -- Sprite 0x17
      12'hB9: dout  = 8'b10000000; //  185 : 128 - 0x80
      12'hBA: dout  = 8'b10000000; //  186 : 128 - 0x80
      12'hBB: dout  = 8'b10000011; //  187 : 131 - 0x83
      12'hBC: dout  = 8'b01001111; //  188 :  79 - 0x4f
      12'hBD: dout  = 8'b00110010; //  189 :  50 - 0x32
      12'hBE: dout  = 8'b00000010; //  190 :   2 - 0x2
      12'hBF: dout  = 8'b00000011; //  191 :   3 - 0x3
      12'hC0: dout  = 8'b00000010; //  192 :   2 - 0x2 -- Sprite 0x18
      12'hC1: dout  = 8'b00000001; //  193 :   1 - 0x1
      12'hC2: dout  = 8'b00000010; //  194 :   2 - 0x2
      12'hC3: dout  = 8'b11111100; //  195 : 252 - 0xfc
      12'hC4: dout  = 8'b11000000; //  196 : 192 - 0xc0
      12'hC5: dout  = 8'b01000000; //  197 :  64 - 0x40
      12'hC6: dout  = 8'b00100000; //  198 :  32 - 0x20
      12'hC7: dout  = 8'b11100000; //  199 : 224 - 0xe0
      12'hC8: dout  = 8'b00001011; //  200 :  11 - 0xb -- Sprite 0x19
      12'hC9: dout  = 8'b00001011; //  201 :  11 - 0xb
      12'hCA: dout  = 8'b00001111; //  202 :  15 - 0xf
      12'hCB: dout  = 8'b00001001; //  203 :   9 - 0x9
      12'hCC: dout  = 8'b00001000; //  204 :   8 - 0x8
      12'hCD: dout  = 8'b00001001; //  205 :   9 - 0x9
      12'hCE: dout  = 8'b00001111; //  206 :  15 - 0xf
      12'hCF: dout  = 8'b00110000; //  207 :  48 - 0x30
      12'hD0: dout  = 8'b11111000; //  208 : 248 - 0xf8 -- Sprite 0x1a
      12'hD1: dout  = 8'b11110000; //  209 : 240 - 0xf0
      12'hD2: dout  = 8'b11100000; //  210 : 224 - 0xe0
      12'hD3: dout  = 8'b11000000; //  211 : 192 - 0xc0
      12'hD4: dout  = 8'b11000000; //  212 : 192 - 0xc0
      12'hD5: dout  = 8'b11000000; //  213 : 192 - 0xc0
      12'hD6: dout  = 8'b11111000; //  214 : 248 - 0xf8
      12'hD7: dout  = 8'b00011111; //  215 :  31 - 0x1f
      12'hD8: dout  = 8'b01000000; //  216 :  64 - 0x40 -- Sprite 0x1b
      12'hD9: dout  = 8'b01000000; //  217 :  64 - 0x40
      12'hDA: dout  = 8'b10000000; //  218 : 128 - 0x80
      12'hDB: dout  = 8'b10000000; //  219 : 128 - 0x80
      12'hDC: dout  = 8'b01000000; //  220 :  64 - 0x40
      12'hDD: dout  = 8'b00111111; //  221 :  63 - 0x3f
      12'hDE: dout  = 8'b00000100; //  222 :   4 - 0x4
      12'hDF: dout  = 8'b00000111; //  223 :   7 - 0x7
      12'hE0: dout  = 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0x1c
      12'hE1: dout  = 8'b00000000; //  225 :   0 - 0x0
      12'hE2: dout  = 8'b00000000; //  226 :   0 - 0x0
      12'hE3: dout  = 8'b00000000; //  227 :   0 - 0x0
      12'hE4: dout  = 8'b00000000; //  228 :   0 - 0x0
      12'hE5: dout  = 8'b11111111; //  229 : 255 - 0xff
      12'hE6: dout  = 8'b01000000; //  230 :  64 - 0x40
      12'hE7: dout  = 8'b11000000; //  231 : 192 - 0xc0
      12'hE8: dout  = 8'b11000000; //  232 : 192 - 0xc0 -- Sprite 0x1d
      12'hE9: dout  = 8'b00100000; //  233 :  32 - 0x20
      12'hEA: dout  = 8'b00100000; //  234 :  32 - 0x20
      12'hEB: dout  = 8'b00100000; //  235 :  32 - 0x20
      12'hEC: dout  = 8'b01000000; //  236 :  64 - 0x40
      12'hED: dout  = 8'b10000000; //  237 : 128 - 0x80
      12'hEE: dout  = 8'b00000000; //  238 :   0 - 0x0
      12'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      12'hF0: dout  = 8'b01111111; //  240 : 127 - 0x7f -- Sprite 0x1e
      12'hF1: dout  = 8'b01100010; //  241 :  98 - 0x62
      12'hF2: dout  = 8'b11000100; //  242 : 196 - 0xc4
      12'hF3: dout  = 8'b00011000; //  243 :  24 - 0x18
      12'hF4: dout  = 8'b00111100; //  244 :  60 - 0x3c
      12'hF5: dout  = 8'b11111110; //  245 : 254 - 0xfe
      12'hF6: dout  = 8'b11111110; //  246 : 254 - 0xfe
      12'hF7: dout  = 8'b11111110; //  247 : 254 - 0xfe
      12'hF8: dout  = 8'b00000000; //  248 :   0 - 0x0 -- Sprite 0x1f
      12'hF9: dout  = 8'b00111000; //  249 :  56 - 0x38
      12'hFA: dout  = 8'b11000110; //  250 : 198 - 0xc6
      12'hFB: dout  = 8'b11001011; //  251 : 203 - 0xcb
      12'hFC: dout  = 8'b11011100; //  252 : 220 - 0xdc
      12'hFD: dout  = 8'b00111010; //  253 :  58 - 0x3a
      12'hFE: dout  = 8'b10011010; //  254 : 154 - 0x9a
      12'hFF: dout  = 8'b11100001; //  255 : 225 - 0xe1
      12'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      12'h101: dout  = 8'b00011100; //  257 :  28 - 0x1c
      12'h102: dout  = 8'b00010011; //  258 :  19 - 0x13
      12'h103: dout  = 8'b00001000; //  259 :   8 - 0x8
      12'h104: dout  = 8'b00010000; //  260 :  16 - 0x10
      12'h105: dout  = 8'b00001000; //  261 :   8 - 0x8
      12'h106: dout  = 8'b00010000; //  262 :  16 - 0x10
      12'h107: dout  = 8'b00010000; //  263 :  16 - 0x10
      12'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- Sprite 0x21
      12'h109: dout  = 8'b00111000; //  265 :  56 - 0x38
      12'h10A: dout  = 8'b11001000; //  266 : 200 - 0xc8
      12'h10B: dout  = 8'b00010000; //  267 :  16 - 0x10
      12'h10C: dout  = 8'b00001000; //  268 :   8 - 0x8
      12'h10D: dout  = 8'b00010000; //  269 :  16 - 0x10
      12'h10E: dout  = 8'b00001000; //  270 :   8 - 0x8
      12'h10F: dout  = 8'b00001000; //  271 :   8 - 0x8
      12'h110: dout  = 8'b00001000; //  272 :   8 - 0x8 -- Sprite 0x22
      12'h111: dout  = 8'b00011100; //  273 :  28 - 0x1c
      12'h112: dout  = 8'b00100111; //  274 :  39 - 0x27
      12'h113: dout  = 8'b00101111; //  275 :  47 - 0x2f
      12'h114: dout  = 8'b00011111; //  276 :  31 - 0x1f
      12'h115: dout  = 8'b00001111; //  277 :  15 - 0xf
      12'h116: dout  = 8'b00001111; //  278 :  15 - 0xf
      12'h117: dout  = 8'b00001111; //  279 :  15 - 0xf
      12'h118: dout  = 8'b00010000; //  280 :  16 - 0x10 -- Sprite 0x23
      12'h119: dout  = 8'b00111100; //  281 :  60 - 0x3c
      12'h11A: dout  = 8'b11000010; //  282 : 194 - 0xc2
      12'h11B: dout  = 8'b10000010; //  283 : 130 - 0x82
      12'h11C: dout  = 8'b10000010; //  284 : 130 - 0x82
      12'h11D: dout  = 8'b10000010; //  285 : 130 - 0x82
      12'h11E: dout  = 8'b00010010; //  286 :  18 - 0x12
      12'h11F: dout  = 8'b00011100; //  287 :  28 - 0x1c
      12'h120: dout  = 8'b00001111; //  288 :  15 - 0xf -- Sprite 0x24
      12'h121: dout  = 8'b00001110; //  289 :  14 - 0xe
      12'h122: dout  = 8'b00010100; //  290 :  20 - 0x14
      12'h123: dout  = 8'b00010100; //  291 :  20 - 0x14
      12'h124: dout  = 8'b00010010; //  292 :  18 - 0x12
      12'h125: dout  = 8'b00100101; //  293 :  37 - 0x25
      12'h126: dout  = 8'b01000100; //  294 :  68 - 0x44
      12'h127: dout  = 8'b00111000; //  295 :  56 - 0x38
      12'h128: dout  = 8'b00010000; //  296 :  16 - 0x10 -- Sprite 0x25
      12'h129: dout  = 8'b00010000; //  297 :  16 - 0x10
      12'h12A: dout  = 8'b00010000; //  298 :  16 - 0x10
      12'h12B: dout  = 8'b00101100; //  299 :  44 - 0x2c
      12'h12C: dout  = 8'b01000100; //  300 :  68 - 0x44
      12'h12D: dout  = 8'b11000100; //  301 : 196 - 0xc4
      12'h12E: dout  = 8'b00111000; //  302 :  56 - 0x38
      12'h12F: dout  = 8'b00000000; //  303 :   0 - 0x0
      12'h130: dout  = 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      12'h131: dout  = 8'b00000000; //  305 :   0 - 0x0
      12'h132: dout  = 8'b00000000; //  306 :   0 - 0x0
      12'h133: dout  = 8'b00000000; //  307 :   0 - 0x0
      12'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      12'h135: dout  = 8'b00000000; //  309 :   0 - 0x0
      12'h136: dout  = 8'b00000000; //  310 :   0 - 0x0
      12'h137: dout  = 8'b00000000; //  311 :   0 - 0x0
      12'h138: dout  = 8'b00000000; //  312 :   0 - 0x0 -- Sprite 0x27
      12'h139: dout  = 8'b00000000; //  313 :   0 - 0x0
      12'h13A: dout  = 8'b00000000; //  314 :   0 - 0x0
      12'h13B: dout  = 8'b00000000; //  315 :   0 - 0x0
      12'h13C: dout  = 8'b00000000; //  316 :   0 - 0x0
      12'h13D: dout  = 8'b00000000; //  317 :   0 - 0x0
      12'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      12'h141: dout  = 8'b00000000; //  321 :   0 - 0x0
      12'h142: dout  = 8'b00000000; //  322 :   0 - 0x0
      12'h143: dout  = 8'b00000000; //  323 :   0 - 0x0
      12'h144: dout  = 8'b00000000; //  324 :   0 - 0x0
      12'h145: dout  = 8'b00000000; //  325 :   0 - 0x0
      12'h146: dout  = 8'b00000000; //  326 :   0 - 0x0
      12'h147: dout  = 8'b00000000; //  327 :   0 - 0x0
      12'h148: dout  = 8'b00100000; //  328 :  32 - 0x20 -- Sprite 0x29
      12'h149: dout  = 8'b00100000; //  329 :  32 - 0x20
      12'h14A: dout  = 8'b00100000; //  330 :  32 - 0x20
      12'h14B: dout  = 8'b00100000; //  331 :  32 - 0x20
      12'h14C: dout  = 8'b00010011; //  332 :  19 - 0x13
      12'h14D: dout  = 8'b00001101; //  333 :  13 - 0xd
      12'h14E: dout  = 8'b00000010; //  334 :   2 - 0x2
      12'h14F: dout  = 8'b00000001; //  335 :   1 - 0x1
      12'h150: dout  = 8'b00100000; //  336 :  32 - 0x20 -- Sprite 0x2a
      12'h151: dout  = 8'b00100000; //  337 :  32 - 0x20
      12'h152: dout  = 8'b00100000; //  338 :  32 - 0x20
      12'h153: dout  = 8'b00100000; //  339 :  32 - 0x20
      12'h154: dout  = 8'b00010011; //  340 :  19 - 0x13
      12'h155: dout  = 8'b00001101; //  341 :  13 - 0xd
      12'h156: dout  = 8'b00000001; //  342 :   1 - 0x1
      12'h157: dout  = 8'b00000001; //  343 :   1 - 0x1
      12'h158: dout  = 8'b00000000; //  344 :   0 - 0x0 -- Sprite 0x2b
      12'h159: dout  = 8'b00000000; //  345 :   0 - 0x0
      12'h15A: dout  = 8'b00000000; //  346 :   0 - 0x0
      12'h15B: dout  = 8'b00000000; //  347 :   0 - 0x0
      12'h15C: dout  = 8'b00000000; //  348 :   0 - 0x0
      12'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      12'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      12'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout  = 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x2c
      12'h161: dout  = 8'b00000000; //  353 :   0 - 0x0
      12'h162: dout  = 8'b00000000; //  354 :   0 - 0x0
      12'h163: dout  = 8'b00000000; //  355 :   0 - 0x0
      12'h164: dout  = 8'b00000000; //  356 :   0 - 0x0
      12'h165: dout  = 8'b00000000; //  357 :   0 - 0x0
      12'h166: dout  = 8'b00000000; //  358 :   0 - 0x0
      12'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout  = 8'b00111100; //  360 :  60 - 0x3c -- Sprite 0x2d
      12'h169: dout  = 8'b00000000; //  361 :   0 - 0x0
      12'h16A: dout  = 8'b10000001; //  362 : 129 - 0x81
      12'h16B: dout  = 8'b10011001; //  363 : 153 - 0x99
      12'h16C: dout  = 8'b10011001; //  364 : 153 - 0x99
      12'h16D: dout  = 8'b10000001; //  365 : 129 - 0x81
      12'h16E: dout  = 8'b00000000; //  366 :   0 - 0x0
      12'h16F: dout  = 8'b00111100; //  367 :  60 - 0x3c
      12'h170: dout  = 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x2e
      12'h171: dout  = 8'b00000000; //  369 :   0 - 0x0
      12'h172: dout  = 8'b00000000; //  370 :   0 - 0x0
      12'h173: dout  = 8'b00000000; //  371 :   0 - 0x0
      12'h174: dout  = 8'b00000000; //  372 :   0 - 0x0
      12'h175: dout  = 8'b00000000; //  373 :   0 - 0x0
      12'h176: dout  = 8'b00000000; //  374 :   0 - 0x0
      12'h177: dout  = 8'b00000000; //  375 :   0 - 0x0
      12'h178: dout  = 8'b10011111; //  376 : 159 - 0x9f -- Sprite 0x2f
      12'h179: dout  = 8'b10011110; //  377 : 158 - 0x9e
      12'h17A: dout  = 8'b10011100; //  378 : 156 - 0x9c
      12'h17B: dout  = 8'b00011000; //  379 :  24 - 0x18
      12'h17C: dout  = 8'b00111000; //  380 :  56 - 0x38
      12'h17D: dout  = 8'b11111100; //  381 : 252 - 0xfc
      12'h17E: dout  = 8'b11111100; //  382 : 252 - 0xfc
      12'h17F: dout  = 8'b11111100; //  383 : 252 - 0xfc
      12'h180: dout  = 8'b01111111; //  384 : 127 - 0x7f -- Sprite 0x30
      12'h181: dout  = 8'b01111110; //  385 : 126 - 0x7e
      12'h182: dout  = 8'b11111100; //  386 : 252 - 0xfc
      12'h183: dout  = 8'b00111000; //  387 :  56 - 0x38
      12'h184: dout  = 8'b00111000; //  388 :  56 - 0x38
      12'h185: dout  = 8'b00000100; //  389 :   4 - 0x4
      12'h186: dout  = 8'b10000100; //  390 : 132 - 0x84
      12'h187: dout  = 8'b11111100; //  391 : 252 - 0xfc
      12'h188: dout  = 8'b01111111; //  392 : 127 - 0x7f -- Sprite 0x31
      12'h189: dout  = 8'b01111110; //  393 : 126 - 0x7e
      12'h18A: dout  = 8'b11111100; //  394 : 252 - 0xfc
      12'h18B: dout  = 8'b00111000; //  395 :  56 - 0x38
      12'h18C: dout  = 8'b00111000; //  396 :  56 - 0x38
      12'h18D: dout  = 8'b00011100; //  397 :  28 - 0x1c
      12'h18E: dout  = 8'b10000100; //  398 : 132 - 0x84
      12'h18F: dout  = 8'b11000100; //  399 : 196 - 0xc4
      12'h190: dout  = 8'b01111111; //  400 : 127 - 0x7f -- Sprite 0x32
      12'h191: dout  = 8'b01111110; //  401 : 126 - 0x7e
      12'h192: dout  = 8'b11111100; //  402 : 252 - 0xfc
      12'h193: dout  = 8'b00111000; //  403 :  56 - 0x38
      12'h194: dout  = 8'b00100100; //  404 :  36 - 0x24
      12'h195: dout  = 8'b00000100; //  405 :   4 - 0x4
      12'h196: dout  = 8'b10011100; //  406 : 156 - 0x9c
      12'h197: dout  = 8'b11111100; //  407 : 252 - 0xfc
      12'h198: dout  = 8'b00100011; //  408 :  35 - 0x23 -- Sprite 0x33
      12'h199: dout  = 8'b00100011; //  409 :  35 - 0x23
      12'h19A: dout  = 8'b00100001; //  410 :  33 - 0x21
      12'h19B: dout  = 8'b00100000; //  411 :  32 - 0x20
      12'h19C: dout  = 8'b00010011; //  412 :  19 - 0x13
      12'h19D: dout  = 8'b00001101; //  413 :  13 - 0xd
      12'h19E: dout  = 8'b00000001; //  414 :   1 - 0x1
      12'h19F: dout  = 8'b00000001; //  415 :   1 - 0x1
      12'h1A0: dout  = 8'b11111100; //  416 : 252 - 0xfc -- Sprite 0x34
      12'h1A1: dout  = 8'b11111100; //  417 : 252 - 0xfc
      12'h1A2: dout  = 8'b11111100; //  418 : 252 - 0xfc
      12'h1A3: dout  = 8'b11111100; //  419 : 252 - 0xfc
      12'h1A4: dout  = 8'b10100100; //  420 : 164 - 0xa4
      12'h1A5: dout  = 8'b00100100; //  421 :  36 - 0x24
      12'h1A6: dout  = 8'b00010010; //  422 :  18 - 0x12
      12'h1A7: dout  = 8'b11101110; //  423 : 238 - 0xee
      12'h1A8: dout  = 8'b00100011; //  424 :  35 - 0x23 -- Sprite 0x35
      12'h1A9: dout  = 8'b00100011; //  425 :  35 - 0x23
      12'h1AA: dout  = 8'b00100001; //  426 :  33 - 0x21
      12'h1AB: dout  = 8'b00100000; //  427 :  32 - 0x20
      12'h1AC: dout  = 8'b00010011; //  428 :  19 - 0x13
      12'h1AD: dout  = 8'b00001110; //  429 :  14 - 0xe
      12'h1AE: dout  = 8'b00000010; //  430 :   2 - 0x2
      12'h1AF: dout  = 8'b00000001; //  431 :   1 - 0x1
      12'h1B0: dout  = 8'b11111100; //  432 : 252 - 0xfc -- Sprite 0x36
      12'h1B1: dout  = 8'b11111100; //  433 : 252 - 0xfc
      12'h1B2: dout  = 8'b11111100; //  434 : 252 - 0xfc
      12'h1B3: dout  = 8'b11111100; //  435 : 252 - 0xfc
      12'h1B4: dout  = 8'b10100110; //  436 : 166 - 0xa6
      12'h1B5: dout  = 8'b00110001; //  437 :  49 - 0x31
      12'h1B6: dout  = 8'b01001001; //  438 :  73 - 0x49
      12'h1B7: dout  = 8'b11000110; //  439 : 198 - 0xc6
      12'h1B8: dout  = 8'b11111100; //  440 : 252 - 0xfc -- Sprite 0x37
      12'h1B9: dout  = 8'b11111100; //  441 : 252 - 0xfc
      12'h1BA: dout  = 8'b11111100; //  442 : 252 - 0xfc
      12'h1BB: dout  = 8'b11111100; //  443 : 252 - 0xfc
      12'h1BC: dout  = 8'b10100100; //  444 : 164 - 0xa4
      12'h1BD: dout  = 8'b00100100; //  445 :  36 - 0x24
      12'h1BE: dout  = 8'b00010010; //  446 :  18 - 0x12
      12'h1BF: dout  = 8'b11101110; //  447 : 238 - 0xee
      12'h1C0: dout  = 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      12'h1C1: dout  = 8'b00000000; //  449 :   0 - 0x0
      12'h1C2: dout  = 8'b00000000; //  450 :   0 - 0x0
      12'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      12'h1C4: dout  = 8'b00000000; //  452 :   0 - 0x0
      12'h1C5: dout  = 8'b00000000; //  453 :   0 - 0x0
      12'h1C6: dout  = 8'b00000000; //  454 :   0 - 0x0
      12'h1C7: dout  = 8'b00000000; //  455 :   0 - 0x0
      12'h1C8: dout  = 8'b00000000; //  456 :   0 - 0x0 -- Sprite 0x39
      12'h1C9: dout  = 8'b00000000; //  457 :   0 - 0x0
      12'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      12'h1CC: dout  = 8'b00000000; //  460 :   0 - 0x0
      12'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      12'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      12'h1D2: dout  = 8'b00000000; //  466 :   0 - 0x0
      12'h1D3: dout  = 8'b00000000; //  467 :   0 - 0x0
      12'h1D4: dout  = 8'b00000000; //  468 :   0 - 0x0
      12'h1D5: dout  = 8'b00000000; //  469 :   0 - 0x0
      12'h1D6: dout  = 8'b00000000; //  470 :   0 - 0x0
      12'h1D7: dout  = 8'b00000000; //  471 :   0 - 0x0
      12'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0 -- Sprite 0x3b
      12'h1D9: dout  = 8'b00000000; //  473 :   0 - 0x0
      12'h1DA: dout  = 8'b00000000; //  474 :   0 - 0x0
      12'h1DB: dout  = 8'b00000000; //  475 :   0 - 0x0
      12'h1DC: dout  = 8'b00000000; //  476 :   0 - 0x0
      12'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      12'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      12'h1E1: dout  = 8'b00000000; //  481 :   0 - 0x0
      12'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      12'h1E3: dout  = 8'b00000000; //  483 :   0 - 0x0
      12'h1E4: dout  = 8'b00000000; //  484 :   0 - 0x0
      12'h1E5: dout  = 8'b00000000; //  485 :   0 - 0x0
      12'h1E6: dout  = 8'b00000000; //  486 :   0 - 0x0
      12'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      12'h1E9: dout  = 8'b00000000; //  489 :   0 - 0x0
      12'h1EA: dout  = 8'b00000000; //  490 :   0 - 0x0
      12'h1EB: dout  = 8'b00000000; //  491 :   0 - 0x0
      12'h1EC: dout  = 8'b00000000; //  492 :   0 - 0x0
      12'h1ED: dout  = 8'b00000000; //  493 :   0 - 0x0
      12'h1EE: dout  = 8'b00000000; //  494 :   0 - 0x0
      12'h1EF: dout  = 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      12'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      12'h1F2: dout  = 8'b00000000; //  498 :   0 - 0x0
      12'h1F3: dout  = 8'b00000000; //  499 :   0 - 0x0
      12'h1F4: dout  = 8'b00000000; //  500 :   0 - 0x0
      12'h1F5: dout  = 8'b00000000; //  501 :   0 - 0x0
      12'h1F6: dout  = 8'b00000000; //  502 :   0 - 0x0
      12'h1F7: dout  = 8'b00000000; //  503 :   0 - 0x0
      12'h1F8: dout  = 8'b00000000; //  504 :   0 - 0x0 -- Sprite 0x3f
      12'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout  = 8'b00000000; //  507 :   0 - 0x0
      12'h1FC: dout  = 8'b00000000; //  508 :   0 - 0x0
      12'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      12'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout  = 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x40
      12'h201: dout  = 8'b00111110; //  513 :  62 - 0x3e
      12'h202: dout  = 8'b01111111; //  514 : 127 - 0x7f
      12'h203: dout  = 8'b01111111; //  515 : 127 - 0x7f
      12'h204: dout  = 8'b01111111; //  516 : 127 - 0x7f
      12'h205: dout  = 8'b01111111; //  517 : 127 - 0x7f
      12'h206: dout  = 8'b01111111; //  518 : 127 - 0x7f
      12'h207: dout  = 8'b00111110; //  519 :  62 - 0x3e
      12'h208: dout  = 8'b00000000; //  520 :   0 - 0x0 -- Sprite 0x41
      12'h209: dout  = 8'b00111100; //  521 :  60 - 0x3c
      12'h20A: dout  = 8'b00011100; //  522 :  28 - 0x1c
      12'h20B: dout  = 8'b00011100; //  523 :  28 - 0x1c
      12'h20C: dout  = 8'b00011100; //  524 :  28 - 0x1c
      12'h20D: dout  = 8'b00011100; //  525 :  28 - 0x1c
      12'h20E: dout  = 8'b00011100; //  526 :  28 - 0x1c
      12'h20F: dout  = 8'b00011100; //  527 :  28 - 0x1c
      12'h210: dout  = 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x42
      12'h211: dout  = 8'b01111100; //  529 : 124 - 0x7c
      12'h212: dout  = 8'b01111111; //  530 : 127 - 0x7f
      12'h213: dout  = 8'b01100111; //  531 : 103 - 0x67
      12'h214: dout  = 8'b00111111; //  532 :  63 - 0x3f
      12'h215: dout  = 8'b01111110; //  533 : 126 - 0x7e
      12'h216: dout  = 8'b01111111; //  534 : 127 - 0x7f
      12'h217: dout  = 8'b01111111; //  535 : 127 - 0x7f
      12'h218: dout  = 8'b00000000; //  536 :   0 - 0x0 -- Sprite 0x43
      12'h219: dout  = 8'b01111110; //  537 : 126 - 0x7e
      12'h21A: dout  = 8'b01111111; //  538 : 127 - 0x7f
      12'h21B: dout  = 8'b01111111; //  539 : 127 - 0x7f
      12'h21C: dout  = 8'b00011111; //  540 :  31 - 0x1f
      12'h21D: dout  = 8'b01110111; //  541 : 119 - 0x77
      12'h21E: dout  = 8'b01111111; //  542 : 127 - 0x7f
      12'h21F: dout  = 8'b01111110; //  543 : 126 - 0x7e
      12'h220: dout  = 8'b00000000; //  544 :   0 - 0x0 -- Sprite 0x44
      12'h221: dout  = 8'b00001110; //  545 :  14 - 0xe
      12'h222: dout  = 8'b00011110; //  546 :  30 - 0x1e
      12'h223: dout  = 8'b00111110; //  547 :  62 - 0x3e
      12'h224: dout  = 8'b01111110; //  548 : 126 - 0x7e
      12'h225: dout  = 8'b01111111; //  549 : 127 - 0x7f
      12'h226: dout  = 8'b01111110; //  550 : 126 - 0x7e
      12'h227: dout  = 8'b00001100; //  551 :  12 - 0xc
      12'h228: dout  = 8'b00000000; //  552 :   0 - 0x0 -- Sprite 0x45
      12'h229: dout  = 8'b01111111; //  553 : 127 - 0x7f
      12'h22A: dout  = 8'b01111111; //  554 : 127 - 0x7f
      12'h22B: dout  = 8'b01111111; //  555 : 127 - 0x7f
      12'h22C: dout  = 8'b01111111; //  556 : 127 - 0x7f
      12'h22D: dout  = 8'b01110111; //  557 : 119 - 0x77
      12'h22E: dout  = 8'b01111111; //  558 : 127 - 0x7f
      12'h22F: dout  = 8'b01111110; //  559 : 126 - 0x7e
      12'h230: dout  = 8'b00000000; //  560 :   0 - 0x0 -- Sprite 0x46
      12'h231: dout  = 8'b00111110; //  561 :  62 - 0x3e
      12'h232: dout  = 8'b01111110; //  562 : 126 - 0x7e
      12'h233: dout  = 8'b01111111; //  563 : 127 - 0x7f
      12'h234: dout  = 8'b01111111; //  564 : 127 - 0x7f
      12'h235: dout  = 8'b01110111; //  565 : 119 - 0x77
      12'h236: dout  = 8'b01111111; //  566 : 127 - 0x7f
      12'h237: dout  = 8'b00111110; //  567 :  62 - 0x3e
      12'h238: dout  = 8'b00000000; //  568 :   0 - 0x0 -- Sprite 0x47
      12'h239: dout  = 8'b01111110; //  569 : 126 - 0x7e
      12'h23A: dout  = 8'b01111110; //  570 : 126 - 0x7e
      12'h23B: dout  = 8'b00011110; //  571 :  30 - 0x1e
      12'h23C: dout  = 8'b00011100; //  572 :  28 - 0x1c
      12'h23D: dout  = 8'b00111100; //  573 :  60 - 0x3c
      12'h23E: dout  = 8'b00111000; //  574 :  56 - 0x38
      12'h23F: dout  = 8'b00111000; //  575 :  56 - 0x38
      12'h240: dout  = 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x48
      12'h241: dout  = 8'b00111110; //  577 :  62 - 0x3e
      12'h242: dout  = 8'b01111111; //  578 : 127 - 0x7f
      12'h243: dout  = 8'b01111111; //  579 : 127 - 0x7f
      12'h244: dout  = 8'b01111111; //  580 : 127 - 0x7f
      12'h245: dout  = 8'b01111111; //  581 : 127 - 0x7f
      12'h246: dout  = 8'b01111111; //  582 : 127 - 0x7f
      12'h247: dout  = 8'b00111110; //  583 :  62 - 0x3e
      12'h248: dout  = 8'b00000000; //  584 :   0 - 0x0 -- Sprite 0x49
      12'h249: dout  = 8'b00111110; //  585 :  62 - 0x3e
      12'h24A: dout  = 8'b01111111; //  586 : 127 - 0x7f
      12'h24B: dout  = 8'b01110111; //  587 : 119 - 0x77
      12'h24C: dout  = 8'b01111111; //  588 : 127 - 0x7f
      12'h24D: dout  = 8'b01111111; //  589 : 127 - 0x7f
      12'h24E: dout  = 8'b00111111; //  590 :  63 - 0x3f
      12'h24F: dout  = 8'b00111110; //  591 :  62 - 0x3e
      12'h250: dout  = 8'b11111111; //  592 : 255 - 0xff -- Sprite 0x4a
      12'h251: dout  = 8'b10011001; //  593 : 153 - 0x99
      12'h252: dout  = 8'b10011001; //  594 : 153 - 0x99
      12'h253: dout  = 8'b10011001; //  595 : 153 - 0x99
      12'h254: dout  = 8'b10011001; //  596 : 153 - 0x99
      12'h255: dout  = 8'b10011001; //  597 : 153 - 0x99
      12'h256: dout  = 8'b10011001; //  598 : 153 - 0x99
      12'h257: dout  = 8'b11111111; //  599 : 255 - 0xff
      12'h258: dout  = 8'b11110000; //  600 : 240 - 0xf0 -- Sprite 0x4b
      12'h259: dout  = 8'b10010000; //  601 : 144 - 0x90
      12'h25A: dout  = 8'b10010000; //  602 : 144 - 0x90
      12'h25B: dout  = 8'b10010000; //  603 : 144 - 0x90
      12'h25C: dout  = 8'b10010000; //  604 : 144 - 0x90
      12'h25D: dout  = 8'b10010000; //  605 : 144 - 0x90
      12'h25E: dout  = 8'b10010000; //  606 : 144 - 0x90
      12'h25F: dout  = 8'b11110000; //  607 : 240 - 0xf0
      12'h260: dout  = 8'b11111111; //  608 : 255 - 0xff -- Sprite 0x4c
      12'h261: dout  = 8'b11111111; //  609 : 255 - 0xff
      12'h262: dout  = 8'b11111111; //  610 : 255 - 0xff
      12'h263: dout  = 8'b11111111; //  611 : 255 - 0xff
      12'h264: dout  = 8'b11111111; //  612 : 255 - 0xff
      12'h265: dout  = 8'b11111111; //  613 : 255 - 0xff
      12'h266: dout  = 8'b11111111; //  614 : 255 - 0xff
      12'h267: dout  = 8'b11111111; //  615 : 255 - 0xff
      12'h268: dout  = 8'b11111111; //  616 : 255 - 0xff -- Sprite 0x4d
      12'h269: dout  = 8'b11111111; //  617 : 255 - 0xff
      12'h26A: dout  = 8'b11111111; //  618 : 255 - 0xff
      12'h26B: dout  = 8'b11111111; //  619 : 255 - 0xff
      12'h26C: dout  = 8'b11111111; //  620 : 255 - 0xff
      12'h26D: dout  = 8'b11111111; //  621 : 255 - 0xff
      12'h26E: dout  = 8'b11111111; //  622 : 255 - 0xff
      12'h26F: dout  = 8'b11111111; //  623 : 255 - 0xff
      12'h270: dout  = 8'b11111111; //  624 : 255 - 0xff -- Sprite 0x4e
      12'h271: dout  = 8'b11111111; //  625 : 255 - 0xff
      12'h272: dout  = 8'b11111111; //  626 : 255 - 0xff
      12'h273: dout  = 8'b11111111; //  627 : 255 - 0xff
      12'h274: dout  = 8'b11111111; //  628 : 255 - 0xff
      12'h275: dout  = 8'b11111111; //  629 : 255 - 0xff
      12'h276: dout  = 8'b11111111; //  630 : 255 - 0xff
      12'h277: dout  = 8'b11111111; //  631 : 255 - 0xff
      12'h278: dout  = 8'b11111111; //  632 : 255 - 0xff -- Sprite 0x4f
      12'h279: dout  = 8'b11111111; //  633 : 255 - 0xff
      12'h27A: dout  = 8'b11111111; //  634 : 255 - 0xff
      12'h27B: dout  = 8'b11111111; //  635 : 255 - 0xff
      12'h27C: dout  = 8'b11111111; //  636 : 255 - 0xff
      12'h27D: dout  = 8'b11111111; //  637 : 255 - 0xff
      12'h27E: dout  = 8'b11111111; //  638 : 255 - 0xff
      12'h27F: dout  = 8'b11111111; //  639 : 255 - 0xff
      12'h280: dout  = 8'b00010000; //  640 :  16 - 0x10 -- Sprite 0x50
      12'h281: dout  = 8'b00101000; //  641 :  40 - 0x28
      12'h282: dout  = 8'b11101110; //  642 : 238 - 0xee
      12'h283: dout  = 8'b10000010; //  643 : 130 - 0x82
      12'h284: dout  = 8'b01000100; //  644 :  68 - 0x44
      12'h285: dout  = 8'b01000100; //  645 :  68 - 0x44
      12'h286: dout  = 8'b10010010; //  646 : 146 - 0x92
      12'h287: dout  = 8'b11101110; //  647 : 238 - 0xee
      12'h288: dout  = 8'b00010000; //  648 :  16 - 0x10 -- Sprite 0x51
      12'h289: dout  = 8'b00101000; //  649 :  40 - 0x28
      12'h28A: dout  = 8'b11101110; //  650 : 238 - 0xee
      12'h28B: dout  = 8'b10000010; //  651 : 130 - 0x82
      12'h28C: dout  = 8'b01000100; //  652 :  68 - 0x44
      12'h28D: dout  = 8'b01000100; //  653 :  68 - 0x44
      12'h28E: dout  = 8'b10010010; //  654 : 146 - 0x92
      12'h28F: dout  = 8'b11101110; //  655 : 238 - 0xee
      12'h290: dout  = 8'b00010000; //  656 :  16 - 0x10 -- Sprite 0x52
      12'h291: dout  = 8'b00111000; //  657 :  56 - 0x38
      12'h292: dout  = 8'b11111110; //  658 : 254 - 0xfe
      12'h293: dout  = 8'b11111110; //  659 : 254 - 0xfe
      12'h294: dout  = 8'b01111100; //  660 : 124 - 0x7c
      12'h295: dout  = 8'b01111100; //  661 : 124 - 0x7c
      12'h296: dout  = 8'b11111110; //  662 : 254 - 0xfe
      12'h297: dout  = 8'b11101110; //  663 : 238 - 0xee
      12'h298: dout  = 8'b11111111; //  664 : 255 - 0xff -- Sprite 0x53
      12'h299: dout  = 8'b11111111; //  665 : 255 - 0xff
      12'h29A: dout  = 8'b11111111; //  666 : 255 - 0xff
      12'h29B: dout  = 8'b11111111; //  667 : 255 - 0xff
      12'h29C: dout  = 8'b11111111; //  668 : 255 - 0xff
      12'h29D: dout  = 8'b11111111; //  669 : 255 - 0xff
      12'h29E: dout  = 8'b11111111; //  670 : 255 - 0xff
      12'h29F: dout  = 8'b11111111; //  671 : 255 - 0xff
      12'h2A0: dout  = 8'b00000000; //  672 :   0 - 0x0 -- Sprite 0x54
      12'h2A1: dout  = 8'b00000000; //  673 :   0 - 0x0
      12'h2A2: dout  = 8'b00000000; //  674 :   0 - 0x0
      12'h2A3: dout  = 8'b00000000; //  675 :   0 - 0x0
      12'h2A4: dout  = 8'b00000000; //  676 :   0 - 0x0
      12'h2A5: dout  = 8'b00000000; //  677 :   0 - 0x0
      12'h2A6: dout  = 8'b00000000; //  678 :   0 - 0x0
      12'h2A7: dout  = 8'b00000000; //  679 :   0 - 0x0
      12'h2A8: dout  = 8'b11111111; //  680 : 255 - 0xff -- Sprite 0x55
      12'h2A9: dout  = 8'b11111111; //  681 : 255 - 0xff
      12'h2AA: dout  = 8'b11111111; //  682 : 255 - 0xff
      12'h2AB: dout  = 8'b11111111; //  683 : 255 - 0xff
      12'h2AC: dout  = 8'b11111111; //  684 : 255 - 0xff
      12'h2AD: dout  = 8'b11111111; //  685 : 255 - 0xff
      12'h2AE: dout  = 8'b11111111; //  686 : 255 - 0xff
      12'h2AF: dout  = 8'b11111111; //  687 : 255 - 0xff
      12'h2B0: dout  = 8'b00101010; //  688 :  42 - 0x2a -- Sprite 0x56
      12'h2B1: dout  = 8'b01000101; //  689 :  69 - 0x45
      12'h2B2: dout  = 8'b00001000; //  690 :   8 - 0x8
      12'h2B3: dout  = 8'b00010101; //  691 :  21 - 0x15
      12'h2B4: dout  = 8'b00100000; //  692 :  32 - 0x20
      12'h2B5: dout  = 8'b01000101; //  693 :  69 - 0x45
      12'h2B6: dout  = 8'b10101000; //  694 : 168 - 0xa8
      12'h2B7: dout  = 8'b00000000; //  695 :   0 - 0x0
      12'h2B8: dout  = 8'b00001000; //  696 :   8 - 0x8 -- Sprite 0x57
      12'h2B9: dout  = 8'b01010101; //  697 :  85 - 0x55
      12'h2BA: dout  = 8'b10100000; //  698 : 160 - 0xa0
      12'h2BB: dout  = 8'b00010000; //  699 :  16 - 0x10
      12'h2BC: dout  = 8'b10000000; //  700 : 128 - 0x80
      12'h2BD: dout  = 8'b00010100; //  701 :  20 - 0x14
      12'h2BE: dout  = 8'b00100010; //  702 :  34 - 0x22
      12'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout  = 8'b11111111; //  704 : 255 - 0xff -- Sprite 0x58
      12'h2C1: dout  = 8'b11010101; //  705 : 213 - 0xd5
      12'h2C2: dout  = 8'b10100000; //  706 : 160 - 0xa0
      12'h2C3: dout  = 8'b11010000; //  707 : 208 - 0xd0
      12'h2C4: dout  = 8'b10001111; //  708 : 143 - 0x8f
      12'h2C5: dout  = 8'b11001000; //  709 : 200 - 0xc8
      12'h2C6: dout  = 8'b10001000; //  710 : 136 - 0x88
      12'h2C7: dout  = 8'b11001000; //  711 : 200 - 0xc8
      12'h2C8: dout  = 8'b10001000; //  712 : 136 - 0x88 -- Sprite 0x59
      12'h2C9: dout  = 8'b11001000; //  713 : 200 - 0xc8
      12'h2CA: dout  = 8'b10001000; //  714 : 136 - 0x88
      12'h2CB: dout  = 8'b11001111; //  715 : 207 - 0xcf
      12'h2CC: dout  = 8'b10010000; //  716 : 144 - 0x90
      12'h2CD: dout  = 8'b11100000; //  717 : 224 - 0xe0
      12'h2CE: dout  = 8'b11101010; //  718 : 234 - 0xea
      12'h2CF: dout  = 8'b11111111; //  719 : 255 - 0xff
      12'h2D0: dout  = 8'b11111111; //  720 : 255 - 0xff -- Sprite 0x5a
      12'h2D1: dout  = 8'b01011011; //  721 :  91 - 0x5b
      12'h2D2: dout  = 8'b00000111; //  722 :   7 - 0x7
      12'h2D3: dout  = 8'b00001001; //  723 :   9 - 0x9
      12'h2D4: dout  = 8'b11110011; //  724 : 243 - 0xf3
      12'h2D5: dout  = 8'b00010001; //  725 :  17 - 0x11
      12'h2D6: dout  = 8'b00010011; //  726 :  19 - 0x13
      12'h2D7: dout  = 8'b00010001; //  727 :  17 - 0x11
      12'h2D8: dout  = 8'b00010011; //  728 :  19 - 0x13 -- Sprite 0x5b
      12'h2D9: dout  = 8'b00010001; //  729 :  17 - 0x11
      12'h2DA: dout  = 8'b00010011; //  730 :  19 - 0x13
      12'h2DB: dout  = 8'b11110001; //  731 : 241 - 0xf1
      12'h2DC: dout  = 8'b00001011; //  732 :  11 - 0xb
      12'h2DD: dout  = 8'b00000101; //  733 :   5 - 0x5
      12'h2DE: dout  = 8'b10101011; //  734 : 171 - 0xab
      12'h2DF: dout  = 8'b11111111; //  735 : 255 - 0xff
      12'h2E0: dout  = 8'b00011100; //  736 :  28 - 0x1c -- Sprite 0x5c
      12'h2E1: dout  = 8'b00100010; //  737 :  34 - 0x22
      12'h2E2: dout  = 8'b01000001; //  738 :  65 - 0x41
      12'h2E3: dout  = 8'b01000001; //  739 :  65 - 0x41
      12'h2E4: dout  = 8'b01000001; //  740 :  65 - 0x41
      12'h2E5: dout  = 8'b00100010; //  741 :  34 - 0x22
      12'h2E6: dout  = 8'b00100010; //  742 :  34 - 0x22
      12'h2E7: dout  = 8'b00011100; //  743 :  28 - 0x1c
      12'h2E8: dout  = 8'b00001000; //  744 :   8 - 0x8 -- Sprite 0x5d
      12'h2E9: dout  = 8'b00010000; //  745 :  16 - 0x10
      12'h2EA: dout  = 8'b00010000; //  746 :  16 - 0x10
      12'h2EB: dout  = 8'b00001000; //  747 :   8 - 0x8
      12'h2EC: dout  = 8'b00000100; //  748 :   4 - 0x4
      12'h2ED: dout  = 8'b00000100; //  749 :   4 - 0x4
      12'h2EE: dout  = 8'b00001000; //  750 :   8 - 0x8
      12'h2EF: dout  = 8'b00010000; //  751 :  16 - 0x10
      12'h2F0: dout  = 8'b00110110; //  752 :  54 - 0x36 -- Sprite 0x5e
      12'h2F1: dout  = 8'b01101011; //  753 : 107 - 0x6b
      12'h2F2: dout  = 8'b01001001; //  754 :  73 - 0x49
      12'h2F3: dout  = 8'b01000001; //  755 :  65 - 0x41
      12'h2F4: dout  = 8'b01000001; //  756 :  65 - 0x41
      12'h2F5: dout  = 8'b00100010; //  757 :  34 - 0x22
      12'h2F6: dout  = 8'b00010100; //  758 :  20 - 0x14
      12'h2F7: dout  = 8'b00001000; //  759 :   8 - 0x8
      12'h2F8: dout  = 8'b00111110; //  760 :  62 - 0x3e -- Sprite 0x5f
      12'h2F9: dout  = 8'b01101011; //  761 : 107 - 0x6b
      12'h2FA: dout  = 8'b00100010; //  762 :  34 - 0x22
      12'h2FB: dout  = 8'b01100011; //  763 :  99 - 0x63
      12'h2FC: dout  = 8'b00100010; //  764 :  34 - 0x22
      12'h2FD: dout  = 8'b01100011; //  765 :  99 - 0x63
      12'h2FE: dout  = 8'b00100010; //  766 :  34 - 0x22
      12'h2FF: dout  = 8'b01111111; //  767 : 127 - 0x7f
      12'h300: dout  = 8'b11111111; //  768 : 255 - 0xff -- Sprite 0x60
      12'h301: dout  = 8'b11111111; //  769 : 255 - 0xff
      12'h302: dout  = 8'b11111111; //  770 : 255 - 0xff
      12'h303: dout  = 8'b11111111; //  771 : 255 - 0xff
      12'h304: dout  = 8'b11010101; //  772 : 213 - 0xd5
      12'h305: dout  = 8'b10101010; //  773 : 170 - 0xaa
      12'h306: dout  = 8'b11010101; //  774 : 213 - 0xd5
      12'h307: dout  = 8'b11111111; //  775 : 255 - 0xff
      12'h308: dout  = 8'b11111111; //  776 : 255 - 0xff -- Sprite 0x61
      12'h309: dout  = 8'b11111111; //  777 : 255 - 0xff
      12'h30A: dout  = 8'b11111111; //  778 : 255 - 0xff
      12'h30B: dout  = 8'b11111111; //  779 : 255 - 0xff
      12'h30C: dout  = 8'b01010101; //  780 :  85 - 0x55
      12'h30D: dout  = 8'b10101010; //  781 : 170 - 0xaa
      12'h30E: dout  = 8'b01010101; //  782 :  85 - 0x55
      12'h30F: dout  = 8'b11111111; //  783 : 255 - 0xff
      12'h310: dout  = 8'b11111111; //  784 : 255 - 0xff -- Sprite 0x62
      12'h311: dout  = 8'b11111111; //  785 : 255 - 0xff
      12'h312: dout  = 8'b11111111; //  786 : 255 - 0xff
      12'h313: dout  = 8'b11111111; //  787 : 255 - 0xff
      12'h314: dout  = 8'b01010101; //  788 :  85 - 0x55
      12'h315: dout  = 8'b10101011; //  789 : 171 - 0xab
      12'h316: dout  = 8'b01010101; //  790 :  85 - 0x55
      12'h317: dout  = 8'b11111111; //  791 : 255 - 0xff
      12'h318: dout  = 8'b00000000; //  792 :   0 - 0x0 -- Sprite 0x63
      12'h319: dout  = 8'b00000000; //  793 :   0 - 0x0
      12'h31A: dout  = 8'b00000000; //  794 :   0 - 0x0
      12'h31B: dout  = 8'b00000000; //  795 :   0 - 0x0
      12'h31C: dout  = 8'b00000000; //  796 :   0 - 0x0
      12'h31D: dout  = 8'b00000000; //  797 :   0 - 0x0
      12'h31E: dout  = 8'b00000000; //  798 :   0 - 0x0
      12'h31F: dout  = 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout  = 8'b00000001; //  800 :   1 - 0x1 -- Sprite 0x64
      12'h321: dout  = 8'b00000001; //  801 :   1 - 0x1
      12'h322: dout  = 8'b00000011; //  802 :   3 - 0x3
      12'h323: dout  = 8'b00000011; //  803 :   3 - 0x3
      12'h324: dout  = 8'b00000110; //  804 :   6 - 0x6
      12'h325: dout  = 8'b00000110; //  805 :   6 - 0x6
      12'h326: dout  = 8'b00001100; //  806 :  12 - 0xc
      12'h327: dout  = 8'b00001100; //  807 :  12 - 0xc
      12'h328: dout  = 8'b00011000; //  808 :  24 - 0x18 -- Sprite 0x65
      12'h329: dout  = 8'b00011000; //  809 :  24 - 0x18
      12'h32A: dout  = 8'b00110000; //  810 :  48 - 0x30
      12'h32B: dout  = 8'b00110000; //  811 :  48 - 0x30
      12'h32C: dout  = 8'b01100000; //  812 :  96 - 0x60
      12'h32D: dout  = 8'b01100000; //  813 :  96 - 0x60
      12'h32E: dout  = 8'b11101010; //  814 : 234 - 0xea
      12'h32F: dout  = 8'b11111111; //  815 : 255 - 0xff
      12'h330: dout  = 8'b10000000; //  816 : 128 - 0x80 -- Sprite 0x66
      12'h331: dout  = 8'b10000000; //  817 : 128 - 0x80
      12'h332: dout  = 8'b11000000; //  818 : 192 - 0xc0
      12'h333: dout  = 8'b01000000; //  819 :  64 - 0x40
      12'h334: dout  = 8'b10100000; //  820 : 160 - 0xa0
      12'h335: dout  = 8'b01100000; //  821 :  96 - 0x60
      12'h336: dout  = 8'b00110000; //  822 :  48 - 0x30
      12'h337: dout  = 8'b00010000; //  823 :  16 - 0x10
      12'h338: dout  = 8'b00101000; //  824 :  40 - 0x28 -- Sprite 0x67
      12'h339: dout  = 8'b00011000; //  825 :  24 - 0x18
      12'h33A: dout  = 8'b00001100; //  826 :  12 - 0xc
      12'h33B: dout  = 8'b00010100; //  827 :  20 - 0x14
      12'h33C: dout  = 8'b00001010; //  828 :  10 - 0xa
      12'h33D: dout  = 8'b00000110; //  829 :   6 - 0x6
      12'h33E: dout  = 8'b10101011; //  830 : 171 - 0xab
      12'h33F: dout  = 8'b11111111; //  831 : 255 - 0xff
      12'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      12'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      12'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      12'h344: dout  = 8'b00000000; //  836 :   0 - 0x0
      12'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout  = 8'b00000000; //  838 :   0 - 0x0
      12'h347: dout  = 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout  = 8'b00000000; //  840 :   0 - 0x0 -- Sprite 0x69
      12'h349: dout  = 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout  = 8'b00000000; //  842 :   0 - 0x0
      12'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout  = 8'b00000000; //  844 :   0 - 0x0
      12'h34D: dout  = 8'b00000000; //  845 :   0 - 0x0
      12'h34E: dout  = 8'b00000000; //  846 :   0 - 0x0
      12'h34F: dout  = 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout  = 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      12'h351: dout  = 8'b00000000; //  849 :   0 - 0x0
      12'h352: dout  = 8'b00000000; //  850 :   0 - 0x0
      12'h353: dout  = 8'b00000000; //  851 :   0 - 0x0
      12'h354: dout  = 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout  = 8'b00000000; //  853 :   0 - 0x0
      12'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout  = 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout  = 8'b00000000; //  856 :   0 - 0x0 -- Sprite 0x6b
      12'h359: dout  = 8'b00000000; //  857 :   0 - 0x0
      12'h35A: dout  = 8'b00000000; //  858 :   0 - 0x0
      12'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout  = 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout  = 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x6c
      12'h361: dout  = 8'b00000000; //  865 :   0 - 0x0
      12'h362: dout  = 8'b00000000; //  866 :   0 - 0x0
      12'h363: dout  = 8'b00000000; //  867 :   0 - 0x0
      12'h364: dout  = 8'b00000000; //  868 :   0 - 0x0
      12'h365: dout  = 8'b00000000; //  869 :   0 - 0x0
      12'h366: dout  = 8'b00000000; //  870 :   0 - 0x0
      12'h367: dout  = 8'b00000000; //  871 :   0 - 0x0
      12'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      12'h369: dout  = 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout  = 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout  = 8'b00000000; //  875 :   0 - 0x0
      12'h36C: dout  = 8'b00000000; //  876 :   0 - 0x0
      12'h36D: dout  = 8'b00000000; //  877 :   0 - 0x0
      12'h36E: dout  = 8'b00000000; //  878 :   0 - 0x0
      12'h36F: dout  = 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      12'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout  = 8'b00000000; //  882 :   0 - 0x0
      12'h373: dout  = 8'b00000000; //  883 :   0 - 0x0
      12'h374: dout  = 8'b00000000; //  884 :   0 - 0x0
      12'h375: dout  = 8'b00000000; //  885 :   0 - 0x0
      12'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout  = 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout  = 8'b00000000; //  888 :   0 - 0x0 -- Sprite 0x6f
      12'h379: dout  = 8'b00000000; //  889 :   0 - 0x0
      12'h37A: dout  = 8'b00000000; //  890 :   0 - 0x0
      12'h37B: dout  = 8'b00000000; //  891 :   0 - 0x0
      12'h37C: dout  = 8'b00000000; //  892 :   0 - 0x0
      12'h37D: dout  = 8'b00000000; //  893 :   0 - 0x0
      12'h37E: dout  = 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout  = 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x70
      12'h381: dout  = 8'b00000000; //  897 :   0 - 0x0
      12'h382: dout  = 8'b00000000; //  898 :   0 - 0x0
      12'h383: dout  = 8'b00000000; //  899 :   0 - 0x0
      12'h384: dout  = 8'b00000000; //  900 :   0 - 0x0
      12'h385: dout  = 8'b00000000; //  901 :   0 - 0x0
      12'h386: dout  = 8'b00000000; //  902 :   0 - 0x0
      12'h387: dout  = 8'b00000000; //  903 :   0 - 0x0
      12'h388: dout  = 8'b00000000; //  904 :   0 - 0x0 -- Sprite 0x71
      12'h389: dout  = 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout  = 8'b00000000; //  906 :   0 - 0x0
      12'h38B: dout  = 8'b00000000; //  907 :   0 - 0x0
      12'h38C: dout  = 8'b00000000; //  908 :   0 - 0x0
      12'h38D: dout  = 8'b00000000; //  909 :   0 - 0x0
      12'h38E: dout  = 8'b00000000; //  910 :   0 - 0x0
      12'h38F: dout  = 8'b00000000; //  911 :   0 - 0x0
      12'h390: dout  = 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x72
      12'h391: dout  = 8'b00000000; //  913 :   0 - 0x0
      12'h392: dout  = 8'b00000000; //  914 :   0 - 0x0
      12'h393: dout  = 8'b00000000; //  915 :   0 - 0x0
      12'h394: dout  = 8'b00000000; //  916 :   0 - 0x0
      12'h395: dout  = 8'b00000000; //  917 :   0 - 0x0
      12'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      12'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout  = 8'b00000000; //  920 :   0 - 0x0 -- Sprite 0x73
      12'h399: dout  = 8'b00000000; //  921 :   0 - 0x0
      12'h39A: dout  = 8'b00000000; //  922 :   0 - 0x0
      12'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      12'h39C: dout  = 8'b00000000; //  924 :   0 - 0x0
      12'h39D: dout  = 8'b00000000; //  925 :   0 - 0x0
      12'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x74
      12'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout  = 8'b00000000; //  930 :   0 - 0x0
      12'h3A3: dout  = 8'b00000000; //  931 :   0 - 0x0
      12'h3A4: dout  = 8'b00000000; //  932 :   0 - 0x0
      12'h3A5: dout  = 8'b00000000; //  933 :   0 - 0x0
      12'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0 -- Sprite 0x75
      12'h3A9: dout  = 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout  = 8'b00000000; //  938 :   0 - 0x0
      12'h3AB: dout  = 8'b00000000; //  939 :   0 - 0x0
      12'h3AC: dout  = 8'b00000000; //  940 :   0 - 0x0
      12'h3AD: dout  = 8'b00000000; //  941 :   0 - 0x0
      12'h3AE: dout  = 8'b00000000; //  942 :   0 - 0x0
      12'h3AF: dout  = 8'b00000000; //  943 :   0 - 0x0
      12'h3B0: dout  = 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x76
      12'h3B1: dout  = 8'b00000000; //  945 :   0 - 0x0
      12'h3B2: dout  = 8'b00000000; //  946 :   0 - 0x0
      12'h3B3: dout  = 8'b00000000; //  947 :   0 - 0x0
      12'h3B4: dout  = 8'b00000000; //  948 :   0 - 0x0
      12'h3B5: dout  = 8'b00000000; //  949 :   0 - 0x0
      12'h3B6: dout  = 8'b00000000; //  950 :   0 - 0x0
      12'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0 -- Sprite 0x77
      12'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      12'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout  = 8'b00000000; //  956 :   0 - 0x0
      12'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout  = 8'b00000000; //  958 :   0 - 0x0
      12'h3BF: dout  = 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x78
      12'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      12'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      12'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      12'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0 -- Sprite 0x79
      12'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x7a
      12'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      12'h3D5: dout  = 8'b00000000; //  981 :   0 - 0x0
      12'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0 -- Sprite 0x7b
      12'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      12'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      12'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      12'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      12'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      12'h3E4: dout  = 8'b00000000; //  996 :   0 - 0x0
      12'h3E5: dout  = 8'b00000000; //  997 :   0 - 0x0
      12'h3E6: dout  = 8'b00000000; //  998 :   0 - 0x0
      12'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      12'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- Sprite 0x7d
      12'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      12'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      12'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      12'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      12'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      12'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x7e
      12'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      12'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0 -- Sprite 0x7f
      12'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      12'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      12'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      12'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      12'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      12'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      12'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout  = 8'b00000011; // 1024 :   3 - 0x3 -- Sprite 0x80
      12'h401: dout  = 8'b00001111; // 1025 :  15 - 0xf
      12'h402: dout  = 8'b00011100; // 1026 :  28 - 0x1c
      12'h403: dout  = 8'b00110000; // 1027 :  48 - 0x30
      12'h404: dout  = 8'b00100000; // 1028 :  32 - 0x20
      12'h405: dout  = 8'b01000000; // 1029 :  64 - 0x40
      12'h406: dout  = 8'b01000000; // 1030 :  64 - 0x40
      12'h407: dout  = 8'b01111111; // 1031 : 127 - 0x7f
      12'h408: dout  = 8'b00000001; // 1032 :   1 - 0x1 -- Sprite 0x81
      12'h409: dout  = 8'b00000001; // 1033 :   1 - 0x1
      12'h40A: dout  = 8'b00000001; // 1034 :   1 - 0x1
      12'h40B: dout  = 8'b00000001; // 1035 :   1 - 0x1
      12'h40C: dout  = 8'b00000001; // 1036 :   1 - 0x1
      12'h40D: dout  = 8'b00000001; // 1037 :   1 - 0x1
      12'h40E: dout  = 8'b00000011; // 1038 :   3 - 0x3
      12'h40F: dout  = 8'b00000011; // 1039 :   3 - 0x3
      12'h410: dout  = 8'b11000000; // 1040 : 192 - 0xc0 -- Sprite 0x82
      12'h411: dout  = 8'b11110000; // 1041 : 240 - 0xf0
      12'h412: dout  = 8'b00111000; // 1042 :  56 - 0x38
      12'h413: dout  = 8'b00001110; // 1043 :  14 - 0xe
      12'h414: dout  = 8'b00011110; // 1044 :  30 - 0x1e
      12'h415: dout  = 8'b00011110; // 1045 :  30 - 0x1e
      12'h416: dout  = 8'b00000010; // 1046 :   2 - 0x2
      12'h417: dout  = 8'b11111110; // 1047 : 254 - 0xfe
      12'h418: dout  = 8'b10000000; // 1048 : 128 - 0x80 -- Sprite 0x83
      12'h419: dout  = 8'b10000000; // 1049 : 128 - 0x80
      12'h41A: dout  = 8'b10000000; // 1050 : 128 - 0x80
      12'h41B: dout  = 8'b10000000; // 1051 : 128 - 0x80
      12'h41C: dout  = 8'b10000000; // 1052 : 128 - 0x80
      12'h41D: dout  = 8'b11100000; // 1053 : 224 - 0xe0
      12'h41E: dout  = 8'b00010000; // 1054 :  16 - 0x10
      12'h41F: dout  = 8'b11110000; // 1055 : 240 - 0xf0
      12'h420: dout  = 8'b00000011; // 1056 :   3 - 0x3 -- Sprite 0x84
      12'h421: dout  = 8'b00001111; // 1057 :  15 - 0xf
      12'h422: dout  = 8'b00011100; // 1058 :  28 - 0x1c
      12'h423: dout  = 8'b00110000; // 1059 :  48 - 0x30
      12'h424: dout  = 8'b00100000; // 1060 :  32 - 0x20
      12'h425: dout  = 8'b01000000; // 1061 :  64 - 0x40
      12'h426: dout  = 8'b01000000; // 1062 :  64 - 0x40
      12'h427: dout  = 8'b01111111; // 1063 : 127 - 0x7f
      12'h428: dout  = 8'b00000011; // 1064 :   3 - 0x3 -- Sprite 0x85
      12'h429: dout  = 8'b00000110; // 1065 :   6 - 0x6
      12'h42A: dout  = 8'b00000110; // 1066 :   6 - 0x6
      12'h42B: dout  = 8'b00011100; // 1067 :  28 - 0x1c
      12'h42C: dout  = 8'b00011000; // 1068 :  24 - 0x18
      12'h42D: dout  = 8'b00110110; // 1069 :  54 - 0x36
      12'h42E: dout  = 8'b00110001; // 1070 :  49 - 0x31
      12'h42F: dout  = 8'b00001111; // 1071 :  15 - 0xf
      12'h430: dout  = 8'b11000000; // 1072 : 192 - 0xc0 -- Sprite 0x86
      12'h431: dout  = 8'b11110000; // 1073 : 240 - 0xf0
      12'h432: dout  = 8'b00111000; // 1074 :  56 - 0x38
      12'h433: dout  = 8'b00001110; // 1075 :  14 - 0xe
      12'h434: dout  = 8'b00011110; // 1076 :  30 - 0x1e
      12'h435: dout  = 8'b00011110; // 1077 :  30 - 0x1e
      12'h436: dout  = 8'b00000010; // 1078 :   2 - 0x2
      12'h437: dout  = 8'b11111110; // 1079 : 254 - 0xfe
      12'h438: dout  = 8'b11000000; // 1080 : 192 - 0xc0 -- Sprite 0x87
      12'h439: dout  = 8'b01100000; // 1081 :  96 - 0x60
      12'h43A: dout  = 8'b01100000; // 1082 :  96 - 0x60
      12'h43B: dout  = 8'b00110000; // 1083 :  48 - 0x30
      12'h43C: dout  = 8'b00111110; // 1084 :  62 - 0x3e
      12'h43D: dout  = 8'b00011001; // 1085 :  25 - 0x19
      12'h43E: dout  = 8'b00110011; // 1086 :  51 - 0x33
      12'h43F: dout  = 8'b00111100; // 1087 :  60 - 0x3c
      12'h440: dout  = 8'b00000011; // 1088 :   3 - 0x3 -- Sprite 0x88
      12'h441: dout  = 8'b00000111; // 1089 :   7 - 0x7
      12'h442: dout  = 8'b00000111; // 1090 :   7 - 0x7
      12'h443: dout  = 8'b00001011; // 1091 :  11 - 0xb
      12'h444: dout  = 8'b00010000; // 1092 :  16 - 0x10
      12'h445: dout  = 8'b01100000; // 1093 :  96 - 0x60
      12'h446: dout  = 8'b11110000; // 1094 : 240 - 0xf0
      12'h447: dout  = 8'b11110000; // 1095 : 240 - 0xf0
      12'h448: dout  = 8'b11110000; // 1096 : 240 - 0xf0 -- Sprite 0x89
      12'h449: dout  = 8'b11110000; // 1097 : 240 - 0xf0
      12'h44A: dout  = 8'b01100000; // 1098 :  96 - 0x60
      12'h44B: dout  = 8'b00010000; // 1099 :  16 - 0x10
      12'h44C: dout  = 8'b00001011; // 1100 :  11 - 0xb
      12'h44D: dout  = 8'b00000111; // 1101 :   7 - 0x7
      12'h44E: dout  = 8'b00000111; // 1102 :   7 - 0x7
      12'h44F: dout  = 8'b00000011; // 1103 :   3 - 0x3
      12'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x8a
      12'h451: dout  = 8'b00011100; // 1105 :  28 - 0x1c
      12'h452: dout  = 8'b00111111; // 1106 :  63 - 0x3f
      12'h453: dout  = 8'b01111000; // 1107 : 120 - 0x78
      12'h454: dout  = 8'b01110000; // 1108 : 112 - 0x70
      12'h455: dout  = 8'b01100000; // 1109 :  96 - 0x60
      12'h456: dout  = 8'b00100000; // 1110 :  32 - 0x20
      12'h457: dout  = 8'b00100000; // 1111 :  32 - 0x20
      12'h458: dout  = 8'b00100000; // 1112 :  32 - 0x20 -- Sprite 0x8b
      12'h459: dout  = 8'b00100000; // 1113 :  32 - 0x20
      12'h45A: dout  = 8'b01100000; // 1114 :  96 - 0x60
      12'h45B: dout  = 8'b01110000; // 1115 : 112 - 0x70
      12'h45C: dout  = 8'b01111000; // 1116 : 120 - 0x78
      12'h45D: dout  = 8'b00111111; // 1117 :  63 - 0x3f
      12'h45E: dout  = 8'b00011100; // 1118 :  28 - 0x1c
      12'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout  = 8'b00000011; // 1120 :   3 - 0x3 -- Sprite 0x8c
      12'h461: dout  = 8'b00001100; // 1121 :  12 - 0xc
      12'h462: dout  = 8'b00011110; // 1122 :  30 - 0x1e
      12'h463: dout  = 8'b00100110; // 1123 :  38 - 0x26
      12'h464: dout  = 8'b01000110; // 1124 :  70 - 0x46
      12'h465: dout  = 8'b01100100; // 1125 : 100 - 0x64
      12'h466: dout  = 8'b01110000; // 1126 : 112 - 0x70
      12'h467: dout  = 8'b11110000; // 1127 : 240 - 0xf0
      12'h468: dout  = 8'b10101010; // 1128 : 170 - 0xaa -- Sprite 0x8d
      12'h469: dout  = 8'b11111111; // 1129 : 255 - 0xff
      12'h46A: dout  = 8'b01111111; // 1130 : 127 - 0x7f
      12'h46B: dout  = 8'b00111001; // 1131 :  57 - 0x39
      12'h46C: dout  = 8'b00011001; // 1132 :  25 - 0x19
      12'h46D: dout  = 8'b00001011; // 1133 :  11 - 0xb
      12'h46E: dout  = 8'b00001000; // 1134 :   8 - 0x8
      12'h46F: dout  = 8'b00000111; // 1135 :   7 - 0x7
      12'h470: dout  = 8'b11000000; // 1136 : 192 - 0xc0 -- Sprite 0x8e
      12'h471: dout  = 8'b00110000; // 1137 :  48 - 0x30
      12'h472: dout  = 8'b00001000; // 1138 :   8 - 0x8
      12'h473: dout  = 8'b01000100; // 1139 :  68 - 0x44
      12'h474: dout  = 8'b01100010; // 1140 :  98 - 0x62
      12'h475: dout  = 8'b01100010; // 1141 :  98 - 0x62
      12'h476: dout  = 8'b00000001; // 1142 :   1 - 0x1
      12'h477: dout  = 8'b00111111; // 1143 :  63 - 0x3f
      12'h478: dout  = 8'b10001011; // 1144 : 139 - 0x8b -- Sprite 0x8f
      12'h479: dout  = 8'b11000001; // 1145 : 193 - 0xc1
      12'h47A: dout  = 8'b11111110; // 1146 : 254 - 0xfe
      12'h47B: dout  = 8'b11111100; // 1147 : 252 - 0xfc
      12'h47C: dout  = 8'b11110000; // 1148 : 240 - 0xf0
      12'h47D: dout  = 8'b11110000; // 1149 : 240 - 0xf0
      12'h47E: dout  = 8'b11111000; // 1150 : 248 - 0xf8
      12'h47F: dout  = 8'b11110000; // 1151 : 240 - 0xf0
      12'h480: dout  = 8'b00000011; // 1152 :   3 - 0x3 -- Sprite 0x90
      12'h481: dout  = 8'b00001110; // 1153 :  14 - 0xe
      12'h482: dout  = 8'b00010110; // 1154 :  22 - 0x16
      12'h483: dout  = 8'b00100110; // 1155 :  38 - 0x26
      12'h484: dout  = 8'b01100011; // 1156 :  99 - 0x63
      12'h485: dout  = 8'b01110010; // 1157 : 114 - 0x72
      12'h486: dout  = 8'b01110000; // 1158 : 112 - 0x70
      12'h487: dout  = 8'b11010000; // 1159 : 208 - 0xd0
      12'h488: dout  = 8'b10101010; // 1160 : 170 - 0xaa -- Sprite 0x91
      12'h489: dout  = 8'b11111111; // 1161 : 255 - 0xff
      12'h48A: dout  = 8'b01111111; // 1162 : 127 - 0x7f
      12'h48B: dout  = 8'b00111100; // 1163 :  60 - 0x3c
      12'h48C: dout  = 8'b00011100; // 1164 :  28 - 0x1c
      12'h48D: dout  = 8'b00000100; // 1165 :   4 - 0x4
      12'h48E: dout  = 8'b00000010; // 1166 :   2 - 0x2
      12'h48F: dout  = 8'b00000001; // 1167 :   1 - 0x1
      12'h490: dout  = 8'b11000000; // 1168 : 192 - 0xc0 -- Sprite 0x92
      12'h491: dout  = 8'b00110000; // 1169 :  48 - 0x30
      12'h492: dout  = 8'b00001000; // 1170 :   8 - 0x8
      12'h493: dout  = 8'b00100100; // 1171 :  36 - 0x24
      12'h494: dout  = 8'b00110010; // 1172 :  50 - 0x32
      12'h495: dout  = 8'b00110010; // 1173 :  50 - 0x32
      12'h496: dout  = 8'b00000001; // 1174 :   1 - 0x1
      12'h497: dout  = 8'b00011111; // 1175 :  31 - 0x1f
      12'h498: dout  = 8'b10001011; // 1176 : 139 - 0x8b -- Sprite 0x93
      12'h499: dout  = 8'b11000001; // 1177 : 193 - 0xc1
      12'h49A: dout  = 8'b11111110; // 1178 : 254 - 0xfe
      12'h49B: dout  = 8'b11111100; // 1179 : 252 - 0xfc
      12'h49C: dout  = 8'b11110000; // 1180 : 240 - 0xf0
      12'h49D: dout  = 8'b11000000; // 1181 : 192 - 0xc0
      12'h49E: dout  = 8'b00100000; // 1182 :  32 - 0x20
      12'h49F: dout  = 8'b11100000; // 1183 : 224 - 0xe0
      12'h4A0: dout  = 8'b00000011; // 1184 :   3 - 0x3 -- Sprite 0x94
      12'h4A1: dout  = 8'b00001111; // 1185 :  15 - 0xf
      12'h4A2: dout  = 8'b00010011; // 1186 :  19 - 0x13
      12'h4A3: dout  = 8'b00110001; // 1187 :  49 - 0x31
      12'h4A4: dout  = 8'b01111001; // 1188 : 121 - 0x79
      12'h4A5: dout  = 8'b01011001; // 1189 :  89 - 0x59
      12'h4A6: dout  = 8'b01001000; // 1190 :  72 - 0x48
      12'h4A7: dout  = 8'b11001100; // 1191 : 204 - 0xcc
      12'h4A8: dout  = 8'b10010101; // 1192 : 149 - 0x95 -- Sprite 0x95
      12'h4A9: dout  = 8'b11111111; // 1193 : 255 - 0xff
      12'h4AA: dout  = 8'b01111111; // 1194 : 127 - 0x7f
      12'h4AB: dout  = 8'b00111110; // 1195 :  62 - 0x3e
      12'h4AC: dout  = 8'b00011111; // 1196 :  31 - 0x1f
      12'h4AD: dout  = 8'b00001111; // 1197 :  15 - 0xf
      12'h4AE: dout  = 8'b00001111; // 1198 :  15 - 0xf
      12'h4AF: dout  = 8'b00000111; // 1199 :   7 - 0x7
      12'h4B0: dout  = 8'b11000000; // 1200 : 192 - 0xc0 -- Sprite 0x96
      12'h4B1: dout  = 8'b00110000; // 1201 :  48 - 0x30
      12'h4B2: dout  = 8'b00001000; // 1202 :   8 - 0x8
      12'h4B3: dout  = 8'b10010100; // 1203 : 148 - 0x94
      12'h4B4: dout  = 8'b10011010; // 1204 : 154 - 0x9a
      12'h4B5: dout  = 8'b00011010; // 1205 :  26 - 0x1a
      12'h4B6: dout  = 8'b00000001; // 1206 :   1 - 0x1
      12'h4B7: dout  = 8'b00001111; // 1207 :  15 - 0xf
      12'h4B8: dout  = 8'b01000101; // 1208 :  69 - 0x45 -- Sprite 0x97
      12'h4B9: dout  = 8'b11100001; // 1209 : 225 - 0xe1
      12'h4BA: dout  = 8'b11111110; // 1210 : 254 - 0xfe
      12'h4BB: dout  = 8'b01111100; // 1211 : 124 - 0x7c
      12'h4BC: dout  = 8'b00110000; // 1212 :  48 - 0x30
      12'h4BD: dout  = 8'b00110000; // 1213 :  48 - 0x30
      12'h4BE: dout  = 8'b10001000; // 1214 : 136 - 0x88
      12'h4BF: dout  = 8'b01111000; // 1215 : 120 - 0x78
      12'h4C0: dout  = 8'b00000001; // 1216 :   1 - 0x1 -- Sprite 0x98
      12'h4C1: dout  = 8'b00000000; // 1217 :   0 - 0x0
      12'h4C2: dout  = 8'b00000000; // 1218 :   0 - 0x0
      12'h4C3: dout  = 8'b00000000; // 1219 :   0 - 0x0
      12'h4C4: dout  = 8'b00000001; // 1220 :   1 - 0x1
      12'h4C5: dout  = 8'b00000001; // 1221 :   1 - 0x1
      12'h4C6: dout  = 8'b00000010; // 1222 :   2 - 0x2
      12'h4C7: dout  = 8'b00000110; // 1223 :   6 - 0x6
      12'h4C8: dout  = 8'b01111000; // 1224 : 120 - 0x78 -- Sprite 0x99
      12'h4C9: dout  = 8'b00101010; // 1225 :  42 - 0x2a
      12'h4CA: dout  = 8'b01010100; // 1226 :  84 - 0x54
      12'h4CB: dout  = 8'b00101001; // 1227 :  41 - 0x29
      12'h4CC: dout  = 8'b00101111; // 1228 :  47 - 0x2f
      12'h4CD: dout  = 8'b00110111; // 1229 :  55 - 0x37
      12'h4CE: dout  = 8'b00000011; // 1230 :   3 - 0x3
      12'h4CF: dout  = 8'b00000111; // 1231 :   7 - 0x7
      12'h4D0: dout  = 8'b10110000; // 1232 : 176 - 0xb0 -- Sprite 0x9a
      12'h4D1: dout  = 8'b11101000; // 1233 : 232 - 0xe8
      12'h4D2: dout  = 8'b10001100; // 1234 : 140 - 0x8c
      12'h4D3: dout  = 8'b10011110; // 1235 : 158 - 0x9e
      12'h4D4: dout  = 8'b00011111; // 1236 :  31 - 0x1f
      12'h4D5: dout  = 8'b00001111; // 1237 :  15 - 0xf
      12'h4D6: dout  = 8'b10010110; // 1238 : 150 - 0x96
      12'h4D7: dout  = 8'b00011100; // 1239 :  28 - 0x1c
      12'h4D8: dout  = 8'b00001100; // 1240 :  12 - 0xc -- Sprite 0x9b
      12'h4D9: dout  = 8'b00111000; // 1241 :  56 - 0x38
      12'h4DA: dout  = 8'b11101000; // 1242 : 232 - 0xe8
      12'h4DB: dout  = 8'b11010000; // 1243 : 208 - 0xd0
      12'h4DC: dout  = 8'b11100000; // 1244 : 224 - 0xe0
      12'h4DD: dout  = 8'b10000000; // 1245 : 128 - 0x80
      12'h4DE: dout  = 8'b00000000; // 1246 :   0 - 0x0
      12'h4DF: dout  = 8'b10000000; // 1247 : 128 - 0x80
      12'h4E0: dout  = 8'b00000001; // 1248 :   1 - 0x1 -- Sprite 0x9c
      12'h4E1: dout  = 8'b00000000; // 1249 :   0 - 0x0
      12'h4E2: dout  = 8'b00000000; // 1250 :   0 - 0x0
      12'h4E3: dout  = 8'b00000000; // 1251 :   0 - 0x0
      12'h4E4: dout  = 8'b00000001; // 1252 :   1 - 0x1
      12'h4E5: dout  = 8'b00000001; // 1253 :   1 - 0x1
      12'h4E6: dout  = 8'b00000010; // 1254 :   2 - 0x2
      12'h4E7: dout  = 8'b00000110; // 1255 :   6 - 0x6
      12'h4E8: dout  = 8'b01111000; // 1256 : 120 - 0x78 -- Sprite 0x9d
      12'h4E9: dout  = 8'b00101010; // 1257 :  42 - 0x2a
      12'h4EA: dout  = 8'b01010100; // 1258 :  84 - 0x54
      12'h4EB: dout  = 8'b00101001; // 1259 :  41 - 0x29
      12'h4EC: dout  = 8'b00101111; // 1260 :  47 - 0x2f
      12'h4ED: dout  = 8'b00111100; // 1261 :  60 - 0x3c
      12'h4EE: dout  = 8'b00011110; // 1262 :  30 - 0x1e
      12'h4EF: dout  = 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout  = 8'b10110000; // 1264 : 176 - 0xb0 -- Sprite 0x9e
      12'h4F1: dout  = 8'b11101000; // 1265 : 232 - 0xe8
      12'h4F2: dout  = 8'b10001100; // 1266 : 140 - 0x8c
      12'h4F3: dout  = 8'b10011110; // 1267 : 158 - 0x9e
      12'h4F4: dout  = 8'b00011111; // 1268 :  31 - 0x1f
      12'h4F5: dout  = 8'b00001111; // 1269 :  15 - 0xf
      12'h4F6: dout  = 8'b10010110; // 1270 : 150 - 0x96
      12'h4F7: dout  = 8'b00011100; // 1271 :  28 - 0x1c
      12'h4F8: dout  = 8'b00001100; // 1272 :  12 - 0xc -- Sprite 0x9f
      12'h4F9: dout  = 8'b00111000; // 1273 :  56 - 0x38
      12'h4FA: dout  = 8'b11101000; // 1274 : 232 - 0xe8
      12'h4FB: dout  = 8'b11110000; // 1275 : 240 - 0xf0
      12'h4FC: dout  = 8'b11000000; // 1276 : 192 - 0xc0
      12'h4FD: dout  = 8'b01110000; // 1277 : 112 - 0x70
      12'h4FE: dout  = 8'b11000000; // 1278 : 192 - 0xc0
      12'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout  = 8'b00000011; // 1280 :   3 - 0x3 -- Sprite 0xa0
      12'h501: dout  = 8'b00001111; // 1281 :  15 - 0xf
      12'h502: dout  = 8'b00011100; // 1282 :  28 - 0x1c
      12'h503: dout  = 8'b00110000; // 1283 :  48 - 0x30
      12'h504: dout  = 8'b01100000; // 1284 :  96 - 0x60
      12'h505: dout  = 8'b01100000; // 1285 :  96 - 0x60
      12'h506: dout  = 8'b11000000; // 1286 : 192 - 0xc0
      12'h507: dout  = 8'b11000000; // 1287 : 192 - 0xc0
      12'h508: dout  = 8'b11000000; // 1288 : 192 - 0xc0 -- Sprite 0xa1
      12'h509: dout  = 8'b11000000; // 1289 : 192 - 0xc0
      12'h50A: dout  = 8'b01100000; // 1290 :  96 - 0x60
      12'h50B: dout  = 8'b01100000; // 1291 :  96 - 0x60
      12'h50C: dout  = 8'b00110000; // 1292 :  48 - 0x30
      12'h50D: dout  = 8'b00011010; // 1293 :  26 - 0x1a
      12'h50E: dout  = 8'b00001101; // 1294 :  13 - 0xd
      12'h50F: dout  = 8'b00000011; // 1295 :   3 - 0x3
      12'h510: dout  = 8'b11000000; // 1296 : 192 - 0xc0 -- Sprite 0xa2
      12'h511: dout  = 8'b11110000; // 1297 : 240 - 0xf0
      12'h512: dout  = 8'b00111000; // 1298 :  56 - 0x38
      12'h513: dout  = 8'b00001100; // 1299 :  12 - 0xc
      12'h514: dout  = 8'b00000110; // 1300 :   6 - 0x6
      12'h515: dout  = 8'b00000010; // 1301 :   2 - 0x2
      12'h516: dout  = 8'b00000101; // 1302 :   5 - 0x5
      12'h517: dout  = 8'b00000011; // 1303 :   3 - 0x3
      12'h518: dout  = 8'b00000101; // 1304 :   5 - 0x5 -- Sprite 0xa3
      12'h519: dout  = 8'b00001011; // 1305 :  11 - 0xb
      12'h51A: dout  = 8'b00010110; // 1306 :  22 - 0x16
      12'h51B: dout  = 8'b00101010; // 1307 :  42 - 0x2a
      12'h51C: dout  = 8'b01010100; // 1308 :  84 - 0x54
      12'h51D: dout  = 8'b10101000; // 1309 : 168 - 0xa8
      12'h51E: dout  = 8'b01110000; // 1310 : 112 - 0x70
      12'h51F: dout  = 8'b11000000; // 1311 : 192 - 0xc0
      12'h520: dout  = 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0xa4
      12'h521: dout  = 8'b00001111; // 1313 :  15 - 0xf
      12'h522: dout  = 8'b00011111; // 1314 :  31 - 0x1f
      12'h523: dout  = 8'b00110001; // 1315 :  49 - 0x31
      12'h524: dout  = 8'b00111111; // 1316 :  63 - 0x3f
      12'h525: dout  = 8'b01111111; // 1317 : 127 - 0x7f
      12'h526: dout  = 8'b11111111; // 1318 : 255 - 0xff
      12'h527: dout  = 8'b11011111; // 1319 : 223 - 0xdf
      12'h528: dout  = 8'b11000000; // 1320 : 192 - 0xc0 -- Sprite 0xa5
      12'h529: dout  = 8'b11000111; // 1321 : 199 - 0xc7
      12'h52A: dout  = 8'b01101111; // 1322 : 111 - 0x6f
      12'h52B: dout  = 8'b01100111; // 1323 : 103 - 0x67
      12'h52C: dout  = 8'b01100011; // 1324 :  99 - 0x63
      12'h52D: dout  = 8'b00110000; // 1325 :  48 - 0x30
      12'h52E: dout  = 8'b00011000; // 1326 :  24 - 0x18
      12'h52F: dout  = 8'b00000111; // 1327 :   7 - 0x7
      12'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0xa6
      12'h531: dout  = 8'b11110000; // 1329 : 240 - 0xf0
      12'h532: dout  = 8'b11111000; // 1330 : 248 - 0xf8
      12'h533: dout  = 8'b10001100; // 1331 : 140 - 0x8c
      12'h534: dout  = 8'b11111100; // 1332 : 252 - 0xfc
      12'h535: dout  = 8'b11111110; // 1333 : 254 - 0xfe
      12'h536: dout  = 8'b11111101; // 1334 : 253 - 0xfd
      12'h537: dout  = 8'b11111001; // 1335 : 249 - 0xf9
      12'h538: dout  = 8'b00000011; // 1336 :   3 - 0x3 -- Sprite 0xa7
      12'h539: dout  = 8'b11100101; // 1337 : 229 - 0xe5
      12'h53A: dout  = 8'b11110010; // 1338 : 242 - 0xf2
      12'h53B: dout  = 8'b11100110; // 1339 : 230 - 0xe6
      12'h53C: dout  = 8'b11001010; // 1340 : 202 - 0xca
      12'h53D: dout  = 8'b00010100; // 1341 :  20 - 0x14
      12'h53E: dout  = 8'b00111000; // 1342 :  56 - 0x38
      12'h53F: dout  = 8'b11100000; // 1343 : 224 - 0xe0
      12'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0xa8
      12'h541: dout  = 8'b00001111; // 1345 :  15 - 0xf
      12'h542: dout  = 8'b00011111; // 1346 :  31 - 0x1f
      12'h543: dout  = 8'b00110001; // 1347 :  49 - 0x31
      12'h544: dout  = 8'b00111111; // 1348 :  63 - 0x3f
      12'h545: dout  = 8'b01111111; // 1349 : 127 - 0x7f
      12'h546: dout  = 8'b11111111; // 1350 : 255 - 0xff
      12'h547: dout  = 8'b11011111; // 1351 : 223 - 0xdf
      12'h548: dout  = 8'b11000000; // 1352 : 192 - 0xc0 -- Sprite 0xa9
      12'h549: dout  = 8'b11000011; // 1353 : 195 - 0xc3
      12'h54A: dout  = 8'b11000111; // 1354 : 199 - 0xc7
      12'h54B: dout  = 8'b11001111; // 1355 : 207 - 0xcf
      12'h54C: dout  = 8'b11000111; // 1356 : 199 - 0xc7
      12'h54D: dout  = 8'b11000000; // 1357 : 192 - 0xc0
      12'h54E: dout  = 8'b11100000; // 1358 : 224 - 0xe0
      12'h54F: dout  = 8'b11111111; // 1359 : 255 - 0xff
      12'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      12'h551: dout  = 8'b11110000; // 1361 : 240 - 0xf0
      12'h552: dout  = 8'b11111000; // 1362 : 248 - 0xf8
      12'h553: dout  = 8'b10001100; // 1363 : 140 - 0x8c
      12'h554: dout  = 8'b11111100; // 1364 : 252 - 0xfc
      12'h555: dout  = 8'b11111110; // 1365 : 254 - 0xfe
      12'h556: dout  = 8'b11111101; // 1366 : 253 - 0xfd
      12'h557: dout  = 8'b11111001; // 1367 : 249 - 0xf9
      12'h558: dout  = 8'b00000011; // 1368 :   3 - 0x3 -- Sprite 0xab
      12'h559: dout  = 8'b11000101; // 1369 : 197 - 0xc5
      12'h55A: dout  = 8'b11100011; // 1370 : 227 - 0xe3
      12'h55B: dout  = 8'b11110101; // 1371 : 245 - 0xf5
      12'h55C: dout  = 8'b11100011; // 1372 : 227 - 0xe3
      12'h55D: dout  = 8'b00000101; // 1373 :   5 - 0x5
      12'h55E: dout  = 8'b00001011; // 1374 :  11 - 0xb
      12'h55F: dout  = 8'b11111111; // 1375 : 255 - 0xff
      12'h560: dout  = 8'b10000011; // 1376 : 131 - 0x83 -- Sprite 0xac
      12'h561: dout  = 8'b10001100; // 1377 : 140 - 0x8c
      12'h562: dout  = 8'b10010000; // 1378 : 144 - 0x90
      12'h563: dout  = 8'b10010000; // 1379 : 144 - 0x90
      12'h564: dout  = 8'b11100000; // 1380 : 224 - 0xe0
      12'h565: dout  = 8'b10100000; // 1381 : 160 - 0xa0
      12'h566: dout  = 8'b10101111; // 1382 : 175 - 0xaf
      12'h567: dout  = 8'b01101111; // 1383 : 111 - 0x6f
      12'h568: dout  = 8'b11111011; // 1384 : 251 - 0xfb -- Sprite 0xad
      12'h569: dout  = 8'b00000101; // 1385 :   5 - 0x5
      12'h56A: dout  = 8'b00000101; // 1386 :   5 - 0x5
      12'h56B: dout  = 8'b00000101; // 1387 :   5 - 0x5
      12'h56C: dout  = 8'b01000101; // 1388 :  69 - 0x45
      12'h56D: dout  = 8'b01100101; // 1389 : 101 - 0x65
      12'h56E: dout  = 8'b11110101; // 1390 : 245 - 0xf5
      12'h56F: dout  = 8'b11111101; // 1391 : 253 - 0xfd
      12'h570: dout  = 8'b10000011; // 1392 : 131 - 0x83 -- Sprite 0xae
      12'h571: dout  = 8'b10001100; // 1393 : 140 - 0x8c
      12'h572: dout  = 8'b10010000; // 1394 : 144 - 0x90
      12'h573: dout  = 8'b10010000; // 1395 : 144 - 0x90
      12'h574: dout  = 8'b11100000; // 1396 : 224 - 0xe0
      12'h575: dout  = 8'b10100000; // 1397 : 160 - 0xa0
      12'h576: dout  = 8'b10101111; // 1398 : 175 - 0xaf
      12'h577: dout  = 8'b01101111; // 1399 : 111 - 0x6f
      12'h578: dout  = 8'b11111011; // 1400 : 251 - 0xfb -- Sprite 0xaf
      12'h579: dout  = 8'b00000101; // 1401 :   5 - 0x5
      12'h57A: dout  = 8'b00000101; // 1402 :   5 - 0x5
      12'h57B: dout  = 8'b00000101; // 1403 :   5 - 0x5
      12'h57C: dout  = 8'b11000101; // 1404 : 197 - 0xc5
      12'h57D: dout  = 8'b11100101; // 1405 : 229 - 0xe5
      12'h57E: dout  = 8'b11110101; // 1406 : 245 - 0xf5
      12'h57F: dout  = 8'b11111101; // 1407 : 253 - 0xfd
      12'h580: dout  = 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      12'h581: dout  = 8'b00000011; // 1409 :   3 - 0x3
      12'h582: dout  = 8'b00001111; // 1410 :  15 - 0xf
      12'h583: dout  = 8'b00111111; // 1411 :  63 - 0x3f
      12'h584: dout  = 8'b01111111; // 1412 : 127 - 0x7f
      12'h585: dout  = 8'b01111111; // 1413 : 127 - 0x7f
      12'h586: dout  = 8'b11111111; // 1414 : 255 - 0xff
      12'h587: dout  = 8'b11111111; // 1415 : 255 - 0xff
      12'h588: dout  = 8'b11111111; // 1416 : 255 - 0xff -- Sprite 0xb1
      12'h589: dout  = 8'b10001111; // 1417 : 143 - 0x8f
      12'h58A: dout  = 8'b10000000; // 1418 : 128 - 0x80
      12'h58B: dout  = 8'b11110000; // 1419 : 240 - 0xf0
      12'h58C: dout  = 8'b11111111; // 1420 : 255 - 0xff
      12'h58D: dout  = 8'b11111111; // 1421 : 255 - 0xff
      12'h58E: dout  = 8'b01111111; // 1422 : 127 - 0x7f
      12'h58F: dout  = 8'b00001111; // 1423 :  15 - 0xf
      12'h590: dout  = 8'b00000000; // 1424 :   0 - 0x0 -- Sprite 0xb2
      12'h591: dout  = 8'b11000000; // 1425 : 192 - 0xc0
      12'h592: dout  = 8'b11110000; // 1426 : 240 - 0xf0
      12'h593: dout  = 8'b11111100; // 1427 : 252 - 0xfc
      12'h594: dout  = 8'b11111110; // 1428 : 254 - 0xfe
      12'h595: dout  = 8'b11111110; // 1429 : 254 - 0xfe
      12'h596: dout  = 8'b11111111; // 1430 : 255 - 0xff
      12'h597: dout  = 8'b11111111; // 1431 : 255 - 0xff
      12'h598: dout  = 8'b11111111; // 1432 : 255 - 0xff -- Sprite 0xb3
      12'h599: dout  = 8'b11110001; // 1433 : 241 - 0xf1
      12'h59A: dout  = 8'b00000001; // 1434 :   1 - 0x1
      12'h59B: dout  = 8'b00001111; // 1435 :  15 - 0xf
      12'h59C: dout  = 8'b11111111; // 1436 : 255 - 0xff
      12'h59D: dout  = 8'b11111111; // 1437 : 255 - 0xff
      12'h59E: dout  = 8'b11111110; // 1438 : 254 - 0xfe
      12'h59F: dout  = 8'b11110000; // 1439 : 240 - 0xf0
      12'h5A0: dout  = 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0xb4
      12'h5A1: dout  = 8'b00000011; // 1441 :   3 - 0x3
      12'h5A2: dout  = 8'b00001110; // 1442 :  14 - 0xe
      12'h5A3: dout  = 8'b00110101; // 1443 :  53 - 0x35
      12'h5A4: dout  = 8'b01101110; // 1444 : 110 - 0x6e
      12'h5A5: dout  = 8'b01010101; // 1445 :  85 - 0x55
      12'h5A6: dout  = 8'b10111010; // 1446 : 186 - 0xba
      12'h5A7: dout  = 8'b11010111; // 1447 : 215 - 0xd7
      12'h5A8: dout  = 8'b11111010; // 1448 : 250 - 0xfa -- Sprite 0xb5
      12'h5A9: dout  = 8'b10001111; // 1449 : 143 - 0x8f
      12'h5AA: dout  = 8'b10000000; // 1450 : 128 - 0x80
      12'h5AB: dout  = 8'b11110000; // 1451 : 240 - 0xf0
      12'h5AC: dout  = 8'b10101111; // 1452 : 175 - 0xaf
      12'h5AD: dout  = 8'b11010101; // 1453 : 213 - 0xd5
      12'h5AE: dout  = 8'b01111010; // 1454 : 122 - 0x7a
      12'h5AF: dout  = 8'b00001111; // 1455 :  15 - 0xf
      12'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0xb6
      12'h5B1: dout  = 8'b11000000; // 1457 : 192 - 0xc0
      12'h5B2: dout  = 8'b10110000; // 1458 : 176 - 0xb0
      12'h5B3: dout  = 8'b01011100; // 1459 :  92 - 0x5c
      12'h5B4: dout  = 8'b11101010; // 1460 : 234 - 0xea
      12'h5B5: dout  = 8'b01011110; // 1461 :  94 - 0x5e
      12'h5B6: dout  = 8'b10101011; // 1462 : 171 - 0xab
      12'h5B7: dout  = 8'b01110101; // 1463 : 117 - 0x75
      12'h5B8: dout  = 8'b10101111; // 1464 : 175 - 0xaf -- Sprite 0xb7
      12'h5B9: dout  = 8'b11110001; // 1465 : 241 - 0xf1
      12'h5BA: dout  = 8'b00000001; // 1466 :   1 - 0x1
      12'h5BB: dout  = 8'b00001111; // 1467 :  15 - 0xf
      12'h5BC: dout  = 8'b11111011; // 1468 : 251 - 0xfb
      12'h5BD: dout  = 8'b01010101; // 1469 :  85 - 0x55
      12'h5BE: dout  = 8'b10101110; // 1470 : 174 - 0xae
      12'h5BF: dout  = 8'b11110000; // 1471 : 240 - 0xf0
      12'h5C0: dout  = 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0xb8
      12'h5C1: dout  = 8'b00000011; // 1473 :   3 - 0x3
      12'h5C2: dout  = 8'b00001100; // 1474 :  12 - 0xc
      12'h5C3: dout  = 8'b00110000; // 1475 :  48 - 0x30
      12'h5C4: dout  = 8'b01000100; // 1476 :  68 - 0x44
      12'h5C5: dout  = 8'b01000000; // 1477 :  64 - 0x40
      12'h5C6: dout  = 8'b10010000; // 1478 : 144 - 0x90
      12'h5C7: dout  = 8'b10000010; // 1479 : 130 - 0x82
      12'h5C8: dout  = 8'b11110000; // 1480 : 240 - 0xf0 -- Sprite 0xb9
      12'h5C9: dout  = 8'b11111111; // 1481 : 255 - 0xff
      12'h5CA: dout  = 8'b11111111; // 1482 : 255 - 0xff
      12'h5CB: dout  = 8'b11111111; // 1483 : 255 - 0xff
      12'h5CC: dout  = 8'b10001111; // 1484 : 143 - 0x8f
      12'h5CD: dout  = 8'b10000000; // 1485 : 128 - 0x80
      12'h5CE: dout  = 8'b01110000; // 1486 : 112 - 0x70
      12'h5CF: dout  = 8'b00001111; // 1487 :  15 - 0xf
      12'h5D0: dout  = 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0xba
      12'h5D1: dout  = 8'b11000000; // 1489 : 192 - 0xc0
      12'h5D2: dout  = 8'b00110000; // 1490 :  48 - 0x30
      12'h5D3: dout  = 8'b00001100; // 1491 :  12 - 0xc
      12'h5D4: dout  = 8'b01000010; // 1492 :  66 - 0x42
      12'h5D5: dout  = 8'b00001010; // 1493 :  10 - 0xa
      12'h5D6: dout  = 8'b00000001; // 1494 :   1 - 0x1
      12'h5D7: dout  = 8'b00100001; // 1495 :  33 - 0x21
      12'h5D8: dout  = 8'b00001111; // 1496 :  15 - 0xf -- Sprite 0xbb
      12'h5D9: dout  = 8'b11111111; // 1497 : 255 - 0xff
      12'h5DA: dout  = 8'b11111111; // 1498 : 255 - 0xff
      12'h5DB: dout  = 8'b11111111; // 1499 : 255 - 0xff
      12'h5DC: dout  = 8'b11110001; // 1500 : 241 - 0xf1
      12'h5DD: dout  = 8'b00000001; // 1501 :   1 - 0x1
      12'h5DE: dout  = 8'b00001110; // 1502 :  14 - 0xe
      12'h5DF: dout  = 8'b11110000; // 1503 : 240 - 0xf0
      12'h5E0: dout  = 8'b11110011; // 1504 : 243 - 0xf3 -- Sprite 0xbc
      12'h5E1: dout  = 8'b11111111; // 1505 : 255 - 0xff
      12'h5E2: dout  = 8'b11000100; // 1506 : 196 - 0xc4
      12'h5E3: dout  = 8'b11000000; // 1507 : 192 - 0xc0
      12'h5E4: dout  = 8'b01000000; // 1508 :  64 - 0x40
      12'h5E5: dout  = 8'b01100011; // 1509 :  99 - 0x63
      12'h5E6: dout  = 8'b11000111; // 1510 : 199 - 0xc7
      12'h5E7: dout  = 8'b11000110; // 1511 : 198 - 0xc6
      12'h5E8: dout  = 8'b11000110; // 1512 : 198 - 0xc6 -- Sprite 0xbd
      12'h5E9: dout  = 8'b11000110; // 1513 : 198 - 0xc6
      12'h5EA: dout  = 8'b01100011; // 1514 :  99 - 0x63
      12'h5EB: dout  = 8'b01000000; // 1515 :  64 - 0x40
      12'h5EC: dout  = 8'b11000000; // 1516 : 192 - 0xc0
      12'h5ED: dout  = 8'b11000100; // 1517 : 196 - 0xc4
      12'h5EE: dout  = 8'b11001100; // 1518 : 204 - 0xcc
      12'h5EF: dout  = 8'b11110011; // 1519 : 243 - 0xf3
      12'h5F0: dout  = 8'b11001111; // 1520 : 207 - 0xcf -- Sprite 0xbe
      12'h5F1: dout  = 8'b11111111; // 1521 : 255 - 0xff
      12'h5F2: dout  = 8'b00100001; // 1522 :  33 - 0x21
      12'h5F3: dout  = 8'b00000001; // 1523 :   1 - 0x1
      12'h5F4: dout  = 8'b00000010; // 1524 :   2 - 0x2
      12'h5F5: dout  = 8'b11000110; // 1525 : 198 - 0xc6
      12'h5F6: dout  = 8'b11100001; // 1526 : 225 - 0xe1
      12'h5F7: dout  = 8'b00100001; // 1527 :  33 - 0x21
      12'h5F8: dout  = 8'b00100001; // 1528 :  33 - 0x21 -- Sprite 0xbf
      12'h5F9: dout  = 8'b00100001; // 1529 :  33 - 0x21
      12'h5FA: dout  = 8'b11000110; // 1530 : 198 - 0xc6
      12'h5FB: dout  = 8'b00000010; // 1531 :   2 - 0x2
      12'h5FC: dout  = 8'b00000001; // 1532 :   1 - 0x1
      12'h5FD: dout  = 8'b00100001; // 1533 :  33 - 0x21
      12'h5FE: dout  = 8'b00110001; // 1534 :  49 - 0x31
      12'h5FF: dout  = 8'b11001111; // 1535 : 207 - 0xcf
      12'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      12'h601: dout  = 8'b01010000; // 1537 :  80 - 0x50
      12'h602: dout  = 8'b10110011; // 1538 : 179 - 0xb3
      12'h603: dout  = 8'b10010111; // 1539 : 151 - 0x97
      12'h604: dout  = 8'b10011111; // 1540 : 159 - 0x9f
      12'h605: dout  = 8'b01101111; // 1541 : 111 - 0x6f
      12'h606: dout  = 8'b00011111; // 1542 :  31 - 0x1f
      12'h607: dout  = 8'b00011111; // 1543 :  31 - 0x1f
      12'h608: dout  = 8'b00011111; // 1544 :  31 - 0x1f -- Sprite 0xc1
      12'h609: dout  = 8'b00011111; // 1545 :  31 - 0x1f
      12'h60A: dout  = 8'b00001111; // 1546 :  15 - 0xf
      12'h60B: dout  = 8'b00000111; // 1547 :   7 - 0x7
      12'h60C: dout  = 8'b00011101; // 1548 :  29 - 0x1d
      12'h60D: dout  = 8'b00101100; // 1549 :  44 - 0x2c
      12'h60E: dout  = 8'b01010100; // 1550 :  84 - 0x54
      12'h60F: dout  = 8'b01111100; // 1551 : 124 - 0x7c
      12'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      12'h611: dout  = 8'b00001010; // 1553 :  10 - 0xa
      12'h612: dout  = 8'b11001101; // 1554 : 205 - 0xcd
      12'h613: dout  = 8'b11101001; // 1555 : 233 - 0xe9
      12'h614: dout  = 8'b11111001; // 1556 : 249 - 0xf9
      12'h615: dout  = 8'b11110110; // 1557 : 246 - 0xf6
      12'h616: dout  = 8'b11110000; // 1558 : 240 - 0xf0
      12'h617: dout  = 8'b11111000; // 1559 : 248 - 0xf8
      12'h618: dout  = 8'b11111000; // 1560 : 248 - 0xf8 -- Sprite 0xc3
      12'h619: dout  = 8'b11111000; // 1561 : 248 - 0xf8
      12'h61A: dout  = 8'b11110000; // 1562 : 240 - 0xf0
      12'h61B: dout  = 8'b11000000; // 1563 : 192 - 0xc0
      12'h61C: dout  = 8'b10111000; // 1564 : 184 - 0xb8
      12'h61D: dout  = 8'b00110100; // 1565 :  52 - 0x34
      12'h61E: dout  = 8'b00101010; // 1566 :  42 - 0x2a
      12'h61F: dout  = 8'b00111110; // 1567 :  62 - 0x3e
      12'h620: dout  = 8'b00000101; // 1568 :   5 - 0x5 -- Sprite 0xc4
      12'h621: dout  = 8'b00001010; // 1569 :  10 - 0xa
      12'h622: dout  = 8'b00001000; // 1570 :   8 - 0x8
      12'h623: dout  = 8'b00001111; // 1571 :  15 - 0xf
      12'h624: dout  = 8'b00000001; // 1572 :   1 - 0x1
      12'h625: dout  = 8'b00000011; // 1573 :   3 - 0x3
      12'h626: dout  = 8'b00000111; // 1574 :   7 - 0x7
      12'h627: dout  = 8'b00001111; // 1575 :  15 - 0xf
      12'h628: dout  = 8'b00001111; // 1576 :  15 - 0xf -- Sprite 0xc5
      12'h629: dout  = 8'b11101111; // 1577 : 239 - 0xef
      12'h62A: dout  = 8'b11011111; // 1578 : 223 - 0xdf
      12'h62B: dout  = 8'b10101111; // 1579 : 175 - 0xaf
      12'h62C: dout  = 8'b01100111; // 1580 : 103 - 0x67
      12'h62D: dout  = 8'b00001101; // 1581 :  13 - 0xd
      12'h62E: dout  = 8'b00001010; // 1582 :  10 - 0xa
      12'h62F: dout  = 8'b00000111; // 1583 :   7 - 0x7
      12'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0xc6
      12'h631: dout  = 8'b10000000; // 1585 : 128 - 0x80
      12'h632: dout  = 8'b10000000; // 1586 : 128 - 0x80
      12'h633: dout  = 8'b11110000; // 1587 : 240 - 0xf0
      12'h634: dout  = 8'b11111000; // 1588 : 248 - 0xf8
      12'h635: dout  = 8'b11111100; // 1589 : 252 - 0xfc
      12'h636: dout  = 8'b11111100; // 1590 : 252 - 0xfc
      12'h637: dout  = 8'b11111100; // 1591 : 252 - 0xfc
      12'h638: dout  = 8'b11111100; // 1592 : 252 - 0xfc -- Sprite 0xc7
      12'h639: dout  = 8'b11111110; // 1593 : 254 - 0xfe
      12'h63A: dout  = 8'b11111001; // 1594 : 249 - 0xf9
      12'h63B: dout  = 8'b11111010; // 1595 : 250 - 0xfa
      12'h63C: dout  = 8'b11101001; // 1596 : 233 - 0xe9
      12'h63D: dout  = 8'b00001110; // 1597 :  14 - 0xe
      12'h63E: dout  = 8'b10000000; // 1598 : 128 - 0x80
      12'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout  = 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      12'h641: dout  = 8'b11000000; // 1601 : 192 - 0xc0
      12'h642: dout  = 8'b10100000; // 1602 : 160 - 0xa0
      12'h643: dout  = 8'b11010011; // 1603 : 211 - 0xd3
      12'h644: dout  = 8'b10110111; // 1604 : 183 - 0xb7
      12'h645: dout  = 8'b11111111; // 1605 : 255 - 0xff
      12'h646: dout  = 8'b00001111; // 1606 :  15 - 0xf
      12'h647: dout  = 8'b00011111; // 1607 :  31 - 0x1f
      12'h648: dout  = 8'b00011111; // 1608 :  31 - 0x1f -- Sprite 0xc9
      12'h649: dout  = 8'b00001111; // 1609 :  15 - 0xf
      12'h64A: dout  = 8'b11110111; // 1610 : 247 - 0xf7
      12'h64B: dout  = 8'b10110111; // 1611 : 183 - 0xb7
      12'h64C: dout  = 8'b11010011; // 1612 : 211 - 0xd3
      12'h64D: dout  = 8'b10100000; // 1613 : 160 - 0xa0
      12'h64E: dout  = 8'b11000000; // 1614 : 192 - 0xc0
      12'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout  = 8'b00011100; // 1616 :  28 - 0x1c -- Sprite 0xca
      12'h651: dout  = 8'b00100010; // 1617 :  34 - 0x22
      12'h652: dout  = 8'b00100100; // 1618 :  36 - 0x24
      12'h653: dout  = 8'b11011110; // 1619 : 222 - 0xde
      12'h654: dout  = 8'b11110000; // 1620 : 240 - 0xf0
      12'h655: dout  = 8'b11111000; // 1621 : 248 - 0xf8
      12'h656: dout  = 8'b11111100; // 1622 : 252 - 0xfc
      12'h657: dout  = 8'b11111100; // 1623 : 252 - 0xfc
      12'h658: dout  = 8'b11111100; // 1624 : 252 - 0xfc -- Sprite 0xcb
      12'h659: dout  = 8'b11111100; // 1625 : 252 - 0xfc
      12'h65A: dout  = 8'b11111000; // 1626 : 248 - 0xf8
      12'h65B: dout  = 8'b11110000; // 1627 : 240 - 0xf0
      12'h65C: dout  = 8'b10011110; // 1628 : 158 - 0x9e
      12'h65D: dout  = 8'b00100100; // 1629 :  36 - 0x24
      12'h65E: dout  = 8'b00100010; // 1630 :  34 - 0x22
      12'h65F: dout  = 8'b00011100; // 1631 :  28 - 0x1c
      12'h660: dout  = 8'b00001110; // 1632 :  14 - 0xe -- Sprite 0xcc
      12'h661: dout  = 8'b00010110; // 1633 :  22 - 0x16
      12'h662: dout  = 8'b00011010; // 1634 :  26 - 0x1a
      12'h663: dout  = 8'b00000100; // 1635 :   4 - 0x4
      12'h664: dout  = 8'b01101111; // 1636 : 111 - 0x6f
      12'h665: dout  = 8'b10111111; // 1637 : 191 - 0xbf
      12'h666: dout  = 8'b11011111; // 1638 : 223 - 0xdf
      12'h667: dout  = 8'b10111111; // 1639 : 191 - 0xbf
      12'h668: dout  = 8'b01011111; // 1640 :  95 - 0x5f -- Sprite 0xcd
      12'h669: dout  = 8'b00011111; // 1641 :  31 - 0x1f
      12'h66A: dout  = 8'b00011111; // 1642 :  31 - 0x1f
      12'h66B: dout  = 8'b00001111; // 1643 :  15 - 0xf
      12'h66C: dout  = 8'b00111111; // 1644 :  63 - 0x3f
      12'h66D: dout  = 8'b00100011; // 1645 :  35 - 0x23
      12'h66E: dout  = 8'b00101010; // 1646 :  42 - 0x2a
      12'h66F: dout  = 8'b00010100; // 1647 :  20 - 0x14
      12'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      12'h671: dout  = 8'b00000000; // 1649 :   0 - 0x0
      12'h672: dout  = 8'b00000000; // 1650 :   0 - 0x0
      12'h673: dout  = 8'b00000000; // 1651 :   0 - 0x0
      12'h674: dout  = 8'b10001110; // 1652 : 142 - 0x8e
      12'h675: dout  = 8'b11001001; // 1653 : 201 - 0xc9
      12'h676: dout  = 8'b11101010; // 1654 : 234 - 0xea
      12'h677: dout  = 8'b11111001; // 1655 : 249 - 0xf9
      12'h678: dout  = 8'b11111110; // 1656 : 254 - 0xfe -- Sprite 0xcf
      12'h679: dout  = 8'b11111000; // 1657 : 248 - 0xf8
      12'h67A: dout  = 8'b11111000; // 1658 : 248 - 0xf8
      12'h67B: dout  = 8'b11111000; // 1659 : 248 - 0xf8
      12'h67C: dout  = 8'b11110000; // 1660 : 240 - 0xf0
      12'h67D: dout  = 8'b11100000; // 1661 : 224 - 0xe0
      12'h67E: dout  = 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      12'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout  = 8'b00000100; // 1666 :   4 - 0x4
      12'h683: dout  = 8'b00100110; // 1667 :  38 - 0x26
      12'h684: dout  = 8'b00101011; // 1668 :  43 - 0x2b
      12'h685: dout  = 8'b01110001; // 1669 : 113 - 0x71
      12'h686: dout  = 8'b01000000; // 1670 :  64 - 0x40
      12'h687: dout  = 8'b01000111; // 1671 :  71 - 0x47
      12'h688: dout  = 8'b10001111; // 1672 : 143 - 0x8f -- Sprite 0xd1
      12'h689: dout  = 8'b10001111; // 1673 : 143 - 0x8f
      12'h68A: dout  = 8'b01001111; // 1674 :  79 - 0x4f
      12'h68B: dout  = 8'b01001111; // 1675 :  79 - 0x4f
      12'h68C: dout  = 8'b00111111; // 1676 :  63 - 0x3f
      12'h68D: dout  = 8'b00010011; // 1677 :  19 - 0x13
      12'h68E: dout  = 8'b00010001; // 1678 :  17 - 0x11
      12'h68F: dout  = 8'b00011111; // 1679 :  31 - 0x1f
      12'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0xd2
      12'h691: dout  = 8'b10000000; // 1681 : 128 - 0x80
      12'h692: dout  = 8'b11001000; // 1682 : 200 - 0xc8
      12'h693: dout  = 8'b11010100; // 1683 : 212 - 0xd4
      12'h694: dout  = 8'b00100100; // 1684 :  36 - 0x24
      12'h695: dout  = 8'b00000010; // 1685 :   2 - 0x2
      12'h696: dout  = 8'b00000010; // 1686 :   2 - 0x2
      12'h697: dout  = 8'b11110010; // 1687 : 242 - 0xf2
      12'h698: dout  = 8'b11110010; // 1688 : 242 - 0xf2 -- Sprite 0xd3
      12'h699: dout  = 8'b11110010; // 1689 : 242 - 0xf2
      12'h69A: dout  = 8'b11110100; // 1690 : 244 - 0xf4
      12'h69B: dout  = 8'b11110100; // 1691 : 244 - 0xf4
      12'h69C: dout  = 8'b11110100; // 1692 : 244 - 0xf4
      12'h69D: dout  = 8'b11001000; // 1693 : 200 - 0xc8
      12'h69E: dout  = 8'b01000100; // 1694 :  68 - 0x44
      12'h69F: dout  = 8'b01111100; // 1695 : 124 - 0x7c
      12'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      12'h6A1: dout  = 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout  = 8'b00000000; // 1698 :   0 - 0x0
      12'h6A3: dout  = 8'b00001001; // 1699 :   9 - 0x9
      12'h6A4: dout  = 8'b00011010; // 1700 :  26 - 0x1a
      12'h6A5: dout  = 8'b00010100; // 1701 :  20 - 0x14
      12'h6A6: dout  = 8'b00100000; // 1702 :  32 - 0x20
      12'h6A7: dout  = 8'b01000111; // 1703 :  71 - 0x47
      12'h6A8: dout  = 8'b10001111; // 1704 : 143 - 0x8f -- Sprite 0xd5
      12'h6A9: dout  = 8'b10001111; // 1705 : 143 - 0x8f
      12'h6AA: dout  = 8'b01001111; // 1706 :  79 - 0x4f
      12'h6AB: dout  = 8'b01001111; // 1707 :  79 - 0x4f
      12'h6AC: dout  = 8'b00111111; // 1708 :  63 - 0x3f
      12'h6AD: dout  = 8'b01000111; // 1709 :  71 - 0x47
      12'h6AE: dout  = 8'b00100010; // 1710 :  34 - 0x22
      12'h6AF: dout  = 8'b00011100; // 1711 :  28 - 0x1c
      12'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      12'h6B1: dout  = 8'b01000000; // 1713 :  64 - 0x40
      12'h6B2: dout  = 8'b11000000; // 1714 : 192 - 0xc0
      12'h6B3: dout  = 8'b00101100; // 1715 :  44 - 0x2c
      12'h6B4: dout  = 8'b00110100; // 1716 :  52 - 0x34
      12'h6B5: dout  = 8'b00000100; // 1717 :   4 - 0x4
      12'h6B6: dout  = 8'b00000010; // 1718 :   2 - 0x2
      12'h6B7: dout  = 8'b11110010; // 1719 : 242 - 0xf2
      12'h6B8: dout  = 8'b11110010; // 1720 : 242 - 0xf2 -- Sprite 0xd7
      12'h6B9: dout  = 8'b11110010; // 1721 : 242 - 0xf2
      12'h6BA: dout  = 8'b11110100; // 1722 : 244 - 0xf4
      12'h6BB: dout  = 8'b11110111; // 1723 : 247 - 0xf7
      12'h6BC: dout  = 8'b11111101; // 1724 : 253 - 0xfd
      12'h6BD: dout  = 8'b11100001; // 1725 : 225 - 0xe1
      12'h6BE: dout  = 8'b00010010; // 1726 :  18 - 0x12
      12'h6BF: dout  = 8'b00001100; // 1727 :  12 - 0xc
      12'h6C0: dout  = 8'b01111000; // 1728 : 120 - 0x78 -- Sprite 0xd8
      12'h6C1: dout  = 8'b01001110; // 1729 :  78 - 0x4e
      12'h6C2: dout  = 8'b11000010; // 1730 : 194 - 0xc2
      12'h6C3: dout  = 8'b10011010; // 1731 : 154 - 0x9a
      12'h6C4: dout  = 8'b10011011; // 1732 : 155 - 0x9b
      12'h6C5: dout  = 8'b11011001; // 1733 : 217 - 0xd9
      12'h6C6: dout  = 8'b01100011; // 1734 :  99 - 0x63
      12'h6C7: dout  = 8'b00111110; // 1735 :  62 - 0x3e
      12'h6C8: dout  = 8'b00011110; // 1736 :  30 - 0x1e -- Sprite 0xd9
      12'h6C9: dout  = 8'b01110001; // 1737 : 113 - 0x71
      12'h6CA: dout  = 8'b01001001; // 1738 :  73 - 0x49
      12'h6CB: dout  = 8'b10111001; // 1739 : 185 - 0xb9
      12'h6CC: dout  = 8'b10011101; // 1740 : 157 - 0x9d
      12'h6CD: dout  = 8'b01010010; // 1741 :  82 - 0x52
      12'h6CE: dout  = 8'b01110010; // 1742 : 114 - 0x72
      12'h6CF: dout  = 8'b00011110; // 1743 :  30 - 0x1e
      12'h6D0: dout  = 8'b01100000; // 1744 :  96 - 0x60 -- Sprite 0xda
      12'h6D1: dout  = 8'b01011110; // 1745 :  94 - 0x5e
      12'h6D2: dout  = 8'b10001001; // 1746 : 137 - 0x89
      12'h6D3: dout  = 8'b10111101; // 1747 : 189 - 0xbd
      12'h6D4: dout  = 8'b10011101; // 1748 : 157 - 0x9d
      12'h6D5: dout  = 8'b11010011; // 1749 : 211 - 0xd3
      12'h6D6: dout  = 8'b01000110; // 1750 :  70 - 0x46
      12'h6D7: dout  = 8'b01111100; // 1751 : 124 - 0x7c
      12'h6D8: dout  = 8'b00011110; // 1752 :  30 - 0x1e -- Sprite 0xdb
      12'h6D9: dout  = 8'b00100011; // 1753 :  35 - 0x23
      12'h6DA: dout  = 8'b01001001; // 1754 :  73 - 0x49
      12'h6DB: dout  = 8'b10111101; // 1755 : 189 - 0xbd
      12'h6DC: dout  = 8'b10011001; // 1756 : 153 - 0x99
      12'h6DD: dout  = 8'b01000011; // 1757 :  67 - 0x43
      12'h6DE: dout  = 8'b01101110; // 1758 : 110 - 0x6e
      12'h6DF: dout  = 8'b00011000; // 1759 :  24 - 0x18
      12'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0xdc
      12'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout  = 8'b00000001; // 1762 :   1 - 0x1
      12'h6E3: dout  = 8'b00000010; // 1763 :   2 - 0x2
      12'h6E4: dout  = 8'b00000100; // 1764 :   4 - 0x4
      12'h6E5: dout  = 8'b00000010; // 1765 :   2 - 0x2
      12'h6E6: dout  = 8'b00011110; // 1766 :  30 - 0x1e
      12'h6E7: dout  = 8'b00010000; // 1767 :  16 - 0x10
      12'h6E8: dout  = 8'b00001000; // 1768 :   8 - 0x8 -- Sprite 0xdd
      12'h6E9: dout  = 8'b00001101; // 1769 :  13 - 0xd
      12'h6EA: dout  = 8'b00111010; // 1770 :  58 - 0x3a
      12'h6EB: dout  = 8'b00100101; // 1771 :  37 - 0x25
      12'h6EC: dout  = 8'b00011011; // 1772 :  27 - 0x1b
      12'h6ED: dout  = 8'b00001111; // 1773 :  15 - 0xf
      12'h6EE: dout  = 8'b00000111; // 1774 :   7 - 0x7
      12'h6EF: dout  = 8'b00000011; // 1775 :   3 - 0x3
      12'h6F0: dout  = 8'b00000000; // 1776 :   0 - 0x0 -- Sprite 0xde
      12'h6F1: dout  = 8'b00000000; // 1777 :   0 - 0x0
      12'h6F2: dout  = 8'b00000000; // 1778 :   0 - 0x0
      12'h6F3: dout  = 8'b11000000; // 1779 : 192 - 0xc0
      12'h6F4: dout  = 8'b01000000; // 1780 :  64 - 0x40
      12'h6F5: dout  = 8'b01011000; // 1781 :  88 - 0x58
      12'h6F6: dout  = 8'b01101000; // 1782 : 104 - 0x68
      12'h6F7: dout  = 8'b00001000; // 1783 :   8 - 0x8
      12'h6F8: dout  = 8'b00010000; // 1784 :  16 - 0x10 -- Sprite 0xdf
      12'h6F9: dout  = 8'b01011100; // 1785 :  92 - 0x5c
      12'h6FA: dout  = 8'b10101000; // 1786 : 168 - 0xa8
      12'h6FB: dout  = 8'b11011000; // 1787 : 216 - 0xd8
      12'h6FC: dout  = 8'b10111000; // 1788 : 184 - 0xb8
      12'h6FD: dout  = 8'b11110000; // 1789 : 240 - 0xf0
      12'h6FE: dout  = 8'b11100000; // 1790 : 224 - 0xe0
      12'h6FF: dout  = 8'b11000000; // 1791 : 192 - 0xc0
      12'h700: dout  = 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0xe0
      12'h701: dout  = 8'b00000000; // 1793 :   0 - 0x0
      12'h702: dout  = 8'b00000000; // 1794 :   0 - 0x0
      12'h703: dout  = 8'b00010011; // 1795 :  19 - 0x13
      12'h704: dout  = 8'b00010011; // 1796 :  19 - 0x13
      12'h705: dout  = 8'b00110111; // 1797 :  55 - 0x37
      12'h706: dout  = 8'b00110111; // 1798 :  55 - 0x37
      12'h707: dout  = 8'b00000111; // 1799 :   7 - 0x7
      12'h708: dout  = 8'b00000111; // 1800 :   7 - 0x7 -- Sprite 0xe1
      12'h709: dout  = 8'b00000100; // 1801 :   4 - 0x4
      12'h70A: dout  = 8'b00000000; // 1802 :   0 - 0x0
      12'h70B: dout  = 8'b00000000; // 1803 :   0 - 0x0
      12'h70C: dout  = 8'b00000000; // 1804 :   0 - 0x0
      12'h70D: dout  = 8'b00100000; // 1805 :  32 - 0x20
      12'h70E: dout  = 8'b01110000; // 1806 : 112 - 0x70
      12'h70F: dout  = 8'b11111000; // 1807 : 248 - 0xf8
      12'h710: dout  = 8'b00000000; // 1808 :   0 - 0x0 -- Sprite 0xe2
      12'h711: dout  = 8'b00000000; // 1809 :   0 - 0x0
      12'h712: dout  = 8'b00000000; // 1810 :   0 - 0x0
      12'h713: dout  = 8'b11111000; // 1811 : 248 - 0xf8
      12'h714: dout  = 8'b11111100; // 1812 : 252 - 0xfc
      12'h715: dout  = 8'b11111100; // 1813 : 252 - 0xfc
      12'h716: dout  = 8'b11111100; // 1814 : 252 - 0xfc
      12'h717: dout  = 8'b11111101; // 1815 : 253 - 0xfd
      12'h718: dout  = 8'b11111100; // 1816 : 252 - 0xfc -- Sprite 0xe3
      12'h719: dout  = 8'b00011100; // 1817 :  28 - 0x1c
      12'h71A: dout  = 8'b11000000; // 1818 : 192 - 0xc0
      12'h71B: dout  = 8'b11100000; // 1819 : 224 - 0xe0
      12'h71C: dout  = 8'b00000000; // 1820 :   0 - 0x0
      12'h71D: dout  = 8'b00000000; // 1821 :   0 - 0x0
      12'h71E: dout  = 8'b00000110; // 1822 :   6 - 0x6
      12'h71F: dout  = 8'b00001111; // 1823 :  15 - 0xf
      12'h720: dout  = 8'b00000000; // 1824 :   0 - 0x0 -- Sprite 0xe4
      12'h721: dout  = 8'b00000000; // 1825 :   0 - 0x0
      12'h722: dout  = 8'b00000000; // 1826 :   0 - 0x0
      12'h723: dout  = 8'b00010011; // 1827 :  19 - 0x13
      12'h724: dout  = 8'b00010011; // 1828 :  19 - 0x13
      12'h725: dout  = 8'b00110111; // 1829 :  55 - 0x37
      12'h726: dout  = 8'b00110111; // 1830 :  55 - 0x37
      12'h727: dout  = 8'b00000111; // 1831 :   7 - 0x7
      12'h728: dout  = 8'b00000111; // 1832 :   7 - 0x7 -- Sprite 0xe5
      12'h729: dout  = 8'b00000100; // 1833 :   4 - 0x4
      12'h72A: dout  = 8'b00000001; // 1834 :   1 - 0x1
      12'h72B: dout  = 8'b00000000; // 1835 :   0 - 0x0
      12'h72C: dout  = 8'b00000000; // 1836 :   0 - 0x0
      12'h72D: dout  = 8'b00100000; // 1837 :  32 - 0x20
      12'h72E: dout  = 8'b01110000; // 1838 : 112 - 0x70
      12'h72F: dout  = 8'b11111000; // 1839 : 248 - 0xf8
      12'h730: dout  = 8'b00000000; // 1840 :   0 - 0x0 -- Sprite 0xe6
      12'h731: dout  = 8'b00000000; // 1841 :   0 - 0x0
      12'h732: dout  = 8'b00000000; // 1842 :   0 - 0x0
      12'h733: dout  = 8'b11111100; // 1843 : 252 - 0xfc
      12'h734: dout  = 8'b11111100; // 1844 : 252 - 0xfc
      12'h735: dout  = 8'b11111100; // 1845 : 252 - 0xfc
      12'h736: dout  = 8'b11111100; // 1846 : 252 - 0xfc
      12'h737: dout  = 8'b11111101; // 1847 : 253 - 0xfd
      12'h738: dout  = 8'b11111100; // 1848 : 252 - 0xfc -- Sprite 0xe7
      12'h739: dout  = 8'b00001100; // 1849 :  12 - 0xc
      12'h73A: dout  = 8'b11000000; // 1850 : 192 - 0xc0
      12'h73B: dout  = 8'b11110000; // 1851 : 240 - 0xf0
      12'h73C: dout  = 8'b11110000; // 1852 : 240 - 0xf0
      12'h73D: dout  = 8'b00000000; // 1853 :   0 - 0x0
      12'h73E: dout  = 8'b00000110; // 1854 :   6 - 0x6
      12'h73F: dout  = 8'b00001111; // 1855 :  15 - 0xf
      12'h740: dout  = 8'b11111111; // 1856 : 255 - 0xff -- Sprite 0xe8
      12'h741: dout  = 8'b11111111; // 1857 : 255 - 0xff
      12'h742: dout  = 8'b01111111; // 1858 : 127 - 0x7f
      12'h743: dout  = 8'b01111111; // 1859 : 127 - 0x7f
      12'h744: dout  = 8'b01111111; // 1860 : 127 - 0x7f
      12'h745: dout  = 8'b00111111; // 1861 :  63 - 0x3f
      12'h746: dout  = 8'b00111111; // 1862 :  63 - 0x3f
      12'h747: dout  = 8'b00111111; // 1863 :  63 - 0x3f
      12'h748: dout  = 8'b00111100; // 1864 :  60 - 0x3c -- Sprite 0xe9
      12'h749: dout  = 8'b00111110; // 1865 :  62 - 0x3e
      12'h74A: dout  = 8'b00011111; // 1866 :  31 - 0x1f
      12'h74B: dout  = 8'b00001111; // 1867 :  15 - 0xf
      12'h74C: dout  = 8'b00000111; // 1868 :   7 - 0x7
      12'h74D: dout  = 8'b00000000; // 1869 :   0 - 0x0
      12'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      12'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout  = 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0xea
      12'h751: dout  = 8'b11111110; // 1873 : 254 - 0xfe
      12'h752: dout  = 8'b11111110; // 1874 : 254 - 0xfe
      12'h753: dout  = 8'b11111100; // 1875 : 252 - 0xfc
      12'h754: dout  = 8'b11111000; // 1876 : 248 - 0xf8
      12'h755: dout  = 8'b11110000; // 1877 : 240 - 0xf0
      12'h756: dout  = 8'b10110000; // 1878 : 176 - 0xb0
      12'h757: dout  = 8'b00111001; // 1879 :  57 - 0x39
      12'h758: dout  = 8'b00011111; // 1880 :  31 - 0x1f -- Sprite 0xeb
      12'h759: dout  = 8'b11001111; // 1881 : 207 - 0xcf
      12'h75A: dout  = 8'b11000110; // 1882 : 198 - 0xc6
      12'h75B: dout  = 8'b10000000; // 1883 : 128 - 0x80
      12'h75C: dout  = 8'b00000000; // 1884 :   0 - 0x0
      12'h75D: dout  = 8'b00000000; // 1885 :   0 - 0x0
      12'h75E: dout  = 8'b00000000; // 1886 :   0 - 0x0
      12'h75F: dout  = 8'b00000000; // 1887 :   0 - 0x0
      12'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      12'h761: dout  = 8'b00000000; // 1889 :   0 - 0x0
      12'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout  = 8'b00000000; // 1891 :   0 - 0x0
      12'h764: dout  = 8'b00000000; // 1892 :   0 - 0x0
      12'h765: dout  = 8'b00000000; // 1893 :   0 - 0x0
      12'h766: dout  = 8'b00001100; // 1894 :  12 - 0xc
      12'h767: dout  = 8'b00001100; // 1895 :  12 - 0xc
      12'h768: dout  = 8'b00110000; // 1896 :  48 - 0x30 -- Sprite 0xed
      12'h769: dout  = 8'b01000011; // 1897 :  67 - 0x43
      12'h76A: dout  = 8'b01000000; // 1898 :  64 - 0x40
      12'h76B: dout  = 8'b01100000; // 1899 :  96 - 0x60
      12'h76C: dout  = 8'b00000011; // 1900 :   3 - 0x3
      12'h76D: dout  = 8'b00000000; // 1901 :   0 - 0x0
      12'h76E: dout  = 8'b01111111; // 1902 : 127 - 0x7f
      12'h76F: dout  = 8'b00000000; // 1903 :   0 - 0x0
      12'h770: dout  = 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0xee
      12'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout  = 8'b00000000; // 1906 :   0 - 0x0
      12'h773: dout  = 8'b00000000; // 1907 :   0 - 0x0
      12'h774: dout  = 8'b00000000; // 1908 :   0 - 0x0
      12'h775: dout  = 8'b00000000; // 1909 :   0 - 0x0
      12'h776: dout  = 8'b00110000; // 1910 :  48 - 0x30
      12'h777: dout  = 8'b00110000; // 1911 :  48 - 0x30
      12'h778: dout  = 8'b00001110; // 1912 :  14 - 0xe -- Sprite 0xef
      12'h779: dout  = 8'b11001011; // 1913 : 203 - 0xcb
      12'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      12'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      12'h77C: dout  = 8'b11000000; // 1916 : 192 - 0xc0
      12'h77D: dout  = 8'b00000000; // 1917 :   0 - 0x0
      12'h77E: dout  = 8'b11111110; // 1918 : 254 - 0xfe
      12'h77F: dout  = 8'b00000000; // 1919 :   0 - 0x0
      12'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      12'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout  = 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout  = 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout  = 8'b00001100; // 1926 :  12 - 0xc
      12'h787: dout  = 8'b00001100; // 1927 :  12 - 0xc
      12'h788: dout  = 8'b00110000; // 1928 :  48 - 0x30 -- Sprite 0xf1
      12'h789: dout  = 8'b00100011; // 1929 :  35 - 0x23
      12'h78A: dout  = 8'b00100000; // 1930 :  32 - 0x20
      12'h78B: dout  = 8'b01100000; // 1931 :  96 - 0x60
      12'h78C: dout  = 8'b00000011; // 1932 :   3 - 0x3
      12'h78D: dout  = 8'b00000000; // 1933 :   0 - 0x0
      12'h78E: dout  = 8'b01111111; // 1934 : 127 - 0x7f
      12'h78F: dout  = 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout  = 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0xf2
      12'h791: dout  = 8'b00000000; // 1937 :   0 - 0x0
      12'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout  = 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout  = 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout  = 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout  = 8'b00110000; // 1942 :  48 - 0x30
      12'h797: dout  = 8'b00110000; // 1943 :  48 - 0x30
      12'h798: dout  = 8'b00001001; // 1944 :   9 - 0x9 -- Sprite 0xf3
      12'h799: dout  = 8'b11001111; // 1945 : 207 - 0xcf
      12'h79A: dout  = 8'b00000000; // 1946 :   0 - 0x0
      12'h79B: dout  = 8'b00000000; // 1947 :   0 - 0x0
      12'h79C: dout  = 8'b11000000; // 1948 : 192 - 0xc0
      12'h79D: dout  = 8'b00000000; // 1949 :   0 - 0x0
      12'h79E: dout  = 8'b11111110; // 1950 : 254 - 0xfe
      12'h79F: dout  = 8'b00000000; // 1951 :   0 - 0x0
      12'h7A0: dout  = 8'b00111111; // 1952 :  63 - 0x3f -- Sprite 0xf4
      12'h7A1: dout  = 8'b00110101; // 1953 :  53 - 0x35
      12'h7A2: dout  = 8'b00011010; // 1954 :  26 - 0x1a
      12'h7A3: dout  = 8'b00001101; // 1955 :  13 - 0xd
      12'h7A4: dout  = 8'b00001010; // 1956 :  10 - 0xa
      12'h7A5: dout  = 8'b00001101; // 1957 :  13 - 0xd
      12'h7A6: dout  = 8'b00001000; // 1958 :   8 - 0x8
      12'h7A7: dout  = 8'b00111000; // 1959 :  56 - 0x38
      12'h7A8: dout  = 8'b01110011; // 1960 : 115 - 0x73 -- Sprite 0xf5
      12'h7A9: dout  = 8'b11000100; // 1961 : 196 - 0xc4
      12'h7AA: dout  = 8'b11000100; // 1962 : 196 - 0xc4
      12'h7AB: dout  = 8'b11000000; // 1963 : 192 - 0xc0
      12'h7AC: dout  = 8'b11000001; // 1964 : 193 - 0xc1
      12'h7AD: dout  = 8'b11000000; // 1965 : 192 - 0xc0
      12'h7AE: dout  = 8'b01100001; // 1966 :  97 - 0x61
      12'h7AF: dout  = 8'b00111111; // 1967 :  63 - 0x3f
      12'h7B0: dout  = 8'b11111100; // 1968 : 252 - 0xfc -- Sprite 0xf6
      12'h7B1: dout  = 8'b01010100; // 1969 :  84 - 0x54
      12'h7B2: dout  = 8'b10101000; // 1970 : 168 - 0xa8
      12'h7B3: dout  = 8'b01010000; // 1971 :  80 - 0x50
      12'h7B4: dout  = 8'b10110000; // 1972 : 176 - 0xb0
      12'h7B5: dout  = 8'b01010000; // 1973 :  80 - 0x50
      12'h7B6: dout  = 8'b10010000; // 1974 : 144 - 0x90
      12'h7B7: dout  = 8'b00011100; // 1975 :  28 - 0x1c
      12'h7B8: dout  = 8'b10000110; // 1976 : 134 - 0x86 -- Sprite 0xf7
      12'h7B9: dout  = 8'b01000010; // 1977 :  66 - 0x42
      12'h7BA: dout  = 8'b01000111; // 1978 :  71 - 0x47
      12'h7BB: dout  = 8'b01000001; // 1979 :  65 - 0x41
      12'h7BC: dout  = 8'b10000011; // 1980 : 131 - 0x83
      12'h7BD: dout  = 8'b00000001; // 1981 :   1 - 0x1
      12'h7BE: dout  = 8'b10000110; // 1982 : 134 - 0x86
      12'h7BF: dout  = 8'b11111100; // 1983 : 252 - 0xfc
      12'h7C0: dout  = 8'b11100100; // 1984 : 228 - 0xe4 -- Sprite 0xf8
      12'h7C1: dout  = 8'b11100100; // 1985 : 228 - 0xe4
      12'h7C2: dout  = 8'b11101111; // 1986 : 239 - 0xef
      12'h7C3: dout  = 8'b11101111; // 1987 : 239 - 0xef
      12'h7C4: dout  = 8'b11111111; // 1988 : 255 - 0xff
      12'h7C5: dout  = 8'b11111111; // 1989 : 255 - 0xff
      12'h7C6: dout  = 8'b01111111; // 1990 : 127 - 0x7f
      12'h7C7: dout  = 8'b01111111; // 1991 : 127 - 0x7f
      12'h7C8: dout  = 8'b00111111; // 1992 :  63 - 0x3f -- Sprite 0xf9
      12'h7C9: dout  = 8'b01111111; // 1993 : 127 - 0x7f
      12'h7CA: dout  = 8'b01111111; // 1994 : 127 - 0x7f
      12'h7CB: dout  = 8'b11111111; // 1995 : 255 - 0xff
      12'h7CC: dout  = 8'b11111111; // 1996 : 255 - 0xff
      12'h7CD: dout  = 8'b11111111; // 1997 : 255 - 0xff
      12'h7CE: dout  = 8'b11111111; // 1998 : 255 - 0xff
      12'h7CF: dout  = 8'b11111111; // 1999 : 255 - 0xff
      12'h7D0: dout  = 8'b00010011; // 2000 :  19 - 0x13 -- Sprite 0xfa
      12'h7D1: dout  = 8'b00010011; // 2001 :  19 - 0x13
      12'h7D2: dout  = 8'b11111011; // 2002 : 251 - 0xfb
      12'h7D3: dout  = 8'b11111011; // 2003 : 251 - 0xfb
      12'h7D4: dout  = 8'b11111111; // 2004 : 255 - 0xff
      12'h7D5: dout  = 8'b11111111; // 2005 : 255 - 0xff
      12'h7D6: dout  = 8'b11111110; // 2006 : 254 - 0xfe
      12'h7D7: dout  = 8'b11111110; // 2007 : 254 - 0xfe
      12'h7D8: dout  = 8'b11111110; // 2008 : 254 - 0xfe -- Sprite 0xfb
      12'h7D9: dout  = 8'b11111111; // 2009 : 255 - 0xff
      12'h7DA: dout  = 8'b11111111; // 2010 : 255 - 0xff
      12'h7DB: dout  = 8'b11111111; // 2011 : 255 - 0xff
      12'h7DC: dout  = 8'b11111111; // 2012 : 255 - 0xff
      12'h7DD: dout  = 8'b11111111; // 2013 : 255 - 0xff
      12'h7DE: dout  = 8'b11111111; // 2014 : 255 - 0xff
      12'h7DF: dout  = 8'b11111111; // 2015 : 255 - 0xff
      12'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      12'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout  = 8'b01111100; // 2018 : 124 - 0x7c
      12'h7E3: dout  = 8'b11111110; // 2019 : 254 - 0xfe
      12'h7E4: dout  = 8'b11111110; // 2020 : 254 - 0xfe
      12'h7E5: dout  = 8'b01111100; // 2021 : 124 - 0x7c
      12'h7E6: dout  = 8'b01000100; // 2022 :  68 - 0x44
      12'h7E7: dout  = 8'b10000010; // 2023 : 130 - 0x82
      12'h7E8: dout  = 8'b10000010; // 2024 : 130 - 0x82 -- Sprite 0xfd
      12'h7E9: dout  = 8'b10000010; // 2025 : 130 - 0x82
      12'h7EA: dout  = 8'b10000010; // 2026 : 130 - 0x82
      12'h7EB: dout  = 8'b11000110; // 2027 : 198 - 0xc6
      12'h7EC: dout  = 8'b11111110; // 2028 : 254 - 0xfe
      12'h7ED: dout  = 8'b11111110; // 2029 : 254 - 0xfe
      12'h7EE: dout  = 8'b10111010; // 2030 : 186 - 0xba
      12'h7EF: dout  = 8'b01111100; // 2031 : 124 - 0x7c
      12'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0xfe
      12'h7F1: dout  = 8'b00011001; // 2033 :  25 - 0x19
      12'h7F2: dout  = 8'b00111110; // 2034 :  62 - 0x3e
      12'h7F3: dout  = 8'b00111100; // 2035 :  60 - 0x3c
      12'h7F4: dout  = 8'b00111100; // 2036 :  60 - 0x3c
      12'h7F5: dout  = 8'b00111100; // 2037 :  60 - 0x3c
      12'h7F6: dout  = 8'b00111110; // 2038 :  62 - 0x3e
      12'h7F7: dout  = 8'b00011001; // 2039 :  25 - 0x19
      12'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      12'h7F9: dout  = 8'b11111110; // 2041 : 254 - 0xfe
      12'h7FA: dout  = 8'b00011101; // 2042 :  29 - 0x1d
      12'h7FB: dout  = 8'b00001111; // 2043 :  15 - 0xf
      12'h7FC: dout  = 8'b00001111; // 2044 :  15 - 0xf
      12'h7FD: dout  = 8'b00001111; // 2045 :  15 - 0xf
      12'h7FE: dout  = 8'b00011101; // 2046 :  29 - 0x1d
      12'h7FF: dout  = 8'b11111110; // 2047 : 254 - 0xfe
          // Background pattern Table
      12'h800: dout  = 8'b11111111; // 2048 : 255 - 0xff -- Background 0x0
      12'h801: dout  = 8'b11111111; // 2049 : 255 - 0xff
      12'h802: dout  = 8'b11000000; // 2050 : 192 - 0xc0
      12'h803: dout  = 8'b11000000; // 2051 : 192 - 0xc0
      12'h804: dout  = 8'b11000000; // 2052 : 192 - 0xc0
      12'h805: dout  = 8'b11000000; // 2053 : 192 - 0xc0
      12'h806: dout  = 8'b11010101; // 2054 : 213 - 0xd5
      12'h807: dout  = 8'b11111111; // 2055 : 255 - 0xff
      12'h808: dout  = 8'b11111111; // 2056 : 255 - 0xff -- Background 0x1
      12'h809: dout  = 8'b11111111; // 2057 : 255 - 0xff
      12'h80A: dout  = 8'b11001110; // 2058 : 206 - 0xce
      12'h80B: dout  = 8'b11000110; // 2059 : 198 - 0xc6
      12'h80C: dout  = 8'b11001110; // 2060 : 206 - 0xce
      12'h80D: dout  = 8'b11000110; // 2061 : 198 - 0xc6
      12'h80E: dout  = 8'b11101110; // 2062 : 238 - 0xee
      12'h80F: dout  = 8'b11111111; // 2063 : 255 - 0xff
      12'h810: dout  = 8'b11111111; // 2064 : 255 - 0xff -- Background 0x2
      12'h811: dout  = 8'b11111111; // 2065 : 255 - 0xff
      12'h812: dout  = 8'b01110001; // 2066 : 113 - 0x71
      12'h813: dout  = 8'b00110011; // 2067 :  51 - 0x33
      12'h814: dout  = 8'b01110001; // 2068 : 113 - 0x71
      12'h815: dout  = 8'b00110011; // 2069 :  51 - 0x33
      12'h816: dout  = 8'b01110101; // 2070 : 117 - 0x75
      12'h817: dout  = 8'b11111111; // 2071 : 255 - 0xff
      12'h818: dout  = 8'b11111111; // 2072 : 255 - 0xff -- Background 0x3
      12'h819: dout  = 8'b11111111; // 2073 : 255 - 0xff
      12'h81A: dout  = 8'b00000011; // 2074 :   3 - 0x3
      12'h81B: dout  = 8'b00000001; // 2075 :   1 - 0x1
      12'h81C: dout  = 8'b00000011; // 2076 :   3 - 0x3
      12'h81D: dout  = 8'b00000001; // 2077 :   1 - 0x1
      12'h81E: dout  = 8'b10101011; // 2078 : 171 - 0xab
      12'h81F: dout  = 8'b11111111; // 2079 : 255 - 0xff
      12'h820: dout  = 8'b11111111; // 2080 : 255 - 0xff -- Background 0x4
      12'h821: dout  = 8'b11111111; // 2081 : 255 - 0xff
      12'h822: dout  = 8'b11100000; // 2082 : 224 - 0xe0
      12'h823: dout  = 8'b11000110; // 2083 : 198 - 0xc6
      12'h824: dout  = 8'b11000110; // 2084 : 198 - 0xc6
      12'h825: dout  = 8'b11110110; // 2085 : 246 - 0xf6
      12'h826: dout  = 8'b11110000; // 2086 : 240 - 0xf0
      12'h827: dout  = 8'b11110001; // 2087 : 241 - 0xf1
      12'h828: dout  = 8'b11000111; // 2088 : 199 - 0xc7 -- Background 0x5
      12'h829: dout  = 8'b11001111; // 2089 : 207 - 0xcf
      12'h82A: dout  = 8'b11011111; // 2090 : 223 - 0xdf
      12'h82B: dout  = 8'b11011111; // 2091 : 223 - 0xdf
      12'h82C: dout  = 8'b11001110; // 2092 : 206 - 0xce
      12'h82D: dout  = 8'b11100000; // 2093 : 224 - 0xe0
      12'h82E: dout  = 8'b11111111; // 2094 : 255 - 0xff
      12'h82F: dout  = 8'b11111111; // 2095 : 255 - 0xff
      12'h830: dout  = 8'b11111111; // 2096 : 255 - 0xff -- Background 0x6
      12'h831: dout  = 8'b11111111; // 2097 : 255 - 0xff
      12'h832: dout  = 8'b00000111; // 2098 :   7 - 0x7
      12'h833: dout  = 8'b01100011; // 2099 :  99 - 0x63
      12'h834: dout  = 8'b01100011; // 2100 :  99 - 0x63
      12'h835: dout  = 8'b01101111; // 2101 : 111 - 0x6f
      12'h836: dout  = 8'b00001111; // 2102 :  15 - 0xf
      12'h837: dout  = 8'b10001111; // 2103 : 143 - 0x8f
      12'h838: dout  = 8'b11100011; // 2104 : 227 - 0xe3 -- Background 0x7
      12'h839: dout  = 8'b11110011; // 2105 : 243 - 0xf3
      12'h83A: dout  = 8'b11111011; // 2106 : 251 - 0xfb
      12'h83B: dout  = 8'b11111011; // 2107 : 251 - 0xfb
      12'h83C: dout  = 8'b01110011; // 2108 : 115 - 0x73
      12'h83D: dout  = 8'b00000111; // 2109 :   7 - 0x7
      12'h83E: dout  = 8'b11111111; // 2110 : 255 - 0xff
      12'h83F: dout  = 8'b11111111; // 2111 : 255 - 0xff
      12'h840: dout  = 8'b11111111; // 2112 : 255 - 0xff -- Background 0x8
      12'h841: dout  = 8'b11010101; // 2113 : 213 - 0xd5
      12'h842: dout  = 8'b10101010; // 2114 : 170 - 0xaa
      12'h843: dout  = 8'b11010101; // 2115 : 213 - 0xd5
      12'h844: dout  = 8'b10101010; // 2116 : 170 - 0xaa
      12'h845: dout  = 8'b11010101; // 2117 : 213 - 0xd5
      12'h846: dout  = 8'b10101010; // 2118 : 170 - 0xaa
      12'h847: dout  = 8'b11010101; // 2119 : 213 - 0xd5
      12'h848: dout  = 8'b10101010; // 2120 : 170 - 0xaa -- Background 0x9
      12'h849: dout  = 8'b11010101; // 2121 : 213 - 0xd5
      12'h84A: dout  = 8'b10101010; // 2122 : 170 - 0xaa
      12'h84B: dout  = 8'b11010101; // 2123 : 213 - 0xd5
      12'h84C: dout  = 8'b10101010; // 2124 : 170 - 0xaa
      12'h84D: dout  = 8'b11110101; // 2125 : 245 - 0xf5
      12'h84E: dout  = 8'b10101010; // 2126 : 170 - 0xaa
      12'h84F: dout  = 8'b11111111; // 2127 : 255 - 0xff
      12'h850: dout  = 8'b11111111; // 2128 : 255 - 0xff -- Background 0xa
      12'h851: dout  = 8'b01010101; // 2129 :  85 - 0x55
      12'h852: dout  = 8'b10101111; // 2130 : 175 - 0xaf
      12'h853: dout  = 8'b01010101; // 2131 :  85 - 0x55
      12'h854: dout  = 8'b10101011; // 2132 : 171 - 0xab
      12'h855: dout  = 8'b01010101; // 2133 :  85 - 0x55
      12'h856: dout  = 8'b10101011; // 2134 : 171 - 0xab
      12'h857: dout  = 8'b01010101; // 2135 :  85 - 0x55
      12'h858: dout  = 8'b10101011; // 2136 : 171 - 0xab -- Background 0xb
      12'h859: dout  = 8'b01010101; // 2137 :  85 - 0x55
      12'h85A: dout  = 8'b10101011; // 2138 : 171 - 0xab
      12'h85B: dout  = 8'b01010101; // 2139 :  85 - 0x55
      12'h85C: dout  = 8'b10101011; // 2140 : 171 - 0xab
      12'h85D: dout  = 8'b01010101; // 2141 :  85 - 0x55
      12'h85E: dout  = 8'b10101011; // 2142 : 171 - 0xab
      12'h85F: dout  = 8'b11111111; // 2143 : 255 - 0xff
      12'h860: dout  = 8'b11111111; // 2144 : 255 - 0xff -- Background 0xc
      12'h861: dout  = 8'b11010101; // 2145 : 213 - 0xd5
      12'h862: dout  = 8'b10100000; // 2146 : 160 - 0xa0
      12'h863: dout  = 8'b11010000; // 2147 : 208 - 0xd0
      12'h864: dout  = 8'b10001111; // 2148 : 143 - 0x8f
      12'h865: dout  = 8'b11001000; // 2149 : 200 - 0xc8
      12'h866: dout  = 8'b10001000; // 2150 : 136 - 0x88
      12'h867: dout  = 8'b11001000; // 2151 : 200 - 0xc8
      12'h868: dout  = 8'b10001000; // 2152 : 136 - 0x88 -- Background 0xd
      12'h869: dout  = 8'b11001000; // 2153 : 200 - 0xc8
      12'h86A: dout  = 8'b10001000; // 2154 : 136 - 0x88
      12'h86B: dout  = 8'b11001111; // 2155 : 207 - 0xcf
      12'h86C: dout  = 8'b10010000; // 2156 : 144 - 0x90
      12'h86D: dout  = 8'b11100000; // 2157 : 224 - 0xe0
      12'h86E: dout  = 8'b11101010; // 2158 : 234 - 0xea
      12'h86F: dout  = 8'b11111111; // 2159 : 255 - 0xff
      12'h870: dout  = 8'b11111111; // 2160 : 255 - 0xff -- Background 0xe
      12'h871: dout  = 8'b01011011; // 2161 :  91 - 0x5b
      12'h872: dout  = 8'b00000111; // 2162 :   7 - 0x7
      12'h873: dout  = 8'b00001001; // 2163 :   9 - 0x9
      12'h874: dout  = 8'b11110011; // 2164 : 243 - 0xf3
      12'h875: dout  = 8'b00010001; // 2165 :  17 - 0x11
      12'h876: dout  = 8'b00010011; // 2166 :  19 - 0x13
      12'h877: dout  = 8'b00010001; // 2167 :  17 - 0x11
      12'h878: dout  = 8'b00010011; // 2168 :  19 - 0x13 -- Background 0xf
      12'h879: dout  = 8'b00010001; // 2169 :  17 - 0x11
      12'h87A: dout  = 8'b00010011; // 2170 :  19 - 0x13
      12'h87B: dout  = 8'b11110001; // 2171 : 241 - 0xf1
      12'h87C: dout  = 8'b00001011; // 2172 :  11 - 0xb
      12'h87D: dout  = 8'b00000101; // 2173 :   5 - 0x5
      12'h87E: dout  = 8'b10101011; // 2174 : 171 - 0xab
      12'h87F: dout  = 8'b11111111; // 2175 : 255 - 0xff
      12'h880: dout  = 8'b11010000; // 2176 : 208 - 0xd0 -- Background 0x10
      12'h881: dout  = 8'b10010000; // 2177 : 144 - 0x90
      12'h882: dout  = 8'b11011111; // 2178 : 223 - 0xdf
      12'h883: dout  = 8'b10011010; // 2179 : 154 - 0x9a
      12'h884: dout  = 8'b11010101; // 2180 : 213 - 0xd5
      12'h885: dout  = 8'b10011111; // 2181 : 159 - 0x9f
      12'h886: dout  = 8'b11010000; // 2182 : 208 - 0xd0
      12'h887: dout  = 8'b10010000; // 2183 : 144 - 0x90
      12'h888: dout  = 8'b00001001; // 2184 :   9 - 0x9 -- Background 0x11
      12'h889: dout  = 8'b00001011; // 2185 :  11 - 0xb
      12'h88A: dout  = 8'b11111001; // 2186 : 249 - 0xf9
      12'h88B: dout  = 8'b10101011; // 2187 : 171 - 0xab
      12'h88C: dout  = 8'b01011001; // 2188 :  89 - 0x59
      12'h88D: dout  = 8'b11111011; // 2189 : 251 - 0xfb
      12'h88E: dout  = 8'b00001001; // 2190 :   9 - 0x9
      12'h88F: dout  = 8'b00001011; // 2191 :  11 - 0xb
      12'h890: dout  = 8'b00011000; // 2192 :  24 - 0x18 -- Background 0x12
      12'h891: dout  = 8'b00010100; // 2193 :  20 - 0x14
      12'h892: dout  = 8'b00010100; // 2194 :  20 - 0x14
      12'h893: dout  = 8'b00111010; // 2195 :  58 - 0x3a
      12'h894: dout  = 8'b00111010; // 2196 :  58 - 0x3a
      12'h895: dout  = 8'b01111010; // 2197 : 122 - 0x7a
      12'h896: dout  = 8'b01111010; // 2198 : 122 - 0x7a
      12'h897: dout  = 8'b01111010; // 2199 : 122 - 0x7a
      12'h898: dout  = 8'b11111011; // 2200 : 251 - 0xfb -- Background 0x13
      12'h899: dout  = 8'b11111101; // 2201 : 253 - 0xfd
      12'h89A: dout  = 8'b11111101; // 2202 : 253 - 0xfd
      12'h89B: dout  = 8'b11111101; // 2203 : 253 - 0xfd
      12'h89C: dout  = 8'b11111101; // 2204 : 253 - 0xfd
      12'h89D: dout  = 8'b11111101; // 2205 : 253 - 0xfd
      12'h89E: dout  = 8'b10000001; // 2206 : 129 - 0x81
      12'h89F: dout  = 8'b11111111; // 2207 : 255 - 0xff
      12'h8A0: dout  = 8'b00000000; // 2208 :   0 - 0x0 -- Background 0x14
      12'h8A1: dout  = 8'b00000111; // 2209 :   7 - 0x7
      12'h8A2: dout  = 8'b00000010; // 2210 :   2 - 0x2
      12'h8A3: dout  = 8'b00000100; // 2211 :   4 - 0x4
      12'h8A4: dout  = 8'b00000011; // 2212 :   3 - 0x3
      12'h8A5: dout  = 8'b00000011; // 2213 :   3 - 0x3
      12'h8A6: dout  = 8'b00001101; // 2214 :  13 - 0xd
      12'h8A7: dout  = 8'b00010111; // 2215 :  23 - 0x17
      12'h8A8: dout  = 8'b00101111; // 2216 :  47 - 0x2f -- Background 0x15
      12'h8A9: dout  = 8'b01001111; // 2217 :  79 - 0x4f
      12'h8AA: dout  = 8'b01001111; // 2218 :  79 - 0x4f
      12'h8AB: dout  = 8'b01001111; // 2219 :  79 - 0x4f
      12'h8AC: dout  = 8'b01001111; // 2220 :  79 - 0x4f
      12'h8AD: dout  = 8'b00100111; // 2221 :  39 - 0x27
      12'h8AE: dout  = 8'b00010000; // 2222 :  16 - 0x10
      12'h8AF: dout  = 8'b00001111; // 2223 :  15 - 0xf
      12'h8B0: dout  = 8'b00000000; // 2224 :   0 - 0x0 -- Background 0x16
      12'h8B1: dout  = 8'b11100000; // 2225 : 224 - 0xe0
      12'h8B2: dout  = 8'b10100000; // 2226 : 160 - 0xa0
      12'h8B3: dout  = 8'b00100000; // 2227 :  32 - 0x20
      12'h8B4: dout  = 8'b11000000; // 2228 : 192 - 0xc0
      12'h8B5: dout  = 8'b01000000; // 2229 :  64 - 0x40
      12'h8B6: dout  = 8'b00110000; // 2230 :  48 - 0x30
      12'h8B7: dout  = 8'b11101000; // 2231 : 232 - 0xe8
      12'h8B8: dout  = 8'b11110100; // 2232 : 244 - 0xf4 -- Background 0x17
      12'h8B9: dout  = 8'b11110010; // 2233 : 242 - 0xf2
      12'h8BA: dout  = 8'b11110010; // 2234 : 242 - 0xf2
      12'h8BB: dout  = 8'b11110010; // 2235 : 242 - 0xf2
      12'h8BC: dout  = 8'b11110010; // 2236 : 242 - 0xf2
      12'h8BD: dout  = 8'b11100100; // 2237 : 228 - 0xe4
      12'h8BE: dout  = 8'b00001000; // 2238 :   8 - 0x8
      12'h8BF: dout  = 8'b11110000; // 2239 : 240 - 0xf0
      12'h8C0: dout  = 8'b00111111; // 2240 :  63 - 0x3f -- Background 0x18
      12'h8C1: dout  = 8'b01000000; // 2241 :  64 - 0x40
      12'h8C2: dout  = 8'b01000000; // 2242 :  64 - 0x40
      12'h8C3: dout  = 8'b10000000; // 2243 : 128 - 0x80
      12'h8C4: dout  = 8'b10000000; // 2244 : 128 - 0x80
      12'h8C5: dout  = 8'b01111111; // 2245 : 127 - 0x7f
      12'h8C6: dout  = 8'b00000001; // 2246 :   1 - 0x1
      12'h8C7: dout  = 8'b01111111; // 2247 : 127 - 0x7f
      12'h8C8: dout  = 8'b11111100; // 2248 : 252 - 0xfc -- Background 0x19
      12'h8C9: dout  = 8'b00000010; // 2249 :   2 - 0x2
      12'h8CA: dout  = 8'b00000010; // 2250 :   2 - 0x2
      12'h8CB: dout  = 8'b00000001; // 2251 :   1 - 0x1
      12'h8CC: dout  = 8'b00000001; // 2252 :   1 - 0x1
      12'h8CD: dout  = 8'b11111110; // 2253 : 254 - 0xfe
      12'h8CE: dout  = 8'b10000000; // 2254 : 128 - 0x80
      12'h8CF: dout  = 8'b11111110; // 2255 : 254 - 0xfe
      12'h8D0: dout  = 8'b00000000; // 2256 :   0 - 0x0 -- Background 0x1a
      12'h8D1: dout  = 8'b00000000; // 2257 :   0 - 0x0
      12'h8D2: dout  = 8'b00111111; // 2258 :  63 - 0x3f
      12'h8D3: dout  = 8'b01000000; // 2259 :  64 - 0x40
      12'h8D4: dout  = 8'b01000000; // 2260 :  64 - 0x40
      12'h8D5: dout  = 8'b10000000; // 2261 : 128 - 0x80
      12'h8D6: dout  = 8'b10000000; // 2262 : 128 - 0x80
      12'h8D7: dout  = 8'b01111111; // 2263 : 127 - 0x7f
      12'h8D8: dout  = 8'b00000000; // 2264 :   0 - 0x0 -- Background 0x1b
      12'h8D9: dout  = 8'b00000000; // 2265 :   0 - 0x0
      12'h8DA: dout  = 8'b11111100; // 2266 : 252 - 0xfc
      12'h8DB: dout  = 8'b00000010; // 2267 :   2 - 0x2
      12'h8DC: dout  = 8'b00000010; // 2268 :   2 - 0x2
      12'h8DD: dout  = 8'b00000001; // 2269 :   1 - 0x1
      12'h8DE: dout  = 8'b00000001; // 2270 :   1 - 0x1
      12'h8DF: dout  = 8'b11111110; // 2271 : 254 - 0xfe
      12'h8E0: dout  = 8'b01111111; // 2272 : 127 - 0x7f -- Background 0x1c
      12'h8E1: dout  = 8'b10000000; // 2273 : 128 - 0x80
      12'h8E2: dout  = 8'b10000000; // 2274 : 128 - 0x80
      12'h8E3: dout  = 8'b10000000; // 2275 : 128 - 0x80
      12'h8E4: dout  = 8'b10011011; // 2276 : 155 - 0x9b
      12'h8E5: dout  = 8'b10100100; // 2277 : 164 - 0xa4
      12'h8E6: dout  = 8'b10100110; // 2278 : 166 - 0xa6
      12'h8E7: dout  = 8'b10000000; // 2279 : 128 - 0x80
      12'h8E8: dout  = 8'b10000000; // 2280 : 128 - 0x80 -- Background 0x1d
      12'h8E9: dout  = 8'b01111111; // 2281 : 127 - 0x7f
      12'h8EA: dout  = 8'b00000010; // 2282 :   2 - 0x2
      12'h8EB: dout  = 8'b00000010; // 2283 :   2 - 0x2
      12'h8EC: dout  = 8'b00000010; // 2284 :   2 - 0x2
      12'h8ED: dout  = 8'b00000010; // 2285 :   2 - 0x2
      12'h8EE: dout  = 8'b00000010; // 2286 :   2 - 0x2
      12'h8EF: dout  = 8'b00001111; // 2287 :  15 - 0xf
      12'h8F0: dout  = 8'b11111110; // 2288 : 254 - 0xfe -- Background 0x1e
      12'h8F1: dout  = 8'b00000001; // 2289 :   1 - 0x1
      12'h8F2: dout  = 8'b00000001; // 2290 :   1 - 0x1
      12'h8F3: dout  = 8'b00000001; // 2291 :   1 - 0x1
      12'h8F4: dout  = 8'b01000001; // 2292 :  65 - 0x41
      12'h8F5: dout  = 8'b11110101; // 2293 : 245 - 0xf5
      12'h8F6: dout  = 8'b00011101; // 2294 :  29 - 0x1d
      12'h8F7: dout  = 8'b00000001; // 2295 :   1 - 0x1
      12'h8F8: dout  = 8'b00000001; // 2296 :   1 - 0x1 -- Background 0x1f
      12'h8F9: dout  = 8'b11111110; // 2297 : 254 - 0xfe
      12'h8FA: dout  = 8'b01000000; // 2298 :  64 - 0x40
      12'h8FB: dout  = 8'b01000000; // 2299 :  64 - 0x40
      12'h8FC: dout  = 8'b01000000; // 2300 :  64 - 0x40
      12'h8FD: dout  = 8'b01000000; // 2301 :  64 - 0x40
      12'h8FE: dout  = 8'b01000000; // 2302 :  64 - 0x40
      12'h8FF: dout  = 8'b11110000; // 2303 : 240 - 0xf0
      12'h900: dout  = 8'b00000111; // 2304 :   7 - 0x7 -- Background 0x20
      12'h901: dout  = 8'b00011111; // 2305 :  31 - 0x1f
      12'h902: dout  = 8'b00111111; // 2306 :  63 - 0x3f
      12'h903: dout  = 8'b01111111; // 2307 : 127 - 0x7f
      12'h904: dout  = 8'b01111111; // 2308 : 127 - 0x7f
      12'h905: dout  = 8'b11111111; // 2309 : 255 - 0xff
      12'h906: dout  = 8'b11111111; // 2310 : 255 - 0xff
      12'h907: dout  = 8'b11111111; // 2311 : 255 - 0xff
      12'h908: dout  = 8'b11100000; // 2312 : 224 - 0xe0 -- Background 0x21
      12'h909: dout  = 8'b11111000; // 2313 : 248 - 0xf8
      12'h90A: dout  = 8'b11111100; // 2314 : 252 - 0xfc
      12'h90B: dout  = 8'b11111110; // 2315 : 254 - 0xfe
      12'h90C: dout  = 8'b11111110; // 2316 : 254 - 0xfe
      12'h90D: dout  = 8'b11111111; // 2317 : 255 - 0xff
      12'h90E: dout  = 8'b11111111; // 2318 : 255 - 0xff
      12'h90F: dout  = 8'b11111111; // 2319 : 255 - 0xff
      12'h910: dout  = 8'b00000111; // 2320 :   7 - 0x7 -- Background 0x22
      12'h911: dout  = 8'b00011111; // 2321 :  31 - 0x1f
      12'h912: dout  = 8'b00111111; // 2322 :  63 - 0x3f
      12'h913: dout  = 8'b01111111; // 2323 : 127 - 0x7f
      12'h914: dout  = 8'b01111111; // 2324 : 127 - 0x7f
      12'h915: dout  = 8'b11111111; // 2325 : 255 - 0xff
      12'h916: dout  = 8'b11111111; // 2326 : 255 - 0xff
      12'h917: dout  = 8'b11111111; // 2327 : 255 - 0xff
      12'h918: dout  = 8'b11100000; // 2328 : 224 - 0xe0 -- Background 0x23
      12'h919: dout  = 8'b11111000; // 2329 : 248 - 0xf8
      12'h91A: dout  = 8'b11111100; // 2330 : 252 - 0xfc
      12'h91B: dout  = 8'b11111110; // 2331 : 254 - 0xfe
      12'h91C: dout  = 8'b11111110; // 2332 : 254 - 0xfe
      12'h91D: dout  = 8'b11111111; // 2333 : 255 - 0xff
      12'h91E: dout  = 8'b11111111; // 2334 : 255 - 0xff
      12'h91F: dout  = 8'b11111111; // 2335 : 255 - 0xff
      12'h920: dout  = 8'b00000000; // 2336 :   0 - 0x0 -- Background 0x24
      12'h921: dout  = 8'b00000000; // 2337 :   0 - 0x0
      12'h922: dout  = 8'b00000000; // 2338 :   0 - 0x0
      12'h923: dout  = 8'b00000000; // 2339 :   0 - 0x0
      12'h924: dout  = 8'b00000000; // 2340 :   0 - 0x0
      12'h925: dout  = 8'b00000000; // 2341 :   0 - 0x0
      12'h926: dout  = 8'b00000000; // 2342 :   0 - 0x0
      12'h927: dout  = 8'b00000000; // 2343 :   0 - 0x0
      12'h928: dout  = 8'b00101111; // 2344 :  47 - 0x2f -- Background 0x25
      12'h929: dout  = 8'b01001111; // 2345 :  79 - 0x4f
      12'h92A: dout  = 8'b01001111; // 2346 :  79 - 0x4f
      12'h92B: dout  = 8'b01001111; // 2347 :  79 - 0x4f
      12'h92C: dout  = 8'b01001111; // 2348 :  79 - 0x4f
      12'h92D: dout  = 8'b00100111; // 2349 :  39 - 0x27
      12'h92E: dout  = 8'b00010000; // 2350 :  16 - 0x10
      12'h92F: dout  = 8'b00001111; // 2351 :  15 - 0xf
      12'h930: dout  = 8'b00000000; // 2352 :   0 - 0x0 -- Background 0x26
      12'h931: dout  = 8'b11100000; // 2353 : 224 - 0xe0
      12'h932: dout  = 8'b10100000; // 2354 : 160 - 0xa0
      12'h933: dout  = 8'b00100000; // 2355 :  32 - 0x20
      12'h934: dout  = 8'b11000000; // 2356 : 192 - 0xc0
      12'h935: dout  = 8'b01000000; // 2357 :  64 - 0x40
      12'h936: dout  = 8'b00110000; // 2358 :  48 - 0x30
      12'h937: dout  = 8'b11101000; // 2359 : 232 - 0xe8
      12'h938: dout  = 8'b11110100; // 2360 : 244 - 0xf4 -- Background 0x27
      12'h939: dout  = 8'b11110010; // 2361 : 242 - 0xf2
      12'h93A: dout  = 8'b11110010; // 2362 : 242 - 0xf2
      12'h93B: dout  = 8'b11110010; // 2363 : 242 - 0xf2
      12'h93C: dout  = 8'b11110010; // 2364 : 242 - 0xf2
      12'h93D: dout  = 8'b11100100; // 2365 : 228 - 0xe4
      12'h93E: dout  = 8'b00001000; // 2366 :   8 - 0x8
      12'h93F: dout  = 8'b11110000; // 2367 : 240 - 0xf0
      12'h940: dout  = 8'b11111111; // 2368 : 255 - 0xff -- Background 0x28
      12'h941: dout  = 8'b11010101; // 2369 : 213 - 0xd5
      12'h942: dout  = 8'b10100011; // 2370 : 163 - 0xa3
      12'h943: dout  = 8'b11010111; // 2371 : 215 - 0xd7
      12'h944: dout  = 8'b10001111; // 2372 : 143 - 0x8f
      12'h945: dout  = 8'b11001111; // 2373 : 207 - 0xcf
      12'h946: dout  = 8'b10001011; // 2374 : 139 - 0x8b
      12'h947: dout  = 8'b11001011; // 2375 : 203 - 0xcb
      12'h948: dout  = 8'b10001111; // 2376 : 143 - 0x8f -- Background 0x29
      12'h949: dout  = 8'b11001111; // 2377 : 207 - 0xcf
      12'h94A: dout  = 8'b10001111; // 2378 : 143 - 0x8f
      12'h94B: dout  = 8'b11001111; // 2379 : 207 - 0xcf
      12'h94C: dout  = 8'b10010000; // 2380 : 144 - 0x90
      12'h94D: dout  = 8'b11100000; // 2381 : 224 - 0xe0
      12'h94E: dout  = 8'b11101010; // 2382 : 234 - 0xea
      12'h94F: dout  = 8'b11111111; // 2383 : 255 - 0xff
      12'h950: dout  = 8'b11111111; // 2384 : 255 - 0xff -- Background 0x2a
      12'h951: dout  = 8'b11011011; // 2385 : 219 - 0xdb
      12'h952: dout  = 8'b11000111; // 2386 : 199 - 0xc7
      12'h953: dout  = 8'b11101001; // 2387 : 233 - 0xe9
      12'h954: dout  = 8'b11110011; // 2388 : 243 - 0xf3
      12'h955: dout  = 8'b11110001; // 2389 : 241 - 0xf1
      12'h956: dout  = 8'b11010011; // 2390 : 211 - 0xd3
      12'h957: dout  = 8'b11010001; // 2391 : 209 - 0xd1
      12'h958: dout  = 8'b11110011; // 2392 : 243 - 0xf3 -- Background 0x2b
      12'h959: dout  = 8'b11110001; // 2393 : 241 - 0xf1
      12'h95A: dout  = 8'b11110011; // 2394 : 243 - 0xf3
      12'h95B: dout  = 8'b11110001; // 2395 : 241 - 0xf1
      12'h95C: dout  = 8'b00001011; // 2396 :  11 - 0xb
      12'h95D: dout  = 8'b00000101; // 2397 :   5 - 0x5
      12'h95E: dout  = 8'b10101011; // 2398 : 171 - 0xab
      12'h95F: dout  = 8'b11111111; // 2399 : 255 - 0xff
      12'h960: dout  = 8'b00000000; // 2400 :   0 - 0x0 -- Background 0x2c
      12'h961: dout  = 8'b00000000; // 2401 :   0 - 0x0
      12'h962: dout  = 8'b00000000; // 2402 :   0 - 0x0
      12'h963: dout  = 8'b00000000; // 2403 :   0 - 0x0
      12'h964: dout  = 8'b00000000; // 2404 :   0 - 0x0
      12'h965: dout  = 8'b00000000; // 2405 :   0 - 0x0
      12'h966: dout  = 8'b00000000; // 2406 :   0 - 0x0
      12'h967: dout  = 8'b00000000; // 2407 :   0 - 0x0
      12'h968: dout  = 8'b00101111; // 2408 :  47 - 0x2f -- Background 0x2d
      12'h969: dout  = 8'b01001111; // 2409 :  79 - 0x4f
      12'h96A: dout  = 8'b01001111; // 2410 :  79 - 0x4f
      12'h96B: dout  = 8'b01001111; // 2411 :  79 - 0x4f
      12'h96C: dout  = 8'b01001111; // 2412 :  79 - 0x4f
      12'h96D: dout  = 8'b00100111; // 2413 :  39 - 0x27
      12'h96E: dout  = 8'b00010000; // 2414 :  16 - 0x10
      12'h96F: dout  = 8'b00001111; // 2415 :  15 - 0xf
      12'h970: dout  = 8'b00000000; // 2416 :   0 - 0x0 -- Background 0x2e
      12'h971: dout  = 8'b00000000; // 2417 :   0 - 0x0
      12'h972: dout  = 8'b00000000; // 2418 :   0 - 0x0
      12'h973: dout  = 8'b00000000; // 2419 :   0 - 0x0
      12'h974: dout  = 8'b00000000; // 2420 :   0 - 0x0
      12'h975: dout  = 8'b00000000; // 2421 :   0 - 0x0
      12'h976: dout  = 8'b00000000; // 2422 :   0 - 0x0
      12'h977: dout  = 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout  = 8'b11110100; // 2424 : 244 - 0xf4 -- Background 0x2f
      12'h979: dout  = 8'b11110010; // 2425 : 242 - 0xf2
      12'h97A: dout  = 8'b11110010; // 2426 : 242 - 0xf2
      12'h97B: dout  = 8'b11110010; // 2427 : 242 - 0xf2
      12'h97C: dout  = 8'b11110010; // 2428 : 242 - 0xf2
      12'h97D: dout  = 8'b11100100; // 2429 : 228 - 0xe4
      12'h97E: dout  = 8'b00001000; // 2430 :   8 - 0x8
      12'h97F: dout  = 8'b11110000; // 2431 : 240 - 0xf0
      12'h980: dout  = 8'b00011000; // 2432 :  24 - 0x18 -- Background 0x30
      12'h981: dout  = 8'b00100100; // 2433 :  36 - 0x24
      12'h982: dout  = 8'b01000010; // 2434 :  66 - 0x42
      12'h983: dout  = 8'b10100101; // 2435 : 165 - 0xa5
      12'h984: dout  = 8'b11100111; // 2436 : 231 - 0xe7
      12'h985: dout  = 8'b00100100; // 2437 :  36 - 0x24
      12'h986: dout  = 8'b00100100; // 2438 :  36 - 0x24
      12'h987: dout  = 8'b00111100; // 2439 :  60 - 0x3c
      12'h988: dout  = 8'b00111100; // 2440 :  60 - 0x3c -- Background 0x31
      12'h989: dout  = 8'b00100100; // 2441 :  36 - 0x24
      12'h98A: dout  = 8'b00100100; // 2442 :  36 - 0x24
      12'h98B: dout  = 8'b01100110; // 2443 : 102 - 0x66
      12'h98C: dout  = 8'b10100101; // 2444 : 165 - 0xa5
      12'h98D: dout  = 8'b01000010; // 2445 :  66 - 0x42
      12'h98E: dout  = 8'b00100100; // 2446 :  36 - 0x24
      12'h98F: dout  = 8'b00011000; // 2447 :  24 - 0x18
      12'h990: dout  = 8'b00000010; // 2448 :   2 - 0x2 -- Background 0x32
      12'h991: dout  = 8'b00000010; // 2449 :   2 - 0x2
      12'h992: dout  = 8'b00000011; // 2450 :   3 - 0x3
      12'h993: dout  = 8'b00000010; // 2451 :   2 - 0x2
      12'h994: dout  = 8'b00000010; // 2452 :   2 - 0x2
      12'h995: dout  = 8'b00000010; // 2453 :   2 - 0x2
      12'h996: dout  = 8'b00000011; // 2454 :   3 - 0x3
      12'h997: dout  = 8'b00000010; // 2455 :   2 - 0x2
      12'h998: dout  = 8'b01000000; // 2456 :  64 - 0x40 -- Background 0x33
      12'h999: dout  = 8'b11000000; // 2457 : 192 - 0xc0
      12'h99A: dout  = 8'b01000000; // 2458 :  64 - 0x40
      12'h99B: dout  = 8'b01000000; // 2459 :  64 - 0x40
      12'h99C: dout  = 8'b01000000; // 2460 :  64 - 0x40
      12'h99D: dout  = 8'b11000000; // 2461 : 192 - 0xc0
      12'h99E: dout  = 8'b01000000; // 2462 :  64 - 0x40
      12'h99F: dout  = 8'b01000000; // 2463 :  64 - 0x40
      12'h9A0: dout  = 8'b00000000; // 2464 :   0 - 0x0 -- Background 0x34
      12'h9A1: dout  = 8'b00011000; // 2465 :  24 - 0x18
      12'h9A2: dout  = 8'b00111100; // 2466 :  60 - 0x3c
      12'h9A3: dout  = 8'b01100010; // 2467 :  98 - 0x62
      12'h9A4: dout  = 8'b01100001; // 2468 :  97 - 0x61
      12'h9A5: dout  = 8'b11000000; // 2469 : 192 - 0xc0
      12'h9A6: dout  = 8'b11000000; // 2470 : 192 - 0xc0
      12'h9A7: dout  = 8'b11000000; // 2471 : 192 - 0xc0
      12'h9A8: dout  = 8'b01100000; // 2472 :  96 - 0x60 -- Background 0x35
      12'h9A9: dout  = 8'b01100000; // 2473 :  96 - 0x60
      12'h9AA: dout  = 8'b00110000; // 2474 :  48 - 0x30
      12'h9AB: dout  = 8'b00011000; // 2475 :  24 - 0x18
      12'h9AC: dout  = 8'b00001100; // 2476 :  12 - 0xc
      12'h9AD: dout  = 8'b00000110; // 2477 :   6 - 0x6
      12'h9AE: dout  = 8'b00000010; // 2478 :   2 - 0x2
      12'h9AF: dout  = 8'b00000001; // 2479 :   1 - 0x1
      12'h9B0: dout  = 8'b00000000; // 2480 :   0 - 0x0 -- Background 0x36
      12'h9B1: dout  = 8'b00011000; // 2481 :  24 - 0x18
      12'h9B2: dout  = 8'b00100100; // 2482 :  36 - 0x24
      12'h9B3: dout  = 8'b01000010; // 2483 :  66 - 0x42
      12'h9B4: dout  = 8'b10000010; // 2484 : 130 - 0x82
      12'h9B5: dout  = 8'b00000001; // 2485 :   1 - 0x1
      12'h9B6: dout  = 8'b00000001; // 2486 :   1 - 0x1
      12'h9B7: dout  = 8'b00000001; // 2487 :   1 - 0x1
      12'h9B8: dout  = 8'b00000010; // 2488 :   2 - 0x2 -- Background 0x37
      12'h9B9: dout  = 8'b00000010; // 2489 :   2 - 0x2
      12'h9BA: dout  = 8'b00000100; // 2490 :   4 - 0x4
      12'h9BB: dout  = 8'b00001000; // 2491 :   8 - 0x8
      12'h9BC: dout  = 8'b00010000; // 2492 :  16 - 0x10
      12'h9BD: dout  = 8'b00100000; // 2493 :  32 - 0x20
      12'h9BE: dout  = 8'b01000000; // 2494 :  64 - 0x40
      12'h9BF: dout  = 8'b10000000; // 2495 : 128 - 0x80
      12'h9C0: dout  = 8'b00000000; // 2496 :   0 - 0x0 -- Background 0x38
      12'h9C1: dout  = 8'b00000110; // 2497 :   6 - 0x6
      12'h9C2: dout  = 8'b00001101; // 2498 :  13 - 0xd
      12'h9C3: dout  = 8'b00001100; // 2499 :  12 - 0xc
      12'h9C4: dout  = 8'b00001100; // 2500 :  12 - 0xc
      12'h9C5: dout  = 8'b00000110; // 2501 :   6 - 0x6
      12'h9C6: dout  = 8'b00000010; // 2502 :   2 - 0x2
      12'h9C7: dout  = 8'b00000001; // 2503 :   1 - 0x1
      12'h9C8: dout  = 8'b11111111; // 2504 : 255 - 0xff -- Background 0x39
      12'h9C9: dout  = 8'b00000000; // 2505 :   0 - 0x0
      12'h9CA: dout  = 8'b00000000; // 2506 :   0 - 0x0
      12'h9CB: dout  = 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout  = 8'b00000000; // 2508 :   0 - 0x0
      12'h9CD: dout  = 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout  = 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout  = 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout  = 8'b00000000; // 2512 :   0 - 0x0 -- Background 0x3a
      12'h9D1: dout  = 8'b01100000; // 2513 :  96 - 0x60
      12'h9D2: dout  = 8'b10010000; // 2514 : 144 - 0x90
      12'h9D3: dout  = 8'b00010000; // 2515 :  16 - 0x10
      12'h9D4: dout  = 8'b00010000; // 2516 :  16 - 0x10
      12'h9D5: dout  = 8'b00100000; // 2517 :  32 - 0x20
      12'h9D6: dout  = 8'b01000000; // 2518 :  64 - 0x40
      12'h9D7: dout  = 8'b10000000; // 2519 : 128 - 0x80
      12'h9D8: dout  = 8'b00000000; // 2520 :   0 - 0x0 -- Background 0x3b
      12'h9D9: dout  = 8'b01010100; // 2521 :  84 - 0x54
      12'h9DA: dout  = 8'b00000010; // 2522 :   2 - 0x2
      12'h9DB: dout  = 8'b01000000; // 2523 :  64 - 0x40
      12'h9DC: dout  = 8'b00000010; // 2524 :   2 - 0x2
      12'h9DD: dout  = 8'b01000000; // 2525 :  64 - 0x40
      12'h9DE: dout  = 8'b00101010; // 2526 :  42 - 0x2a
      12'h9DF: dout  = 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout  = 8'b11111111; // 2528 : 255 - 0xff -- Background 0x3c
      12'h9E1: dout  = 8'b11111111; // 2529 : 255 - 0xff
      12'h9E2: dout  = 8'b11111111; // 2530 : 255 - 0xff
      12'h9E3: dout  = 8'b11111111; // 2531 : 255 - 0xff
      12'h9E4: dout  = 8'b11111111; // 2532 : 255 - 0xff
      12'h9E5: dout  = 8'b11111111; // 2533 : 255 - 0xff
      12'h9E6: dout  = 8'b11111111; // 2534 : 255 - 0xff
      12'h9E7: dout  = 8'b11111111; // 2535 : 255 - 0xff
      12'h9E8: dout  = 8'b00000000; // 2536 :   0 - 0x0 -- Background 0x3d
      12'h9E9: dout  = 8'b00000000; // 2537 :   0 - 0x0
      12'h9EA: dout  = 8'b00000000; // 2538 :   0 - 0x0
      12'h9EB: dout  = 8'b00000000; // 2539 :   0 - 0x0
      12'h9EC: dout  = 8'b00000000; // 2540 :   0 - 0x0
      12'h9ED: dout  = 8'b00000000; // 2541 :   0 - 0x0
      12'h9EE: dout  = 8'b00000000; // 2542 :   0 - 0x0
      12'h9EF: dout  = 8'b00000000; // 2543 :   0 - 0x0
      12'h9F0: dout  = 8'b11111111; // 2544 : 255 - 0xff -- Background 0x3e
      12'h9F1: dout  = 8'b11111111; // 2545 : 255 - 0xff
      12'h9F2: dout  = 8'b11111111; // 2546 : 255 - 0xff
      12'h9F3: dout  = 8'b11111111; // 2547 : 255 - 0xff
      12'h9F4: dout  = 8'b11111111; // 2548 : 255 - 0xff
      12'h9F5: dout  = 8'b11111111; // 2549 : 255 - 0xff
      12'h9F6: dout  = 8'b11111111; // 2550 : 255 - 0xff
      12'h9F7: dout  = 8'b11111111; // 2551 : 255 - 0xff
      12'h9F8: dout  = 8'b00000000; // 2552 :   0 - 0x0 -- Background 0x3f
      12'h9F9: dout  = 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout  = 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout  = 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout  = 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout  = 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout  = 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout  = 8'b00111100; // 2560 :  60 - 0x3c -- Background 0x40
      12'hA01: dout  = 8'b01000010; // 2561 :  66 - 0x42
      12'hA02: dout  = 8'b10011001; // 2562 : 153 - 0x99
      12'hA03: dout  = 8'b10100101; // 2563 : 165 - 0xa5
      12'hA04: dout  = 8'b10100101; // 2564 : 165 - 0xa5
      12'hA05: dout  = 8'b10011010; // 2565 : 154 - 0x9a
      12'hA06: dout  = 8'b01000000; // 2566 :  64 - 0x40
      12'hA07: dout  = 8'b00111100; // 2567 :  60 - 0x3c
      12'hA08: dout  = 8'b00001100; // 2568 :  12 - 0xc -- Background 0x41
      12'hA09: dout  = 8'b00010010; // 2569 :  18 - 0x12
      12'hA0A: dout  = 8'b00100010; // 2570 :  34 - 0x22
      12'hA0B: dout  = 8'b00100010; // 2571 :  34 - 0x22
      12'hA0C: dout  = 8'b01111110; // 2572 : 126 - 0x7e
      12'hA0D: dout  = 8'b00100010; // 2573 :  34 - 0x22
      12'hA0E: dout  = 8'b00100100; // 2574 :  36 - 0x24
      12'hA0F: dout  = 8'b00000000; // 2575 :   0 - 0x0
      12'hA10: dout  = 8'b00111100; // 2576 :  60 - 0x3c -- Background 0x42
      12'hA11: dout  = 8'b01000010; // 2577 :  66 - 0x42
      12'hA12: dout  = 8'b01010010; // 2578 :  82 - 0x52
      12'hA13: dout  = 8'b00011100; // 2579 :  28 - 0x1c
      12'hA14: dout  = 8'b00010010; // 2580 :  18 - 0x12
      12'hA15: dout  = 8'b00110010; // 2581 :  50 - 0x32
      12'hA16: dout  = 8'b00011100; // 2582 :  28 - 0x1c
      12'hA17: dout  = 8'b00000000; // 2583 :   0 - 0x0
      12'hA18: dout  = 8'b00011000; // 2584 :  24 - 0x18 -- Background 0x43
      12'hA19: dout  = 8'b00100100; // 2585 :  36 - 0x24
      12'hA1A: dout  = 8'b01010100; // 2586 :  84 - 0x54
      12'hA1B: dout  = 8'b01001000; // 2587 :  72 - 0x48
      12'hA1C: dout  = 8'b01000010; // 2588 :  66 - 0x42
      12'hA1D: dout  = 8'b00100100; // 2589 :  36 - 0x24
      12'hA1E: dout  = 8'b00011000; // 2590 :  24 - 0x18
      12'hA1F: dout  = 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout  = 8'b01011000; // 2592 :  88 - 0x58 -- Background 0x44
      12'hA21: dout  = 8'b11100100; // 2593 : 228 - 0xe4
      12'hA22: dout  = 8'b01000010; // 2594 :  66 - 0x42
      12'hA23: dout  = 8'b01000010; // 2595 :  66 - 0x42
      12'hA24: dout  = 8'b00100010; // 2596 :  34 - 0x22
      12'hA25: dout  = 8'b01100100; // 2597 : 100 - 0x64
      12'hA26: dout  = 8'b00111000; // 2598 :  56 - 0x38
      12'hA27: dout  = 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout  = 8'b00011100; // 2600 :  28 - 0x1c -- Background 0x45
      12'hA29: dout  = 8'b00100000; // 2601 :  32 - 0x20
      12'hA2A: dout  = 8'b00100000; // 2602 :  32 - 0x20
      12'hA2B: dout  = 8'b00101100; // 2603 :  44 - 0x2c
      12'hA2C: dout  = 8'b01110000; // 2604 : 112 - 0x70
      12'hA2D: dout  = 8'b00100010; // 2605 :  34 - 0x22
      12'hA2E: dout  = 8'b00011100; // 2606 :  28 - 0x1c
      12'hA2F: dout  = 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout  = 8'b00011100; // 2608 :  28 - 0x1c -- Background 0x46
      12'hA31: dout  = 8'b00100000; // 2609 :  32 - 0x20
      12'hA32: dout  = 8'b00100000; // 2610 :  32 - 0x20
      12'hA33: dout  = 8'b00101100; // 2611 :  44 - 0x2c
      12'hA34: dout  = 8'b01110000; // 2612 : 112 - 0x70
      12'hA35: dout  = 8'b00010000; // 2613 :  16 - 0x10
      12'hA36: dout  = 8'b00010000; // 2614 :  16 - 0x10
      12'hA37: dout  = 8'b00000000; // 2615 :   0 - 0x0
      12'hA38: dout  = 8'b00011000; // 2616 :  24 - 0x18 -- Background 0x47
      12'hA39: dout  = 8'b00100100; // 2617 :  36 - 0x24
      12'hA3A: dout  = 8'b01000000; // 2618 :  64 - 0x40
      12'hA3B: dout  = 8'b01001110; // 2619 :  78 - 0x4e
      12'hA3C: dout  = 8'b01000010; // 2620 :  66 - 0x42
      12'hA3D: dout  = 8'b00100100; // 2621 :  36 - 0x24
      12'hA3E: dout  = 8'b00011000; // 2622 :  24 - 0x18
      12'hA3F: dout  = 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout  = 8'b00100000; // 2624 :  32 - 0x20 -- Background 0x48
      12'hA41: dout  = 8'b01000100; // 2625 :  68 - 0x44
      12'hA42: dout  = 8'b01000100; // 2626 :  68 - 0x44
      12'hA43: dout  = 8'b01000100; // 2627 :  68 - 0x44
      12'hA44: dout  = 8'b11111100; // 2628 : 252 - 0xfc
      12'hA45: dout  = 8'b01000100; // 2629 :  68 - 0x44
      12'hA46: dout  = 8'b01001000; // 2630 :  72 - 0x48
      12'hA47: dout  = 8'b00000000; // 2631 :   0 - 0x0
      12'hA48: dout  = 8'b00010000; // 2632 :  16 - 0x10 -- Background 0x49
      12'hA49: dout  = 8'b00010000; // 2633 :  16 - 0x10
      12'hA4A: dout  = 8'b00010000; // 2634 :  16 - 0x10
      12'hA4B: dout  = 8'b00010000; // 2635 :  16 - 0x10
      12'hA4C: dout  = 8'b00010000; // 2636 :  16 - 0x10
      12'hA4D: dout  = 8'b00001000; // 2637 :   8 - 0x8
      12'hA4E: dout  = 8'b00001000; // 2638 :   8 - 0x8
      12'hA4F: dout  = 8'b00000000; // 2639 :   0 - 0x0
      12'hA50: dout  = 8'b00001000; // 2640 :   8 - 0x8 -- Background 0x4a
      12'hA51: dout  = 8'b00001000; // 2641 :   8 - 0x8
      12'hA52: dout  = 8'b00000100; // 2642 :   4 - 0x4
      12'hA53: dout  = 8'b00000100; // 2643 :   4 - 0x4
      12'hA54: dout  = 8'b01000100; // 2644 :  68 - 0x44
      12'hA55: dout  = 8'b01001000; // 2645 :  72 - 0x48
      12'hA56: dout  = 8'b00110000; // 2646 :  48 - 0x30
      12'hA57: dout  = 8'b00000000; // 2647 :   0 - 0x0
      12'hA58: dout  = 8'b01000100; // 2648 :  68 - 0x44 -- Background 0x4b
      12'hA59: dout  = 8'b01000100; // 2649 :  68 - 0x44
      12'hA5A: dout  = 8'b01001000; // 2650 :  72 - 0x48
      12'hA5B: dout  = 8'b01110000; // 2651 : 112 - 0x70
      12'hA5C: dout  = 8'b01001000; // 2652 :  72 - 0x48
      12'hA5D: dout  = 8'b00100100; // 2653 :  36 - 0x24
      12'hA5E: dout  = 8'b00100010; // 2654 :  34 - 0x22
      12'hA5F: dout  = 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout  = 8'b00010000; // 2656 :  16 - 0x10 -- Background 0x4c
      12'hA61: dout  = 8'b00100000; // 2657 :  32 - 0x20
      12'hA62: dout  = 8'b00100000; // 2658 :  32 - 0x20
      12'hA63: dout  = 8'b00100000; // 2659 :  32 - 0x20
      12'hA64: dout  = 8'b01000000; // 2660 :  64 - 0x40
      12'hA65: dout  = 8'b01000000; // 2661 :  64 - 0x40
      12'hA66: dout  = 8'b01000110; // 2662 :  70 - 0x46
      12'hA67: dout  = 8'b00111000; // 2663 :  56 - 0x38
      12'hA68: dout  = 8'b00100100; // 2664 :  36 - 0x24 -- Background 0x4d
      12'hA69: dout  = 8'b01011010; // 2665 :  90 - 0x5a
      12'hA6A: dout  = 8'b01011010; // 2666 :  90 - 0x5a
      12'hA6B: dout  = 8'b01011010; // 2667 :  90 - 0x5a
      12'hA6C: dout  = 8'b01000010; // 2668 :  66 - 0x42
      12'hA6D: dout  = 8'b01000010; // 2669 :  66 - 0x42
      12'hA6E: dout  = 8'b00100010; // 2670 :  34 - 0x22
      12'hA6F: dout  = 8'b00000000; // 2671 :   0 - 0x0
      12'hA70: dout  = 8'b00100100; // 2672 :  36 - 0x24 -- Background 0x4e
      12'hA71: dout  = 8'b01010010; // 2673 :  82 - 0x52
      12'hA72: dout  = 8'b01010010; // 2674 :  82 - 0x52
      12'hA73: dout  = 8'b01010010; // 2675 :  82 - 0x52
      12'hA74: dout  = 8'b01010010; // 2676 :  82 - 0x52
      12'hA75: dout  = 8'b01010010; // 2677 :  82 - 0x52
      12'hA76: dout  = 8'b01001100; // 2678 :  76 - 0x4c
      12'hA77: dout  = 8'b00000000; // 2679 :   0 - 0x0
      12'hA78: dout  = 8'b00111000; // 2680 :  56 - 0x38 -- Background 0x4f
      12'hA79: dout  = 8'b01000100; // 2681 :  68 - 0x44
      12'hA7A: dout  = 8'b10000010; // 2682 : 130 - 0x82
      12'hA7B: dout  = 8'b10000010; // 2683 : 130 - 0x82
      12'hA7C: dout  = 8'b10000010; // 2684 : 130 - 0x82
      12'hA7D: dout  = 8'b01000100; // 2685 :  68 - 0x44
      12'hA7E: dout  = 8'b00111000; // 2686 :  56 - 0x38
      12'hA7F: dout  = 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout  = 8'b01111111; // 2688 : 127 - 0x7f -- Background 0x50
      12'hA81: dout  = 8'b11000000; // 2689 : 192 - 0xc0
      12'hA82: dout  = 8'b10000000; // 2690 : 128 - 0x80
      12'hA83: dout  = 8'b10000000; // 2691 : 128 - 0x80
      12'hA84: dout  = 8'b10000000; // 2692 : 128 - 0x80
      12'hA85: dout  = 8'b11000011; // 2693 : 195 - 0xc3
      12'hA86: dout  = 8'b11111111; // 2694 : 255 - 0xff
      12'hA87: dout  = 8'b11111111; // 2695 : 255 - 0xff
      12'hA88: dout  = 8'b11111110; // 2696 : 254 - 0xfe -- Background 0x51
      12'hA89: dout  = 8'b00000011; // 2697 :   3 - 0x3
      12'hA8A: dout  = 8'b00000001; // 2698 :   1 - 0x1
      12'hA8B: dout  = 8'b00000001; // 2699 :   1 - 0x1
      12'hA8C: dout  = 8'b00000001; // 2700 :   1 - 0x1
      12'hA8D: dout  = 8'b11000011; // 2701 : 195 - 0xc3
      12'hA8E: dout  = 8'b11111111; // 2702 : 255 - 0xff
      12'hA8F: dout  = 8'b11111111; // 2703 : 255 - 0xff
      12'hA90: dout  = 8'b00000000; // 2704 :   0 - 0x0 -- Background 0x52
      12'hA91: dout  = 8'b00000111; // 2705 :   7 - 0x7
      12'hA92: dout  = 8'b00001100; // 2706 :  12 - 0xc
      12'hA93: dout  = 8'b00011000; // 2707 :  24 - 0x18
      12'hA94: dout  = 8'b00110000; // 2708 :  48 - 0x30
      12'hA95: dout  = 8'b01100000; // 2709 :  96 - 0x60
      12'hA96: dout  = 8'b01000000; // 2710 :  64 - 0x40
      12'hA97: dout  = 8'b01001111; // 2711 :  79 - 0x4f
      12'hA98: dout  = 8'b00000000; // 2712 :   0 - 0x0 -- Background 0x53
      12'hA99: dout  = 8'b11110000; // 2713 : 240 - 0xf0
      12'hA9A: dout  = 8'b01010000; // 2714 :  80 - 0x50
      12'hA9B: dout  = 8'b01001000; // 2715 :  72 - 0x48
      12'hA9C: dout  = 8'b01001100; // 2716 :  76 - 0x4c
      12'hA9D: dout  = 8'b01000100; // 2717 :  68 - 0x44
      12'hA9E: dout  = 8'b10000010; // 2718 : 130 - 0x82
      12'hA9F: dout  = 8'b10000011; // 2719 : 131 - 0x83
      12'hAA0: dout  = 8'b01111111; // 2720 : 127 - 0x7f -- Background 0x54
      12'hAA1: dout  = 8'b11011110; // 2721 : 222 - 0xde
      12'hAA2: dout  = 8'b10001110; // 2722 : 142 - 0x8e
      12'hAA3: dout  = 8'b11000101; // 2723 : 197 - 0xc5
      12'hAA4: dout  = 8'b10010010; // 2724 : 146 - 0x92
      12'hAA5: dout  = 8'b11000111; // 2725 : 199 - 0xc7
      12'hAA6: dout  = 8'b11100010; // 2726 : 226 - 0xe2
      12'hAA7: dout  = 8'b11010000; // 2727 : 208 - 0xd0
      12'hAA8: dout  = 8'b11111111; // 2728 : 255 - 0xff -- Background 0x55
      12'hAA9: dout  = 8'b11011110; // 2729 : 222 - 0xde
      12'hAAA: dout  = 8'b10001110; // 2730 : 142 - 0x8e
      12'hAAB: dout  = 8'b11000101; // 2731 : 197 - 0xc5
      12'hAAC: dout  = 8'b10010010; // 2732 : 146 - 0x92
      12'hAAD: dout  = 8'b01000111; // 2733 :  71 - 0x47
      12'hAAE: dout  = 8'b11100010; // 2734 : 226 - 0xe2
      12'hAAF: dout  = 8'b01010000; // 2735 :  80 - 0x50
      12'hAB0: dout  = 8'b11111110; // 2736 : 254 - 0xfe -- Background 0x56
      12'hAB1: dout  = 8'b11011111; // 2737 : 223 - 0xdf
      12'hAB2: dout  = 8'b10001111; // 2738 : 143 - 0x8f
      12'hAB3: dout  = 8'b11000101; // 2739 : 197 - 0xc5
      12'hAB4: dout  = 8'b10010011; // 2740 : 147 - 0x93
      12'hAB5: dout  = 8'b01000111; // 2741 :  71 - 0x47
      12'hAB6: dout  = 8'b11100011; // 2742 : 227 - 0xe3
      12'hAB7: dout  = 8'b01010001; // 2743 :  81 - 0x51
      12'hAB8: dout  = 8'b01111111; // 2744 : 127 - 0x7f -- Background 0x57
      12'hAB9: dout  = 8'b10000000; // 2745 : 128 - 0x80
      12'hABA: dout  = 8'b10110011; // 2746 : 179 - 0xb3
      12'hABB: dout  = 8'b01001100; // 2747 :  76 - 0x4c
      12'hABC: dout  = 8'b00111111; // 2748 :  63 - 0x3f
      12'hABD: dout  = 8'b00000011; // 2749 :   3 - 0x3
      12'hABE: dout  = 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout  = 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout  = 8'b11111111; // 2752 : 255 - 0xff -- Background 0x58
      12'hAC1: dout  = 8'b00000000; // 2753 :   0 - 0x0
      12'hAC2: dout  = 8'b00110011; // 2754 :  51 - 0x33
      12'hAC3: dout  = 8'b11001100; // 2755 : 204 - 0xcc
      12'hAC4: dout  = 8'b00110011; // 2756 :  51 - 0x33
      12'hAC5: dout  = 8'b11111111; // 2757 : 255 - 0xff
      12'hAC6: dout  = 8'b00000000; // 2758 :   0 - 0x0
      12'hAC7: dout  = 8'b00000000; // 2759 :   0 - 0x0
      12'hAC8: dout  = 8'b11111110; // 2760 : 254 - 0xfe -- Background 0x59
      12'hAC9: dout  = 8'b00000001; // 2761 :   1 - 0x1
      12'hACA: dout  = 8'b00110011; // 2762 :  51 - 0x33
      12'hACB: dout  = 8'b11001110; // 2763 : 206 - 0xce
      12'hACC: dout  = 8'b00111100; // 2764 :  60 - 0x3c
      12'hACD: dout  = 8'b11000000; // 2765 : 192 - 0xc0
      12'hACE: dout  = 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout  = 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout  = 8'b00000000; // 2768 :   0 - 0x0 -- Background 0x5a
      12'hAD1: dout  = 8'b00000000; // 2769 :   0 - 0x0
      12'hAD2: dout  = 8'b00000000; // 2770 :   0 - 0x0
      12'hAD3: dout  = 8'b00000000; // 2771 :   0 - 0x0
      12'hAD4: dout  = 8'b00000000; // 2772 :   0 - 0x0
      12'hAD5: dout  = 8'b00000000; // 2773 :   0 - 0x0
      12'hAD6: dout  = 8'b00000000; // 2774 :   0 - 0x0
      12'hAD7: dout  = 8'b00000000; // 2775 :   0 - 0x0
      12'hAD8: dout  = 8'b00000000; // 2776 :   0 - 0x0 -- Background 0x5b
      12'hAD9: dout  = 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout  = 8'b00000000; // 2778 :   0 - 0x0
      12'hADB: dout  = 8'b00000001; // 2779 :   1 - 0x1
      12'hADC: dout  = 8'b00000011; // 2780 :   3 - 0x3
      12'hADD: dout  = 8'b00000011; // 2781 :   3 - 0x3
      12'hADE: dout  = 8'b00000111; // 2782 :   7 - 0x7
      12'hADF: dout  = 8'b00111111; // 2783 :  63 - 0x3f
      12'hAE0: dout  = 8'b00000000; // 2784 :   0 - 0x0 -- Background 0x5c
      12'hAE1: dout  = 8'b00000001; // 2785 :   1 - 0x1
      12'hAE2: dout  = 8'b01111111; // 2786 : 127 - 0x7f
      12'hAE3: dout  = 8'b11111111; // 2787 : 255 - 0xff
      12'hAE4: dout  = 8'b11111111; // 2788 : 255 - 0xff
      12'hAE5: dout  = 8'b11111111; // 2789 : 255 - 0xff
      12'hAE6: dout  = 8'b11111111; // 2790 : 255 - 0xff
      12'hAE7: dout  = 8'b11111111; // 2791 : 255 - 0xff
      12'hAE8: dout  = 8'b11111111; // 2792 : 255 - 0xff -- Background 0x5d
      12'hAE9: dout  = 8'b11111111; // 2793 : 255 - 0xff
      12'hAEA: dout  = 8'b11111111; // 2794 : 255 - 0xff
      12'hAEB: dout  = 8'b11111111; // 2795 : 255 - 0xff
      12'hAEC: dout  = 8'b11111111; // 2796 : 255 - 0xff
      12'hAED: dout  = 8'b11111111; // 2797 : 255 - 0xff
      12'hAEE: dout  = 8'b11111111; // 2798 : 255 - 0xff
      12'hAEF: dout  = 8'b11111111; // 2799 : 255 - 0xff
      12'hAF0: dout  = 8'b00000000; // 2800 :   0 - 0x0 -- Background 0x5e
      12'hAF1: dout  = 8'b10000000; // 2801 : 128 - 0x80
      12'hAF2: dout  = 8'b11111110; // 2802 : 254 - 0xfe
      12'hAF3: dout  = 8'b11111111; // 2803 : 255 - 0xff
      12'hAF4: dout  = 8'b11111111; // 2804 : 255 - 0xff
      12'hAF5: dout  = 8'b11111111; // 2805 : 255 - 0xff
      12'hAF6: dout  = 8'b11111111; // 2806 : 255 - 0xff
      12'hAF7: dout  = 8'b11111111; // 2807 : 255 - 0xff
      12'hAF8: dout  = 8'b00000000; // 2808 :   0 - 0x0 -- Background 0x5f
      12'hAF9: dout  = 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout  = 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout  = 8'b10000000; // 2811 : 128 - 0x80
      12'hAFC: dout  = 8'b11000000; // 2812 : 192 - 0xc0
      12'hAFD: dout  = 8'b11000000; // 2813 : 192 - 0xc0
      12'hAFE: dout  = 8'b11100000; // 2814 : 224 - 0xe0
      12'hAFF: dout  = 8'b11111000; // 2815 : 248 - 0xf8
      12'hB00: dout  = 8'b11111111; // 2816 : 255 - 0xff -- Background 0x60
      12'hB01: dout  = 8'b11111111; // 2817 : 255 - 0xff
      12'hB02: dout  = 8'b11111111; // 2818 : 255 - 0xff
      12'hB03: dout  = 8'b11111111; // 2819 : 255 - 0xff
      12'hB04: dout  = 8'b11111111; // 2820 : 255 - 0xff
      12'hB05: dout  = 8'b11111111; // 2821 : 255 - 0xff
      12'hB06: dout  = 8'b11111111; // 2822 : 255 - 0xff
      12'hB07: dout  = 8'b11111111; // 2823 : 255 - 0xff
      12'hB08: dout  = 8'b11111111; // 2824 : 255 - 0xff -- Background 0x61
      12'hB09: dout  = 8'b11111111; // 2825 : 255 - 0xff
      12'hB0A: dout  = 8'b11111111; // 2826 : 255 - 0xff
      12'hB0B: dout  = 8'b11111111; // 2827 : 255 - 0xff
      12'hB0C: dout  = 8'b11111111; // 2828 : 255 - 0xff
      12'hB0D: dout  = 8'b11111111; // 2829 : 255 - 0xff
      12'hB0E: dout  = 8'b11111111; // 2830 : 255 - 0xff
      12'hB0F: dout  = 8'b11111111; // 2831 : 255 - 0xff
      12'hB10: dout  = 8'b01111000; // 2832 : 120 - 0x78 -- Background 0x62
      12'hB11: dout  = 8'b01100000; // 2833 :  96 - 0x60
      12'hB12: dout  = 8'b01000000; // 2834 :  64 - 0x40
      12'hB13: dout  = 8'b01000000; // 2835 :  64 - 0x40
      12'hB14: dout  = 8'b01000000; // 2836 :  64 - 0x40
      12'hB15: dout  = 8'b01100000; // 2837 :  96 - 0x60
      12'hB16: dout  = 8'b00110000; // 2838 :  48 - 0x30
      12'hB17: dout  = 8'b00011111; // 2839 :  31 - 0x1f
      12'hB18: dout  = 8'b10000001; // 2840 : 129 - 0x81 -- Background 0x63
      12'hB19: dout  = 8'b10000011; // 2841 : 131 - 0x83
      12'hB1A: dout  = 8'b11000001; // 2842 : 193 - 0xc1
      12'hB1B: dout  = 8'b01000011; // 2843 :  67 - 0x43
      12'hB1C: dout  = 8'b01000001; // 2844 :  65 - 0x41
      12'hB1D: dout  = 8'b01100011; // 2845 :  99 - 0x63
      12'hB1E: dout  = 8'b00100110; // 2846 :  38 - 0x26
      12'hB1F: dout  = 8'b11111000; // 2847 : 248 - 0xf8
      12'hB20: dout  = 8'b10111001; // 2848 : 185 - 0xb9 -- Background 0x64
      12'hB21: dout  = 8'b10010100; // 2849 : 148 - 0x94
      12'hB22: dout  = 8'b10001110; // 2850 : 142 - 0x8e
      12'hB23: dout  = 8'b11000101; // 2851 : 197 - 0xc5
      12'hB24: dout  = 8'b10010010; // 2852 : 146 - 0x92
      12'hB25: dout  = 8'b11000111; // 2853 : 199 - 0xc7
      12'hB26: dout  = 8'b11100010; // 2854 : 226 - 0xe2
      12'hB27: dout  = 8'b11010000; // 2855 : 208 - 0xd0
      12'hB28: dout  = 8'b10111001; // 2856 : 185 - 0xb9 -- Background 0x65
      12'hB29: dout  = 8'b00010100; // 2857 :  20 - 0x14
      12'hB2A: dout  = 8'b10001110; // 2858 : 142 - 0x8e
      12'hB2B: dout  = 8'b11000101; // 2859 : 197 - 0xc5
      12'hB2C: dout  = 8'b10010010; // 2860 : 146 - 0x92
      12'hB2D: dout  = 8'b01000111; // 2861 :  71 - 0x47
      12'hB2E: dout  = 8'b11100010; // 2862 : 226 - 0xe2
      12'hB2F: dout  = 8'b01010000; // 2863 :  80 - 0x50
      12'hB30: dout  = 8'b10111001; // 2864 : 185 - 0xb9 -- Background 0x66
      12'hB31: dout  = 8'b00010101; // 2865 :  21 - 0x15
      12'hB32: dout  = 8'b10001111; // 2866 : 143 - 0x8f
      12'hB33: dout  = 8'b11000101; // 2867 : 197 - 0xc5
      12'hB34: dout  = 8'b10010011; // 2868 : 147 - 0x93
      12'hB35: dout  = 8'b01000111; // 2869 :  71 - 0x47
      12'hB36: dout  = 8'b11100011; // 2870 : 227 - 0xe3
      12'hB37: dout  = 8'b01010001; // 2871 :  81 - 0x51
      12'hB38: dout  = 8'b01111111; // 2872 : 127 - 0x7f -- Background 0x67
      12'hB39: dout  = 8'b10000000; // 2873 : 128 - 0x80
      12'hB3A: dout  = 8'b11001100; // 2874 : 204 - 0xcc
      12'hB3B: dout  = 8'b01111111; // 2875 : 127 - 0x7f
      12'hB3C: dout  = 8'b00111111; // 2876 :  63 - 0x3f
      12'hB3D: dout  = 8'b00000011; // 2877 :   3 - 0x3
      12'hB3E: dout  = 8'b00000000; // 2878 :   0 - 0x0
      12'hB3F: dout  = 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout  = 8'b11111111; // 2880 : 255 - 0xff -- Background 0x68
      12'hB41: dout  = 8'b00000000; // 2881 :   0 - 0x0
      12'hB42: dout  = 8'b11001100; // 2882 : 204 - 0xcc
      12'hB43: dout  = 8'b00110011; // 2883 :  51 - 0x33
      12'hB44: dout  = 8'b11111111; // 2884 : 255 - 0xff
      12'hB45: dout  = 8'b11111111; // 2885 : 255 - 0xff
      12'hB46: dout  = 8'b00000000; // 2886 :   0 - 0x0
      12'hB47: dout  = 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout  = 8'b11111110; // 2888 : 254 - 0xfe -- Background 0x69
      12'hB49: dout  = 8'b00000001; // 2889 :   1 - 0x1
      12'hB4A: dout  = 8'b11001101; // 2890 : 205 - 0xcd
      12'hB4B: dout  = 8'b00111110; // 2891 :  62 - 0x3e
      12'hB4C: dout  = 8'b11111100; // 2892 : 252 - 0xfc
      12'hB4D: dout  = 8'b11000000; // 2893 : 192 - 0xc0
      12'hB4E: dout  = 8'b00000000; // 2894 :   0 - 0x0
      12'hB4F: dout  = 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout  = 8'b00000000; // 2896 :   0 - 0x0 -- Background 0x6a
      12'hB51: dout  = 8'b00000000; // 2897 :   0 - 0x0
      12'hB52: dout  = 8'b00000000; // 2898 :   0 - 0x0
      12'hB53: dout  = 8'b00000000; // 2899 :   0 - 0x0
      12'hB54: dout  = 8'b00000000; // 2900 :   0 - 0x0
      12'hB55: dout  = 8'b00000000; // 2901 :   0 - 0x0
      12'hB56: dout  = 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout  = 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout  = 8'b01111111; // 2904 : 127 - 0x7f -- Background 0x6b
      12'hB59: dout  = 8'b11111111; // 2905 : 255 - 0xff
      12'hB5A: dout  = 8'b11111111; // 2906 : 255 - 0xff
      12'hB5B: dout  = 8'b11111111; // 2907 : 255 - 0xff
      12'hB5C: dout  = 8'b01111111; // 2908 : 127 - 0x7f
      12'hB5D: dout  = 8'b00110000; // 2909 :  48 - 0x30
      12'hB5E: dout  = 8'b00001111; // 2910 :  15 - 0xf
      12'hB5F: dout  = 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout  = 8'b11111111; // 2912 : 255 - 0xff -- Background 0x6c
      12'hB61: dout  = 8'b11111111; // 2913 : 255 - 0xff
      12'hB62: dout  = 8'b11111111; // 2914 : 255 - 0xff
      12'hB63: dout  = 8'b11111111; // 2915 : 255 - 0xff
      12'hB64: dout  = 8'b11111111; // 2916 : 255 - 0xff
      12'hB65: dout  = 8'b11111110; // 2917 : 254 - 0xfe
      12'hB66: dout  = 8'b00000001; // 2918 :   1 - 0x1
      12'hB67: dout  = 8'b11111110; // 2919 : 254 - 0xfe
      12'hB68: dout  = 8'b00000000; // 2920 :   0 - 0x0 -- Background 0x6d
      12'hB69: dout  = 8'b00000000; // 2921 :   0 - 0x0
      12'hB6A: dout  = 8'b00000000; // 2922 :   0 - 0x0
      12'hB6B: dout  = 8'b00000000; // 2923 :   0 - 0x0
      12'hB6C: dout  = 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout  = 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout  = 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout  = 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout  = 8'b00000000; // 2928 :   0 - 0x0 -- Background 0x6e
      12'hB71: dout  = 8'b00000000; // 2929 :   0 - 0x0
      12'hB72: dout  = 8'b00000000; // 2930 :   0 - 0x0
      12'hB73: dout  = 8'b00000000; // 2931 :   0 - 0x0
      12'hB74: dout  = 8'b00000000; // 2932 :   0 - 0x0
      12'hB75: dout  = 8'b00000000; // 2933 :   0 - 0x0
      12'hB76: dout  = 8'b00000000; // 2934 :   0 - 0x0
      12'hB77: dout  = 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout  = 8'b11111100; // 2936 : 252 - 0xfc -- Background 0x6f
      12'hB79: dout  = 8'b11111110; // 2937 : 254 - 0xfe
      12'hB7A: dout  = 8'b11111111; // 2938 : 255 - 0xff
      12'hB7B: dout  = 8'b11111111; // 2939 : 255 - 0xff
      12'hB7C: dout  = 8'b11110010; // 2940 : 242 - 0xf2
      12'hB7D: dout  = 8'b00001100; // 2941 :  12 - 0xc
      12'hB7E: dout  = 8'b11110000; // 2942 : 240 - 0xf0
      12'hB7F: dout  = 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout  = 8'b01111111; // 2944 : 127 - 0x7f -- Background 0x70
      12'hB81: dout  = 8'b11000000; // 2945 : 192 - 0xc0
      12'hB82: dout  = 8'b10000000; // 2946 : 128 - 0x80
      12'hB83: dout  = 8'b10000000; // 2947 : 128 - 0x80
      12'hB84: dout  = 8'b11100011; // 2948 : 227 - 0xe3
      12'hB85: dout  = 8'b11111111; // 2949 : 255 - 0xff
      12'hB86: dout  = 8'b11111111; // 2950 : 255 - 0xff
      12'hB87: dout  = 8'b11111111; // 2951 : 255 - 0xff
      12'hB88: dout  = 8'b11111111; // 2952 : 255 - 0xff -- Background 0x71
      12'hB89: dout  = 8'b00000000; // 2953 :   0 - 0x0
      12'hB8A: dout  = 8'b00000000; // 2954 :   0 - 0x0
      12'hB8B: dout  = 8'b00000000; // 2955 :   0 - 0x0
      12'hB8C: dout  = 8'b00000000; // 2956 :   0 - 0x0
      12'hB8D: dout  = 8'b11000011; // 2957 : 195 - 0xc3
      12'hB8E: dout  = 8'b11111111; // 2958 : 255 - 0xff
      12'hB8F: dout  = 8'b11111111; // 2959 : 255 - 0xff
      12'hB90: dout  = 8'b11111110; // 2960 : 254 - 0xfe -- Background 0x72
      12'hB91: dout  = 8'b00000011; // 2961 :   3 - 0x3
      12'hB92: dout  = 8'b00000001; // 2962 :   1 - 0x1
      12'hB93: dout  = 8'b00000001; // 2963 :   1 - 0x1
      12'hB94: dout  = 8'b11000111; // 2964 : 199 - 0xc7
      12'hB95: dout  = 8'b11111111; // 2965 : 255 - 0xff
      12'hB96: dout  = 8'b11111111; // 2966 : 255 - 0xff
      12'hB97: dout  = 8'b11111111; // 2967 : 255 - 0xff
      12'hB98: dout  = 8'b11111111; // 2968 : 255 - 0xff -- Background 0x73
      12'hB99: dout  = 8'b11111111; // 2969 : 255 - 0xff
      12'hB9A: dout  = 8'b11111111; // 2970 : 255 - 0xff
      12'hB9B: dout  = 8'b11111111; // 2971 : 255 - 0xff
      12'hB9C: dout  = 8'b11111111; // 2972 : 255 - 0xff
      12'hB9D: dout  = 8'b11111111; // 2973 : 255 - 0xff
      12'hB9E: dout  = 8'b11111111; // 2974 : 255 - 0xff
      12'hB9F: dout  = 8'b11111111; // 2975 : 255 - 0xff
      12'hBA0: dout  = 8'b10111001; // 2976 : 185 - 0xb9 -- Background 0x74
      12'hBA1: dout  = 8'b10010100; // 2977 : 148 - 0x94
      12'hBA2: dout  = 8'b10001110; // 2978 : 142 - 0x8e
      12'hBA3: dout  = 8'b11000101; // 2979 : 197 - 0xc5
      12'hBA4: dout  = 8'b10010010; // 2980 : 146 - 0x92
      12'hBA5: dout  = 8'b11000111; // 2981 : 199 - 0xc7
      12'hBA6: dout  = 8'b11100010; // 2982 : 226 - 0xe2
      12'hBA7: dout  = 8'b01111111; // 2983 : 127 - 0x7f
      12'hBA8: dout  = 8'b10111001; // 2984 : 185 - 0xb9 -- Background 0x75
      12'hBA9: dout  = 8'b00010100; // 2985 :  20 - 0x14
      12'hBAA: dout  = 8'b10001110; // 2986 : 142 - 0x8e
      12'hBAB: dout  = 8'b11000101; // 2987 : 197 - 0xc5
      12'hBAC: dout  = 8'b10010010; // 2988 : 146 - 0x92
      12'hBAD: dout  = 8'b01000111; // 2989 :  71 - 0x47
      12'hBAE: dout  = 8'b11100010; // 2990 : 226 - 0xe2
      12'hBAF: dout  = 8'b11111111; // 2991 : 255 - 0xff
      12'hBB0: dout  = 8'b10111001; // 2992 : 185 - 0xb9 -- Background 0x76
      12'hBB1: dout  = 8'b00010101; // 2993 :  21 - 0x15
      12'hBB2: dout  = 8'b10001111; // 2994 : 143 - 0x8f
      12'hBB3: dout  = 8'b11000101; // 2995 : 197 - 0xc5
      12'hBB4: dout  = 8'b10010011; // 2996 : 147 - 0x93
      12'hBB5: dout  = 8'b01000111; // 2997 :  71 - 0x47
      12'hBB6: dout  = 8'b11100011; // 2998 : 227 - 0xe3
      12'hBB7: dout  = 8'b11111110; // 2999 : 254 - 0xfe
      12'hBB8: dout  = 8'b11111111; // 3000 : 255 - 0xff -- Background 0x77
      12'hBB9: dout  = 8'b11111111; // 3001 : 255 - 0xff
      12'hBBA: dout  = 8'b11111111; // 3002 : 255 - 0xff
      12'hBBB: dout  = 8'b11111111; // 3003 : 255 - 0xff
      12'hBBC: dout  = 8'b11111111; // 3004 : 255 - 0xff
      12'hBBD: dout  = 8'b11111111; // 3005 : 255 - 0xff
      12'hBBE: dout  = 8'b11111111; // 3006 : 255 - 0xff
      12'hBBF: dout  = 8'b11111111; // 3007 : 255 - 0xff
      12'hBC0: dout  = 8'b00000000; // 3008 :   0 - 0x0 -- Background 0x78
      12'hBC1: dout  = 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout  = 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout  = 8'b00000000; // 3011 :   0 - 0x0
      12'hBC4: dout  = 8'b00000000; // 3012 :   0 - 0x0
      12'hBC5: dout  = 8'b00000000; // 3013 :   0 - 0x0
      12'hBC6: dout  = 8'b00000000; // 3014 :   0 - 0x0
      12'hBC7: dout  = 8'b00000000; // 3015 :   0 - 0x0
      12'hBC8: dout  = 8'b00000000; // 3016 :   0 - 0x0 -- Background 0x79
      12'hBC9: dout  = 8'b00000000; // 3017 :   0 - 0x0
      12'hBCA: dout  = 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout  = 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout  = 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout  = 8'b00000000; // 3021 :   0 - 0x0
      12'hBCE: dout  = 8'b00000000; // 3022 :   0 - 0x0
      12'hBCF: dout  = 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout  = 8'b00000000; // 3024 :   0 - 0x0 -- Background 0x7a
      12'hBD1: dout  = 8'b00000000; // 3025 :   0 - 0x0
      12'hBD2: dout  = 8'b00000000; // 3026 :   0 - 0x0
      12'hBD3: dout  = 8'b00000000; // 3027 :   0 - 0x0
      12'hBD4: dout  = 8'b00000000; // 3028 :   0 - 0x0
      12'hBD5: dout  = 8'b00000000; // 3029 :   0 - 0x0
      12'hBD6: dout  = 8'b00000000; // 3030 :   0 - 0x0
      12'hBD7: dout  = 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout  = 8'b00000000; // 3032 :   0 - 0x0 -- Background 0x7b
      12'hBD9: dout  = 8'b00000000; // 3033 :   0 - 0x0
      12'hBDA: dout  = 8'b00000000; // 3034 :   0 - 0x0
      12'hBDB: dout  = 8'b00000000; // 3035 :   0 - 0x0
      12'hBDC: dout  = 8'b00000000; // 3036 :   0 - 0x0
      12'hBDD: dout  = 8'b00000000; // 3037 :   0 - 0x0
      12'hBDE: dout  = 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout  = 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout  = 8'b00100010; // 3040 :  34 - 0x22 -- Background 0x7c
      12'hBE1: dout  = 8'b01010101; // 3041 :  85 - 0x55
      12'hBE2: dout  = 8'b10101010; // 3042 : 170 - 0xaa
      12'hBE3: dout  = 8'b00000101; // 3043 :   5 - 0x5
      12'hBE4: dout  = 8'b00000100; // 3044 :   4 - 0x4
      12'hBE5: dout  = 8'b00001010; // 3045 :  10 - 0xa
      12'hBE6: dout  = 8'b01010000; // 3046 :  80 - 0x50
      12'hBE7: dout  = 8'b00000010; // 3047 :   2 - 0x2
      12'hBE8: dout  = 8'b01110011; // 3048 : 115 - 0x73 -- Background 0x7d
      12'hBE9: dout  = 8'b11111111; // 3049 : 255 - 0xff
      12'hBEA: dout  = 8'b11111111; // 3050 : 255 - 0xff
      12'hBEB: dout  = 8'b10111101; // 3051 : 189 - 0xbd
      12'hBEC: dout  = 8'b01101110; // 3052 : 110 - 0x6e
      12'hBED: dout  = 8'b00001010; // 3053 :  10 - 0xa
      12'hBEE: dout  = 8'b01010000; // 3054 :  80 - 0x50
      12'hBEF: dout  = 8'b00000010; // 3055 :   2 - 0x2
      12'hBF0: dout  = 8'b00100000; // 3056 :  32 - 0x20 -- Background 0x7e
      12'hBF1: dout  = 8'b01010000; // 3057 :  80 - 0x50
      12'hBF2: dout  = 8'b10000100; // 3058 : 132 - 0x84
      12'hBF3: dout  = 8'b00000000; // 3059 :   0 - 0x0
      12'hBF4: dout  = 8'b00100100; // 3060 :  36 - 0x24
      12'hBF5: dout  = 8'b01011010; // 3061 :  90 - 0x5a
      12'hBF6: dout  = 8'b00010000; // 3062 :  16 - 0x10
      12'hBF7: dout  = 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout  = 8'b11111111; // 3064 : 255 - 0xff -- Background 0x7f
      12'hBF9: dout  = 8'b01010000; // 3065 :  80 - 0x50
      12'hBFA: dout  = 8'b10000100; // 3066 : 132 - 0x84
      12'hBFB: dout  = 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout  = 8'b00100100; // 3068 :  36 - 0x24
      12'hBFD: dout  = 8'b01011010; // 3069 :  90 - 0x5a
      12'hBFE: dout  = 8'b00010000; // 3070 :  16 - 0x10
      12'hBFF: dout  = 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout  = 8'b11111111; // 3072 : 255 - 0xff -- Background 0x80
      12'hC01: dout  = 8'b10000000; // 3073 : 128 - 0x80
      12'hC02: dout  = 8'b11001111; // 3074 : 207 - 0xcf
      12'hC03: dout  = 8'b01001000; // 3075 :  72 - 0x48
      12'hC04: dout  = 8'b11001111; // 3076 : 207 - 0xcf
      12'hC05: dout  = 8'b10000000; // 3077 : 128 - 0x80
      12'hC06: dout  = 8'b11001111; // 3078 : 207 - 0xcf
      12'hC07: dout  = 8'b01001000; // 3079 :  72 - 0x48
      12'hC08: dout  = 8'b11111111; // 3080 : 255 - 0xff -- Background 0x81
      12'hC09: dout  = 8'b10000000; // 3081 : 128 - 0x80
      12'hC0A: dout  = 8'b11111111; // 3082 : 255 - 0xff
      12'hC0B: dout  = 8'b10000000; // 3083 : 128 - 0x80
      12'hC0C: dout  = 8'b10000000; // 3084 : 128 - 0x80
      12'hC0D: dout  = 8'b11011111; // 3085 : 223 - 0xdf
      12'hC0E: dout  = 8'b10110000; // 3086 : 176 - 0xb0
      12'hC0F: dout  = 8'b11000000; // 3087 : 192 - 0xc0
      12'hC10: dout  = 8'b11111111; // 3088 : 255 - 0xff -- Background 0x82
      12'hC11: dout  = 8'b00000001; // 3089 :   1 - 0x1
      12'hC12: dout  = 8'b11110011; // 3090 : 243 - 0xf3
      12'hC13: dout  = 8'b00010010; // 3091 :  18 - 0x12
      12'hC14: dout  = 8'b11110011; // 3092 : 243 - 0xf3
      12'hC15: dout  = 8'b00000001; // 3093 :   1 - 0x1
      12'hC16: dout  = 8'b11110011; // 3094 : 243 - 0xf3
      12'hC17: dout  = 8'b00010010; // 3095 :  18 - 0x12
      12'hC18: dout  = 8'b11111111; // 3096 : 255 - 0xff -- Background 0x83
      12'hC19: dout  = 8'b00000000; // 3097 :   0 - 0x0
      12'hC1A: dout  = 8'b11111111; // 3098 : 255 - 0xff
      12'hC1B: dout  = 8'b00000000; // 3099 :   0 - 0x0
      12'hC1C: dout  = 8'b00000000; // 3100 :   0 - 0x0
      12'hC1D: dout  = 8'b11111111; // 3101 : 255 - 0xff
      12'hC1E: dout  = 8'b00000000; // 3102 :   0 - 0x0
      12'hC1F: dout  = 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout  = 8'b11111111; // 3104 : 255 - 0xff -- Background 0x84
      12'hC21: dout  = 8'b10000010; // 3105 : 130 - 0x82
      12'hC22: dout  = 8'b00010000; // 3106 :  16 - 0x10
      12'hC23: dout  = 8'b00000000; // 3107 :   0 - 0x0
      12'hC24: dout  = 8'b00000000; // 3108 :   0 - 0x0
      12'hC25: dout  = 8'b00010000; // 3109 :  16 - 0x10
      12'hC26: dout  = 8'b01000100; // 3110 :  68 - 0x44
      12'hC27: dout  = 8'b11111111; // 3111 : 255 - 0xff
      12'hC28: dout  = 8'b11111111; // 3112 : 255 - 0xff -- Background 0x85
      12'hC29: dout  = 8'b00000001; // 3113 :   1 - 0x1
      12'hC2A: dout  = 8'b11111111; // 3114 : 255 - 0xff
      12'hC2B: dout  = 8'b00000001; // 3115 :   1 - 0x1
      12'hC2C: dout  = 8'b00000001; // 3116 :   1 - 0x1
      12'hC2D: dout  = 8'b11110011; // 3117 : 243 - 0xf3
      12'hC2E: dout  = 8'b00001101; // 3118 :  13 - 0xd
      12'hC2F: dout  = 8'b00000011; // 3119 :   3 - 0x3
      12'hC30: dout  = 8'b00000000; // 3120 :   0 - 0x0 -- Background 0x86
      12'hC31: dout  = 8'b00000000; // 3121 :   0 - 0x0
      12'hC32: dout  = 8'b00000000; // 3122 :   0 - 0x0
      12'hC33: dout  = 8'b00000000; // 3123 :   0 - 0x0
      12'hC34: dout  = 8'b00000000; // 3124 :   0 - 0x0
      12'hC35: dout  = 8'b00000000; // 3125 :   0 - 0x0
      12'hC36: dout  = 8'b00000000; // 3126 :   0 - 0x0
      12'hC37: dout  = 8'b00000000; // 3127 :   0 - 0x0
      12'hC38: dout  = 8'b00000000; // 3128 :   0 - 0x0 -- Background 0x87
      12'hC39: dout  = 8'b00000000; // 3129 :   0 - 0x0
      12'hC3A: dout  = 8'b00000000; // 3130 :   0 - 0x0
      12'hC3B: dout  = 8'b00000000; // 3131 :   0 - 0x0
      12'hC3C: dout  = 8'b00000000; // 3132 :   0 - 0x0
      12'hC3D: dout  = 8'b00000000; // 3133 :   0 - 0x0
      12'hC3E: dout  = 8'b00000000; // 3134 :   0 - 0x0
      12'hC3F: dout  = 8'b00000000; // 3135 :   0 - 0x0
      12'hC40: dout  = 8'b00000111; // 3136 :   7 - 0x7 -- Background 0x88
      12'hC41: dout  = 8'b00011110; // 3137 :  30 - 0x1e
      12'hC42: dout  = 8'b00101111; // 3138 :  47 - 0x2f
      12'hC43: dout  = 8'b01010011; // 3139 :  83 - 0x53
      12'hC44: dout  = 8'b01101110; // 3140 : 110 - 0x6e
      12'hC45: dout  = 8'b11011011; // 3141 : 219 - 0xdb
      12'hC46: dout  = 8'b11111010; // 3142 : 250 - 0xfa
      12'hC47: dout  = 8'b11010101; // 3143 : 213 - 0xd5
      12'hC48: dout  = 8'b10111011; // 3144 : 187 - 0xbb -- Background 0x89
      12'hC49: dout  = 8'b11110010; // 3145 : 242 - 0xf2
      12'hC4A: dout  = 8'b11011101; // 3146 : 221 - 0xdd
      12'hC4B: dout  = 8'b01001111; // 3147 :  79 - 0x4f
      12'hC4C: dout  = 8'b01111011; // 3148 : 123 - 0x7b
      12'hC4D: dout  = 8'b00110010; // 3149 :  50 - 0x32
      12'hC4E: dout  = 8'b00011111; // 3150 :  31 - 0x1f
      12'hC4F: dout  = 8'b00000111; // 3151 :   7 - 0x7
      12'hC50: dout  = 8'b11100000; // 3152 : 224 - 0xe0 -- Background 0x8a
      12'hC51: dout  = 8'b11011000; // 3153 : 216 - 0xd8
      12'hC52: dout  = 8'b01010100; // 3154 :  84 - 0x54
      12'hC53: dout  = 8'b11101010; // 3155 : 234 - 0xea
      12'hC54: dout  = 8'b10111010; // 3156 : 186 - 0xba
      12'hC55: dout  = 8'b10010011; // 3157 : 147 - 0x93
      12'hC56: dout  = 8'b11011111; // 3158 : 223 - 0xdf
      12'hC57: dout  = 8'b10111101; // 3159 : 189 - 0xbd
      12'hC58: dout  = 8'b01101011; // 3160 : 107 - 0x6b -- Background 0x8b
      12'hC59: dout  = 8'b10011111; // 3161 : 159 - 0x9f
      12'hC5A: dout  = 8'b01011101; // 3162 :  93 - 0x5d
      12'hC5B: dout  = 8'b10110110; // 3163 : 182 - 0xb6
      12'hC5C: dout  = 8'b11101010; // 3164 : 234 - 0xea
      12'hC5D: dout  = 8'b11001100; // 3165 : 204 - 0xcc
      12'hC5E: dout  = 8'b01111000; // 3166 : 120 - 0x78
      12'hC5F: dout  = 8'b11100000; // 3167 : 224 - 0xe0
      12'hC60: dout  = 8'b00000111; // 3168 :   7 - 0x7 -- Background 0x8c
      12'hC61: dout  = 8'b00011000; // 3169 :  24 - 0x18
      12'hC62: dout  = 8'b00100011; // 3170 :  35 - 0x23
      12'hC63: dout  = 8'b01001100; // 3171 :  76 - 0x4c
      12'hC64: dout  = 8'b01110000; // 3172 : 112 - 0x70
      12'hC65: dout  = 8'b10100001; // 3173 : 161 - 0xa1
      12'hC66: dout  = 8'b10100110; // 3174 : 166 - 0xa6
      12'hC67: dout  = 8'b10101000; // 3175 : 168 - 0xa8
      12'hC68: dout  = 8'b10100101; // 3176 : 165 - 0xa5 -- Background 0x8d
      12'hC69: dout  = 8'b10100010; // 3177 : 162 - 0xa2
      12'hC6A: dout  = 8'b10010000; // 3178 : 144 - 0x90
      12'hC6B: dout  = 8'b01001000; // 3179 :  72 - 0x48
      12'hC6C: dout  = 8'b01000111; // 3180 :  71 - 0x47
      12'hC6D: dout  = 8'b00100000; // 3181 :  32 - 0x20
      12'hC6E: dout  = 8'b00011001; // 3182 :  25 - 0x19
      12'hC6F: dout  = 8'b00000111; // 3183 :   7 - 0x7
      12'hC70: dout  = 8'b11100000; // 3184 : 224 - 0xe0 -- Background 0x8e
      12'hC71: dout  = 8'b00011000; // 3185 :  24 - 0x18
      12'hC72: dout  = 8'b00000100; // 3186 :   4 - 0x4
      12'hC73: dout  = 8'b11000010; // 3187 : 194 - 0xc2
      12'hC74: dout  = 8'b00110010; // 3188 :  50 - 0x32
      12'hC75: dout  = 8'b00001001; // 3189 :   9 - 0x9
      12'hC76: dout  = 8'b11000101; // 3190 : 197 - 0xc5
      12'hC77: dout  = 8'b00100101; // 3191 :  37 - 0x25
      12'hC78: dout  = 8'b10100101; // 3192 : 165 - 0xa5 -- Background 0x8f
      12'hC79: dout  = 8'b01100101; // 3193 : 101 - 0x65
      12'hC7A: dout  = 8'b01000101; // 3194 :  69 - 0x45
      12'hC7B: dout  = 8'b10001010; // 3195 : 138 - 0x8a
      12'hC7C: dout  = 8'b10010010; // 3196 : 146 - 0x92
      12'hC7D: dout  = 8'b00100100; // 3197 :  36 - 0x24
      12'hC7E: dout  = 8'b11011000; // 3198 : 216 - 0xd8
      12'hC7F: dout  = 8'b11100000; // 3199 : 224 - 0xe0
      12'hC80: dout  = 8'b00000000; // 3200 :   0 - 0x0 -- Background 0x90
      12'hC81: dout  = 8'b00000000; // 3201 :   0 - 0x0
      12'hC82: dout  = 8'b00100000; // 3202 :  32 - 0x20
      12'hC83: dout  = 8'b00110000; // 3203 :  48 - 0x30
      12'hC84: dout  = 8'b00101100; // 3204 :  44 - 0x2c
      12'hC85: dout  = 8'b00100010; // 3205 :  34 - 0x22
      12'hC86: dout  = 8'b00010001; // 3206 :  17 - 0x11
      12'hC87: dout  = 8'b00001000; // 3207 :   8 - 0x8
      12'hC88: dout  = 8'b00000100; // 3208 :   4 - 0x4 -- Background 0x91
      12'hC89: dout  = 8'b11110010; // 3209 : 242 - 0xf2
      12'hC8A: dout  = 8'b11001111; // 3210 : 207 - 0xcf
      12'hC8B: dout  = 8'b00110000; // 3211 :  48 - 0x30
      12'hC8C: dout  = 8'b00001100; // 3212 :  12 - 0xc
      12'hC8D: dout  = 8'b11111111; // 3213 : 255 - 0xff
      12'hC8E: dout  = 8'b10000000; // 3214 : 128 - 0x80
      12'hC8F: dout  = 8'b11111111; // 3215 : 255 - 0xff
      12'hC90: dout  = 8'b01000010; // 3216 :  66 - 0x42 -- Background 0x92
      12'hC91: dout  = 8'b10100101; // 3217 : 165 - 0xa5
      12'hC92: dout  = 8'b10100101; // 3218 : 165 - 0xa5
      12'hC93: dout  = 8'b10011001; // 3219 : 153 - 0x99
      12'hC94: dout  = 8'b10011001; // 3220 : 153 - 0x99
      12'hC95: dout  = 8'b10011001; // 3221 : 153 - 0x99
      12'hC96: dout  = 8'b00000001; // 3222 :   1 - 0x1
      12'hC97: dout  = 8'b00000000; // 3223 :   0 - 0x0
      12'hC98: dout  = 8'b11111111; // 3224 : 255 - 0xff -- Background 0x93
      12'hC99: dout  = 8'b11111111; // 3225 : 255 - 0xff
      12'hC9A: dout  = 8'b11111111; // 3226 : 255 - 0xff
      12'hC9B: dout  = 8'b10000001; // 3227 : 129 - 0x81
      12'hC9C: dout  = 8'b11111111; // 3228 : 255 - 0xff
      12'hC9D: dout  = 8'b11111111; // 3229 : 255 - 0xff
      12'hC9E: dout  = 8'b11111111; // 3230 : 255 - 0xff
      12'hC9F: dout  = 8'b10000001; // 3231 : 129 - 0x81
      12'hCA0: dout  = 8'b00000000; // 3232 :   0 - 0x0 -- Background 0x94
      12'hCA1: dout  = 8'b00000000; // 3233 :   0 - 0x0
      12'hCA2: dout  = 8'b00000100; // 3234 :   4 - 0x4
      12'hCA3: dout  = 8'b00001100; // 3235 :  12 - 0xc
      12'hCA4: dout  = 8'b00110100; // 3236 :  52 - 0x34
      12'hCA5: dout  = 8'b01000100; // 3237 :  68 - 0x44
      12'hCA6: dout  = 8'b10001000; // 3238 : 136 - 0x88
      12'hCA7: dout  = 8'b00010000; // 3239 :  16 - 0x10
      12'hCA8: dout  = 8'b00100000; // 3240 :  32 - 0x20 -- Background 0x95
      12'hCA9: dout  = 8'b01001111; // 3241 :  79 - 0x4f
      12'hCAA: dout  = 8'b11110011; // 3242 : 243 - 0xf3
      12'hCAB: dout  = 8'b00001100; // 3243 :  12 - 0xc
      12'hCAC: dout  = 8'b00110000; // 3244 :  48 - 0x30
      12'hCAD: dout  = 8'b11111111; // 3245 : 255 - 0xff
      12'hCAE: dout  = 8'b00000001; // 3246 :   1 - 0x1
      12'hCAF: dout  = 8'b11111111; // 3247 : 255 - 0xff
      12'hCB0: dout  = 8'b01111111; // 3248 : 127 - 0x7f -- Background 0x96
      12'hCB1: dout  = 8'b11111111; // 3249 : 255 - 0xff
      12'hCB2: dout  = 8'b11111111; // 3250 : 255 - 0xff
      12'hCB3: dout  = 8'b11111111; // 3251 : 255 - 0xff
      12'hCB4: dout  = 8'b11111011; // 3252 : 251 - 0xfb
      12'hCB5: dout  = 8'b11111111; // 3253 : 255 - 0xff
      12'hCB6: dout  = 8'b11111111; // 3254 : 255 - 0xff
      12'hCB7: dout  = 8'b11111111; // 3255 : 255 - 0xff
      12'hCB8: dout  = 8'b11111111; // 3256 : 255 - 0xff -- Background 0x97
      12'hCB9: dout  = 8'b11111111; // 3257 : 255 - 0xff
      12'hCBA: dout  = 8'b11111111; // 3258 : 255 - 0xff
      12'hCBB: dout  = 8'b11111111; // 3259 : 255 - 0xff
      12'hCBC: dout  = 8'b11111111; // 3260 : 255 - 0xff
      12'hCBD: dout  = 8'b11111111; // 3261 : 255 - 0xff
      12'hCBE: dout  = 8'b11111110; // 3262 : 254 - 0xfe
      12'hCBF: dout  = 8'b11111111; // 3263 : 255 - 0xff
      12'hCC0: dout  = 8'b11111111; // 3264 : 255 - 0xff -- Background 0x98
      12'hCC1: dout  = 8'b10111111; // 3265 : 191 - 0xbf
      12'hCC2: dout  = 8'b11111111; // 3266 : 255 - 0xff
      12'hCC3: dout  = 8'b11111111; // 3267 : 255 - 0xff
      12'hCC4: dout  = 8'b11111011; // 3268 : 251 - 0xfb
      12'hCC5: dout  = 8'b11111111; // 3269 : 255 - 0xff
      12'hCC6: dout  = 8'b11111111; // 3270 : 255 - 0xff
      12'hCC7: dout  = 8'b11111111; // 3271 : 255 - 0xff
      12'hCC8: dout  = 8'b11111111; // 3272 : 255 - 0xff -- Background 0x99
      12'hCC9: dout  = 8'b11111111; // 3273 : 255 - 0xff
      12'hCCA: dout  = 8'b11111111; // 3274 : 255 - 0xff
      12'hCCB: dout  = 8'b11111111; // 3275 : 255 - 0xff
      12'hCCC: dout  = 8'b11111111; // 3276 : 255 - 0xff
      12'hCCD: dout  = 8'b11111111; // 3277 : 255 - 0xff
      12'hCCE: dout  = 8'b11111110; // 3278 : 254 - 0xfe
      12'hCCF: dout  = 8'b11111111; // 3279 : 255 - 0xff
      12'hCD0: dout  = 8'b11111110; // 3280 : 254 - 0xfe -- Background 0x9a
      12'hCD1: dout  = 8'b11111111; // 3281 : 255 - 0xff
      12'hCD2: dout  = 8'b11111111; // 3282 : 255 - 0xff
      12'hCD3: dout  = 8'b11111111; // 3283 : 255 - 0xff
      12'hCD4: dout  = 8'b11111011; // 3284 : 251 - 0xfb
      12'hCD5: dout  = 8'b11111111; // 3285 : 255 - 0xff
      12'hCD6: dout  = 8'b11111111; // 3286 : 255 - 0xff
      12'hCD7: dout  = 8'b11111111; // 3287 : 255 - 0xff
      12'hCD8: dout  = 8'b11111111; // 3288 : 255 - 0xff -- Background 0x9b
      12'hCD9: dout  = 8'b11111111; // 3289 : 255 - 0xff
      12'hCDA: dout  = 8'b11111111; // 3290 : 255 - 0xff
      12'hCDB: dout  = 8'b11111111; // 3291 : 255 - 0xff
      12'hCDC: dout  = 8'b11111111; // 3292 : 255 - 0xff
      12'hCDD: dout  = 8'b11111111; // 3293 : 255 - 0xff
      12'hCDE: dout  = 8'b11111111; // 3294 : 255 - 0xff
      12'hCDF: dout  = 8'b11111111; // 3295 : 255 - 0xff
      12'hCE0: dout  = 8'b11111111; // 3296 : 255 - 0xff -- Background 0x9c
      12'hCE1: dout  = 8'b11111111; // 3297 : 255 - 0xff
      12'hCE2: dout  = 8'b10100000; // 3298 : 160 - 0xa0
      12'hCE3: dout  = 8'b10010000; // 3299 : 144 - 0x90
      12'hCE4: dout  = 8'b10001000; // 3300 : 136 - 0x88
      12'hCE5: dout  = 8'b10000100; // 3301 : 132 - 0x84
      12'hCE6: dout  = 8'b01101010; // 3302 : 106 - 0x6a
      12'hCE7: dout  = 8'b00111111; // 3303 :  63 - 0x3f
      12'hCE8: dout  = 8'b11111111; // 3304 : 255 - 0xff -- Background 0x9d
      12'hCE9: dout  = 8'b11111111; // 3305 : 255 - 0xff
      12'hCEA: dout  = 8'b00100001; // 3306 :  33 - 0x21
      12'hCEB: dout  = 8'b00010001; // 3307 :  17 - 0x11
      12'hCEC: dout  = 8'b00001001; // 3308 :   9 - 0x9
      12'hCED: dout  = 8'b00000101; // 3309 :   5 - 0x5
      12'hCEE: dout  = 8'b10101010; // 3310 : 170 - 0xaa
      12'hCEF: dout  = 8'b11111100; // 3311 : 252 - 0xfc
      12'hCF0: dout  = 8'b11111111; // 3312 : 255 - 0xff -- Background 0x9e
      12'hCF1: dout  = 8'b11111111; // 3313 : 255 - 0xff
      12'hCF2: dout  = 8'b00100000; // 3314 :  32 - 0x20
      12'hCF3: dout  = 8'b00010000; // 3315 :  16 - 0x10
      12'hCF4: dout  = 8'b00001000; // 3316 :   8 - 0x8
      12'hCF5: dout  = 8'b00000100; // 3317 :   4 - 0x4
      12'hCF6: dout  = 8'b10101010; // 3318 : 170 - 0xaa
      12'hCF7: dout  = 8'b11111111; // 3319 : 255 - 0xff
      12'hCF8: dout  = 8'b00000000; // 3320 :   0 - 0x0 -- Background 0x9f
      12'hCF9: dout  = 8'b00000000; // 3321 :   0 - 0x0
      12'hCFA: dout  = 8'b00000000; // 3322 :   0 - 0x0
      12'hCFB: dout  = 8'b00000000; // 3323 :   0 - 0x0
      12'hCFC: dout  = 8'b00000000; // 3324 :   0 - 0x0
      12'hCFD: dout  = 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout  = 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout  = 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout  = 8'b11111111; // 3328 : 255 - 0xff -- Background 0xa0
      12'hD01: dout  = 8'b11010101; // 3329 : 213 - 0xd5
      12'hD02: dout  = 8'b11111111; // 3330 : 255 - 0xff
      12'hD03: dout  = 8'b00000010; // 3331 :   2 - 0x2
      12'hD04: dout  = 8'b00000010; // 3332 :   2 - 0x2
      12'hD05: dout  = 8'b00000010; // 3333 :   2 - 0x2
      12'hD06: dout  = 8'b00000010; // 3334 :   2 - 0x2
      12'hD07: dout  = 8'b00000010; // 3335 :   2 - 0x2
      12'hD08: dout  = 8'b00000010; // 3336 :   2 - 0x2 -- Background 0xa1
      12'hD09: dout  = 8'b00000010; // 3337 :   2 - 0x2
      12'hD0A: dout  = 8'b00000010; // 3338 :   2 - 0x2
      12'hD0B: dout  = 8'b00000010; // 3339 :   2 - 0x2
      12'hD0C: dout  = 8'b00000010; // 3340 :   2 - 0x2
      12'hD0D: dout  = 8'b00000010; // 3341 :   2 - 0x2
      12'hD0E: dout  = 8'b00000010; // 3342 :   2 - 0x2
      12'hD0F: dout  = 8'b00000010; // 3343 :   2 - 0x2
      12'hD10: dout  = 8'b11111111; // 3344 : 255 - 0xff -- Background 0xa2
      12'hD11: dout  = 8'b01010101; // 3345 :  85 - 0x55
      12'hD12: dout  = 8'b11111111; // 3346 : 255 - 0xff
      12'hD13: dout  = 8'b01000000; // 3347 :  64 - 0x40
      12'hD14: dout  = 8'b01000000; // 3348 :  64 - 0x40
      12'hD15: dout  = 8'b01000000; // 3349 :  64 - 0x40
      12'hD16: dout  = 8'b01000000; // 3350 :  64 - 0x40
      12'hD17: dout  = 8'b01000000; // 3351 :  64 - 0x40
      12'hD18: dout  = 8'b01000000; // 3352 :  64 - 0x40 -- Background 0xa3
      12'hD19: dout  = 8'b01000000; // 3353 :  64 - 0x40
      12'hD1A: dout  = 8'b01000000; // 3354 :  64 - 0x40
      12'hD1B: dout  = 8'b01000000; // 3355 :  64 - 0x40
      12'hD1C: dout  = 8'b01000000; // 3356 :  64 - 0x40
      12'hD1D: dout  = 8'b01000000; // 3357 :  64 - 0x40
      12'hD1E: dout  = 8'b01000000; // 3358 :  64 - 0x40
      12'hD1F: dout  = 8'b01000000; // 3359 :  64 - 0x40
      12'hD20: dout  = 8'b00110001; // 3360 :  49 - 0x31 -- Background 0xa4
      12'hD21: dout  = 8'b01001000; // 3361 :  72 - 0x48
      12'hD22: dout  = 8'b01000101; // 3362 :  69 - 0x45
      12'hD23: dout  = 8'b10000101; // 3363 : 133 - 0x85
      12'hD24: dout  = 8'b10000011; // 3364 : 131 - 0x83
      12'hD25: dout  = 8'b10000010; // 3365 : 130 - 0x82
      12'hD26: dout  = 8'b01100010; // 3366 :  98 - 0x62
      12'hD27: dout  = 8'b00010010; // 3367 :  18 - 0x12
      12'hD28: dout  = 8'b00110010; // 3368 :  50 - 0x32 -- Background 0xa5
      12'hD29: dout  = 8'b00100010; // 3369 :  34 - 0x22
      12'hD2A: dout  = 8'b01000010; // 3370 :  66 - 0x42
      12'hD2B: dout  = 8'b01000000; // 3371 :  64 - 0x40
      12'hD2C: dout  = 8'b01000000; // 3372 :  64 - 0x40
      12'hD2D: dout  = 8'b00100000; // 3373 :  32 - 0x20
      12'hD2E: dout  = 8'b00011110; // 3374 :  30 - 0x1e
      12'hD2F: dout  = 8'b00000111; // 3375 :   7 - 0x7
      12'hD30: dout  = 8'b10000000; // 3376 : 128 - 0x80 -- Background 0xa6
      12'hD31: dout  = 8'b11100000; // 3377 : 224 - 0xe0
      12'hD32: dout  = 8'b00111000; // 3378 :  56 - 0x38
      12'hD33: dout  = 8'b00100100; // 3379 :  36 - 0x24
      12'hD34: dout  = 8'b00000100; // 3380 :   4 - 0x4
      12'hD35: dout  = 8'b00001000; // 3381 :   8 - 0x8
      12'hD36: dout  = 8'b00110000; // 3382 :  48 - 0x30
      12'hD37: dout  = 8'b00100000; // 3383 :  32 - 0x20
      12'hD38: dout  = 8'b00110000; // 3384 :  48 - 0x30 -- Background 0xa7
      12'hD39: dout  = 8'b00001000; // 3385 :   8 - 0x8
      12'hD3A: dout  = 8'b00001000; // 3386 :   8 - 0x8
      12'hD3B: dout  = 8'b00110000; // 3387 :  48 - 0x30
      12'hD3C: dout  = 8'b00100000; // 3388 :  32 - 0x20
      12'hD3D: dout  = 8'b00100000; // 3389 :  32 - 0x20
      12'hD3E: dout  = 8'b00110000; // 3390 :  48 - 0x30
      12'hD3F: dout  = 8'b11110000; // 3391 : 240 - 0xf0
      12'hD40: dout  = 8'b11111111; // 3392 : 255 - 0xff -- Background 0xa8
      12'hD41: dout  = 8'b11010010; // 3393 : 210 - 0xd2
      12'hD42: dout  = 8'b11110100; // 3394 : 244 - 0xf4
      12'hD43: dout  = 8'b11011000; // 3395 : 216 - 0xd8
      12'hD44: dout  = 8'b11111000; // 3396 : 248 - 0xf8
      12'hD45: dout  = 8'b11010100; // 3397 : 212 - 0xd4
      12'hD46: dout  = 8'b11110010; // 3398 : 242 - 0xf2
      12'hD47: dout  = 8'b11010001; // 3399 : 209 - 0xd1
      12'hD48: dout  = 8'b11110001; // 3400 : 241 - 0xf1 -- Background 0xa9
      12'hD49: dout  = 8'b11010010; // 3401 : 210 - 0xd2
      12'hD4A: dout  = 8'b11110100; // 3402 : 244 - 0xf4
      12'hD4B: dout  = 8'b11011000; // 3403 : 216 - 0xd8
      12'hD4C: dout  = 8'b11111000; // 3404 : 248 - 0xf8
      12'hD4D: dout  = 8'b11010100; // 3405 : 212 - 0xd4
      12'hD4E: dout  = 8'b11110010; // 3406 : 242 - 0xf2
      12'hD4F: dout  = 8'b11111111; // 3407 : 255 - 0xff
      12'hD50: dout  = 8'b11111111; // 3408 : 255 - 0xff -- Background 0xaa
      12'hD51: dout  = 8'b01000010; // 3409 :  66 - 0x42
      12'hD52: dout  = 8'b00100100; // 3410 :  36 - 0x24
      12'hD53: dout  = 8'b00011000; // 3411 :  24 - 0x18
      12'hD54: dout  = 8'b00011000; // 3412 :  24 - 0x18
      12'hD55: dout  = 8'b00100100; // 3413 :  36 - 0x24
      12'hD56: dout  = 8'b01000010; // 3414 :  66 - 0x42
      12'hD57: dout  = 8'b10000001; // 3415 : 129 - 0x81
      12'hD58: dout  = 8'b10000001; // 3416 : 129 - 0x81 -- Background 0xab
      12'hD59: dout  = 8'b01000010; // 3417 :  66 - 0x42
      12'hD5A: dout  = 8'b00100100; // 3418 :  36 - 0x24
      12'hD5B: dout  = 8'b00011000; // 3419 :  24 - 0x18
      12'hD5C: dout  = 8'b00011000; // 3420 :  24 - 0x18
      12'hD5D: dout  = 8'b00100100; // 3421 :  36 - 0x24
      12'hD5E: dout  = 8'b01000010; // 3422 :  66 - 0x42
      12'hD5F: dout  = 8'b11111111; // 3423 : 255 - 0xff
      12'hD60: dout  = 8'b11111111; // 3424 : 255 - 0xff -- Background 0xac
      12'hD61: dout  = 8'b01001101; // 3425 :  77 - 0x4d
      12'hD62: dout  = 8'b00101111; // 3426 :  47 - 0x2f
      12'hD63: dout  = 8'b00011101; // 3427 :  29 - 0x1d
      12'hD64: dout  = 8'b00011111; // 3428 :  31 - 0x1f
      12'hD65: dout  = 8'b00101101; // 3429 :  45 - 0x2d
      12'hD66: dout  = 8'b01001111; // 3430 :  79 - 0x4f
      12'hD67: dout  = 8'b10001101; // 3431 : 141 - 0x8d
      12'hD68: dout  = 8'b10001111; // 3432 : 143 - 0x8f -- Background 0xad
      12'hD69: dout  = 8'b01001101; // 3433 :  77 - 0x4d
      12'hD6A: dout  = 8'b00101111; // 3434 :  47 - 0x2f
      12'hD6B: dout  = 8'b00011101; // 3435 :  29 - 0x1d
      12'hD6C: dout  = 8'b00011111; // 3436 :  31 - 0x1f
      12'hD6D: dout  = 8'b00101101; // 3437 :  45 - 0x2d
      12'hD6E: dout  = 8'b01001111; // 3438 :  79 - 0x4f
      12'hD6F: dout  = 8'b11111111; // 3439 : 255 - 0xff
      12'hD70: dout  = 8'b00000001; // 3440 :   1 - 0x1 -- Background 0xae
      12'hD71: dout  = 8'b00000011; // 3441 :   3 - 0x3
      12'hD72: dout  = 8'b00000110; // 3442 :   6 - 0x6
      12'hD73: dout  = 8'b00000111; // 3443 :   7 - 0x7
      12'hD74: dout  = 8'b00000111; // 3444 :   7 - 0x7
      12'hD75: dout  = 8'b00000111; // 3445 :   7 - 0x7
      12'hD76: dout  = 8'b00000110; // 3446 :   6 - 0x6
      12'hD77: dout  = 8'b00000111; // 3447 :   7 - 0x7
      12'hD78: dout  = 8'b00000110; // 3448 :   6 - 0x6 -- Background 0xaf
      12'hD79: dout  = 8'b00000110; // 3449 :   6 - 0x6
      12'hD7A: dout  = 8'b00001110; // 3450 :  14 - 0xe
      12'hD7B: dout  = 8'b00001111; // 3451 :  15 - 0xf
      12'hD7C: dout  = 8'b00001110; // 3452 :  14 - 0xe
      12'hD7D: dout  = 8'b00011010; // 3453 :  26 - 0x1a
      12'hD7E: dout  = 8'b00011011; // 3454 :  27 - 0x1b
      12'hD7F: dout  = 8'b00001111; // 3455 :  15 - 0xf
      12'hD80: dout  = 8'b00000000; // 3456 :   0 - 0x0 -- Background 0xb0
      12'hD81: dout  = 8'b11000000; // 3457 : 192 - 0xc0
      12'hD82: dout  = 8'b11110000; // 3458 : 240 - 0xf0
      12'hD83: dout  = 8'b10001000; // 3459 : 136 - 0x88
      12'hD84: dout  = 8'b00010100; // 3460 :  20 - 0x14
      12'hD85: dout  = 8'b01101000; // 3461 : 104 - 0x68
      12'hD86: dout  = 8'b10101000; // 3462 : 168 - 0xa8
      12'hD87: dout  = 8'b00101100; // 3463 :  44 - 0x2c
      12'hD88: dout  = 8'b00000100; // 3464 :   4 - 0x4 -- Background 0xb1
      12'hD89: dout  = 8'b00111000; // 3465 :  56 - 0x38
      12'hD8A: dout  = 8'b00010000; // 3466 :  16 - 0x10
      12'hD8B: dout  = 8'b10100000; // 3467 : 160 - 0xa0
      12'hD8C: dout  = 8'b01100000; // 3468 :  96 - 0x60
      12'hD8D: dout  = 8'b00100000; // 3469 :  32 - 0x20
      12'hD8E: dout  = 8'b00010000; // 3470 :  16 - 0x10
      12'hD8F: dout  = 8'b10001000; // 3471 : 136 - 0x88
      12'hD90: dout  = 8'b00001111; // 3472 :  15 - 0xf -- Background 0xb2
      12'hD91: dout  = 8'b00011011; // 3473 :  27 - 0x1b
      12'hD92: dout  = 8'b00011011; // 3474 :  27 - 0x1b
      12'hD93: dout  = 8'b00001110; // 3475 :  14 - 0xe
      12'hD94: dout  = 8'b00000110; // 3476 :   6 - 0x6
      12'hD95: dout  = 8'b00001100; // 3477 :  12 - 0xc
      12'hD96: dout  = 8'b00001100; // 3478 :  12 - 0xc
      12'hD97: dout  = 8'b00111111; // 3479 :  63 - 0x3f
      12'hD98: dout  = 8'b01111111; // 3480 : 127 - 0x7f -- Background 0xb3
      12'hD99: dout  = 8'b01100000; // 3481 :  96 - 0x60
      12'hD9A: dout  = 8'b01100000; // 3482 :  96 - 0x60
      12'hD9B: dout  = 8'b01100000; // 3483 :  96 - 0x60
      12'hD9C: dout  = 8'b01100000; // 3484 :  96 - 0x60
      12'hD9D: dout  = 8'b01100000; // 3485 :  96 - 0x60
      12'hD9E: dout  = 8'b01101010; // 3486 : 106 - 0x6a
      12'hD9F: dout  = 8'b01111111; // 3487 : 127 - 0x7f
      12'hDA0: dout  = 8'b01001000; // 3488 :  72 - 0x48 -- Background 0xb4
      12'hDA1: dout  = 8'b00110000; // 3489 :  48 - 0x30
      12'hDA2: dout  = 8'b00010000; // 3490 :  16 - 0x10
      12'hDA3: dout  = 8'b00010000; // 3491 :  16 - 0x10
      12'hDA4: dout  = 8'b00001000; // 3492 :   8 - 0x8
      12'hDA5: dout  = 8'b00001000; // 3493 :   8 - 0x8
      12'hDA6: dout  = 8'b00001000; // 3494 :   8 - 0x8
      12'hDA7: dout  = 8'b11111100; // 3495 : 252 - 0xfc
      12'hDA8: dout  = 8'b11111110; // 3496 : 254 - 0xfe -- Background 0xb5
      12'hDA9: dout  = 8'b00000110; // 3497 :   6 - 0x6
      12'hDAA: dout  = 8'b00000010; // 3498 :   2 - 0x2
      12'hDAB: dout  = 8'b00000110; // 3499 :   6 - 0x6
      12'hDAC: dout  = 8'b00000010; // 3500 :   2 - 0x2
      12'hDAD: dout  = 8'b00000110; // 3501 :   6 - 0x6
      12'hDAE: dout  = 8'b10101010; // 3502 : 170 - 0xaa
      12'hDAF: dout  = 8'b11111110; // 3503 : 254 - 0xfe
      12'hDB0: dout  = 8'b11111111; // 3504 : 255 - 0xff -- Background 0xb6
      12'hDB1: dout  = 8'b10000000; // 3505 : 128 - 0x80
      12'hDB2: dout  = 8'b10000000; // 3506 : 128 - 0x80
      12'hDB3: dout  = 8'b10000000; // 3507 : 128 - 0x80
      12'hDB4: dout  = 8'b10000000; // 3508 : 128 - 0x80
      12'hDB5: dout  = 8'b10000000; // 3509 : 128 - 0x80
      12'hDB6: dout  = 8'b10010101; // 3510 : 149 - 0x95
      12'hDB7: dout  = 8'b11111111; // 3511 : 255 - 0xff
      12'hDB8: dout  = 8'b11111111; // 3512 : 255 - 0xff -- Background 0xb7
      12'hDB9: dout  = 8'b10000100; // 3513 : 132 - 0x84
      12'hDBA: dout  = 8'b10001100; // 3514 : 140 - 0x8c
      12'hDBB: dout  = 8'b10000100; // 3515 : 132 - 0x84
      12'hDBC: dout  = 8'b10001100; // 3516 : 140 - 0x8c
      12'hDBD: dout  = 8'b10000100; // 3517 : 132 - 0x84
      12'hDBE: dout  = 8'b10101100; // 3518 : 172 - 0xac
      12'hDBF: dout  = 8'b11111111; // 3519 : 255 - 0xff
      12'hDC0: dout  = 8'b11111111; // 3520 : 255 - 0xff -- Background 0xb8
      12'hDC1: dout  = 8'b00100001; // 3521 :  33 - 0x21
      12'hDC2: dout  = 8'b01100001; // 3522 :  97 - 0x61
      12'hDC3: dout  = 8'b00100011; // 3523 :  35 - 0x23
      12'hDC4: dout  = 8'b01100001; // 3524 :  97 - 0x61
      12'hDC5: dout  = 8'b00100011; // 3525 :  35 - 0x23
      12'hDC6: dout  = 8'b01100101; // 3526 : 101 - 0x65
      12'hDC7: dout  = 8'b11111111; // 3527 : 255 - 0xff
      12'hDC8: dout  = 8'b11111111; // 3528 : 255 - 0xff -- Background 0xb9
      12'hDC9: dout  = 8'b00000001; // 3529 :   1 - 0x1
      12'hDCA: dout  = 8'b00000011; // 3530 :   3 - 0x3
      12'hDCB: dout  = 8'b00000001; // 3531 :   1 - 0x1
      12'hDCC: dout  = 8'b00000011; // 3532 :   3 - 0x3
      12'hDCD: dout  = 8'b00000001; // 3533 :   1 - 0x1
      12'hDCE: dout  = 8'b10101011; // 3534 : 171 - 0xab
      12'hDCF: dout  = 8'b11111111; // 3535 : 255 - 0xff
      12'hDD0: dout  = 8'b11111111; // 3536 : 255 - 0xff -- Background 0xba
      12'hDD1: dout  = 8'b11010101; // 3537 : 213 - 0xd5
      12'hDD2: dout  = 8'b10101010; // 3538 : 170 - 0xaa
      12'hDD3: dout  = 8'b11111111; // 3539 : 255 - 0xff
      12'hDD4: dout  = 8'b10000000; // 3540 : 128 - 0x80
      12'hDD5: dout  = 8'b10000000; // 3541 : 128 - 0x80
      12'hDD6: dout  = 8'b10010101; // 3542 : 149 - 0x95
      12'hDD7: dout  = 8'b11111111; // 3543 : 255 - 0xff
      12'hDD8: dout  = 8'b00000000; // 3544 :   0 - 0x0 -- Background 0xbb
      12'hDD9: dout  = 8'b00000000; // 3545 :   0 - 0x0
      12'hDDA: dout  = 8'b00000000; // 3546 :   0 - 0x0
      12'hDDB: dout  = 8'b00000000; // 3547 :   0 - 0x0
      12'hDDC: dout  = 8'b00000000; // 3548 :   0 - 0x0
      12'hDDD: dout  = 8'b00000000; // 3549 :   0 - 0x0
      12'hDDE: dout  = 8'b00000000; // 3550 :   0 - 0x0
      12'hDDF: dout  = 8'b00000000; // 3551 :   0 - 0x0
      12'hDE0: dout  = 8'b11111111; // 3552 : 255 - 0xff -- Background 0xbc
      12'hDE1: dout  = 8'b01010101; // 3553 :  85 - 0x55
      12'hDE2: dout  = 8'b10101011; // 3554 : 171 - 0xab
      12'hDE3: dout  = 8'b11111111; // 3555 : 255 - 0xff
      12'hDE4: dout  = 8'b01100001; // 3556 :  97 - 0x61
      12'hDE5: dout  = 8'b00100011; // 3557 :  35 - 0x23
      12'hDE6: dout  = 8'b01100101; // 3558 : 101 - 0x65
      12'hDE7: dout  = 8'b11111111; // 3559 : 255 - 0xff
      12'hDE8: dout  = 8'b00000000; // 3560 :   0 - 0x0 -- Background 0xbd
      12'hDE9: dout  = 8'b00000000; // 3561 :   0 - 0x0
      12'hDEA: dout  = 8'b00000000; // 3562 :   0 - 0x0
      12'hDEB: dout  = 8'b00000000; // 3563 :   0 - 0x0
      12'hDEC: dout  = 8'b00000000; // 3564 :   0 - 0x0
      12'hDED: dout  = 8'b00000000; // 3565 :   0 - 0x0
      12'hDEE: dout  = 8'b00000000; // 3566 :   0 - 0x0
      12'hDEF: dout  = 8'b00000000; // 3567 :   0 - 0x0
      12'hDF0: dout  = 8'b00000000; // 3568 :   0 - 0x0 -- Background 0xbe
      12'hDF1: dout  = 8'b00000000; // 3569 :   0 - 0x0
      12'hDF2: dout  = 8'b00000000; // 3570 :   0 - 0x0
      12'hDF3: dout  = 8'b00000000; // 3571 :   0 - 0x0
      12'hDF4: dout  = 8'b00000000; // 3572 :   0 - 0x0
      12'hDF5: dout  = 8'b00000000; // 3573 :   0 - 0x0
      12'hDF6: dout  = 8'b00000000; // 3574 :   0 - 0x0
      12'hDF7: dout  = 8'b00000000; // 3575 :   0 - 0x0
      12'hDF8: dout  = 8'b00000000; // 3576 :   0 - 0x0 -- Background 0xbf
      12'hDF9: dout  = 8'b00000000; // 3577 :   0 - 0x0
      12'hDFA: dout  = 8'b00000000; // 3578 :   0 - 0x0
      12'hDFB: dout  = 8'b00000000; // 3579 :   0 - 0x0
      12'hDFC: dout  = 8'b00000000; // 3580 :   0 - 0x0
      12'hDFD: dout  = 8'b00000000; // 3581 :   0 - 0x0
      12'hDFE: dout  = 8'b00000000; // 3582 :   0 - 0x0
      12'hDFF: dout  = 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout  = 8'b00000000; // 3584 :   0 - 0x0 -- Background 0xc0
      12'hE01: dout  = 8'b00000000; // 3585 :   0 - 0x0
      12'hE02: dout  = 8'b00000000; // 3586 :   0 - 0x0
      12'hE03: dout  = 8'b00000000; // 3587 :   0 - 0x0
      12'hE04: dout  = 8'b00000000; // 3588 :   0 - 0x0
      12'hE05: dout  = 8'b00000000; // 3589 :   0 - 0x0
      12'hE06: dout  = 8'b00000000; // 3590 :   0 - 0x0
      12'hE07: dout  = 8'b00000000; // 3591 :   0 - 0x0
      12'hE08: dout  = 8'b00000000; // 3592 :   0 - 0x0 -- Background 0xc1
      12'hE09: dout  = 8'b00000000; // 3593 :   0 - 0x0
      12'hE0A: dout  = 8'b00000000; // 3594 :   0 - 0x0
      12'hE0B: dout  = 8'b00000000; // 3595 :   0 - 0x0
      12'hE0C: dout  = 8'b00000000; // 3596 :   0 - 0x0
      12'hE0D: dout  = 8'b00000000; // 3597 :   0 - 0x0
      12'hE0E: dout  = 8'b00000000; // 3598 :   0 - 0x0
      12'hE0F: dout  = 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout  = 8'b00000000; // 3600 :   0 - 0x0 -- Background 0xc2
      12'hE11: dout  = 8'b00000000; // 3601 :   0 - 0x0
      12'hE12: dout  = 8'b00000000; // 3602 :   0 - 0x0
      12'hE13: dout  = 8'b00000000; // 3603 :   0 - 0x0
      12'hE14: dout  = 8'b00000000; // 3604 :   0 - 0x0
      12'hE15: dout  = 8'b00000000; // 3605 :   0 - 0x0
      12'hE16: dout  = 8'b00000000; // 3606 :   0 - 0x0
      12'hE17: dout  = 8'b00000000; // 3607 :   0 - 0x0
      12'hE18: dout  = 8'b00000000; // 3608 :   0 - 0x0 -- Background 0xc3
      12'hE19: dout  = 8'b00000000; // 3609 :   0 - 0x0
      12'hE1A: dout  = 8'b00000000; // 3610 :   0 - 0x0
      12'hE1B: dout  = 8'b00000000; // 3611 :   0 - 0x0
      12'hE1C: dout  = 8'b00000000; // 3612 :   0 - 0x0
      12'hE1D: dout  = 8'b00000000; // 3613 :   0 - 0x0
      12'hE1E: dout  = 8'b00000000; // 3614 :   0 - 0x0
      12'hE1F: dout  = 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout  = 8'b00000000; // 3616 :   0 - 0x0 -- Background 0xc4
      12'hE21: dout  = 8'b00000000; // 3617 :   0 - 0x0
      12'hE22: dout  = 8'b00000000; // 3618 :   0 - 0x0
      12'hE23: dout  = 8'b00000000; // 3619 :   0 - 0x0
      12'hE24: dout  = 8'b00000000; // 3620 :   0 - 0x0
      12'hE25: dout  = 8'b00000000; // 3621 :   0 - 0x0
      12'hE26: dout  = 8'b00000000; // 3622 :   0 - 0x0
      12'hE27: dout  = 8'b00000000; // 3623 :   0 - 0x0
      12'hE28: dout  = 8'b00000000; // 3624 :   0 - 0x0 -- Background 0xc5
      12'hE29: dout  = 8'b00000000; // 3625 :   0 - 0x0
      12'hE2A: dout  = 8'b00000001; // 3626 :   1 - 0x1
      12'hE2B: dout  = 8'b00000110; // 3627 :   6 - 0x6
      12'hE2C: dout  = 8'b00001010; // 3628 :  10 - 0xa
      12'hE2D: dout  = 8'b00010100; // 3629 :  20 - 0x14
      12'hE2E: dout  = 8'b00010000; // 3630 :  16 - 0x10
      12'hE2F: dout  = 8'b00101000; // 3631 :  40 - 0x28
      12'hE30: dout  = 8'b00011111; // 3632 :  31 - 0x1f -- Background 0xc6
      12'hE31: dout  = 8'b01100000; // 3633 :  96 - 0x60
      12'hE32: dout  = 8'b10100000; // 3634 : 160 - 0xa0
      12'hE33: dout  = 8'b01000000; // 3635 :  64 - 0x40
      12'hE34: dout  = 8'b00000000; // 3636 :   0 - 0x0
      12'hE35: dout  = 8'b00000000; // 3637 :   0 - 0x0
      12'hE36: dout  = 8'b00000000; // 3638 :   0 - 0x0
      12'hE37: dout  = 8'b00000000; // 3639 :   0 - 0x0
      12'hE38: dout  = 8'b00110000; // 3640 :  48 - 0x30 -- Background 0xc7
      12'hE39: dout  = 8'b01000000; // 3641 :  64 - 0x40
      12'hE3A: dout  = 8'b01100000; // 3642 :  96 - 0x60
      12'hE3B: dout  = 8'b11000000; // 3643 : 192 - 0xc0
      12'hE3C: dout  = 8'b10000000; // 3644 : 128 - 0x80
      12'hE3D: dout  = 8'b10100000; // 3645 : 160 - 0xa0
      12'hE3E: dout  = 8'b11000000; // 3646 : 192 - 0xc0
      12'hE3F: dout  = 8'b10000000; // 3647 : 128 - 0x80
      12'hE40: dout  = 8'b11111111; // 3648 : 255 - 0xff -- Background 0xc8
      12'hE41: dout  = 8'b00000000; // 3649 :   0 - 0x0
      12'hE42: dout  = 8'b00000000; // 3650 :   0 - 0x0
      12'hE43: dout  = 8'b00000000; // 3651 :   0 - 0x0
      12'hE44: dout  = 8'b00000000; // 3652 :   0 - 0x0
      12'hE45: dout  = 8'b00000000; // 3653 :   0 - 0x0
      12'hE46: dout  = 8'b00000000; // 3654 :   0 - 0x0
      12'hE47: dout  = 8'b00000000; // 3655 :   0 - 0x0
      12'hE48: dout  = 8'b00010100; // 3656 :  20 - 0x14 -- Background 0xc9
      12'hE49: dout  = 8'b00101010; // 3657 :  42 - 0x2a
      12'hE4A: dout  = 8'b00010110; // 3658 :  22 - 0x16
      12'hE4B: dout  = 8'b00101011; // 3659 :  43 - 0x2b
      12'hE4C: dout  = 8'b00010101; // 3660 :  21 - 0x15
      12'hE4D: dout  = 8'b00101011; // 3661 :  43 - 0x2b
      12'hE4E: dout  = 8'b00010101; // 3662 :  21 - 0x15
      12'hE4F: dout  = 8'b00101011; // 3663 :  43 - 0x2b
      12'hE50: dout  = 8'b00000000; // 3664 :   0 - 0x0 -- Background 0xca
      12'hE51: dout  = 8'b00000100; // 3665 :   4 - 0x4
      12'hE52: dout  = 8'b00000100; // 3666 :   4 - 0x4
      12'hE53: dout  = 8'b00000101; // 3667 :   5 - 0x5
      12'hE54: dout  = 8'b00010101; // 3668 :  21 - 0x15
      12'hE55: dout  = 8'b00010101; // 3669 :  21 - 0x15
      12'hE56: dout  = 8'b01010101; // 3670 :  85 - 0x55
      12'hE57: dout  = 8'b01010101; // 3671 :  85 - 0x55
      12'hE58: dout  = 8'b00000000; // 3672 :   0 - 0x0 -- Background 0xcb
      12'hE59: dout  = 8'b00000000; // 3673 :   0 - 0x0
      12'hE5A: dout  = 8'b00010000; // 3674 :  16 - 0x10
      12'hE5B: dout  = 8'b00010000; // 3675 :  16 - 0x10
      12'hE5C: dout  = 8'b01010001; // 3676 :  81 - 0x51
      12'hE5D: dout  = 8'b01010101; // 3677 :  85 - 0x55
      12'hE5E: dout  = 8'b01010101; // 3678 :  85 - 0x55
      12'hE5F: dout  = 8'b01010101; // 3679 :  85 - 0x55
      12'hE60: dout  = 8'b00000000; // 3680 :   0 - 0x0 -- Background 0xcc
      12'hE61: dout  = 8'b00000000; // 3681 :   0 - 0x0
      12'hE62: dout  = 8'b00000000; // 3682 :   0 - 0x0
      12'hE63: dout  = 8'b00000101; // 3683 :   5 - 0x5
      12'hE64: dout  = 8'b00001111; // 3684 :  15 - 0xf
      12'hE65: dout  = 8'b00000111; // 3685 :   7 - 0x7
      12'hE66: dout  = 8'b00000011; // 3686 :   3 - 0x3
      12'hE67: dout  = 8'b00000001; // 3687 :   1 - 0x1
      12'hE68: dout  = 8'b00000000; // 3688 :   0 - 0x0 -- Background 0xcd
      12'hE69: dout  = 8'b00000000; // 3689 :   0 - 0x0
      12'hE6A: dout  = 8'b10000000; // 3690 : 128 - 0x80
      12'hE6B: dout  = 8'b11010000; // 3691 : 208 - 0xd0
      12'hE6C: dout  = 8'b11111000; // 3692 : 248 - 0xf8
      12'hE6D: dout  = 8'b11110000; // 3693 : 240 - 0xf0
      12'hE6E: dout  = 8'b11100000; // 3694 : 224 - 0xe0
      12'hE6F: dout  = 8'b11000000; // 3695 : 192 - 0xc0
      12'hE70: dout  = 8'b00000000; // 3696 :   0 - 0x0 -- Background 0xce
      12'hE71: dout  = 8'b00000000; // 3697 :   0 - 0x0
      12'hE72: dout  = 8'b00000000; // 3698 :   0 - 0x0
      12'hE73: dout  = 8'b01111000; // 3699 : 120 - 0x78
      12'hE74: dout  = 8'b11001111; // 3700 : 207 - 0xcf
      12'hE75: dout  = 8'b10000000; // 3701 : 128 - 0x80
      12'hE76: dout  = 8'b11001111; // 3702 : 207 - 0xcf
      12'hE77: dout  = 8'b01001000; // 3703 :  72 - 0x48
      12'hE78: dout  = 8'b00000000; // 3704 :   0 - 0x0 -- Background 0xcf
      12'hE79: dout  = 8'b00000000; // 3705 :   0 - 0x0
      12'hE7A: dout  = 8'b00000000; // 3706 :   0 - 0x0
      12'hE7B: dout  = 8'b00011110; // 3707 :  30 - 0x1e
      12'hE7C: dout  = 8'b11110011; // 3708 : 243 - 0xf3
      12'hE7D: dout  = 8'b00000001; // 3709 :   1 - 0x1
      12'hE7E: dout  = 8'b11110011; // 3710 : 243 - 0xf3
      12'hE7F: dout  = 8'b00010010; // 3711 :  18 - 0x12
      12'hE80: dout  = 8'b00000000; // 3712 :   0 - 0x0 -- Background 0xd0
      12'hE81: dout  = 8'b00000000; // 3713 :   0 - 0x0
      12'hE82: dout  = 8'b00000000; // 3714 :   0 - 0x0
      12'hE83: dout  = 8'b00000000; // 3715 :   0 - 0x0
      12'hE84: dout  = 8'b00000000; // 3716 :   0 - 0x0
      12'hE85: dout  = 8'b00000000; // 3717 :   0 - 0x0
      12'hE86: dout  = 8'b00000000; // 3718 :   0 - 0x0
      12'hE87: dout  = 8'b00000000; // 3719 :   0 - 0x0
      12'hE88: dout  = 8'b00000000; // 3720 :   0 - 0x0 -- Background 0xd1
      12'hE89: dout  = 8'b00000000; // 3721 :   0 - 0x0
      12'hE8A: dout  = 8'b00000000; // 3722 :   0 - 0x0
      12'hE8B: dout  = 8'b00000000; // 3723 :   0 - 0x0
      12'hE8C: dout  = 8'b00000000; // 3724 :   0 - 0x0
      12'hE8D: dout  = 8'b00000000; // 3725 :   0 - 0x0
      12'hE8E: dout  = 8'b00000000; // 3726 :   0 - 0x0
      12'hE8F: dout  = 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout  = 8'b00001000; // 3728 :   8 - 0x8 -- Background 0xd2
      12'hE91: dout  = 8'b00001100; // 3729 :  12 - 0xc
      12'hE92: dout  = 8'b00001000; // 3730 :   8 - 0x8
      12'hE93: dout  = 8'b00001000; // 3731 :   8 - 0x8
      12'hE94: dout  = 8'b00001010; // 3732 :  10 - 0xa
      12'hE95: dout  = 8'b00001000; // 3733 :   8 - 0x8
      12'hE96: dout  = 8'b00001000; // 3734 :   8 - 0x8
      12'hE97: dout  = 8'b00001100; // 3735 :  12 - 0xc
      12'hE98: dout  = 8'b00010000; // 3736 :  16 - 0x10 -- Background 0xd3
      12'hE99: dout  = 8'b00010000; // 3737 :  16 - 0x10
      12'hE9A: dout  = 8'b00110000; // 3738 :  48 - 0x30
      12'hE9B: dout  = 8'b00010000; // 3739 :  16 - 0x10
      12'hE9C: dout  = 8'b01010000; // 3740 :  80 - 0x50
      12'hE9D: dout  = 8'b00010000; // 3741 :  16 - 0x10
      12'hE9E: dout  = 8'b00110000; // 3742 :  48 - 0x30
      12'hE9F: dout  = 8'b00010000; // 3743 :  16 - 0x10
      12'hEA0: dout  = 8'b00000000; // 3744 :   0 - 0x0 -- Background 0xd4
      12'hEA1: dout  = 8'b00000000; // 3745 :   0 - 0x0
      12'hEA2: dout  = 8'b00000000; // 3746 :   0 - 0x0
      12'hEA3: dout  = 8'b00000000; // 3747 :   0 - 0x0
      12'hEA4: dout  = 8'b00000000; // 3748 :   0 - 0x0
      12'hEA5: dout  = 8'b00000000; // 3749 :   0 - 0x0
      12'hEA6: dout  = 8'b00000000; // 3750 :   0 - 0x0
      12'hEA7: dout  = 8'b00000000; // 3751 :   0 - 0x0
      12'hEA8: dout  = 8'b11111000; // 3752 : 248 - 0xf8 -- Background 0xd5
      12'hEA9: dout  = 8'b00000110; // 3753 :   6 - 0x6
      12'hEAA: dout  = 8'b00000001; // 3754 :   1 - 0x1
      12'hEAB: dout  = 8'b00000000; // 3755 :   0 - 0x0
      12'hEAC: dout  = 8'b00000000; // 3756 :   0 - 0x0
      12'hEAD: dout  = 8'b00000000; // 3757 :   0 - 0x0
      12'hEAE: dout  = 8'b00000000; // 3758 :   0 - 0x0
      12'hEAF: dout  = 8'b00000000; // 3759 :   0 - 0x0
      12'hEB0: dout  = 8'b00000000; // 3760 :   0 - 0x0 -- Background 0xd6
      12'hEB1: dout  = 8'b00000000; // 3761 :   0 - 0x0
      12'hEB2: dout  = 8'b10000000; // 3762 : 128 - 0x80
      12'hEB3: dout  = 8'b01100000; // 3763 :  96 - 0x60
      12'hEB4: dout  = 8'b01010000; // 3764 :  80 - 0x50
      12'hEB5: dout  = 8'b10101000; // 3765 : 168 - 0xa8
      12'hEB6: dout  = 8'b01011000; // 3766 :  88 - 0x58
      12'hEB7: dout  = 8'b00101100; // 3767 :  44 - 0x2c
      12'hEB8: dout  = 8'b10100000; // 3768 : 160 - 0xa0 -- Background 0xd7
      12'hEB9: dout  = 8'b11000000; // 3769 : 192 - 0xc0
      12'hEBA: dout  = 8'b10000000; // 3770 : 128 - 0x80
      12'hEBB: dout  = 8'b01010000; // 3771 :  80 - 0x50
      12'hEBC: dout  = 8'b01100000; // 3772 :  96 - 0x60
      12'hEBD: dout  = 8'b00111000; // 3773 :  56 - 0x38
      12'hEBE: dout  = 8'b00001000; // 3774 :   8 - 0x8
      12'hEBF: dout  = 8'b00000111; // 3775 :   7 - 0x7
      12'hEC0: dout  = 8'b00000000; // 3776 :   0 - 0x0 -- Background 0xd8
      12'hEC1: dout  = 8'b00000000; // 3777 :   0 - 0x0
      12'hEC2: dout  = 8'b00000000; // 3778 :   0 - 0x0
      12'hEC3: dout  = 8'b00000000; // 3779 :   0 - 0x0
      12'hEC4: dout  = 8'b00000000; // 3780 :   0 - 0x0
      12'hEC5: dout  = 8'b00000000; // 3781 :   0 - 0x0
      12'hEC6: dout  = 8'b00000000; // 3782 :   0 - 0x0
      12'hEC7: dout  = 8'b11111111; // 3783 : 255 - 0xff
      12'hEC8: dout  = 8'b00010101; // 3784 :  21 - 0x15 -- Background 0xd9
      12'hEC9: dout  = 8'b00101011; // 3785 :  43 - 0x2b
      12'hECA: dout  = 8'b00010101; // 3786 :  21 - 0x15
      12'hECB: dout  = 8'b00101010; // 3787 :  42 - 0x2a
      12'hECC: dout  = 8'b01010110; // 3788 :  86 - 0x56
      12'hECD: dout  = 8'b10101100; // 3789 : 172 - 0xac
      12'hECE: dout  = 8'b01010000; // 3790 :  80 - 0x50
      12'hECF: dout  = 8'b11100000; // 3791 : 224 - 0xe0
      12'hED0: dout  = 8'b00000001; // 3792 :   1 - 0x1 -- Background 0xda
      12'hED1: dout  = 8'b00001101; // 3793 :  13 - 0xd
      12'hED2: dout  = 8'b00010011; // 3794 :  19 - 0x13
      12'hED3: dout  = 8'b00001101; // 3795 :  13 - 0xd
      12'hED4: dout  = 8'b00000001; // 3796 :   1 - 0x1
      12'hED5: dout  = 8'b00000001; // 3797 :   1 - 0x1
      12'hED6: dout  = 8'b00000001; // 3798 :   1 - 0x1
      12'hED7: dout  = 8'b00000001; // 3799 :   1 - 0x1
      12'hED8: dout  = 8'b11000000; // 3800 : 192 - 0xc0 -- Background 0xdb
      12'hED9: dout  = 8'b01000000; // 3801 :  64 - 0x40
      12'hEDA: dout  = 8'b01000000; // 3802 :  64 - 0x40
      12'hEDB: dout  = 8'b01011000; // 3803 :  88 - 0x58
      12'hEDC: dout  = 8'b01100100; // 3804 : 100 - 0x64
      12'hEDD: dout  = 8'b01011000; // 3805 :  88 - 0x58
      12'hEDE: dout  = 8'b01000000; // 3806 :  64 - 0x40
      12'hEDF: dout  = 8'b01000000; // 3807 :  64 - 0x40
      12'hEE0: dout  = 8'b00000000; // 3808 :   0 - 0x0 -- Background 0xdc
      12'hEE1: dout  = 8'b00000000; // 3809 :   0 - 0x0
      12'hEE2: dout  = 8'b00000000; // 3810 :   0 - 0x0
      12'hEE3: dout  = 8'b00000110; // 3811 :   6 - 0x6
      12'hEE4: dout  = 8'b00000111; // 3812 :   7 - 0x7
      12'hEE5: dout  = 8'b00000111; // 3813 :   7 - 0x7
      12'hEE6: dout  = 8'b00000111; // 3814 :   7 - 0x7
      12'hEE7: dout  = 8'b00000011; // 3815 :   3 - 0x3
      12'hEE8: dout  = 8'b00000000; // 3816 :   0 - 0x0 -- Background 0xdd
      12'hEE9: dout  = 8'b00000000; // 3817 :   0 - 0x0
      12'hEEA: dout  = 8'b00000000; // 3818 :   0 - 0x0
      12'hEEB: dout  = 8'b10110000; // 3819 : 176 - 0xb0
      12'hEEC: dout  = 8'b11110000; // 3820 : 240 - 0xf0
      12'hEED: dout  = 8'b11110000; // 3821 : 240 - 0xf0
      12'hEEE: dout  = 8'b11110000; // 3822 : 240 - 0xf0
      12'hEEF: dout  = 8'b11100000; // 3823 : 224 - 0xe0
      12'hEF0: dout  = 8'b11001111; // 3824 : 207 - 0xcf -- Background 0xde
      12'hEF1: dout  = 8'b10000000; // 3825 : 128 - 0x80
      12'hEF2: dout  = 8'b11001111; // 3826 : 207 - 0xcf
      12'hEF3: dout  = 8'b01001000; // 3827 :  72 - 0x48
      12'hEF4: dout  = 8'b01001000; // 3828 :  72 - 0x48
      12'hEF5: dout  = 8'b01001000; // 3829 :  72 - 0x48
      12'hEF6: dout  = 8'b01001000; // 3830 :  72 - 0x48
      12'hEF7: dout  = 8'b01001000; // 3831 :  72 - 0x48
      12'hEF8: dout  = 8'b11110011; // 3832 : 243 - 0xf3 -- Background 0xdf
      12'hEF9: dout  = 8'b00000001; // 3833 :   1 - 0x1
      12'hEFA: dout  = 8'b11110011; // 3834 : 243 - 0xf3
      12'hEFB: dout  = 8'b00010010; // 3835 :  18 - 0x12
      12'hEFC: dout  = 8'b00010010; // 3836 :  18 - 0x12
      12'hEFD: dout  = 8'b00010010; // 3837 :  18 - 0x12
      12'hEFE: dout  = 8'b00010010; // 3838 :  18 - 0x12
      12'hEFF: dout  = 8'b00010010; // 3839 :  18 - 0x12
      12'hF00: dout  = 8'b00000000; // 3840 :   0 - 0x0 -- Background 0xe0
      12'hF01: dout  = 8'b00000000; // 3841 :   0 - 0x0
      12'hF02: dout  = 8'b00000000; // 3842 :   0 - 0x0
      12'hF03: dout  = 8'b00000000; // 3843 :   0 - 0x0
      12'hF04: dout  = 8'b00000000; // 3844 :   0 - 0x0
      12'hF05: dout  = 8'b00000000; // 3845 :   0 - 0x0
      12'hF06: dout  = 8'b00000000; // 3846 :   0 - 0x0
      12'hF07: dout  = 8'b00000000; // 3847 :   0 - 0x0
      12'hF08: dout  = 8'b00000000; // 3848 :   0 - 0x0 -- Background 0xe1
      12'hF09: dout  = 8'b00000000; // 3849 :   0 - 0x0
      12'hF0A: dout  = 8'b00000000; // 3850 :   0 - 0x0
      12'hF0B: dout  = 8'b00000000; // 3851 :   0 - 0x0
      12'hF0C: dout  = 8'b00000000; // 3852 :   0 - 0x0
      12'hF0D: dout  = 8'b00000000; // 3853 :   0 - 0x0
      12'hF0E: dout  = 8'b00000000; // 3854 :   0 - 0x0
      12'hF0F: dout  = 8'b00000000; // 3855 :   0 - 0x0
      12'hF10: dout  = 8'b00000000; // 3856 :   0 - 0x0 -- Background 0xe2
      12'hF11: dout  = 8'b00000000; // 3857 :   0 - 0x0
      12'hF12: dout  = 8'b00000000; // 3858 :   0 - 0x0
      12'hF13: dout  = 8'b00000000; // 3859 :   0 - 0x0
      12'hF14: dout  = 8'b00000000; // 3860 :   0 - 0x0
      12'hF15: dout  = 8'b00000000; // 3861 :   0 - 0x0
      12'hF16: dout  = 8'b00000000; // 3862 :   0 - 0x0
      12'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout  = 8'b00000000; // 3864 :   0 - 0x0 -- Background 0xe3
      12'hF19: dout  = 8'b00000000; // 3865 :   0 - 0x0
      12'hF1A: dout  = 8'b00000000; // 3866 :   0 - 0x0
      12'hF1B: dout  = 8'b00000000; // 3867 :   0 - 0x0
      12'hF1C: dout  = 8'b00000000; // 3868 :   0 - 0x0
      12'hF1D: dout  = 8'b00000000; // 3869 :   0 - 0x0
      12'hF1E: dout  = 8'b00000000; // 3870 :   0 - 0x0
      12'hF1F: dout  = 8'b00000000; // 3871 :   0 - 0x0
      12'hF20: dout  = 8'b00000000; // 3872 :   0 - 0x0 -- Background 0xe4
      12'hF21: dout  = 8'b00000000; // 3873 :   0 - 0x0
      12'hF22: dout  = 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout  = 8'b00000000; // 3875 :   0 - 0x0
      12'hF24: dout  = 8'b00000000; // 3876 :   0 - 0x0
      12'hF25: dout  = 8'b00000000; // 3877 :   0 - 0x0
      12'hF26: dout  = 8'b00000000; // 3878 :   0 - 0x0
      12'hF27: dout  = 8'b00000000; // 3879 :   0 - 0x0
      12'hF28: dout  = 8'b00000000; // 3880 :   0 - 0x0 -- Background 0xe5
      12'hF29: dout  = 8'b00000000; // 3881 :   0 - 0x0
      12'hF2A: dout  = 8'b00000000; // 3882 :   0 - 0x0
      12'hF2B: dout  = 8'b00000000; // 3883 :   0 - 0x0
      12'hF2C: dout  = 8'b00000000; // 3884 :   0 - 0x0
      12'hF2D: dout  = 8'b00000000; // 3885 :   0 - 0x0
      12'hF2E: dout  = 8'b00000000; // 3886 :   0 - 0x0
      12'hF2F: dout  = 8'b00000000; // 3887 :   0 - 0x0
      12'hF30: dout  = 8'b00000000; // 3888 :   0 - 0x0 -- Background 0xe6
      12'hF31: dout  = 8'b00000000; // 3889 :   0 - 0x0
      12'hF32: dout  = 8'b00000000; // 3890 :   0 - 0x0
      12'hF33: dout  = 8'b00000000; // 3891 :   0 - 0x0
      12'hF34: dout  = 8'b00000000; // 3892 :   0 - 0x0
      12'hF35: dout  = 8'b00000000; // 3893 :   0 - 0x0
      12'hF36: dout  = 8'b00000000; // 3894 :   0 - 0x0
      12'hF37: dout  = 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout  = 8'b00000000; // 3896 :   0 - 0x0 -- Background 0xe7
      12'hF39: dout  = 8'b00000000; // 3897 :   0 - 0x0
      12'hF3A: dout  = 8'b00000000; // 3898 :   0 - 0x0
      12'hF3B: dout  = 8'b00000000; // 3899 :   0 - 0x0
      12'hF3C: dout  = 8'b00000000; // 3900 :   0 - 0x0
      12'hF3D: dout  = 8'b00000000; // 3901 :   0 - 0x0
      12'hF3E: dout  = 8'b00000000; // 3902 :   0 - 0x0
      12'hF3F: dout  = 8'b00000000; // 3903 :   0 - 0x0
      12'hF40: dout  = 8'b00000000; // 3904 :   0 - 0x0 -- Background 0xe8
      12'hF41: dout  = 8'b00000000; // 3905 :   0 - 0x0
      12'hF42: dout  = 8'b00000000; // 3906 :   0 - 0x0
      12'hF43: dout  = 8'b00000000; // 3907 :   0 - 0x0
      12'hF44: dout  = 8'b00000000; // 3908 :   0 - 0x0
      12'hF45: dout  = 8'b00000000; // 3909 :   0 - 0x0
      12'hF46: dout  = 8'b00000000; // 3910 :   0 - 0x0
      12'hF47: dout  = 8'b00000000; // 3911 :   0 - 0x0
      12'hF48: dout  = 8'b00000000; // 3912 :   0 - 0x0 -- Background 0xe9
      12'hF49: dout  = 8'b00000000; // 3913 :   0 - 0x0
      12'hF4A: dout  = 8'b00000000; // 3914 :   0 - 0x0
      12'hF4B: dout  = 8'b00000000; // 3915 :   0 - 0x0
      12'hF4C: dout  = 8'b00000000; // 3916 :   0 - 0x0
      12'hF4D: dout  = 8'b00000000; // 3917 :   0 - 0x0
      12'hF4E: dout  = 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout  = 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout  = 8'b00000000; // 3920 :   0 - 0x0 -- Background 0xea
      12'hF51: dout  = 8'b00000000; // 3921 :   0 - 0x0
      12'hF52: dout  = 8'b00000000; // 3922 :   0 - 0x0
      12'hF53: dout  = 8'b00000000; // 3923 :   0 - 0x0
      12'hF54: dout  = 8'b00000000; // 3924 :   0 - 0x0
      12'hF55: dout  = 8'b00000000; // 3925 :   0 - 0x0
      12'hF56: dout  = 8'b00000000; // 3926 :   0 - 0x0
      12'hF57: dout  = 8'b00000000; // 3927 :   0 - 0x0
      12'hF58: dout  = 8'b00000000; // 3928 :   0 - 0x0 -- Background 0xeb
      12'hF59: dout  = 8'b00000000; // 3929 :   0 - 0x0
      12'hF5A: dout  = 8'b00000000; // 3930 :   0 - 0x0
      12'hF5B: dout  = 8'b00000000; // 3931 :   0 - 0x0
      12'hF5C: dout  = 8'b00000000; // 3932 :   0 - 0x0
      12'hF5D: dout  = 8'b00000000; // 3933 :   0 - 0x0
      12'hF5E: dout  = 8'b00000000; // 3934 :   0 - 0x0
      12'hF5F: dout  = 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout  = 8'b00000000; // 3936 :   0 - 0x0 -- Background 0xec
      12'hF61: dout  = 8'b00000000; // 3937 :   0 - 0x0
      12'hF62: dout  = 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout  = 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout  = 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout  = 8'b00000000; // 3941 :   0 - 0x0
      12'hF66: dout  = 8'b00000000; // 3942 :   0 - 0x0
      12'hF67: dout  = 8'b00000000; // 3943 :   0 - 0x0
      12'hF68: dout  = 8'b00000000; // 3944 :   0 - 0x0 -- Background 0xed
      12'hF69: dout  = 8'b00000000; // 3945 :   0 - 0x0
      12'hF6A: dout  = 8'b00000000; // 3946 :   0 - 0x0
      12'hF6B: dout  = 8'b00000000; // 3947 :   0 - 0x0
      12'hF6C: dout  = 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout  = 8'b00000000; // 3949 :   0 - 0x0
      12'hF6E: dout  = 8'b00000000; // 3950 :   0 - 0x0
      12'hF6F: dout  = 8'b00000000; // 3951 :   0 - 0x0
      12'hF70: dout  = 8'b00000000; // 3952 :   0 - 0x0 -- Background 0xee
      12'hF71: dout  = 8'b00000000; // 3953 :   0 - 0x0
      12'hF72: dout  = 8'b00000000; // 3954 :   0 - 0x0
      12'hF73: dout  = 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout  = 8'b00000000; // 3956 :   0 - 0x0
      12'hF75: dout  = 8'b00000000; // 3957 :   0 - 0x0
      12'hF76: dout  = 8'b00000000; // 3958 :   0 - 0x0
      12'hF77: dout  = 8'b00000000; // 3959 :   0 - 0x0
      12'hF78: dout  = 8'b00000000; // 3960 :   0 - 0x0 -- Background 0xef
      12'hF79: dout  = 8'b00000000; // 3961 :   0 - 0x0
      12'hF7A: dout  = 8'b00000000; // 3962 :   0 - 0x0
      12'hF7B: dout  = 8'b00000000; // 3963 :   0 - 0x0
      12'hF7C: dout  = 8'b00000000; // 3964 :   0 - 0x0
      12'hF7D: dout  = 8'b00000000; // 3965 :   0 - 0x0
      12'hF7E: dout  = 8'b00000000; // 3966 :   0 - 0x0
      12'hF7F: dout  = 8'b00000000; // 3967 :   0 - 0x0
      12'hF80: dout  = 8'b00000000; // 3968 :   0 - 0x0 -- Background 0xf0
      12'hF81: dout  = 8'b00000000; // 3969 :   0 - 0x0
      12'hF82: dout  = 8'b00000000; // 3970 :   0 - 0x0
      12'hF83: dout  = 8'b00000000; // 3971 :   0 - 0x0
      12'hF84: dout  = 8'b00000000; // 3972 :   0 - 0x0
      12'hF85: dout  = 8'b00000000; // 3973 :   0 - 0x0
      12'hF86: dout  = 8'b00000000; // 3974 :   0 - 0x0
      12'hF87: dout  = 8'b00000000; // 3975 :   0 - 0x0
      12'hF88: dout  = 8'b00000000; // 3976 :   0 - 0x0 -- Background 0xf1
      12'hF89: dout  = 8'b00000000; // 3977 :   0 - 0x0
      12'hF8A: dout  = 8'b00000000; // 3978 :   0 - 0x0
      12'hF8B: dout  = 8'b00000000; // 3979 :   0 - 0x0
      12'hF8C: dout  = 8'b00000000; // 3980 :   0 - 0x0
      12'hF8D: dout  = 8'b00000000; // 3981 :   0 - 0x0
      12'hF8E: dout  = 8'b00000000; // 3982 :   0 - 0x0
      12'hF8F: dout  = 8'b00000000; // 3983 :   0 - 0x0
      12'hF90: dout  = 8'b00000000; // 3984 :   0 - 0x0 -- Background 0xf2
      12'hF91: dout  = 8'b00000000; // 3985 :   0 - 0x0
      12'hF92: dout  = 8'b00000000; // 3986 :   0 - 0x0
      12'hF93: dout  = 8'b00000000; // 3987 :   0 - 0x0
      12'hF94: dout  = 8'b00000000; // 3988 :   0 - 0x0
      12'hF95: dout  = 8'b00000000; // 3989 :   0 - 0x0
      12'hF96: dout  = 8'b00000000; // 3990 :   0 - 0x0
      12'hF97: dout  = 8'b00000000; // 3991 :   0 - 0x0
      12'hF98: dout  = 8'b00000000; // 3992 :   0 - 0x0 -- Background 0xf3
      12'hF99: dout  = 8'b00000000; // 3993 :   0 - 0x0
      12'hF9A: dout  = 8'b00000000; // 3994 :   0 - 0x0
      12'hF9B: dout  = 8'b00000000; // 3995 :   0 - 0x0
      12'hF9C: dout  = 8'b00000000; // 3996 :   0 - 0x0
      12'hF9D: dout  = 8'b00000000; // 3997 :   0 - 0x0
      12'hF9E: dout  = 8'b00000000; // 3998 :   0 - 0x0
      12'hF9F: dout  = 8'b00000000; // 3999 :   0 - 0x0
      12'hFA0: dout  = 8'b00000000; // 4000 :   0 - 0x0 -- Background 0xf4
      12'hFA1: dout  = 8'b00000000; // 4001 :   0 - 0x0
      12'hFA2: dout  = 8'b00000000; // 4002 :   0 - 0x0
      12'hFA3: dout  = 8'b00000000; // 4003 :   0 - 0x0
      12'hFA4: dout  = 8'b00000000; // 4004 :   0 - 0x0
      12'hFA5: dout  = 8'b00000000; // 4005 :   0 - 0x0
      12'hFA6: dout  = 8'b00000000; // 4006 :   0 - 0x0
      12'hFA7: dout  = 8'b00000000; // 4007 :   0 - 0x0
      12'hFA8: dout  = 8'b00000000; // 4008 :   0 - 0x0 -- Background 0xf5
      12'hFA9: dout  = 8'b00000000; // 4009 :   0 - 0x0
      12'hFAA: dout  = 8'b00000000; // 4010 :   0 - 0x0
      12'hFAB: dout  = 8'b00000000; // 4011 :   0 - 0x0
      12'hFAC: dout  = 8'b00000000; // 4012 :   0 - 0x0
      12'hFAD: dout  = 8'b00000000; // 4013 :   0 - 0x0
      12'hFAE: dout  = 8'b00000000; // 4014 :   0 - 0x0
      12'hFAF: dout  = 8'b00000000; // 4015 :   0 - 0x0
      12'hFB0: dout  = 8'b00000000; // 4016 :   0 - 0x0 -- Background 0xf6
      12'hFB1: dout  = 8'b00000000; // 4017 :   0 - 0x0
      12'hFB2: dout  = 8'b00000000; // 4018 :   0 - 0x0
      12'hFB3: dout  = 8'b00000000; // 4019 :   0 - 0x0
      12'hFB4: dout  = 8'b00000000; // 4020 :   0 - 0x0
      12'hFB5: dout  = 8'b00000000; // 4021 :   0 - 0x0
      12'hFB6: dout  = 8'b00000000; // 4022 :   0 - 0x0
      12'hFB7: dout  = 8'b00000000; // 4023 :   0 - 0x0
      12'hFB8: dout  = 8'b00000000; // 4024 :   0 - 0x0 -- Background 0xf7
      12'hFB9: dout  = 8'b00000000; // 4025 :   0 - 0x0
      12'hFBA: dout  = 8'b00000000; // 4026 :   0 - 0x0
      12'hFBB: dout  = 8'b00000000; // 4027 :   0 - 0x0
      12'hFBC: dout  = 8'b00000000; // 4028 :   0 - 0x0
      12'hFBD: dout  = 8'b00000000; // 4029 :   0 - 0x0
      12'hFBE: dout  = 8'b00000000; // 4030 :   0 - 0x0
      12'hFBF: dout  = 8'b00000000; // 4031 :   0 - 0x0
      12'hFC0: dout  = 8'b00000000; // 4032 :   0 - 0x0 -- Background 0xf8
      12'hFC1: dout  = 8'b00000000; // 4033 :   0 - 0x0
      12'hFC2: dout  = 8'b00000000; // 4034 :   0 - 0x0
      12'hFC3: dout  = 8'b00000000; // 4035 :   0 - 0x0
      12'hFC4: dout  = 8'b00000000; // 4036 :   0 - 0x0
      12'hFC5: dout  = 8'b00000000; // 4037 :   0 - 0x0
      12'hFC6: dout  = 8'b00000000; // 4038 :   0 - 0x0
      12'hFC7: dout  = 8'b00000000; // 4039 :   0 - 0x0
      12'hFC8: dout  = 8'b00000000; // 4040 :   0 - 0x0 -- Background 0xf9
      12'hFC9: dout  = 8'b00000000; // 4041 :   0 - 0x0
      12'hFCA: dout  = 8'b00000000; // 4042 :   0 - 0x0
      12'hFCB: dout  = 8'b00000000; // 4043 :   0 - 0x0
      12'hFCC: dout  = 8'b00000000; // 4044 :   0 - 0x0
      12'hFCD: dout  = 8'b00000000; // 4045 :   0 - 0x0
      12'hFCE: dout  = 8'b00000000; // 4046 :   0 - 0x0
      12'hFCF: dout  = 8'b00000000; // 4047 :   0 - 0x0
      12'hFD0: dout  = 8'b00000000; // 4048 :   0 - 0x0 -- Background 0xfa
      12'hFD1: dout  = 8'b00000000; // 4049 :   0 - 0x0
      12'hFD2: dout  = 8'b00000000; // 4050 :   0 - 0x0
      12'hFD3: dout  = 8'b00000000; // 4051 :   0 - 0x0
      12'hFD4: dout  = 8'b00000000; // 4052 :   0 - 0x0
      12'hFD5: dout  = 8'b00000000; // 4053 :   0 - 0x0
      12'hFD6: dout  = 8'b00000000; // 4054 :   0 - 0x0
      12'hFD7: dout  = 8'b00000000; // 4055 :   0 - 0x0
      12'hFD8: dout  = 8'b00000000; // 4056 :   0 - 0x0 -- Background 0xfb
      12'hFD9: dout  = 8'b00000000; // 4057 :   0 - 0x0
      12'hFDA: dout  = 8'b00000000; // 4058 :   0 - 0x0
      12'hFDB: dout  = 8'b00000000; // 4059 :   0 - 0x0
      12'hFDC: dout  = 8'b00000000; // 4060 :   0 - 0x0
      12'hFDD: dout  = 8'b00000000; // 4061 :   0 - 0x0
      12'hFDE: dout  = 8'b00000000; // 4062 :   0 - 0x0
      12'hFDF: dout  = 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout  = 8'b00000000; // 4064 :   0 - 0x0 -- Background 0xfc
      12'hFE1: dout  = 8'b00000000; // 4065 :   0 - 0x0
      12'hFE2: dout  = 8'b10001110; // 4066 : 142 - 0x8e
      12'hFE3: dout  = 8'b10001010; // 4067 : 138 - 0x8a
      12'hFE4: dout  = 8'b10001010; // 4068 : 138 - 0x8a
      12'hFE5: dout  = 8'b10001010; // 4069 : 138 - 0x8a
      12'hFE6: dout  = 8'b10001010; // 4070 : 138 - 0x8a
      12'hFE7: dout  = 8'b11101110; // 4071 : 238 - 0xee
      12'hFE8: dout  = 8'b00000000; // 4072 :   0 - 0x0 -- Background 0xfd
      12'hFE9: dout  = 8'b00000000; // 4073 :   0 - 0x0
      12'hFEA: dout  = 8'b01001100; // 4074 :  76 - 0x4c
      12'hFEB: dout  = 8'b10101010; // 4075 : 170 - 0xaa
      12'hFEC: dout  = 8'b10101010; // 4076 : 170 - 0xaa
      12'hFED: dout  = 8'b11101010; // 4077 : 234 - 0xea
      12'hFEE: dout  = 8'b10101010; // 4078 : 170 - 0xaa
      12'hFEF: dout  = 8'b10101100; // 4079 : 172 - 0xac
      12'hFF0: dout  = 8'b00000000; // 4080 :   0 - 0x0 -- Background 0xfe
      12'hFF1: dout  = 8'b00000000; // 4081 :   0 - 0x0
      12'hFF2: dout  = 8'b11101100; // 4082 : 236 - 0xec
      12'hFF3: dout  = 8'b01001010; // 4083 :  74 - 0x4a
      12'hFF4: dout  = 8'b01001010; // 4084 :  74 - 0x4a
      12'hFF5: dout  = 8'b01001010; // 4085 :  74 - 0x4a
      12'hFF6: dout  = 8'b01001010; // 4086 :  74 - 0x4a
      12'hFF7: dout  = 8'b11101010; // 4087 : 234 - 0xea
      12'hFF8: dout  = 8'b00000000; // 4088 :   0 - 0x0 -- Background 0xff
      12'hFF9: dout  = 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout  = 8'b01100000; // 4090 :  96 - 0x60
      12'hFFB: dout  = 8'b10001000; // 4091 : 136 - 0x88
      12'hFFC: dout  = 8'b10100000; // 4092 : 160 - 0xa0
      12'hFFD: dout  = 8'b10100000; // 4093 : 160 - 0xa0
      12'hFFE: dout  = 8'b10101000; // 4094 : 168 - 0xa8
      12'hFFF: dout  = 8'b01000000; // 4095 :  64 - 0x40
    endcase
  end

endmodule
