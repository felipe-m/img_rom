--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables


---  Original memory dump file name: smario_ntable_01.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_SMARIO_01 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_SMARIO_01;

architecture BEHAVIORAL of ROM_NTABLE_SMARIO_01 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "00100100", --    0 -  0x0  :   36 - 0x24
    "00100100", --    1 -  0x1  :   36 - 0x24
    "00100100", --    2 -  0x2  :   36 - 0x24
    "00100100", --    3 -  0x3  :   36 - 0x24
    "00100100", --    4 -  0x4  :   36 - 0x24
    "00100100", --    5 -  0x5  :   36 - 0x24
    "00100100", --    6 -  0x6  :   36 - 0x24
    "00100100", --    7 -  0x7  :   36 - 0x24
    "00100100", --    8 -  0x8  :   36 - 0x24
    "00100100", --    9 -  0x9  :   36 - 0x24
    "00100100", --   10 -  0xa  :   36 - 0x24
    "00100100", --   11 -  0xb  :   36 - 0x24
    "00100100", --   12 -  0xc  :   36 - 0x24
    "00100100", --   13 -  0xd  :   36 - 0x24
    "00100100", --   14 -  0xe  :   36 - 0x24
    "00100100", --   15 -  0xf  :   36 - 0x24
    "00100100", --   16 - 0x10  :   36 - 0x24
    "00100100", --   17 - 0x11  :   36 - 0x24
    "00100100", --   18 - 0x12  :   36 - 0x24
    "00100100", --   19 - 0x13  :   36 - 0x24
    "00100100", --   20 - 0x14  :   36 - 0x24
    "00100100", --   21 - 0x15  :   36 - 0x24
    "00100100", --   22 - 0x16  :   36 - 0x24
    "00100100", --   23 - 0x17  :   36 - 0x24
    "00100100", --   24 - 0x18  :   36 - 0x24
    "00100100", --   25 - 0x19  :   36 - 0x24
    "00100100", --   26 - 0x1a  :   36 - 0x24
    "00100100", --   27 - 0x1b  :   36 - 0x24
    "00100100", --   28 - 0x1c  :   36 - 0x24
    "00100100", --   29 - 0x1d  :   36 - 0x24
    "00100100", --   30 - 0x1e  :   36 - 0x24
    "00100100", --   31 - 0x1f  :   36 - 0x24
    "00100100", --   32 - 0x20  :   36 - 0x24
    "00100100", --   33 - 0x21  :   36 - 0x24
    "00100100", --   34 - 0x22  :   36 - 0x24
    "00100100", --   35 - 0x23  :   36 - 0x24
    "00100100", --   36 - 0x24  :   36 - 0x24
    "00100100", --   37 - 0x25  :   36 - 0x24
    "00100100", --   38 - 0x26  :   36 - 0x24
    "00100100", --   39 - 0x27  :   36 - 0x24
    "00100100", --   40 - 0x28  :   36 - 0x24
    "00100100", --   41 - 0x29  :   36 - 0x24
    "00100100", --   42 - 0x2a  :   36 - 0x24
    "00100100", --   43 - 0x2b  :   36 - 0x24
    "00100100", --   44 - 0x2c  :   36 - 0x24
    "00100100", --   45 - 0x2d  :   36 - 0x24
    "00100100", --   46 - 0x2e  :   36 - 0x24
    "00100100", --   47 - 0x2f  :   36 - 0x24
    "00100100", --   48 - 0x30  :   36 - 0x24
    "00100100", --   49 - 0x31  :   36 - 0x24
    "00100100", --   50 - 0x32  :   36 - 0x24
    "00100100", --   51 - 0x33  :   36 - 0x24
    "00100100", --   52 - 0x34  :   36 - 0x24
    "00100100", --   53 - 0x35  :   36 - 0x24
    "00100100", --   54 - 0x36  :   36 - 0x24
    "00100100", --   55 - 0x37  :   36 - 0x24
    "00100100", --   56 - 0x38  :   36 - 0x24
    "00100100", --   57 - 0x39  :   36 - 0x24
    "00100100", --   58 - 0x3a  :   36 - 0x24
    "00100100", --   59 - 0x3b  :   36 - 0x24
    "00100100", --   60 - 0x3c  :   36 - 0x24
    "00100100", --   61 - 0x3d  :   36 - 0x24
    "00100100", --   62 - 0x3e  :   36 - 0x24
    "00100100", --   63 - 0x3f  :   36 - 0x24
    "00100100", --   64 - 0x40  :   36 - 0x24
    "00100100", --   65 - 0x41  :   36 - 0x24
    "00100100", --   66 - 0x42  :   36 - 0x24
    "00010110", --   67 - 0x43  :   22 - 0x16
    "00001010", --   68 - 0x44  :   10 - 0xa
    "00011011", --   69 - 0x45  :   27 - 0x1b
    "00010010", --   70 - 0x46  :   18 - 0x12
    "00011000", --   71 - 0x47  :   24 - 0x18
    "00100100", --   72 - 0x48  :   36 - 0x24
    "00100100", --   73 - 0x49  :   36 - 0x24
    "00100100", --   74 - 0x4a  :   36 - 0x24
    "00100100", --   75 - 0x4b  :   36 - 0x24
    "00100100", --   76 - 0x4c  :   36 - 0x24
    "00100100", --   77 - 0x4d  :   36 - 0x24
    "00100100", --   78 - 0x4e  :   36 - 0x24
    "00100100", --   79 - 0x4f  :   36 - 0x24
    "00100100", --   80 - 0x50  :   36 - 0x24
    "00100100", --   81 - 0x51  :   36 - 0x24
    "00100000", --   82 - 0x52  :   32 - 0x20
    "00011000", --   83 - 0x53  :   24 - 0x18
    "00011011", --   84 - 0x54  :   27 - 0x1b
    "00010101", --   85 - 0x55  :   21 - 0x15
    "00001101", --   86 - 0x56  :   13 - 0xd
    "00100100", --   87 - 0x57  :   36 - 0x24
    "00100100", --   88 - 0x58  :   36 - 0x24
    "00011101", --   89 - 0x59  :   29 - 0x1d
    "00010010", --   90 - 0x5a  :   18 - 0x12
    "00010110", --   91 - 0x5b  :   22 - 0x16
    "00001110", --   92 - 0x5c  :   14 - 0xe
    "00100100", --   93 - 0x5d  :   36 - 0x24
    "00100100", --   94 - 0x5e  :   36 - 0x24
    "00100100", --   95 - 0x5f  :   36 - 0x24
    "00100100", --   96 - 0x60  :   36 - 0x24
    "00100100", --   97 - 0x61  :   36 - 0x24
    "00100100", --   98 - 0x62  :   36 - 0x24
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0
    "00100100", --  105 - 0x69  :   36 - 0x24
    "00100100", --  106 - 0x6a  :   36 - 0x24
    "00101110", --  107 - 0x6b  :   46 - 0x2e
    "00101001", --  108 - 0x6c  :   41 - 0x29
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00100100", --  111 - 0x6f  :   36 - 0x24
    "00100100", --  112 - 0x70  :   36 - 0x24
    "00100100", --  113 - 0x71  :   36 - 0x24
    "00100100", --  114 - 0x72  :   36 - 0x24
    "00000001", --  115 - 0x73  :    1 - 0x1
    "00101000", --  116 - 0x74  :   40 - 0x28
    "00000001", --  117 - 0x75  :    1 - 0x1
    "00100100", --  118 - 0x76  :   36 - 0x24
    "00100100", --  119 - 0x77  :   36 - 0x24
    "00100100", --  120 - 0x78  :   36 - 0x24
    "00100100", --  121 - 0x79  :   36 - 0x24
    "00100100", --  122 - 0x7a  :   36 - 0x24
    "00100100", --  123 - 0x7b  :   36 - 0x24
    "00100100", --  124 - 0x7c  :   36 - 0x24
    "00100100", --  125 - 0x7d  :   36 - 0x24
    "00100100", --  126 - 0x7e  :   36 - 0x24
    "00100100", --  127 - 0x7f  :   36 - 0x24
    "00100100", --  128 - 0x80  :   36 - 0x24
    "00100100", --  129 - 0x81  :   36 - 0x24
    "00100100", --  130 - 0x82  :   36 - 0x24
    "00100100", --  131 - 0x83  :   36 - 0x24
    "00100100", --  132 - 0x84  :   36 - 0x24
    "01000100", --  133 - 0x85  :   68 - 0x44
    "01001000", --  134 - 0x86  :   72 - 0x48
    "01001000", --  135 - 0x87  :   72 - 0x48
    "01001000", --  136 - 0x88  :   72 - 0x48
    "01001000", --  137 - 0x89  :   72 - 0x48
    "01001000", --  138 - 0x8a  :   72 - 0x48
    "01001000", --  139 - 0x8b  :   72 - 0x48
    "01001000", --  140 - 0x8c  :   72 - 0x48
    "01001000", --  141 - 0x8d  :   72 - 0x48
    "01001000", --  142 - 0x8e  :   72 - 0x48
    "01001000", --  143 - 0x8f  :   72 - 0x48
    "01001000", --  144 - 0x90  :   72 - 0x48
    "01001000", --  145 - 0x91  :   72 - 0x48
    "01001000", --  146 - 0x92  :   72 - 0x48
    "01001000", --  147 - 0x93  :   72 - 0x48
    "01001000", --  148 - 0x94  :   72 - 0x48
    "01001000", --  149 - 0x95  :   72 - 0x48
    "01001000", --  150 - 0x96  :   72 - 0x48
    "01001000", --  151 - 0x97  :   72 - 0x48
    "01001000", --  152 - 0x98  :   72 - 0x48
    "01001000", --  153 - 0x99  :   72 - 0x48
    "01001001", --  154 - 0x9a  :   73 - 0x49
    "00100100", --  155 - 0x9b  :   36 - 0x24
    "00100100", --  156 - 0x9c  :   36 - 0x24
    "00100100", --  157 - 0x9d  :   36 - 0x24
    "00100100", --  158 - 0x9e  :   36 - 0x24
    "00100100", --  159 - 0x9f  :   36 - 0x24
    "00100100", --  160 - 0xa0  :   36 - 0x24
    "00100100", --  161 - 0xa1  :   36 - 0x24
    "00100100", --  162 - 0xa2  :   36 - 0x24
    "00100100", --  163 - 0xa3  :   36 - 0x24
    "00100100", --  164 - 0xa4  :   36 - 0x24
    "01000110", --  165 - 0xa5  :   70 - 0x46
    "11010000", --  166 - 0xa6  :  208 - 0xd0
    "11010001", --  167 - 0xa7  :  209 - 0xd1
    "11011000", --  168 - 0xa8  :  216 - 0xd8
    "11011000", --  169 - 0xa9  :  216 - 0xd8
    "11011110", --  170 - 0xaa  :  222 - 0xde
    "11010001", --  171 - 0xab  :  209 - 0xd1
    "11010000", --  172 - 0xac  :  208 - 0xd0
    "11011010", --  173 - 0xad  :  218 - 0xda
    "11011110", --  174 - 0xae  :  222 - 0xde
    "11010001", --  175 - 0xaf  :  209 - 0xd1
    "00100110", --  176 - 0xb0  :   38 - 0x26
    "00100110", --  177 - 0xb1  :   38 - 0x26
    "00100110", --  178 - 0xb2  :   38 - 0x26
    "00100110", --  179 - 0xb3  :   38 - 0x26
    "00100110", --  180 - 0xb4  :   38 - 0x26
    "00100110", --  181 - 0xb5  :   38 - 0x26
    "00100110", --  182 - 0xb6  :   38 - 0x26
    "00100110", --  183 - 0xb7  :   38 - 0x26
    "00100110", --  184 - 0xb8  :   38 - 0x26
    "00100110", --  185 - 0xb9  :   38 - 0x26
    "01001010", --  186 - 0xba  :   74 - 0x4a
    "00100100", --  187 - 0xbb  :   36 - 0x24
    "00100100", --  188 - 0xbc  :   36 - 0x24
    "00100100", --  189 - 0xbd  :   36 - 0x24
    "00100100", --  190 - 0xbe  :   36 - 0x24
    "00100100", --  191 - 0xbf  :   36 - 0x24
    "00100100", --  192 - 0xc0  :   36 - 0x24
    "00100100", --  193 - 0xc1  :   36 - 0x24
    "00100100", --  194 - 0xc2  :   36 - 0x24
    "00100100", --  195 - 0xc3  :   36 - 0x24
    "00100100", --  196 - 0xc4  :   36 - 0x24
    "01000110", --  197 - 0xc5  :   70 - 0x46
    "11010010", --  198 - 0xc6  :  210 - 0xd2
    "11010011", --  199 - 0xc7  :  211 - 0xd3
    "11011011", --  200 - 0xc8  :  219 - 0xdb
    "11011011", --  201 - 0xc9  :  219 - 0xdb
    "11011011", --  202 - 0xca  :  219 - 0xdb
    "11011001", --  203 - 0xcb  :  217 - 0xd9
    "11011011", --  204 - 0xcc  :  219 - 0xdb
    "11011100", --  205 - 0xcd  :  220 - 0xdc
    "11011011", --  206 - 0xce  :  219 - 0xdb
    "11011111", --  207 - 0xcf  :  223 - 0xdf
    "00100110", --  208 - 0xd0  :   38 - 0x26
    "00100110", --  209 - 0xd1  :   38 - 0x26
    "00100110", --  210 - 0xd2  :   38 - 0x26
    "00100110", --  211 - 0xd3  :   38 - 0x26
    "00100110", --  212 - 0xd4  :   38 - 0x26
    "00100110", --  213 - 0xd5  :   38 - 0x26
    "00100110", --  214 - 0xd6  :   38 - 0x26
    "00100110", --  215 - 0xd7  :   38 - 0x26
    "00100110", --  216 - 0xd8  :   38 - 0x26
    "00100110", --  217 - 0xd9  :   38 - 0x26
    "01001010", --  218 - 0xda  :   74 - 0x4a
    "00100100", --  219 - 0xdb  :   36 - 0x24
    "00100100", --  220 - 0xdc  :   36 - 0x24
    "00100100", --  221 - 0xdd  :   36 - 0x24
    "00100100", --  222 - 0xde  :   36 - 0x24
    "00100100", --  223 - 0xdf  :   36 - 0x24
    "00100100", --  224 - 0xe0  :   36 - 0x24
    "00100100", --  225 - 0xe1  :   36 - 0x24
    "00100100", --  226 - 0xe2  :   36 - 0x24
    "00100100", --  227 - 0xe3  :   36 - 0x24
    "00100100", --  228 - 0xe4  :   36 - 0x24
    "01000110", --  229 - 0xe5  :   70 - 0x46
    "11010100", --  230 - 0xe6  :  212 - 0xd4
    "11010101", --  231 - 0xe7  :  213 - 0xd5
    "11010100", --  232 - 0xe8  :  212 - 0xd4
    "11011001", --  233 - 0xe9  :  217 - 0xd9
    "11011011", --  234 - 0xea  :  219 - 0xdb
    "11100010", --  235 - 0xeb  :  226 - 0xe2
    "11010100", --  236 - 0xec  :  212 - 0xd4
    "11011010", --  237 - 0xed  :  218 - 0xda
    "11011011", --  238 - 0xee  :  219 - 0xdb
    "11100000", --  239 - 0xef  :  224 - 0xe0
    "00100110", --  240 - 0xf0  :   38 - 0x26
    "00100110", --  241 - 0xf1  :   38 - 0x26
    "00100110", --  242 - 0xf2  :   38 - 0x26
    "00100110", --  243 - 0xf3  :   38 - 0x26
    "00100110", --  244 - 0xf4  :   38 - 0x26
    "00100110", --  245 - 0xf5  :   38 - 0x26
    "00100110", --  246 - 0xf6  :   38 - 0x26
    "00100110", --  247 - 0xf7  :   38 - 0x26
    "00100110", --  248 - 0xf8  :   38 - 0x26
    "00100110", --  249 - 0xf9  :   38 - 0x26
    "01001010", --  250 - 0xfa  :   74 - 0x4a
    "00100100", --  251 - 0xfb  :   36 - 0x24
    "00100100", --  252 - 0xfc  :   36 - 0x24
    "00100100", --  253 - 0xfd  :   36 - 0x24
    "00100100", --  254 - 0xfe  :   36 - 0x24
    "00100100", --  255 - 0xff  :   36 - 0x24
    "00100100", --  256 - 0x100  :   36 - 0x24
    "00100100", --  257 - 0x101  :   36 - 0x24
    "00100100", --  258 - 0x102  :   36 - 0x24
    "00100100", --  259 - 0x103  :   36 - 0x24
    "00100100", --  260 - 0x104  :   36 - 0x24
    "01000110", --  261 - 0x105  :   70 - 0x46
    "11010110", --  262 - 0x106  :  214 - 0xd6
    "11010111", --  263 - 0x107  :  215 - 0xd7
    "11010110", --  264 - 0x108  :  214 - 0xd6
    "11010111", --  265 - 0x109  :  215 - 0xd7
    "11100001", --  266 - 0x10a  :  225 - 0xe1
    "00100110", --  267 - 0x10b  :   38 - 0x26
    "11010110", --  268 - 0x10c  :  214 - 0xd6
    "11011101", --  269 - 0x10d  :  221 - 0xdd
    "11100001", --  270 - 0x10e  :  225 - 0xe1
    "11100001", --  271 - 0x10f  :  225 - 0xe1
    "00100110", --  272 - 0x110  :   38 - 0x26
    "00100110", --  273 - 0x111  :   38 - 0x26
    "00100110", --  274 - 0x112  :   38 - 0x26
    "00100110", --  275 - 0x113  :   38 - 0x26
    "00100110", --  276 - 0x114  :   38 - 0x26
    "00100110", --  277 - 0x115  :   38 - 0x26
    "00100110", --  278 - 0x116  :   38 - 0x26
    "00100110", --  279 - 0x117  :   38 - 0x26
    "00100110", --  280 - 0x118  :   38 - 0x26
    "00100110", --  281 - 0x119  :   38 - 0x26
    "01001010", --  282 - 0x11a  :   74 - 0x4a
    "00100100", --  283 - 0x11b  :   36 - 0x24
    "00100100", --  284 - 0x11c  :   36 - 0x24
    "00100100", --  285 - 0x11d  :   36 - 0x24
    "00100100", --  286 - 0x11e  :   36 - 0x24
    "00100100", --  287 - 0x11f  :   36 - 0x24
    "00100100", --  288 - 0x120  :   36 - 0x24
    "00100100", --  289 - 0x121  :   36 - 0x24
    "00100100", --  290 - 0x122  :   36 - 0x24
    "00100100", --  291 - 0x123  :   36 - 0x24
    "00100100", --  292 - 0x124  :   36 - 0x24
    "01000110", --  293 - 0x125  :   70 - 0x46
    "11010000", --  294 - 0x126  :  208 - 0xd0
    "11101000", --  295 - 0x127  :  232 - 0xe8
    "11010001", --  296 - 0x128  :  209 - 0xd1
    "11010000", --  297 - 0x129  :  208 - 0xd0
    "11010001", --  298 - 0x12a  :  209 - 0xd1
    "11011110", --  299 - 0x12b  :  222 - 0xde
    "11010001", --  300 - 0x12c  :  209 - 0xd1
    "11011000", --  301 - 0x12d  :  216 - 0xd8
    "11010000", --  302 - 0x12e  :  208 - 0xd0
    "11010001", --  303 - 0x12f  :  209 - 0xd1
    "00100110", --  304 - 0x130  :   38 - 0x26
    "11011110", --  305 - 0x131  :  222 - 0xde
    "11010001", --  306 - 0x132  :  209 - 0xd1
    "11011110", --  307 - 0x133  :  222 - 0xde
    "11010001", --  308 - 0x134  :  209 - 0xd1
    "11010000", --  309 - 0x135  :  208 - 0xd0
    "11010001", --  310 - 0x136  :  209 - 0xd1
    "11010000", --  311 - 0x137  :  208 - 0xd0
    "11010001", --  312 - 0x138  :  209 - 0xd1
    "00100110", --  313 - 0x139  :   38 - 0x26
    "01001010", --  314 - 0x13a  :   74 - 0x4a
    "00100100", --  315 - 0x13b  :   36 - 0x24
    "00100100", --  316 - 0x13c  :   36 - 0x24
    "00100100", --  317 - 0x13d  :   36 - 0x24
    "00100100", --  318 - 0x13e  :   36 - 0x24
    "00100100", --  319 - 0x13f  :   36 - 0x24
    "00100100", --  320 - 0x140  :   36 - 0x24
    "00100100", --  321 - 0x141  :   36 - 0x24
    "00100100", --  322 - 0x142  :   36 - 0x24
    "00100100", --  323 - 0x143  :   36 - 0x24
    "00100100", --  324 - 0x144  :   36 - 0x24
    "01000110", --  325 - 0x145  :   70 - 0x46
    "11011011", --  326 - 0x146  :  219 - 0xdb
    "01000010", --  327 - 0x147  :   66 - 0x42
    "01000010", --  328 - 0x148  :   66 - 0x42
    "11011011", --  329 - 0x149  :  219 - 0xdb
    "01000010", --  330 - 0x14a  :   66 - 0x42
    "11011011", --  331 - 0x14b  :  219 - 0xdb
    "01000010", --  332 - 0x14c  :   66 - 0x42
    "11011011", --  333 - 0x14d  :  219 - 0xdb
    "11011011", --  334 - 0x14e  :  219 - 0xdb
    "01000010", --  335 - 0x14f  :   66 - 0x42
    "00100110", --  336 - 0x150  :   38 - 0x26
    "11011011", --  337 - 0x151  :  219 - 0xdb
    "01000010", --  338 - 0x152  :   66 - 0x42
    "11011011", --  339 - 0x153  :  219 - 0xdb
    "01000010", --  340 - 0x154  :   66 - 0x42
    "11011011", --  341 - 0x155  :  219 - 0xdb
    "01000010", --  342 - 0x156  :   66 - 0x42
    "11011011", --  343 - 0x157  :  219 - 0xdb
    "01000010", --  344 - 0x158  :   66 - 0x42
    "00100110", --  345 - 0x159  :   38 - 0x26
    "01001010", --  346 - 0x15a  :   74 - 0x4a
    "00100100", --  347 - 0x15b  :   36 - 0x24
    "00100100", --  348 - 0x15c  :   36 - 0x24
    "00100100", --  349 - 0x15d  :   36 - 0x24
    "00100100", --  350 - 0x15e  :   36 - 0x24
    "00100100", --  351 - 0x15f  :   36 - 0x24
    "00100100", --  352 - 0x160  :   36 - 0x24
    "00100100", --  353 - 0x161  :   36 - 0x24
    "00100100", --  354 - 0x162  :   36 - 0x24
    "00100100", --  355 - 0x163  :   36 - 0x24
    "00100100", --  356 - 0x164  :   36 - 0x24
    "01000110", --  357 - 0x165  :   70 - 0x46
    "11011011", --  358 - 0x166  :  219 - 0xdb
    "11011011", --  359 - 0x167  :  219 - 0xdb
    "11011011", --  360 - 0x168  :  219 - 0xdb
    "11011011", --  361 - 0x169  :  219 - 0xdb
    "11011011", --  362 - 0x16a  :  219 - 0xdb
    "11011011", --  363 - 0x16b  :  219 - 0xdb
    "11011111", --  364 - 0x16c  :  223 - 0xdf
    "11011011", --  365 - 0x16d  :  219 - 0xdb
    "11011011", --  366 - 0x16e  :  219 - 0xdb
    "11011011", --  367 - 0x16f  :  219 - 0xdb
    "00100110", --  368 - 0x170  :   38 - 0x26
    "11011011", --  369 - 0x171  :  219 - 0xdb
    "11011111", --  370 - 0x172  :  223 - 0xdf
    "11011011", --  371 - 0x173  :  219 - 0xdb
    "11011111", --  372 - 0x174  :  223 - 0xdf
    "11011011", --  373 - 0x175  :  219 - 0xdb
    "11011011", --  374 - 0x176  :  219 - 0xdb
    "11100100", --  375 - 0x177  :  228 - 0xe4
    "11100101", --  376 - 0x178  :  229 - 0xe5
    "00100110", --  377 - 0x179  :   38 - 0x26
    "01001010", --  378 - 0x17a  :   74 - 0x4a
    "00100100", --  379 - 0x17b  :   36 - 0x24
    "00100100", --  380 - 0x17c  :   36 - 0x24
    "00100100", --  381 - 0x17d  :   36 - 0x24
    "00100100", --  382 - 0x17e  :   36 - 0x24
    "00100100", --  383 - 0x17f  :   36 - 0x24
    "00100100", --  384 - 0x180  :   36 - 0x24
    "00100100", --  385 - 0x181  :   36 - 0x24
    "00100100", --  386 - 0x182  :   36 - 0x24
    "00100100", --  387 - 0x183  :   36 - 0x24
    "00100100", --  388 - 0x184  :   36 - 0x24
    "01000110", --  389 - 0x185  :   70 - 0x46
    "11011011", --  390 - 0x186  :  219 - 0xdb
    "11011011", --  391 - 0x187  :  219 - 0xdb
    "11011011", --  392 - 0x188  :  219 - 0xdb
    "11011110", --  393 - 0x189  :  222 - 0xde
    "01000011", --  394 - 0x18a  :   67 - 0x43
    "11011011", --  395 - 0x18b  :  219 - 0xdb
    "11100000", --  396 - 0x18c  :  224 - 0xe0
    "11011011", --  397 - 0x18d  :  219 - 0xdb
    "11011011", --  398 - 0x18e  :  219 - 0xdb
    "11011011", --  399 - 0x18f  :  219 - 0xdb
    "00100110", --  400 - 0x190  :   38 - 0x26
    "11011011", --  401 - 0x191  :  219 - 0xdb
    "11100011", --  402 - 0x192  :  227 - 0xe3
    "11011011", --  403 - 0x193  :  219 - 0xdb
    "11100000", --  404 - 0x194  :  224 - 0xe0
    "11011011", --  405 - 0x195  :  219 - 0xdb
    "11011011", --  406 - 0x196  :  219 - 0xdb
    "11100110", --  407 - 0x197  :  230 - 0xe6
    "11100011", --  408 - 0x198  :  227 - 0xe3
    "00100110", --  409 - 0x199  :   38 - 0x26
    "01001010", --  410 - 0x19a  :   74 - 0x4a
    "00100100", --  411 - 0x19b  :   36 - 0x24
    "00100100", --  412 - 0x19c  :   36 - 0x24
    "00100100", --  413 - 0x19d  :   36 - 0x24
    "00100100", --  414 - 0x19e  :   36 - 0x24
    "00100100", --  415 - 0x19f  :   36 - 0x24
    "00100100", --  416 - 0x1a0  :   36 - 0x24
    "00100100", --  417 - 0x1a1  :   36 - 0x24
    "00100100", --  418 - 0x1a2  :   36 - 0x24
    "00100100", --  419 - 0x1a3  :   36 - 0x24
    "00100100", --  420 - 0x1a4  :   36 - 0x24
    "01000110", --  421 - 0x1a5  :   70 - 0x46
    "11011011", --  422 - 0x1a6  :  219 - 0xdb
    "11011011", --  423 - 0x1a7  :  219 - 0xdb
    "11011011", --  424 - 0x1a8  :  219 - 0xdb
    "11011011", --  425 - 0x1a9  :  219 - 0xdb
    "01000010", --  426 - 0x1aa  :   66 - 0x42
    "11011011", --  427 - 0x1ab  :  219 - 0xdb
    "11011011", --  428 - 0x1ac  :  219 - 0xdb
    "11011011", --  429 - 0x1ad  :  219 - 0xdb
    "11010100", --  430 - 0x1ae  :  212 - 0xd4
    "11011001", --  431 - 0x1af  :  217 - 0xd9
    "00100110", --  432 - 0x1b0  :   38 - 0x26
    "11011011", --  433 - 0x1b1  :  219 - 0xdb
    "11011001", --  434 - 0x1b2  :  217 - 0xd9
    "11011011", --  435 - 0x1b3  :  219 - 0xdb
    "11011011", --  436 - 0x1b4  :  219 - 0xdb
    "11010100", --  437 - 0x1b5  :  212 - 0xd4
    "11011001", --  438 - 0x1b6  :  217 - 0xd9
    "11010100", --  439 - 0x1b7  :  212 - 0xd4
    "11011001", --  440 - 0x1b8  :  217 - 0xd9
    "11100111", --  441 - 0x1b9  :  231 - 0xe7
    "01001010", --  442 - 0x1ba  :   74 - 0x4a
    "00100100", --  443 - 0x1bb  :   36 - 0x24
    "00100100", --  444 - 0x1bc  :   36 - 0x24
    "00100100", --  445 - 0x1bd  :   36 - 0x24
    "00100100", --  446 - 0x1be  :   36 - 0x24
    "00100100", --  447 - 0x1bf  :   36 - 0x24
    "00100100", --  448 - 0x1c0  :   36 - 0x24
    "00100100", --  449 - 0x1c1  :   36 - 0x24
    "00100100", --  450 - 0x1c2  :   36 - 0x24
    "00100100", --  451 - 0x1c3  :   36 - 0x24
    "00100100", --  452 - 0x1c4  :   36 - 0x24
    "01011111", --  453 - 0x1c5  :   95 - 0x5f
    "10010101", --  454 - 0x1c6  :  149 - 0x95
    "10010101", --  455 - 0x1c7  :  149 - 0x95
    "10010101", --  456 - 0x1c8  :  149 - 0x95
    "10010101", --  457 - 0x1c9  :  149 - 0x95
    "10010101", --  458 - 0x1ca  :  149 - 0x95
    "10010101", --  459 - 0x1cb  :  149 - 0x95
    "10010101", --  460 - 0x1cc  :  149 - 0x95
    "10010101", --  461 - 0x1cd  :  149 - 0x95
    "10010111", --  462 - 0x1ce  :  151 - 0x97
    "10011000", --  463 - 0x1cf  :  152 - 0x98
    "01111000", --  464 - 0x1d0  :  120 - 0x78
    "10010101", --  465 - 0x1d1  :  149 - 0x95
    "10010110", --  466 - 0x1d2  :  150 - 0x96
    "10010101", --  467 - 0x1d3  :  149 - 0x95
    "10010101", --  468 - 0x1d4  :  149 - 0x95
    "10010111", --  469 - 0x1d5  :  151 - 0x97
    "10011000", --  470 - 0x1d6  :  152 - 0x98
    "10010111", --  471 - 0x1d7  :  151 - 0x97
    "10011000", --  472 - 0x1d8  :  152 - 0x98
    "10010101", --  473 - 0x1d9  :  149 - 0x95
    "01111010", --  474 - 0x1da  :  122 - 0x7a
    "00100100", --  475 - 0x1db  :   36 - 0x24
    "00100100", --  476 - 0x1dc  :   36 - 0x24
    "00100100", --  477 - 0x1dd  :   36 - 0x24
    "00100100", --  478 - 0x1de  :   36 - 0x24
    "00100100", --  479 - 0x1df  :   36 - 0x24
    "00100100", --  480 - 0x1e0  :   36 - 0x24
    "00100100", --  481 - 0x1e1  :   36 - 0x24
    "00100100", --  482 - 0x1e2  :   36 - 0x24
    "00100100", --  483 - 0x1e3  :   36 - 0x24
    "00100100", --  484 - 0x1e4  :   36 - 0x24
    "00100100", --  485 - 0x1e5  :   36 - 0x24
    "00100100", --  486 - 0x1e6  :   36 - 0x24
    "00100100", --  487 - 0x1e7  :   36 - 0x24
    "00100100", --  488 - 0x1e8  :   36 - 0x24
    "00100100", --  489 - 0x1e9  :   36 - 0x24
    "00100100", --  490 - 0x1ea  :   36 - 0x24
    "00100100", --  491 - 0x1eb  :   36 - 0x24
    "00100100", --  492 - 0x1ec  :   36 - 0x24
    "11001111", --  493 - 0x1ed  :  207 - 0xcf
    "00000001", --  494 - 0x1ee  :    1 - 0x1
    "00001001", --  495 - 0x1ef  :    9 - 0x9
    "00001000", --  496 - 0x1f0  :    8 - 0x8
    "00000101", --  497 - 0x1f1  :    5 - 0x5
    "00100100", --  498 - 0x1f2  :   36 - 0x24
    "00010111", --  499 - 0x1f3  :   23 - 0x17
    "00010010", --  500 - 0x1f4  :   18 - 0x12
    "00010111", --  501 - 0x1f5  :   23 - 0x17
    "00011101", --  502 - 0x1f6  :   29 - 0x1d
    "00001110", --  503 - 0x1f7  :   14 - 0xe
    "00010111", --  504 - 0x1f8  :   23 - 0x17
    "00001101", --  505 - 0x1f9  :   13 - 0xd
    "00011000", --  506 - 0x1fa  :   24 - 0x18
    "00100100", --  507 - 0x1fb  :   36 - 0x24
    "00100100", --  508 - 0x1fc  :   36 - 0x24
    "00100100", --  509 - 0x1fd  :   36 - 0x24
    "00100100", --  510 - 0x1fe  :   36 - 0x24
    "00100100", --  511 - 0x1ff  :   36 - 0x24
    "00100100", --  512 - 0x200  :   36 - 0x24
    "00100100", --  513 - 0x201  :   36 - 0x24
    "00100100", --  514 - 0x202  :   36 - 0x24
    "00100100", --  515 - 0x203  :   36 - 0x24
    "00100100", --  516 - 0x204  :   36 - 0x24
    "00100100", --  517 - 0x205  :   36 - 0x24
    "00100100", --  518 - 0x206  :   36 - 0x24
    "00100100", --  519 - 0x207  :   36 - 0x24
    "00100100", --  520 - 0x208  :   36 - 0x24
    "00100100", --  521 - 0x209  :   36 - 0x24
    "00100100", --  522 - 0x20a  :   36 - 0x24
    "00100100", --  523 - 0x20b  :   36 - 0x24
    "00100100", --  524 - 0x20c  :   36 - 0x24
    "00100100", --  525 - 0x20d  :   36 - 0x24
    "00100100", --  526 - 0x20e  :   36 - 0x24
    "00100100", --  527 - 0x20f  :   36 - 0x24
    "00100100", --  528 - 0x210  :   36 - 0x24
    "00100100", --  529 - 0x211  :   36 - 0x24
    "00100100", --  530 - 0x212  :   36 - 0x24
    "00100100", --  531 - 0x213  :   36 - 0x24
    "00100100", --  532 - 0x214  :   36 - 0x24
    "00100100", --  533 - 0x215  :   36 - 0x24
    "00100100", --  534 - 0x216  :   36 - 0x24
    "00100100", --  535 - 0x217  :   36 - 0x24
    "00100100", --  536 - 0x218  :   36 - 0x24
    "00100100", --  537 - 0x219  :   36 - 0x24
    "00100100", --  538 - 0x21a  :   36 - 0x24
    "00100100", --  539 - 0x21b  :   36 - 0x24
    "00100100", --  540 - 0x21c  :   36 - 0x24
    "00100100", --  541 - 0x21d  :   36 - 0x24
    "00100100", --  542 - 0x21e  :   36 - 0x24
    "00100100", --  543 - 0x21f  :   36 - 0x24
    "00100100", --  544 - 0x220  :   36 - 0x24
    "00100100", --  545 - 0x221  :   36 - 0x24
    "00100100", --  546 - 0x222  :   36 - 0x24
    "00100100", --  547 - 0x223  :   36 - 0x24
    "00100100", --  548 - 0x224  :   36 - 0x24
    "00100100", --  549 - 0x225  :   36 - 0x24
    "00100100", --  550 - 0x226  :   36 - 0x24
    "00100100", --  551 - 0x227  :   36 - 0x24
    "00100100", --  552 - 0x228  :   36 - 0x24
    "00100100", --  553 - 0x229  :   36 - 0x24
    "00100100", --  554 - 0x22a  :   36 - 0x24
    "00100100", --  555 - 0x22b  :   36 - 0x24
    "00100100", --  556 - 0x22c  :   36 - 0x24
    "00100100", --  557 - 0x22d  :   36 - 0x24
    "00100100", --  558 - 0x22e  :   36 - 0x24
    "00100100", --  559 - 0x22f  :   36 - 0x24
    "00100100", --  560 - 0x230  :   36 - 0x24
    "00100100", --  561 - 0x231  :   36 - 0x24
    "00100100", --  562 - 0x232  :   36 - 0x24
    "00100100", --  563 - 0x233  :   36 - 0x24
    "00100100", --  564 - 0x234  :   36 - 0x24
    "00100100", --  565 - 0x235  :   36 - 0x24
    "00100100", --  566 - 0x236  :   36 - 0x24
    "00100100", --  567 - 0x237  :   36 - 0x24
    "00100100", --  568 - 0x238  :   36 - 0x24
    "00100100", --  569 - 0x239  :   36 - 0x24
    "00100100", --  570 - 0x23a  :   36 - 0x24
    "00100100", --  571 - 0x23b  :   36 - 0x24
    "00100100", --  572 - 0x23c  :   36 - 0x24
    "00100100", --  573 - 0x23d  :   36 - 0x24
    "00100100", --  574 - 0x23e  :   36 - 0x24
    "00100100", --  575 - 0x23f  :   36 - 0x24
    "00100100", --  576 - 0x240  :   36 - 0x24
    "00100100", --  577 - 0x241  :   36 - 0x24
    "00100100", --  578 - 0x242  :   36 - 0x24
    "00100100", --  579 - 0x243  :   36 - 0x24
    "00100100", --  580 - 0x244  :   36 - 0x24
    "00100100", --  581 - 0x245  :   36 - 0x24
    "00100100", --  582 - 0x246  :   36 - 0x24
    "00100100", --  583 - 0x247  :   36 - 0x24
    "00100100", --  584 - 0x248  :   36 - 0x24
    "11001110", --  585 - 0x249  :  206 - 0xce
    "00100100", --  586 - 0x24a  :   36 - 0x24
    "00000001", --  587 - 0x24b  :    1 - 0x1
    "00100100", --  588 - 0x24c  :   36 - 0x24
    "00011001", --  589 - 0x24d  :   25 - 0x19
    "00010101", --  590 - 0x24e  :   21 - 0x15
    "00001010", --  591 - 0x24f  :   10 - 0xa
    "00100010", --  592 - 0x250  :   34 - 0x22
    "00001110", --  593 - 0x251  :   14 - 0xe
    "00011011", --  594 - 0x252  :   27 - 0x1b
    "00100100", --  595 - 0x253  :   36 - 0x24
    "00010000", --  596 - 0x254  :   16 - 0x10
    "00001010", --  597 - 0x255  :   10 - 0xa
    "00010110", --  598 - 0x256  :   22 - 0x16
    "00001110", --  599 - 0x257  :   14 - 0xe
    "00100100", --  600 - 0x258  :   36 - 0x24
    "00100100", --  601 - 0x259  :   36 - 0x24
    "00100100", --  602 - 0x25a  :   36 - 0x24
    "00100100", --  603 - 0x25b  :   36 - 0x24
    "00100100", --  604 - 0x25c  :   36 - 0x24
    "00100100", --  605 - 0x25d  :   36 - 0x24
    "00100100", --  606 - 0x25e  :   36 - 0x24
    "00100100", --  607 - 0x25f  :   36 - 0x24
    "00100100", --  608 - 0x260  :   36 - 0x24
    "00100100", --  609 - 0x261  :   36 - 0x24
    "00100100", --  610 - 0x262  :   36 - 0x24
    "00100100", --  611 - 0x263  :   36 - 0x24
    "00100100", --  612 - 0x264  :   36 - 0x24
    "00100100", --  613 - 0x265  :   36 - 0x24
    "00100100", --  614 - 0x266  :   36 - 0x24
    "00100100", --  615 - 0x267  :   36 - 0x24
    "00100100", --  616 - 0x268  :   36 - 0x24
    "00100100", --  617 - 0x269  :   36 - 0x24
    "00100100", --  618 - 0x26a  :   36 - 0x24
    "00100100", --  619 - 0x26b  :   36 - 0x24
    "00100100", --  620 - 0x26c  :   36 - 0x24
    "00100100", --  621 - 0x26d  :   36 - 0x24
    "00100100", --  622 - 0x26e  :   36 - 0x24
    "00100100", --  623 - 0x26f  :   36 - 0x24
    "00100100", --  624 - 0x270  :   36 - 0x24
    "00100100", --  625 - 0x271  :   36 - 0x24
    "00100100", --  626 - 0x272  :   36 - 0x24
    "00100100", --  627 - 0x273  :   36 - 0x24
    "00100100", --  628 - 0x274  :   36 - 0x24
    "00100100", --  629 - 0x275  :   36 - 0x24
    "00100100", --  630 - 0x276  :   36 - 0x24
    "00100100", --  631 - 0x277  :   36 - 0x24
    "00100100", --  632 - 0x278  :   36 - 0x24
    "00100100", --  633 - 0x279  :   36 - 0x24
    "00100100", --  634 - 0x27a  :   36 - 0x24
    "00100100", --  635 - 0x27b  :   36 - 0x24
    "00100100", --  636 - 0x27c  :   36 - 0x24
    "00100100", --  637 - 0x27d  :   36 - 0x24
    "00100100", --  638 - 0x27e  :   36 - 0x24
    "00100100", --  639 - 0x27f  :   36 - 0x24
    "00100100", --  640 - 0x280  :   36 - 0x24
    "00100100", --  641 - 0x281  :   36 - 0x24
    "00100100", --  642 - 0x282  :   36 - 0x24
    "00100100", --  643 - 0x283  :   36 - 0x24
    "00100100", --  644 - 0x284  :   36 - 0x24
    "00100100", --  645 - 0x285  :   36 - 0x24
    "00100100", --  646 - 0x286  :   36 - 0x24
    "00100100", --  647 - 0x287  :   36 - 0x24
    "00100100", --  648 - 0x288  :   36 - 0x24
    "00100100", --  649 - 0x289  :   36 - 0x24
    "00100100", --  650 - 0x28a  :   36 - 0x24
    "00000010", --  651 - 0x28b  :    2 - 0x2
    "00100100", --  652 - 0x28c  :   36 - 0x24
    "00011001", --  653 - 0x28d  :   25 - 0x19
    "00010101", --  654 - 0x28e  :   21 - 0x15
    "00001010", --  655 - 0x28f  :   10 - 0xa
    "00100010", --  656 - 0x290  :   34 - 0x22
    "00001110", --  657 - 0x291  :   14 - 0xe
    "00011011", --  658 - 0x292  :   27 - 0x1b
    "00100100", --  659 - 0x293  :   36 - 0x24
    "00010000", --  660 - 0x294  :   16 - 0x10
    "00001010", --  661 - 0x295  :   10 - 0xa
    "00010110", --  662 - 0x296  :   22 - 0x16
    "00001110", --  663 - 0x297  :   14 - 0xe
    "00100100", --  664 - 0x298  :   36 - 0x24
    "00100100", --  665 - 0x299  :   36 - 0x24
    "00100100", --  666 - 0x29a  :   36 - 0x24
    "00100100", --  667 - 0x29b  :   36 - 0x24
    "00100100", --  668 - 0x29c  :   36 - 0x24
    "00100100", --  669 - 0x29d  :   36 - 0x24
    "00100100", --  670 - 0x29e  :   36 - 0x24
    "00100100", --  671 - 0x29f  :   36 - 0x24
    "00100100", --  672 - 0x2a0  :   36 - 0x24
    "00100100", --  673 - 0x2a1  :   36 - 0x24
    "00100100", --  674 - 0x2a2  :   36 - 0x24
    "00100100", --  675 - 0x2a3  :   36 - 0x24
    "00110001", --  676 - 0x2a4  :   49 - 0x31
    "00110010", --  677 - 0x2a5  :   50 - 0x32
    "00100100", --  678 - 0x2a6  :   36 - 0x24
    "00100100", --  679 - 0x2a7  :   36 - 0x24
    "00100100", --  680 - 0x2a8  :   36 - 0x24
    "00100100", --  681 - 0x2a9  :   36 - 0x24
    "00100100", --  682 - 0x2aa  :   36 - 0x24
    "00100100", --  683 - 0x2ab  :   36 - 0x24
    "00100100", --  684 - 0x2ac  :   36 - 0x24
    "00100100", --  685 - 0x2ad  :   36 - 0x24
    "00100100", --  686 - 0x2ae  :   36 - 0x24
    "00100100", --  687 - 0x2af  :   36 - 0x24
    "00100100", --  688 - 0x2b0  :   36 - 0x24
    "00100100", --  689 - 0x2b1  :   36 - 0x24
    "00100100", --  690 - 0x2b2  :   36 - 0x24
    "00100100", --  691 - 0x2b3  :   36 - 0x24
    "00100100", --  692 - 0x2b4  :   36 - 0x24
    "00100100", --  693 - 0x2b5  :   36 - 0x24
    "00100100", --  694 - 0x2b6  :   36 - 0x24
    "00100100", --  695 - 0x2b7  :   36 - 0x24
    "00100100", --  696 - 0x2b8  :   36 - 0x24
    "00100100", --  697 - 0x2b9  :   36 - 0x24
    "00100100", --  698 - 0x2ba  :   36 - 0x24
    "00100100", --  699 - 0x2bb  :   36 - 0x24
    "00100100", --  700 - 0x2bc  :   36 - 0x24
    "00100100", --  701 - 0x2bd  :   36 - 0x24
    "00100100", --  702 - 0x2be  :   36 - 0x24
    "00100100", --  703 - 0x2bf  :   36 - 0x24
    "00100100", --  704 - 0x2c0  :   36 - 0x24
    "00100100", --  705 - 0x2c1  :   36 - 0x24
    "00100100", --  706 - 0x2c2  :   36 - 0x24
    "00110000", --  707 - 0x2c3  :   48 - 0x30
    "00100110", --  708 - 0x2c4  :   38 - 0x26
    "00110100", --  709 - 0x2c5  :   52 - 0x34
    "00110011", --  710 - 0x2c6  :   51 - 0x33
    "00100100", --  711 - 0x2c7  :   36 - 0x24
    "00100100", --  712 - 0x2c8  :   36 - 0x24
    "00100100", --  713 - 0x2c9  :   36 - 0x24
    "00100100", --  714 - 0x2ca  :   36 - 0x24
    "00100100", --  715 - 0x2cb  :   36 - 0x24
    "00100100", --  716 - 0x2cc  :   36 - 0x24
    "00100100", --  717 - 0x2cd  :   36 - 0x24
    "00100100", --  718 - 0x2ce  :   36 - 0x24
    "00100100", --  719 - 0x2cf  :   36 - 0x24
    "00100100", --  720 - 0x2d0  :   36 - 0x24
    "00100100", --  721 - 0x2d1  :   36 - 0x24
    "00100100", --  722 - 0x2d2  :   36 - 0x24
    "00100100", --  723 - 0x2d3  :   36 - 0x24
    "00100100", --  724 - 0x2d4  :   36 - 0x24
    "00100100", --  725 - 0x2d5  :   36 - 0x24
    "00100100", --  726 - 0x2d6  :   36 - 0x24
    "00100100", --  727 - 0x2d7  :   36 - 0x24
    "00100100", --  728 - 0x2d8  :   36 - 0x24
    "00100100", --  729 - 0x2d9  :   36 - 0x24
    "00100100", --  730 - 0x2da  :   36 - 0x24
    "00100100", --  731 - 0x2db  :   36 - 0x24
    "00100100", --  732 - 0x2dc  :   36 - 0x24
    "00100100", --  733 - 0x2dd  :   36 - 0x24
    "00100100", --  734 - 0x2de  :   36 - 0x24
    "00100100", --  735 - 0x2df  :   36 - 0x24
    "00100100", --  736 - 0x2e0  :   36 - 0x24
    "00100100", --  737 - 0x2e1  :   36 - 0x24
    "00110000", --  738 - 0x2e2  :   48 - 0x30
    "00100110", --  739 - 0x2e3  :   38 - 0x26
    "00100110", --  740 - 0x2e4  :   38 - 0x26
    "00100110", --  741 - 0x2e5  :   38 - 0x26
    "00100110", --  742 - 0x2e6  :   38 - 0x26
    "00110011", --  743 - 0x2e7  :   51 - 0x33
    "00100100", --  744 - 0x2e8  :   36 - 0x24
    "00100100", --  745 - 0x2e9  :   36 - 0x24
    "00100100", --  746 - 0x2ea  :   36 - 0x24
    "00100100", --  747 - 0x2eb  :   36 - 0x24
    "00011101", --  748 - 0x2ec  :   29 - 0x1d
    "00011000", --  749 - 0x2ed  :   24 - 0x18
    "00011001", --  750 - 0x2ee  :   25 - 0x19
    "00101000", --  751 - 0x2ef  :   40 - 0x28
    "00100100", --  752 - 0x2f0  :   36 - 0x24
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00000000", --  754 - 0x2f2  :    0 - 0x0
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "00000000", --  756 - 0x2f4  :    0 - 0x0
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00100100", --  759 - 0x2f7  :   36 - 0x24
    "00100100", --  760 - 0x2f8  :   36 - 0x24
    "00100100", --  761 - 0x2f9  :   36 - 0x24
    "00100100", --  762 - 0x2fa  :   36 - 0x24
    "00100100", --  763 - 0x2fb  :   36 - 0x24
    "00100100", --  764 - 0x2fc  :   36 - 0x24
    "00100100", --  765 - 0x2fd  :   36 - 0x24
    "00100100", --  766 - 0x2fe  :   36 - 0x24
    "00100100", --  767 - 0x2ff  :   36 - 0x24
    "00100100", --  768 - 0x300  :   36 - 0x24
    "00110000", --  769 - 0x301  :   48 - 0x30
    "00100110", --  770 - 0x302  :   38 - 0x26
    "00110100", --  771 - 0x303  :   52 - 0x34
    "00100110", --  772 - 0x304  :   38 - 0x26
    "00100110", --  773 - 0x305  :   38 - 0x26
    "00110100", --  774 - 0x306  :   52 - 0x34
    "00100110", --  775 - 0x307  :   38 - 0x26
    "00110011", --  776 - 0x308  :   51 - 0x33
    "00100100", --  777 - 0x309  :   36 - 0x24
    "00100100", --  778 - 0x30a  :   36 - 0x24
    "00100100", --  779 - 0x30b  :   36 - 0x24
    "00100100", --  780 - 0x30c  :   36 - 0x24
    "00100100", --  781 - 0x30d  :   36 - 0x24
    "00100100", --  782 - 0x30e  :   36 - 0x24
    "00100100", --  783 - 0x30f  :   36 - 0x24
    "00100100", --  784 - 0x310  :   36 - 0x24
    "00100100", --  785 - 0x311  :   36 - 0x24
    "00100100", --  786 - 0x312  :   36 - 0x24
    "00100100", --  787 - 0x313  :   36 - 0x24
    "00100100", --  788 - 0x314  :   36 - 0x24
    "00100100", --  789 - 0x315  :   36 - 0x24
    "00100100", --  790 - 0x316  :   36 - 0x24
    "00100100", --  791 - 0x317  :   36 - 0x24
    "00110110", --  792 - 0x318  :   54 - 0x36
    "00110111", --  793 - 0x319  :   55 - 0x37
    "00110110", --  794 - 0x31a  :   54 - 0x36
    "00110111", --  795 - 0x31b  :   55 - 0x37
    "00110110", --  796 - 0x31c  :   54 - 0x36
    "00110111", --  797 - 0x31d  :   55 - 0x37
    "00100100", --  798 - 0x31e  :   36 - 0x24
    "00100100", --  799 - 0x31f  :   36 - 0x24
    "00110000", --  800 - 0x320  :   48 - 0x30
    "00100110", --  801 - 0x321  :   38 - 0x26
    "00100110", --  802 - 0x322  :   38 - 0x26
    "00100110", --  803 - 0x323  :   38 - 0x26
    "00100110", --  804 - 0x324  :   38 - 0x26
    "00100110", --  805 - 0x325  :   38 - 0x26
    "00100110", --  806 - 0x326  :   38 - 0x26
    "00100110", --  807 - 0x327  :   38 - 0x26
    "00100110", --  808 - 0x328  :   38 - 0x26
    "00110011", --  809 - 0x329  :   51 - 0x33
    "00100100", --  810 - 0x32a  :   36 - 0x24
    "00100100", --  811 - 0x32b  :   36 - 0x24
    "00100100", --  812 - 0x32c  :   36 - 0x24
    "00100100", --  813 - 0x32d  :   36 - 0x24
    "00100100", --  814 - 0x32e  :   36 - 0x24
    "00100100", --  815 - 0x32f  :   36 - 0x24
    "00100100", --  816 - 0x330  :   36 - 0x24
    "00100100", --  817 - 0x331  :   36 - 0x24
    "00100100", --  818 - 0x332  :   36 - 0x24
    "00100100", --  819 - 0x333  :   36 - 0x24
    "00100100", --  820 - 0x334  :   36 - 0x24
    "00100100", --  821 - 0x335  :   36 - 0x24
    "00100100", --  822 - 0x336  :   36 - 0x24
    "00110101", --  823 - 0x337  :   53 - 0x35
    "00100101", --  824 - 0x338  :   37 - 0x25
    "00100101", --  825 - 0x339  :   37 - 0x25
    "00100101", --  826 - 0x33a  :   37 - 0x25
    "00100101", --  827 - 0x33b  :   37 - 0x25
    "00100101", --  828 - 0x33c  :   37 - 0x25
    "00100101", --  829 - 0x33d  :   37 - 0x25
    "00111000", --  830 - 0x33e  :   56 - 0x38
    "00100100", --  831 - 0x33f  :   36 - 0x24
    "10110100", --  832 - 0x340  :  180 - 0xb4
    "10110101", --  833 - 0x341  :  181 - 0xb5
    "10110100", --  834 - 0x342  :  180 - 0xb4
    "10110101", --  835 - 0x343  :  181 - 0xb5
    "10110100", --  836 - 0x344  :  180 - 0xb4
    "10110101", --  837 - 0x345  :  181 - 0xb5
    "10110100", --  838 - 0x346  :  180 - 0xb4
    "10110101", --  839 - 0x347  :  181 - 0xb5
    "10110100", --  840 - 0x348  :  180 - 0xb4
    "10110101", --  841 - 0x349  :  181 - 0xb5
    "10110100", --  842 - 0x34a  :  180 - 0xb4
    "10110101", --  843 - 0x34b  :  181 - 0xb5
    "10110100", --  844 - 0x34c  :  180 - 0xb4
    "10110101", --  845 - 0x34d  :  181 - 0xb5
    "10110100", --  846 - 0x34e  :  180 - 0xb4
    "10110101", --  847 - 0x34f  :  181 - 0xb5
    "10110100", --  848 - 0x350  :  180 - 0xb4
    "10110101", --  849 - 0x351  :  181 - 0xb5
    "10110100", --  850 - 0x352  :  180 - 0xb4
    "10110101", --  851 - 0x353  :  181 - 0xb5
    "10110100", --  852 - 0x354  :  180 - 0xb4
    "10110101", --  853 - 0x355  :  181 - 0xb5
    "10110100", --  854 - 0x356  :  180 - 0xb4
    "10110101", --  855 - 0x357  :  181 - 0xb5
    "10110100", --  856 - 0x358  :  180 - 0xb4
    "10110101", --  857 - 0x359  :  181 - 0xb5
    "10110100", --  858 - 0x35a  :  180 - 0xb4
    "10110101", --  859 - 0x35b  :  181 - 0xb5
    "10110100", --  860 - 0x35c  :  180 - 0xb4
    "10110101", --  861 - 0x35d  :  181 - 0xb5
    "10110100", --  862 - 0x35e  :  180 - 0xb4
    "10110101", --  863 - 0x35f  :  181 - 0xb5
    "10110110", --  864 - 0x360  :  182 - 0xb6
    "10110111", --  865 - 0x361  :  183 - 0xb7
    "10110110", --  866 - 0x362  :  182 - 0xb6
    "10110111", --  867 - 0x363  :  183 - 0xb7
    "10110110", --  868 - 0x364  :  182 - 0xb6
    "10110111", --  869 - 0x365  :  183 - 0xb7
    "10110110", --  870 - 0x366  :  182 - 0xb6
    "10110111", --  871 - 0x367  :  183 - 0xb7
    "10110110", --  872 - 0x368  :  182 - 0xb6
    "10110111", --  873 - 0x369  :  183 - 0xb7
    "10110110", --  874 - 0x36a  :  182 - 0xb6
    "10110111", --  875 - 0x36b  :  183 - 0xb7
    "10110110", --  876 - 0x36c  :  182 - 0xb6
    "10110111", --  877 - 0x36d  :  183 - 0xb7
    "10110110", --  878 - 0x36e  :  182 - 0xb6
    "10110111", --  879 - 0x36f  :  183 - 0xb7
    "10110110", --  880 - 0x370  :  182 - 0xb6
    "10110111", --  881 - 0x371  :  183 - 0xb7
    "10110110", --  882 - 0x372  :  182 - 0xb6
    "10110111", --  883 - 0x373  :  183 - 0xb7
    "10110110", --  884 - 0x374  :  182 - 0xb6
    "10110111", --  885 - 0x375  :  183 - 0xb7
    "10110110", --  886 - 0x376  :  182 - 0xb6
    "10110111", --  887 - 0x377  :  183 - 0xb7
    "10110110", --  888 - 0x378  :  182 - 0xb6
    "10110111", --  889 - 0x379  :  183 - 0xb7
    "10110110", --  890 - 0x37a  :  182 - 0xb6
    "10110111", --  891 - 0x37b  :  183 - 0xb7
    "10110110", --  892 - 0x37c  :  182 - 0xb6
    "10110111", --  893 - 0x37d  :  183 - 0xb7
    "10110110", --  894 - 0x37e  :  182 - 0xb6
    "10110111", --  895 - 0x37f  :  183 - 0xb7
    "10110100", --  896 - 0x380  :  180 - 0xb4
    "10110101", --  897 - 0x381  :  181 - 0xb5
    "10110100", --  898 - 0x382  :  180 - 0xb4
    "10110101", --  899 - 0x383  :  181 - 0xb5
    "10110100", --  900 - 0x384  :  180 - 0xb4
    "10110101", --  901 - 0x385  :  181 - 0xb5
    "10110100", --  902 - 0x386  :  180 - 0xb4
    "10110101", --  903 - 0x387  :  181 - 0xb5
    "10110100", --  904 - 0x388  :  180 - 0xb4
    "10110101", --  905 - 0x389  :  181 - 0xb5
    "10110100", --  906 - 0x38a  :  180 - 0xb4
    "10110101", --  907 - 0x38b  :  181 - 0xb5
    "10110100", --  908 - 0x38c  :  180 - 0xb4
    "10110101", --  909 - 0x38d  :  181 - 0xb5
    "10110100", --  910 - 0x38e  :  180 - 0xb4
    "10110101", --  911 - 0x38f  :  181 - 0xb5
    "10110100", --  912 - 0x390  :  180 - 0xb4
    "10110101", --  913 - 0x391  :  181 - 0xb5
    "10110100", --  914 - 0x392  :  180 - 0xb4
    "10110101", --  915 - 0x393  :  181 - 0xb5
    "10110100", --  916 - 0x394  :  180 - 0xb4
    "10110101", --  917 - 0x395  :  181 - 0xb5
    "10110100", --  918 - 0x396  :  180 - 0xb4
    "10110101", --  919 - 0x397  :  181 - 0xb5
    "10110100", --  920 - 0x398  :  180 - 0xb4
    "10110101", --  921 - 0x399  :  181 - 0xb5
    "10110100", --  922 - 0x39a  :  180 - 0xb4
    "10110101", --  923 - 0x39b  :  181 - 0xb5
    "10110100", --  924 - 0x39c  :  180 - 0xb4
    "10110101", --  925 - 0x39d  :  181 - 0xb5
    "10110100", --  926 - 0x39e  :  180 - 0xb4
    "10110101", --  927 - 0x39f  :  181 - 0xb5
    "10110110", --  928 - 0x3a0  :  182 - 0xb6
    "10110111", --  929 - 0x3a1  :  183 - 0xb7
    "10110110", --  930 - 0x3a2  :  182 - 0xb6
    "10110111", --  931 - 0x3a3  :  183 - 0xb7
    "10110110", --  932 - 0x3a4  :  182 - 0xb6
    "10110111", --  933 - 0x3a5  :  183 - 0xb7
    "10110110", --  934 - 0x3a6  :  182 - 0xb6
    "10110111", --  935 - 0x3a7  :  183 - 0xb7
    "10110110", --  936 - 0x3a8  :  182 - 0xb6
    "10110111", --  937 - 0x3a9  :  183 - 0xb7
    "10110110", --  938 - 0x3aa  :  182 - 0xb6
    "10110111", --  939 - 0x3ab  :  183 - 0xb7
    "10110110", --  940 - 0x3ac  :  182 - 0xb6
    "10110111", --  941 - 0x3ad  :  183 - 0xb7
    "10110110", --  942 - 0x3ae  :  182 - 0xb6
    "10110111", --  943 - 0x3af  :  183 - 0xb7
    "10110110", --  944 - 0x3b0  :  182 - 0xb6
    "10110111", --  945 - 0x3b1  :  183 - 0xb7
    "10110110", --  946 - 0x3b2  :  182 - 0xb6
    "10110111", --  947 - 0x3b3  :  183 - 0xb7
    "10110110", --  948 - 0x3b4  :  182 - 0xb6
    "10110111", --  949 - 0x3b5  :  183 - 0xb7
    "10110110", --  950 - 0x3b6  :  182 - 0xb6
    "10110111", --  951 - 0x3b7  :  183 - 0xb7
    "10110110", --  952 - 0x3b8  :  182 - 0xb6
    "10110111", --  953 - 0x3b9  :  183 - 0xb7
    "10110110", --  954 - 0x3ba  :  182 - 0xb6
    "10110111", --  955 - 0x3bb  :  183 - 0xb7
    "10110110", --  956 - 0x3bc  :  182 - 0xb6
    "10110111", --  957 - 0x3bd  :  183 - 0xb7
    "10110110", --  958 - 0x3be  :  182 - 0xb6
    "10110111", --  959 - 0x3bf  :  183 - 0xb7
        ---- Attribute Table 0----
    "10101010", --  960 - 0x3c0  :  170 - 0xaa
    "10101010", --  961 - 0x3c1  :  170 - 0xaa
    "11101010", --  962 - 0x3c2  :  234 - 0xea
    "10101010", --  963 - 0x3c3  :  170 - 0xaa
    "10101010", --  964 - 0x3c4  :  170 - 0xaa
    "10101010", --  965 - 0x3c5  :  170 - 0xaa
    "10101010", --  966 - 0x3c6  :  170 - 0xaa
    "10101010", --  967 - 0x3c7  :  170 - 0xaa
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "01010101", --  969 - 0x3c9  :   85 - 0x55
    "01010101", --  970 - 0x3ca  :   85 - 0x55
    "01010101", --  971 - 0x3cb  :   85 - 0x55
    "01010101", --  972 - 0x3cc  :   85 - 0x55
    "01010101", --  973 - 0x3cd  :   85 - 0x55
    "01010101", --  974 - 0x3ce  :   85 - 0x55
    "01010101", --  975 - 0x3cf  :   85 - 0x55
    "01010101", --  976 - 0x3d0  :   85 - 0x55
    "01010101", --  977 - 0x3d1  :   85 - 0x55
    "01010101", --  978 - 0x3d2  :   85 - 0x55
    "01010101", --  979 - 0x3d3  :   85 - 0x55
    "01010101", --  980 - 0x3d4  :   85 - 0x55
    "01010101", --  981 - 0x3d5  :   85 - 0x55
    "01010101", --  982 - 0x3d6  :   85 - 0x55
    "01010101", --  983 - 0x3d7  :   85 - 0x55
    "01010101", --  984 - 0x3d8  :   85 - 0x55
    "01010101", --  985 - 0x3d9  :   85 - 0x55
    "01010101", --  986 - 0x3da  :   85 - 0x55
    "01010101", --  987 - 0x3db  :   85 - 0x55
    "01010101", --  988 - 0x3dc  :   85 - 0x55
    "01010101", --  989 - 0x3dd  :   85 - 0x55
    "01010101", --  990 - 0x3de  :   85 - 0x55
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "10011001", --  994 - 0x3e2  :  153 - 0x99
    "10101010", --  995 - 0x3e3  :  170 - 0xaa
    "10101010", --  996 - 0x3e4  :  170 - 0xaa
    "10101010", --  997 - 0x3e5  :  170 - 0xaa
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "10011001", -- 1002 - 0x3ea  :  153 - 0x99
    "10101010", -- 1003 - 0x3eb  :  170 - 0xaa
    "10101010", -- 1004 - 0x3ec  :  170 - 0xaa
    "10101010", -- 1005 - 0x3ed  :  170 - 0xaa
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "01010000", -- 1008 - 0x3f0  :   80 - 0x50
    "01010000", -- 1009 - 0x3f1  :   80 - 0x50
    "01010000", -- 1010 - 0x3f2  :   80 - 0x50
    "01010000", -- 1011 - 0x3f3  :   80 - 0x50
    "01010000", -- 1012 - 0x3f4  :   80 - 0x50
    "01010000", -- 1013 - 0x3f5  :   80 - 0x50
    "01010000", -- 1014 - 0x3f6  :   80 - 0x50
    "01010000", -- 1015 - 0x3f7  :   80 - 0x50
    "00000101", -- 1016 - 0x3f8  :    5 - 0x5
    "00000101", -- 1017 - 0x3f9  :    5 - 0x5
    "00000101", -- 1018 - 0x3fa  :    5 - 0x5
    "00000101", -- 1019 - 0x3fb  :    5 - 0x5
    "00000101", -- 1020 - 0x3fc  :    5 - 0x5
    "00000101", -- 1021 - 0x3fd  :    5 - 0x5
    "00000101", -- 1022 - 0x3fe  :    5 - 0x5
    "00000101", -- 1023 - 0x3ff  :    5 - 0x5
     ------- Name Table 1---------
    "00100100", -- 1024 - 0x400  :   36 - 0x24
    "00100100", -- 1025 - 0x401  :   36 - 0x24
    "00100100", -- 1026 - 0x402  :   36 - 0x24
    "00100100", -- 1027 - 0x403  :   36 - 0x24
    "00100100", -- 1028 - 0x404  :   36 - 0x24
    "00100100", -- 1029 - 0x405  :   36 - 0x24
    "00100100", -- 1030 - 0x406  :   36 - 0x24
    "00100100", -- 1031 - 0x407  :   36 - 0x24
    "00100100", -- 1032 - 0x408  :   36 - 0x24
    "00100100", -- 1033 - 0x409  :   36 - 0x24
    "00100100", -- 1034 - 0x40a  :   36 - 0x24
    "00100100", -- 1035 - 0x40b  :   36 - 0x24
    "00100100", -- 1036 - 0x40c  :   36 - 0x24
    "00100100", -- 1037 - 0x40d  :   36 - 0x24
    "00100100", -- 1038 - 0x40e  :   36 - 0x24
    "00100100", -- 1039 - 0x40f  :   36 - 0x24
    "00100100", -- 1040 - 0x410  :   36 - 0x24
    "00100100", -- 1041 - 0x411  :   36 - 0x24
    "00100100", -- 1042 - 0x412  :   36 - 0x24
    "00100100", -- 1043 - 0x413  :   36 - 0x24
    "00100100", -- 1044 - 0x414  :   36 - 0x24
    "00100100", -- 1045 - 0x415  :   36 - 0x24
    "00100100", -- 1046 - 0x416  :   36 - 0x24
    "00100100", -- 1047 - 0x417  :   36 - 0x24
    "00100100", -- 1048 - 0x418  :   36 - 0x24
    "00100100", -- 1049 - 0x419  :   36 - 0x24
    "00100100", -- 1050 - 0x41a  :   36 - 0x24
    "00100100", -- 1051 - 0x41b  :   36 - 0x24
    "00100100", -- 1052 - 0x41c  :   36 - 0x24
    "00100100", -- 1053 - 0x41d  :   36 - 0x24
    "00100100", -- 1054 - 0x41e  :   36 - 0x24
    "00100100", -- 1055 - 0x41f  :   36 - 0x24
    "00100100", -- 1056 - 0x420  :   36 - 0x24
    "00100100", -- 1057 - 0x421  :   36 - 0x24
    "00100100", -- 1058 - 0x422  :   36 - 0x24
    "00100100", -- 1059 - 0x423  :   36 - 0x24
    "00100100", -- 1060 - 0x424  :   36 - 0x24
    "00100100", -- 1061 - 0x425  :   36 - 0x24
    "00100100", -- 1062 - 0x426  :   36 - 0x24
    "00100100", -- 1063 - 0x427  :   36 - 0x24
    "00100100", -- 1064 - 0x428  :   36 - 0x24
    "00100100", -- 1065 - 0x429  :   36 - 0x24
    "00100100", -- 1066 - 0x42a  :   36 - 0x24
    "00100100", -- 1067 - 0x42b  :   36 - 0x24
    "00100100", -- 1068 - 0x42c  :   36 - 0x24
    "00100100", -- 1069 - 0x42d  :   36 - 0x24
    "00100100", -- 1070 - 0x42e  :   36 - 0x24
    "00100100", -- 1071 - 0x42f  :   36 - 0x24
    "00100100", -- 1072 - 0x430  :   36 - 0x24
    "00100100", -- 1073 - 0x431  :   36 - 0x24
    "00100100", -- 1074 - 0x432  :   36 - 0x24
    "00100100", -- 1075 - 0x433  :   36 - 0x24
    "00100100", -- 1076 - 0x434  :   36 - 0x24
    "00100100", -- 1077 - 0x435  :   36 - 0x24
    "00100100", -- 1078 - 0x436  :   36 - 0x24
    "00100100", -- 1079 - 0x437  :   36 - 0x24
    "00100100", -- 1080 - 0x438  :   36 - 0x24
    "00100100", -- 1081 - 0x439  :   36 - 0x24
    "00100100", -- 1082 - 0x43a  :   36 - 0x24
    "00100100", -- 1083 - 0x43b  :   36 - 0x24
    "00100100", -- 1084 - 0x43c  :   36 - 0x24
    "00100100", -- 1085 - 0x43d  :   36 - 0x24
    "00100100", -- 1086 - 0x43e  :   36 - 0x24
    "00100100", -- 1087 - 0x43f  :   36 - 0x24
    "00100100", -- 1088 - 0x440  :   36 - 0x24
    "00100100", -- 1089 - 0x441  :   36 - 0x24
    "00100100", -- 1090 - 0x442  :   36 - 0x24
    "00100100", -- 1091 - 0x443  :   36 - 0x24
    "00100100", -- 1092 - 0x444  :   36 - 0x24
    "00100100", -- 1093 - 0x445  :   36 - 0x24
    "00100100", -- 1094 - 0x446  :   36 - 0x24
    "00100100", -- 1095 - 0x447  :   36 - 0x24
    "00100100", -- 1096 - 0x448  :   36 - 0x24
    "00100100", -- 1097 - 0x449  :   36 - 0x24
    "00100100", -- 1098 - 0x44a  :   36 - 0x24
    "00100100", -- 1099 - 0x44b  :   36 - 0x24
    "00100100", -- 1100 - 0x44c  :   36 - 0x24
    "00100100", -- 1101 - 0x44d  :   36 - 0x24
    "00100100", -- 1102 - 0x44e  :   36 - 0x24
    "00100100", -- 1103 - 0x44f  :   36 - 0x24
    "00100100", -- 1104 - 0x450  :   36 - 0x24
    "00100100", -- 1105 - 0x451  :   36 - 0x24
    "00100100", -- 1106 - 0x452  :   36 - 0x24
    "00100100", -- 1107 - 0x453  :   36 - 0x24
    "00100100", -- 1108 - 0x454  :   36 - 0x24
    "00100100", -- 1109 - 0x455  :   36 - 0x24
    "00100100", -- 1110 - 0x456  :   36 - 0x24
    "00100100", -- 1111 - 0x457  :   36 - 0x24
    "00100100", -- 1112 - 0x458  :   36 - 0x24
    "00100100", -- 1113 - 0x459  :   36 - 0x24
    "00100100", -- 1114 - 0x45a  :   36 - 0x24
    "00100100", -- 1115 - 0x45b  :   36 - 0x24
    "00100100", -- 1116 - 0x45c  :   36 - 0x24
    "00100100", -- 1117 - 0x45d  :   36 - 0x24
    "00100100", -- 1118 - 0x45e  :   36 - 0x24
    "00100100", -- 1119 - 0x45f  :   36 - 0x24
    "00100100", -- 1120 - 0x460  :   36 - 0x24
    "00100100", -- 1121 - 0x461  :   36 - 0x24
    "00100100", -- 1122 - 0x462  :   36 - 0x24
    "00100100", -- 1123 - 0x463  :   36 - 0x24
    "00100100", -- 1124 - 0x464  :   36 - 0x24
    "00100100", -- 1125 - 0x465  :   36 - 0x24
    "00100100", -- 1126 - 0x466  :   36 - 0x24
    "00100100", -- 1127 - 0x467  :   36 - 0x24
    "00100100", -- 1128 - 0x468  :   36 - 0x24
    "00100100", -- 1129 - 0x469  :   36 - 0x24
    "00100100", -- 1130 - 0x46a  :   36 - 0x24
    "00100100", -- 1131 - 0x46b  :   36 - 0x24
    "00100100", -- 1132 - 0x46c  :   36 - 0x24
    "00100100", -- 1133 - 0x46d  :   36 - 0x24
    "00100100", -- 1134 - 0x46e  :   36 - 0x24
    "00100100", -- 1135 - 0x46f  :   36 - 0x24
    "00100100", -- 1136 - 0x470  :   36 - 0x24
    "00100100", -- 1137 - 0x471  :   36 - 0x24
    "00100100", -- 1138 - 0x472  :   36 - 0x24
    "00100100", -- 1139 - 0x473  :   36 - 0x24
    "00100100", -- 1140 - 0x474  :   36 - 0x24
    "00100100", -- 1141 - 0x475  :   36 - 0x24
    "00100100", -- 1142 - 0x476  :   36 - 0x24
    "00100100", -- 1143 - 0x477  :   36 - 0x24
    "00100100", -- 1144 - 0x478  :   36 - 0x24
    "00100100", -- 1145 - 0x479  :   36 - 0x24
    "00100100", -- 1146 - 0x47a  :   36 - 0x24
    "00100100", -- 1147 - 0x47b  :   36 - 0x24
    "00100100", -- 1148 - 0x47c  :   36 - 0x24
    "00100100", -- 1149 - 0x47d  :   36 - 0x24
    "00100100", -- 1150 - 0x47e  :   36 - 0x24
    "00100100", -- 1151 - 0x47f  :   36 - 0x24
    "00100100", -- 1152 - 0x480  :   36 - 0x24
    "00100100", -- 1153 - 0x481  :   36 - 0x24
    "00100100", -- 1154 - 0x482  :   36 - 0x24
    "00100100", -- 1155 - 0x483  :   36 - 0x24
    "00100100", -- 1156 - 0x484  :   36 - 0x24
    "00100100", -- 1157 - 0x485  :   36 - 0x24
    "00100100", -- 1158 - 0x486  :   36 - 0x24
    "00100100", -- 1159 - 0x487  :   36 - 0x24
    "00110110", -- 1160 - 0x488  :   54 - 0x36
    "00110111", -- 1161 - 0x489  :   55 - 0x37
    "00100100", -- 1162 - 0x48a  :   36 - 0x24
    "00100100", -- 1163 - 0x48b  :   36 - 0x24
    "00100100", -- 1164 - 0x48c  :   36 - 0x24
    "00100100", -- 1165 - 0x48d  :   36 - 0x24
    "00100100", -- 1166 - 0x48e  :   36 - 0x24
    "00100100", -- 1167 - 0x48f  :   36 - 0x24
    "00100100", -- 1168 - 0x490  :   36 - 0x24
    "00100100", -- 1169 - 0x491  :   36 - 0x24
    "00100100", -- 1170 - 0x492  :   36 - 0x24
    "00100100", -- 1171 - 0x493  :   36 - 0x24
    "00100100", -- 1172 - 0x494  :   36 - 0x24
    "00100100", -- 1173 - 0x495  :   36 - 0x24
    "00100100", -- 1174 - 0x496  :   36 - 0x24
    "00100100", -- 1175 - 0x497  :   36 - 0x24
    "00100100", -- 1176 - 0x498  :   36 - 0x24
    "00100100", -- 1177 - 0x499  :   36 - 0x24
    "00100100", -- 1178 - 0x49a  :   36 - 0x24
    "00100100", -- 1179 - 0x49b  :   36 - 0x24
    "00100100", -- 1180 - 0x49c  :   36 - 0x24
    "00100100", -- 1181 - 0x49d  :   36 - 0x24
    "00100100", -- 1182 - 0x49e  :   36 - 0x24
    "00100100", -- 1183 - 0x49f  :   36 - 0x24
    "00100100", -- 1184 - 0x4a0  :   36 - 0x24
    "00100100", -- 1185 - 0x4a1  :   36 - 0x24
    "00100100", -- 1186 - 0x4a2  :   36 - 0x24
    "00100100", -- 1187 - 0x4a3  :   36 - 0x24
    "00100100", -- 1188 - 0x4a4  :   36 - 0x24
    "00100100", -- 1189 - 0x4a5  :   36 - 0x24
    "00100100", -- 1190 - 0x4a6  :   36 - 0x24
    "00110101", -- 1191 - 0x4a7  :   53 - 0x35
    "00100101", -- 1192 - 0x4a8  :   37 - 0x25
    "00100101", -- 1193 - 0x4a9  :   37 - 0x25
    "00111000", -- 1194 - 0x4aa  :   56 - 0x38
    "00100100", -- 1195 - 0x4ab  :   36 - 0x24
    "00100100", -- 1196 - 0x4ac  :   36 - 0x24
    "00100100", -- 1197 - 0x4ad  :   36 - 0x24
    "00100100", -- 1198 - 0x4ae  :   36 - 0x24
    "00100100", -- 1199 - 0x4af  :   36 - 0x24
    "00100100", -- 1200 - 0x4b0  :   36 - 0x24
    "00100100", -- 1201 - 0x4b1  :   36 - 0x24
    "00100100", -- 1202 - 0x4b2  :   36 - 0x24
    "00100100", -- 1203 - 0x4b3  :   36 - 0x24
    "00100100", -- 1204 - 0x4b4  :   36 - 0x24
    "00100100", -- 1205 - 0x4b5  :   36 - 0x24
    "00100100", -- 1206 - 0x4b6  :   36 - 0x24
    "00100100", -- 1207 - 0x4b7  :   36 - 0x24
    "00100100", -- 1208 - 0x4b8  :   36 - 0x24
    "00100100", -- 1209 - 0x4b9  :   36 - 0x24
    "00100100", -- 1210 - 0x4ba  :   36 - 0x24
    "00100100", -- 1211 - 0x4bb  :   36 - 0x24
    "00100100", -- 1212 - 0x4bc  :   36 - 0x24
    "00100100", -- 1213 - 0x4bd  :   36 - 0x24
    "00100100", -- 1214 - 0x4be  :   36 - 0x24
    "00100100", -- 1215 - 0x4bf  :   36 - 0x24
    "00100100", -- 1216 - 0x4c0  :   36 - 0x24
    "00100100", -- 1217 - 0x4c1  :   36 - 0x24
    "00100100", -- 1218 - 0x4c2  :   36 - 0x24
    "00100100", -- 1219 - 0x4c3  :   36 - 0x24
    "00100100", -- 1220 - 0x4c4  :   36 - 0x24
    "00100100", -- 1221 - 0x4c5  :   36 - 0x24
    "00100100", -- 1222 - 0x4c6  :   36 - 0x24
    "00111001", -- 1223 - 0x4c7  :   57 - 0x39
    "00111010", -- 1224 - 0x4c8  :   58 - 0x3a
    "00111011", -- 1225 - 0x4c9  :   59 - 0x3b
    "00111100", -- 1226 - 0x4ca  :   60 - 0x3c
    "00100100", -- 1227 - 0x4cb  :   36 - 0x24
    "00100100", -- 1228 - 0x4cc  :   36 - 0x24
    "00100100", -- 1229 - 0x4cd  :   36 - 0x24
    "00100100", -- 1230 - 0x4ce  :   36 - 0x24
    "00100100", -- 1231 - 0x4cf  :   36 - 0x24
    "00100100", -- 1232 - 0x4d0  :   36 - 0x24
    "00100100", -- 1233 - 0x4d1  :   36 - 0x24
    "00100100", -- 1234 - 0x4d2  :   36 - 0x24
    "00100100", -- 1235 - 0x4d3  :   36 - 0x24
    "00100100", -- 1236 - 0x4d4  :   36 - 0x24
    "00100100", -- 1237 - 0x4d5  :   36 - 0x24
    "00100100", -- 1238 - 0x4d6  :   36 - 0x24
    "00100100", -- 1239 - 0x4d7  :   36 - 0x24
    "00100100", -- 1240 - 0x4d8  :   36 - 0x24
    "00100100", -- 1241 - 0x4d9  :   36 - 0x24
    "00100100", -- 1242 - 0x4da  :   36 - 0x24
    "00100100", -- 1243 - 0x4db  :   36 - 0x24
    "00100100", -- 1244 - 0x4dc  :   36 - 0x24
    "00100100", -- 1245 - 0x4dd  :   36 - 0x24
    "00100100", -- 1246 - 0x4de  :   36 - 0x24
    "00100100", -- 1247 - 0x4df  :   36 - 0x24
    "00100100", -- 1248 - 0x4e0  :   36 - 0x24
    "00100100", -- 1249 - 0x4e1  :   36 - 0x24
    "00100100", -- 1250 - 0x4e2  :   36 - 0x24
    "00100100", -- 1251 - 0x4e3  :   36 - 0x24
    "00100100", -- 1252 - 0x4e4  :   36 - 0x24
    "00100100", -- 1253 - 0x4e5  :   36 - 0x24
    "00100100", -- 1254 - 0x4e6  :   36 - 0x24
    "00100100", -- 1255 - 0x4e7  :   36 - 0x24
    "00100100", -- 1256 - 0x4e8  :   36 - 0x24
    "00100100", -- 1257 - 0x4e9  :   36 - 0x24
    "00100100", -- 1258 - 0x4ea  :   36 - 0x24
    "00100100", -- 1259 - 0x4eb  :   36 - 0x24
    "00100100", -- 1260 - 0x4ec  :   36 - 0x24
    "00100100", -- 1261 - 0x4ed  :   36 - 0x24
    "00100100", -- 1262 - 0x4ee  :   36 - 0x24
    "00100100", -- 1263 - 0x4ef  :   36 - 0x24
    "00100100", -- 1264 - 0x4f0  :   36 - 0x24
    "00100100", -- 1265 - 0x4f1  :   36 - 0x24
    "00100100", -- 1266 - 0x4f2  :   36 - 0x24
    "00100100", -- 1267 - 0x4f3  :   36 - 0x24
    "00100100", -- 1268 - 0x4f4  :   36 - 0x24
    "00100100", -- 1269 - 0x4f5  :   36 - 0x24
    "00100100", -- 1270 - 0x4f6  :   36 - 0x24
    "00100100", -- 1271 - 0x4f7  :   36 - 0x24
    "00100100", -- 1272 - 0x4f8  :   36 - 0x24
    "00100100", -- 1273 - 0x4f9  :   36 - 0x24
    "00100100", -- 1274 - 0x4fa  :   36 - 0x24
    "00100100", -- 1275 - 0x4fb  :   36 - 0x24
    "00100100", -- 1276 - 0x4fc  :   36 - 0x24
    "00100100", -- 1277 - 0x4fd  :   36 - 0x24
    "00100100", -- 1278 - 0x4fe  :   36 - 0x24
    "00100100", -- 1279 - 0x4ff  :   36 - 0x24
    "00100100", -- 1280 - 0x500  :   36 - 0x24
    "00100100", -- 1281 - 0x501  :   36 - 0x24
    "00100100", -- 1282 - 0x502  :   36 - 0x24
    "00100100", -- 1283 - 0x503  :   36 - 0x24
    "00100100", -- 1284 - 0x504  :   36 - 0x24
    "00100100", -- 1285 - 0x505  :   36 - 0x24
    "00100100", -- 1286 - 0x506  :   36 - 0x24
    "00100100", -- 1287 - 0x507  :   36 - 0x24
    "00100100", -- 1288 - 0x508  :   36 - 0x24
    "00100100", -- 1289 - 0x509  :   36 - 0x24
    "00100100", -- 1290 - 0x50a  :   36 - 0x24
    "00100100", -- 1291 - 0x50b  :   36 - 0x24
    "00100100", -- 1292 - 0x50c  :   36 - 0x24
    "00100100", -- 1293 - 0x50d  :   36 - 0x24
    "00100100", -- 1294 - 0x50e  :   36 - 0x24
    "00100100", -- 1295 - 0x50f  :   36 - 0x24
    "00100100", -- 1296 - 0x510  :   36 - 0x24
    "00100100", -- 1297 - 0x511  :   36 - 0x24
    "00100100", -- 1298 - 0x512  :   36 - 0x24
    "00100100", -- 1299 - 0x513  :   36 - 0x24
    "00100100", -- 1300 - 0x514  :   36 - 0x24
    "00100100", -- 1301 - 0x515  :   36 - 0x24
    "00100100", -- 1302 - 0x516  :   36 - 0x24
    "00100100", -- 1303 - 0x517  :   36 - 0x24
    "00100100", -- 1304 - 0x518  :   36 - 0x24
    "00100100", -- 1305 - 0x519  :   36 - 0x24
    "00100100", -- 1306 - 0x51a  :   36 - 0x24
    "00100100", -- 1307 - 0x51b  :   36 - 0x24
    "00100100", -- 1308 - 0x51c  :   36 - 0x24
    "00100100", -- 1309 - 0x51d  :   36 - 0x24
    "00100100", -- 1310 - 0x51e  :   36 - 0x24
    "00100100", -- 1311 - 0x51f  :   36 - 0x24
    "00100100", -- 1312 - 0x520  :   36 - 0x24
    "00100100", -- 1313 - 0x521  :   36 - 0x24
    "00100100", -- 1314 - 0x522  :   36 - 0x24
    "00100100", -- 1315 - 0x523  :   36 - 0x24
    "00100100", -- 1316 - 0x524  :   36 - 0x24
    "00100100", -- 1317 - 0x525  :   36 - 0x24
    "00100100", -- 1318 - 0x526  :   36 - 0x24
    "00100100", -- 1319 - 0x527  :   36 - 0x24
    "00100100", -- 1320 - 0x528  :   36 - 0x24
    "00100100", -- 1321 - 0x529  :   36 - 0x24
    "00100100", -- 1322 - 0x52a  :   36 - 0x24
    "00100100", -- 1323 - 0x52b  :   36 - 0x24
    "00100100", -- 1324 - 0x52c  :   36 - 0x24
    "00100100", -- 1325 - 0x52d  :   36 - 0x24
    "00100100", -- 1326 - 0x52e  :   36 - 0x24
    "00100100", -- 1327 - 0x52f  :   36 - 0x24
    "00100100", -- 1328 - 0x530  :   36 - 0x24
    "00100100", -- 1329 - 0x531  :   36 - 0x24
    "00100100", -- 1330 - 0x532  :   36 - 0x24
    "00100100", -- 1331 - 0x533  :   36 - 0x24
    "00100100", -- 1332 - 0x534  :   36 - 0x24
    "00100100", -- 1333 - 0x535  :   36 - 0x24
    "00100100", -- 1334 - 0x536  :   36 - 0x24
    "00100100", -- 1335 - 0x537  :   36 - 0x24
    "00100100", -- 1336 - 0x538  :   36 - 0x24
    "00100100", -- 1337 - 0x539  :   36 - 0x24
    "00100100", -- 1338 - 0x53a  :   36 - 0x24
    "00100100", -- 1339 - 0x53b  :   36 - 0x24
    "00100100", -- 1340 - 0x53c  :   36 - 0x24
    "00100100", -- 1341 - 0x53d  :   36 - 0x24
    "00100100", -- 1342 - 0x53e  :   36 - 0x24
    "00100100", -- 1343 - 0x53f  :   36 - 0x24
    "00100100", -- 1344 - 0x540  :   36 - 0x24
    "00100100", -- 1345 - 0x541  :   36 - 0x24
    "00100100", -- 1346 - 0x542  :   36 - 0x24
    "00100100", -- 1347 - 0x543  :   36 - 0x24
    "00100100", -- 1348 - 0x544  :   36 - 0x24
    "00100100", -- 1349 - 0x545  :   36 - 0x24
    "00100100", -- 1350 - 0x546  :   36 - 0x24
    "00100100", -- 1351 - 0x547  :   36 - 0x24
    "00100100", -- 1352 - 0x548  :   36 - 0x24
    "00100100", -- 1353 - 0x549  :   36 - 0x24
    "00100100", -- 1354 - 0x54a  :   36 - 0x24
    "00100100", -- 1355 - 0x54b  :   36 - 0x24
    "01010011", -- 1356 - 0x54c  :   83 - 0x53
    "01010100", -- 1357 - 0x54d  :   84 - 0x54
    "00100100", -- 1358 - 0x54e  :   36 - 0x24
    "00100100", -- 1359 - 0x54f  :   36 - 0x24
    "00100100", -- 1360 - 0x550  :   36 - 0x24
    "00100100", -- 1361 - 0x551  :   36 - 0x24
    "00100100", -- 1362 - 0x552  :   36 - 0x24
    "00100100", -- 1363 - 0x553  :   36 - 0x24
    "00100100", -- 1364 - 0x554  :   36 - 0x24
    "00100100", -- 1365 - 0x555  :   36 - 0x24
    "00100100", -- 1366 - 0x556  :   36 - 0x24
    "00100100", -- 1367 - 0x557  :   36 - 0x24
    "00100100", -- 1368 - 0x558  :   36 - 0x24
    "00100100", -- 1369 - 0x559  :   36 - 0x24
    "00100100", -- 1370 - 0x55a  :   36 - 0x24
    "00100100", -- 1371 - 0x55b  :   36 - 0x24
    "00100100", -- 1372 - 0x55c  :   36 - 0x24
    "00100100", -- 1373 - 0x55d  :   36 - 0x24
    "00100100", -- 1374 - 0x55e  :   36 - 0x24
    "00100100", -- 1375 - 0x55f  :   36 - 0x24
    "00100100", -- 1376 - 0x560  :   36 - 0x24
    "00100100", -- 1377 - 0x561  :   36 - 0x24
    "00100100", -- 1378 - 0x562  :   36 - 0x24
    "00100100", -- 1379 - 0x563  :   36 - 0x24
    "00100100", -- 1380 - 0x564  :   36 - 0x24
    "00100100", -- 1381 - 0x565  :   36 - 0x24
    "00100100", -- 1382 - 0x566  :   36 - 0x24
    "00100100", -- 1383 - 0x567  :   36 - 0x24
    "00100100", -- 1384 - 0x568  :   36 - 0x24
    "00100100", -- 1385 - 0x569  :   36 - 0x24
    "00100100", -- 1386 - 0x56a  :   36 - 0x24
    "00100100", -- 1387 - 0x56b  :   36 - 0x24
    "01010101", -- 1388 - 0x56c  :   85 - 0x55
    "01010110", -- 1389 - 0x56d  :   86 - 0x56
    "00100100", -- 1390 - 0x56e  :   36 - 0x24
    "00100100", -- 1391 - 0x56f  :   36 - 0x24
    "00100100", -- 1392 - 0x570  :   36 - 0x24
    "00100100", -- 1393 - 0x571  :   36 - 0x24
    "00100100", -- 1394 - 0x572  :   36 - 0x24
    "00100100", -- 1395 - 0x573  :   36 - 0x24
    "00100100", -- 1396 - 0x574  :   36 - 0x24
    "00100100", -- 1397 - 0x575  :   36 - 0x24
    "00100100", -- 1398 - 0x576  :   36 - 0x24
    "00100100", -- 1399 - 0x577  :   36 - 0x24
    "00100100", -- 1400 - 0x578  :   36 - 0x24
    "00100100", -- 1401 - 0x579  :   36 - 0x24
    "00100100", -- 1402 - 0x57a  :   36 - 0x24
    "00100100", -- 1403 - 0x57b  :   36 - 0x24
    "00100100", -- 1404 - 0x57c  :   36 - 0x24
    "00100100", -- 1405 - 0x57d  :   36 - 0x24
    "00100100", -- 1406 - 0x57e  :   36 - 0x24
    "00100100", -- 1407 - 0x57f  :   36 - 0x24
    "00100100", -- 1408 - 0x580  :   36 - 0x24
    "00100100", -- 1409 - 0x581  :   36 - 0x24
    "00100100", -- 1410 - 0x582  :   36 - 0x24
    "00100100", -- 1411 - 0x583  :   36 - 0x24
    "00100100", -- 1412 - 0x584  :   36 - 0x24
    "00100100", -- 1413 - 0x585  :   36 - 0x24
    "00100100", -- 1414 - 0x586  :   36 - 0x24
    "00100100", -- 1415 - 0x587  :   36 - 0x24
    "00100100", -- 1416 - 0x588  :   36 - 0x24
    "00100100", -- 1417 - 0x589  :   36 - 0x24
    "00100100", -- 1418 - 0x58a  :   36 - 0x24
    "00100100", -- 1419 - 0x58b  :   36 - 0x24
    "00100100", -- 1420 - 0x58c  :   36 - 0x24
    "00100100", -- 1421 - 0x58d  :   36 - 0x24
    "00100100", -- 1422 - 0x58e  :   36 - 0x24
    "00100100", -- 1423 - 0x58f  :   36 - 0x24
    "00100100", -- 1424 - 0x590  :   36 - 0x24
    "00100100", -- 1425 - 0x591  :   36 - 0x24
    "00100100", -- 1426 - 0x592  :   36 - 0x24
    "00100100", -- 1427 - 0x593  :   36 - 0x24
    "00100100", -- 1428 - 0x594  :   36 - 0x24
    "00100100", -- 1429 - 0x595  :   36 - 0x24
    "00100100", -- 1430 - 0x596  :   36 - 0x24
    "00100100", -- 1431 - 0x597  :   36 - 0x24
    "00100100", -- 1432 - 0x598  :   36 - 0x24
    "00100100", -- 1433 - 0x599  :   36 - 0x24
    "00100100", -- 1434 - 0x59a  :   36 - 0x24
    "00100100", -- 1435 - 0x59b  :   36 - 0x24
    "00100100", -- 1436 - 0x59c  :   36 - 0x24
    "00100100", -- 1437 - 0x59d  :   36 - 0x24
    "00100100", -- 1438 - 0x59e  :   36 - 0x24
    "00100100", -- 1439 - 0x59f  :   36 - 0x24
    "00100100", -- 1440 - 0x5a0  :   36 - 0x24
    "00100100", -- 1441 - 0x5a1  :   36 - 0x24
    "00100100", -- 1442 - 0x5a2  :   36 - 0x24
    "00100100", -- 1443 - 0x5a3  :   36 - 0x24
    "00100100", -- 1444 - 0x5a4  :   36 - 0x24
    "00100100", -- 1445 - 0x5a5  :   36 - 0x24
    "00100100", -- 1446 - 0x5a6  :   36 - 0x24
    "00100100", -- 1447 - 0x5a7  :   36 - 0x24
    "00100100", -- 1448 - 0x5a8  :   36 - 0x24
    "00100100", -- 1449 - 0x5a9  :   36 - 0x24
    "00100100", -- 1450 - 0x5aa  :   36 - 0x24
    "00100100", -- 1451 - 0x5ab  :   36 - 0x24
    "00100100", -- 1452 - 0x5ac  :   36 - 0x24
    "00100100", -- 1453 - 0x5ad  :   36 - 0x24
    "00100100", -- 1454 - 0x5ae  :   36 - 0x24
    "00100100", -- 1455 - 0x5af  :   36 - 0x24
    "00100100", -- 1456 - 0x5b0  :   36 - 0x24
    "00100100", -- 1457 - 0x5b1  :   36 - 0x24
    "00100100", -- 1458 - 0x5b2  :   36 - 0x24
    "00100100", -- 1459 - 0x5b3  :   36 - 0x24
    "00100100", -- 1460 - 0x5b4  :   36 - 0x24
    "00100100", -- 1461 - 0x5b5  :   36 - 0x24
    "00100100", -- 1462 - 0x5b6  :   36 - 0x24
    "00100100", -- 1463 - 0x5b7  :   36 - 0x24
    "00100100", -- 1464 - 0x5b8  :   36 - 0x24
    "00100100", -- 1465 - 0x5b9  :   36 - 0x24
    "00100100", -- 1466 - 0x5ba  :   36 - 0x24
    "00100100", -- 1467 - 0x5bb  :   36 - 0x24
    "00100100", -- 1468 - 0x5bc  :   36 - 0x24
    "00100100", -- 1469 - 0x5bd  :   36 - 0x24
    "00100100", -- 1470 - 0x5be  :   36 - 0x24
    "00100100", -- 1471 - 0x5bf  :   36 - 0x24
    "00100100", -- 1472 - 0x5c0  :   36 - 0x24
    "00100100", -- 1473 - 0x5c1  :   36 - 0x24
    "00100100", -- 1474 - 0x5c2  :   36 - 0x24
    "00100100", -- 1475 - 0x5c3  :   36 - 0x24
    "00100100", -- 1476 - 0x5c4  :   36 - 0x24
    "00100100", -- 1477 - 0x5c5  :   36 - 0x24
    "00100100", -- 1478 - 0x5c6  :   36 - 0x24
    "00100100", -- 1479 - 0x5c7  :   36 - 0x24
    "00100100", -- 1480 - 0x5c8  :   36 - 0x24
    "00100100", -- 1481 - 0x5c9  :   36 - 0x24
    "00100100", -- 1482 - 0x5ca  :   36 - 0x24
    "00100100", -- 1483 - 0x5cb  :   36 - 0x24
    "00100100", -- 1484 - 0x5cc  :   36 - 0x24
    "00100100", -- 1485 - 0x5cd  :   36 - 0x24
    "00100100", -- 1486 - 0x5ce  :   36 - 0x24
    "00100100", -- 1487 - 0x5cf  :   36 - 0x24
    "00100100", -- 1488 - 0x5d0  :   36 - 0x24
    "00100100", -- 1489 - 0x5d1  :   36 - 0x24
    "00100100", -- 1490 - 0x5d2  :   36 - 0x24
    "00100100", -- 1491 - 0x5d3  :   36 - 0x24
    "00100100", -- 1492 - 0x5d4  :   36 - 0x24
    "00100100", -- 1493 - 0x5d5  :   36 - 0x24
    "00100100", -- 1494 - 0x5d6  :   36 - 0x24
    "00100100", -- 1495 - 0x5d7  :   36 - 0x24
    "00100100", -- 1496 - 0x5d8  :   36 - 0x24
    "00100100", -- 1497 - 0x5d9  :   36 - 0x24
    "00100100", -- 1498 - 0x5da  :   36 - 0x24
    "00100100", -- 1499 - 0x5db  :   36 - 0x24
    "00100100", -- 1500 - 0x5dc  :   36 - 0x24
    "00100100", -- 1501 - 0x5dd  :   36 - 0x24
    "00100100", -- 1502 - 0x5de  :   36 - 0x24
    "00100100", -- 1503 - 0x5df  :   36 - 0x24
    "00100100", -- 1504 - 0x5e0  :   36 - 0x24
    "00100100", -- 1505 - 0x5e1  :   36 - 0x24
    "00100100", -- 1506 - 0x5e2  :   36 - 0x24
    "00100100", -- 1507 - 0x5e3  :   36 - 0x24
    "00100100", -- 1508 - 0x5e4  :   36 - 0x24
    "00100100", -- 1509 - 0x5e5  :   36 - 0x24
    "00100100", -- 1510 - 0x5e6  :   36 - 0x24
    "00100100", -- 1511 - 0x5e7  :   36 - 0x24
    "00100100", -- 1512 - 0x5e8  :   36 - 0x24
    "00100100", -- 1513 - 0x5e9  :   36 - 0x24
    "00100100", -- 1514 - 0x5ea  :   36 - 0x24
    "00100100", -- 1515 - 0x5eb  :   36 - 0x24
    "00100100", -- 1516 - 0x5ec  :   36 - 0x24
    "00100100", -- 1517 - 0x5ed  :   36 - 0x24
    "00100100", -- 1518 - 0x5ee  :   36 - 0x24
    "00100100", -- 1519 - 0x5ef  :   36 - 0x24
    "00100100", -- 1520 - 0x5f0  :   36 - 0x24
    "00100100", -- 1521 - 0x5f1  :   36 - 0x24
    "00100100", -- 1522 - 0x5f2  :   36 - 0x24
    "00100100", -- 1523 - 0x5f3  :   36 - 0x24
    "00100100", -- 1524 - 0x5f4  :   36 - 0x24
    "00100100", -- 1525 - 0x5f5  :   36 - 0x24
    "00100100", -- 1526 - 0x5f6  :   36 - 0x24
    "00100100", -- 1527 - 0x5f7  :   36 - 0x24
    "00100100", -- 1528 - 0x5f8  :   36 - 0x24
    "00100100", -- 1529 - 0x5f9  :   36 - 0x24
    "00100100", -- 1530 - 0x5fa  :   36 - 0x24
    "00100100", -- 1531 - 0x5fb  :   36 - 0x24
    "00100100", -- 1532 - 0x5fc  :   36 - 0x24
    "00100100", -- 1533 - 0x5fd  :   36 - 0x24
    "00100100", -- 1534 - 0x5fe  :   36 - 0x24
    "00100100", -- 1535 - 0x5ff  :   36 - 0x24
    "00100100", -- 1536 - 0x600  :   36 - 0x24
    "00100100", -- 1537 - 0x601  :   36 - 0x24
    "00100100", -- 1538 - 0x602  :   36 - 0x24
    "00100100", -- 1539 - 0x603  :   36 - 0x24
    "00100100", -- 1540 - 0x604  :   36 - 0x24
    "00100100", -- 1541 - 0x605  :   36 - 0x24
    "00100100", -- 1542 - 0x606  :   36 - 0x24
    "00100100", -- 1543 - 0x607  :   36 - 0x24
    "00100100", -- 1544 - 0x608  :   36 - 0x24
    "00100100", -- 1545 - 0x609  :   36 - 0x24
    "00100100", -- 1546 - 0x60a  :   36 - 0x24
    "00100100", -- 1547 - 0x60b  :   36 - 0x24
    "00100100", -- 1548 - 0x60c  :   36 - 0x24
    "00100100", -- 1549 - 0x60d  :   36 - 0x24
    "00100100", -- 1550 - 0x60e  :   36 - 0x24
    "00100100", -- 1551 - 0x60f  :   36 - 0x24
    "00100100", -- 1552 - 0x610  :   36 - 0x24
    "00100100", -- 1553 - 0x611  :   36 - 0x24
    "00100100", -- 1554 - 0x612  :   36 - 0x24
    "00100100", -- 1555 - 0x613  :   36 - 0x24
    "00100100", -- 1556 - 0x614  :   36 - 0x24
    "00100100", -- 1557 - 0x615  :   36 - 0x24
    "00100100", -- 1558 - 0x616  :   36 - 0x24
    "00100100", -- 1559 - 0x617  :   36 - 0x24
    "00100100", -- 1560 - 0x618  :   36 - 0x24
    "00100100", -- 1561 - 0x619  :   36 - 0x24
    "00100100", -- 1562 - 0x61a  :   36 - 0x24
    "00100100", -- 1563 - 0x61b  :   36 - 0x24
    "00100100", -- 1564 - 0x61c  :   36 - 0x24
    "00100100", -- 1565 - 0x61d  :   36 - 0x24
    "00100100", -- 1566 - 0x61e  :   36 - 0x24
    "00100100", -- 1567 - 0x61f  :   36 - 0x24
    "00100100", -- 1568 - 0x620  :   36 - 0x24
    "00100100", -- 1569 - 0x621  :   36 - 0x24
    "00100100", -- 1570 - 0x622  :   36 - 0x24
    "00100100", -- 1571 - 0x623  :   36 - 0x24
    "00100100", -- 1572 - 0x624  :   36 - 0x24
    "00100100", -- 1573 - 0x625  :   36 - 0x24
    "00100100", -- 1574 - 0x626  :   36 - 0x24
    "00100100", -- 1575 - 0x627  :   36 - 0x24
    "00100100", -- 1576 - 0x628  :   36 - 0x24
    "00100100", -- 1577 - 0x629  :   36 - 0x24
    "00100100", -- 1578 - 0x62a  :   36 - 0x24
    "00100100", -- 1579 - 0x62b  :   36 - 0x24
    "00100100", -- 1580 - 0x62c  :   36 - 0x24
    "00100100", -- 1581 - 0x62d  :   36 - 0x24
    "00100100", -- 1582 - 0x62e  :   36 - 0x24
    "00100100", -- 1583 - 0x62f  :   36 - 0x24
    "00100100", -- 1584 - 0x630  :   36 - 0x24
    "00100100", -- 1585 - 0x631  :   36 - 0x24
    "00100100", -- 1586 - 0x632  :   36 - 0x24
    "00100100", -- 1587 - 0x633  :   36 - 0x24
    "00100100", -- 1588 - 0x634  :   36 - 0x24
    "00100100", -- 1589 - 0x635  :   36 - 0x24
    "00100100", -- 1590 - 0x636  :   36 - 0x24
    "00100100", -- 1591 - 0x637  :   36 - 0x24
    "00100100", -- 1592 - 0x638  :   36 - 0x24
    "00100100", -- 1593 - 0x639  :   36 - 0x24
    "00100100", -- 1594 - 0x63a  :   36 - 0x24
    "00100100", -- 1595 - 0x63b  :   36 - 0x24
    "00100100", -- 1596 - 0x63c  :   36 - 0x24
    "00100100", -- 1597 - 0x63d  :   36 - 0x24
    "00100100", -- 1598 - 0x63e  :   36 - 0x24
    "00100100", -- 1599 - 0x63f  :   36 - 0x24
    "01010011", -- 1600 - 0x640  :   83 - 0x53
    "01010100", -- 1601 - 0x641  :   84 - 0x54
    "00100100", -- 1602 - 0x642  :   36 - 0x24
    "00100100", -- 1603 - 0x643  :   36 - 0x24
    "00100100", -- 1604 - 0x644  :   36 - 0x24
    "00100100", -- 1605 - 0x645  :   36 - 0x24
    "00100100", -- 1606 - 0x646  :   36 - 0x24
    "00100100", -- 1607 - 0x647  :   36 - 0x24
    "01000101", -- 1608 - 0x648  :   69 - 0x45
    "01000101", -- 1609 - 0x649  :   69 - 0x45
    "01010011", -- 1610 - 0x64a  :   83 - 0x53
    "01010100", -- 1611 - 0x64b  :   84 - 0x54
    "01000101", -- 1612 - 0x64c  :   69 - 0x45
    "01000101", -- 1613 - 0x64d  :   69 - 0x45
    "01010011", -- 1614 - 0x64e  :   83 - 0x53
    "01010100", -- 1615 - 0x64f  :   84 - 0x54
    "00100100", -- 1616 - 0x650  :   36 - 0x24
    "00100100", -- 1617 - 0x651  :   36 - 0x24
    "00100100", -- 1618 - 0x652  :   36 - 0x24
    "00100100", -- 1619 - 0x653  :   36 - 0x24
    "00100100", -- 1620 - 0x654  :   36 - 0x24
    "00100100", -- 1621 - 0x655  :   36 - 0x24
    "00100100", -- 1622 - 0x656  :   36 - 0x24
    "00100100", -- 1623 - 0x657  :   36 - 0x24
    "00100100", -- 1624 - 0x658  :   36 - 0x24
    "00100100", -- 1625 - 0x659  :   36 - 0x24
    "00100100", -- 1626 - 0x65a  :   36 - 0x24
    "00100100", -- 1627 - 0x65b  :   36 - 0x24
    "00100100", -- 1628 - 0x65c  :   36 - 0x24
    "00100100", -- 1629 - 0x65d  :   36 - 0x24
    "00100100", -- 1630 - 0x65e  :   36 - 0x24
    "00100100", -- 1631 - 0x65f  :   36 - 0x24
    "01010101", -- 1632 - 0x660  :   85 - 0x55
    "01010110", -- 1633 - 0x661  :   86 - 0x56
    "00100100", -- 1634 - 0x662  :   36 - 0x24
    "00100100", -- 1635 - 0x663  :   36 - 0x24
    "00100100", -- 1636 - 0x664  :   36 - 0x24
    "00100100", -- 1637 - 0x665  :   36 - 0x24
    "00100100", -- 1638 - 0x666  :   36 - 0x24
    "00100100", -- 1639 - 0x667  :   36 - 0x24
    "01000111", -- 1640 - 0x668  :   71 - 0x47
    "01000111", -- 1641 - 0x669  :   71 - 0x47
    "01010101", -- 1642 - 0x66a  :   85 - 0x55
    "01010110", -- 1643 - 0x66b  :   86 - 0x56
    "01000111", -- 1644 - 0x66c  :   71 - 0x47
    "01000111", -- 1645 - 0x66d  :   71 - 0x47
    "01010101", -- 1646 - 0x66e  :   85 - 0x55
    "01010110", -- 1647 - 0x66f  :   86 - 0x56
    "00100100", -- 1648 - 0x670  :   36 - 0x24
    "00100100", -- 1649 - 0x671  :   36 - 0x24
    "00100100", -- 1650 - 0x672  :   36 - 0x24
    "00100100", -- 1651 - 0x673  :   36 - 0x24
    "00100100", -- 1652 - 0x674  :   36 - 0x24
    "00100100", -- 1653 - 0x675  :   36 - 0x24
    "00100100", -- 1654 - 0x676  :   36 - 0x24
    "00100100", -- 1655 - 0x677  :   36 - 0x24
    "00100100", -- 1656 - 0x678  :   36 - 0x24
    "00100100", -- 1657 - 0x679  :   36 - 0x24
    "00100100", -- 1658 - 0x67a  :   36 - 0x24
    "00100100", -- 1659 - 0x67b  :   36 - 0x24
    "00100100", -- 1660 - 0x67c  :   36 - 0x24
    "00100100", -- 1661 - 0x67d  :   36 - 0x24
    "00100100", -- 1662 - 0x67e  :   36 - 0x24
    "00100100", -- 1663 - 0x67f  :   36 - 0x24
    "00100100", -- 1664 - 0x680  :   36 - 0x24
    "00100100", -- 1665 - 0x681  :   36 - 0x24
    "00100100", -- 1666 - 0x682  :   36 - 0x24
    "00100100", -- 1667 - 0x683  :   36 - 0x24
    "00100100", -- 1668 - 0x684  :   36 - 0x24
    "00100100", -- 1669 - 0x685  :   36 - 0x24
    "00100100", -- 1670 - 0x686  :   36 - 0x24
    "00100100", -- 1671 - 0x687  :   36 - 0x24
    "00100100", -- 1672 - 0x688  :   36 - 0x24
    "00100100", -- 1673 - 0x689  :   36 - 0x24
    "00100100", -- 1674 - 0x68a  :   36 - 0x24
    "00100100", -- 1675 - 0x68b  :   36 - 0x24
    "00100100", -- 1676 - 0x68c  :   36 - 0x24
    "00100100", -- 1677 - 0x68d  :   36 - 0x24
    "00100100", -- 1678 - 0x68e  :   36 - 0x24
    "00100100", -- 1679 - 0x68f  :   36 - 0x24
    "00100100", -- 1680 - 0x690  :   36 - 0x24
    "00100100", -- 1681 - 0x691  :   36 - 0x24
    "00100100", -- 1682 - 0x692  :   36 - 0x24
    "00100100", -- 1683 - 0x693  :   36 - 0x24
    "00100100", -- 1684 - 0x694  :   36 - 0x24
    "00100100", -- 1685 - 0x695  :   36 - 0x24
    "00100100", -- 1686 - 0x696  :   36 - 0x24
    "00100100", -- 1687 - 0x697  :   36 - 0x24
    "00100100", -- 1688 - 0x698  :   36 - 0x24
    "00100100", -- 1689 - 0x699  :   36 - 0x24
    "00100100", -- 1690 - 0x69a  :   36 - 0x24
    "00100100", -- 1691 - 0x69b  :   36 - 0x24
    "00100100", -- 1692 - 0x69c  :   36 - 0x24
    "00100100", -- 1693 - 0x69d  :   36 - 0x24
    "00100100", -- 1694 - 0x69e  :   36 - 0x24
    "00100100", -- 1695 - 0x69f  :   36 - 0x24
    "00100100", -- 1696 - 0x6a0  :   36 - 0x24
    "00100100", -- 1697 - 0x6a1  :   36 - 0x24
    "00100100", -- 1698 - 0x6a2  :   36 - 0x24
    "00100100", -- 1699 - 0x6a3  :   36 - 0x24
    "00100100", -- 1700 - 0x6a4  :   36 - 0x24
    "00100100", -- 1701 - 0x6a5  :   36 - 0x24
    "00100100", -- 1702 - 0x6a6  :   36 - 0x24
    "00100100", -- 1703 - 0x6a7  :   36 - 0x24
    "00100100", -- 1704 - 0x6a8  :   36 - 0x24
    "00100100", -- 1705 - 0x6a9  :   36 - 0x24
    "00100100", -- 1706 - 0x6aa  :   36 - 0x24
    "00100100", -- 1707 - 0x6ab  :   36 - 0x24
    "00100100", -- 1708 - 0x6ac  :   36 - 0x24
    "00100100", -- 1709 - 0x6ad  :   36 - 0x24
    "00100100", -- 1710 - 0x6ae  :   36 - 0x24
    "00100100", -- 1711 - 0x6af  :   36 - 0x24
    "00100100", -- 1712 - 0x6b0  :   36 - 0x24
    "00100100", -- 1713 - 0x6b1  :   36 - 0x24
    "00100100", -- 1714 - 0x6b2  :   36 - 0x24
    "00100100", -- 1715 - 0x6b3  :   36 - 0x24
    "00100100", -- 1716 - 0x6b4  :   36 - 0x24
    "00100100", -- 1717 - 0x6b5  :   36 - 0x24
    "00100100", -- 1718 - 0x6b6  :   36 - 0x24
    "00100100", -- 1719 - 0x6b7  :   36 - 0x24
    "00100100", -- 1720 - 0x6b8  :   36 - 0x24
    "00100100", -- 1721 - 0x6b9  :   36 - 0x24
    "00100100", -- 1722 - 0x6ba  :   36 - 0x24
    "00100100", -- 1723 - 0x6bb  :   36 - 0x24
    "00100100", -- 1724 - 0x6bc  :   36 - 0x24
    "00100100", -- 1725 - 0x6bd  :   36 - 0x24
    "00100100", -- 1726 - 0x6be  :   36 - 0x24
    "00100100", -- 1727 - 0x6bf  :   36 - 0x24
    "00100100", -- 1728 - 0x6c0  :   36 - 0x24
    "00100100", -- 1729 - 0x6c1  :   36 - 0x24
    "00100100", -- 1730 - 0x6c2  :   36 - 0x24
    "00100100", -- 1731 - 0x6c3  :   36 - 0x24
    "00100100", -- 1732 - 0x6c4  :   36 - 0x24
    "00100100", -- 1733 - 0x6c5  :   36 - 0x24
    "00100100", -- 1734 - 0x6c6  :   36 - 0x24
    "00100100", -- 1735 - 0x6c7  :   36 - 0x24
    "00100100", -- 1736 - 0x6c8  :   36 - 0x24
    "00100100", -- 1737 - 0x6c9  :   36 - 0x24
    "00100100", -- 1738 - 0x6ca  :   36 - 0x24
    "00100100", -- 1739 - 0x6cb  :   36 - 0x24
    "00100100", -- 1740 - 0x6cc  :   36 - 0x24
    "00100100", -- 1741 - 0x6cd  :   36 - 0x24
    "00100100", -- 1742 - 0x6ce  :   36 - 0x24
    "00100100", -- 1743 - 0x6cf  :   36 - 0x24
    "00100100", -- 1744 - 0x6d0  :   36 - 0x24
    "00100100", -- 1745 - 0x6d1  :   36 - 0x24
    "00100100", -- 1746 - 0x6d2  :   36 - 0x24
    "00100100", -- 1747 - 0x6d3  :   36 - 0x24
    "00100100", -- 1748 - 0x6d4  :   36 - 0x24
    "00100100", -- 1749 - 0x6d5  :   36 - 0x24
    "00100100", -- 1750 - 0x6d6  :   36 - 0x24
    "00100100", -- 1751 - 0x6d7  :   36 - 0x24
    "00100100", -- 1752 - 0x6d8  :   36 - 0x24
    "00100100", -- 1753 - 0x6d9  :   36 - 0x24
    "00100100", -- 1754 - 0x6da  :   36 - 0x24
    "00100100", -- 1755 - 0x6db  :   36 - 0x24
    "00100100", -- 1756 - 0x6dc  :   36 - 0x24
    "00100100", -- 1757 - 0x6dd  :   36 - 0x24
    "00100100", -- 1758 - 0x6de  :   36 - 0x24
    "00100100", -- 1759 - 0x6df  :   36 - 0x24
    "00100100", -- 1760 - 0x6e0  :   36 - 0x24
    "00100100", -- 1761 - 0x6e1  :   36 - 0x24
    "00110001", -- 1762 - 0x6e2  :   49 - 0x31
    "00110010", -- 1763 - 0x6e3  :   50 - 0x32
    "00100100", -- 1764 - 0x6e4  :   36 - 0x24
    "00100100", -- 1765 - 0x6e5  :   36 - 0x24
    "00100100", -- 1766 - 0x6e6  :   36 - 0x24
    "00100100", -- 1767 - 0x6e7  :   36 - 0x24
    "00100100", -- 1768 - 0x6e8  :   36 - 0x24
    "00100100", -- 1769 - 0x6e9  :   36 - 0x24
    "00100100", -- 1770 - 0x6ea  :   36 - 0x24
    "00100100", -- 1771 - 0x6eb  :   36 - 0x24
    "00100100", -- 1772 - 0x6ec  :   36 - 0x24
    "00100100", -- 1773 - 0x6ed  :   36 - 0x24
    "00100100", -- 1774 - 0x6ee  :   36 - 0x24
    "00100100", -- 1775 - 0x6ef  :   36 - 0x24
    "00100100", -- 1776 - 0x6f0  :   36 - 0x24
    "00100100", -- 1777 - 0x6f1  :   36 - 0x24
    "00100100", -- 1778 - 0x6f2  :   36 - 0x24
    "00100100", -- 1779 - 0x6f3  :   36 - 0x24
    "00100100", -- 1780 - 0x6f4  :   36 - 0x24
    "00100100", -- 1781 - 0x6f5  :   36 - 0x24
    "00100100", -- 1782 - 0x6f6  :   36 - 0x24
    "00100100", -- 1783 - 0x6f7  :   36 - 0x24
    "00100100", -- 1784 - 0x6f8  :   36 - 0x24
    "00100100", -- 1785 - 0x6f9  :   36 - 0x24
    "00100100", -- 1786 - 0x6fa  :   36 - 0x24
    "00100100", -- 1787 - 0x6fb  :   36 - 0x24
    "00100100", -- 1788 - 0x6fc  :   36 - 0x24
    "00100100", -- 1789 - 0x6fd  :   36 - 0x24
    "00100100", -- 1790 - 0x6fe  :   36 - 0x24
    "00100100", -- 1791 - 0x6ff  :   36 - 0x24
    "00100100", -- 1792 - 0x700  :   36 - 0x24
    "00110000", -- 1793 - 0x701  :   48 - 0x30
    "00100110", -- 1794 - 0x702  :   38 - 0x26
    "00110100", -- 1795 - 0x703  :   52 - 0x34
    "00110011", -- 1796 - 0x704  :   51 - 0x33
    "00100100", -- 1797 - 0x705  :   36 - 0x24
    "00100100", -- 1798 - 0x706  :   36 - 0x24
    "00100100", -- 1799 - 0x707  :   36 - 0x24
    "00100100", -- 1800 - 0x708  :   36 - 0x24
    "00100100", -- 1801 - 0x709  :   36 - 0x24
    "00100100", -- 1802 - 0x70a  :   36 - 0x24
    "00100100", -- 1803 - 0x70b  :   36 - 0x24
    "00100100", -- 1804 - 0x70c  :   36 - 0x24
    "00100100", -- 1805 - 0x70d  :   36 - 0x24
    "00100100", -- 1806 - 0x70e  :   36 - 0x24
    "00100100", -- 1807 - 0x70f  :   36 - 0x24
    "00100100", -- 1808 - 0x710  :   36 - 0x24
    "00100100", -- 1809 - 0x711  :   36 - 0x24
    "00100100", -- 1810 - 0x712  :   36 - 0x24
    "00100100", -- 1811 - 0x713  :   36 - 0x24
    "00100100", -- 1812 - 0x714  :   36 - 0x24
    "00100100", -- 1813 - 0x715  :   36 - 0x24
    "00100100", -- 1814 - 0x716  :   36 - 0x24
    "00100100", -- 1815 - 0x717  :   36 - 0x24
    "00100100", -- 1816 - 0x718  :   36 - 0x24
    "00100100", -- 1817 - 0x719  :   36 - 0x24
    "00100100", -- 1818 - 0x71a  :   36 - 0x24
    "00100100", -- 1819 - 0x71b  :   36 - 0x24
    "00100100", -- 1820 - 0x71c  :   36 - 0x24
    "00100100", -- 1821 - 0x71d  :   36 - 0x24
    "00100100", -- 1822 - 0x71e  :   36 - 0x24
    "00100100", -- 1823 - 0x71f  :   36 - 0x24
    "00110000", -- 1824 - 0x720  :   48 - 0x30
    "00100110", -- 1825 - 0x721  :   38 - 0x26
    "00100110", -- 1826 - 0x722  :   38 - 0x26
    "00100110", -- 1827 - 0x723  :   38 - 0x26
    "00100110", -- 1828 - 0x724  :   38 - 0x26
    "00110011", -- 1829 - 0x725  :   51 - 0x33
    "00100100", -- 1830 - 0x726  :   36 - 0x24
    "00100100", -- 1831 - 0x727  :   36 - 0x24
    "00100100", -- 1832 - 0x728  :   36 - 0x24
    "00100100", -- 1833 - 0x729  :   36 - 0x24
    "00100100", -- 1834 - 0x72a  :   36 - 0x24
    "00100100", -- 1835 - 0x72b  :   36 - 0x24
    "00100100", -- 1836 - 0x72c  :   36 - 0x24
    "00100100", -- 1837 - 0x72d  :   36 - 0x24
    "00100100", -- 1838 - 0x72e  :   36 - 0x24
    "00110101", -- 1839 - 0x72f  :   53 - 0x35
    "00100100", -- 1840 - 0x730  :   36 - 0x24
    "00100100", -- 1841 - 0x731  :   36 - 0x24
    "00100100", -- 1842 - 0x732  :   36 - 0x24
    "00100100", -- 1843 - 0x733  :   36 - 0x24
    "00100100", -- 1844 - 0x734  :   36 - 0x24
    "00100100", -- 1845 - 0x735  :   36 - 0x24
    "00100100", -- 1846 - 0x736  :   36 - 0x24
    "00100100", -- 1847 - 0x737  :   36 - 0x24
    "00100100", -- 1848 - 0x738  :   36 - 0x24
    "00100100", -- 1849 - 0x739  :   36 - 0x24
    "00100100", -- 1850 - 0x73a  :   36 - 0x24
    "00100100", -- 1851 - 0x73b  :   36 - 0x24
    "00100100", -- 1852 - 0x73c  :   36 - 0x24
    "00100100", -- 1853 - 0x73d  :   36 - 0x24
    "00100100", -- 1854 - 0x73e  :   36 - 0x24
    "00100100", -- 1855 - 0x73f  :   36 - 0x24
    "10110100", -- 1856 - 0x740  :  180 - 0xb4
    "10110101", -- 1857 - 0x741  :  181 - 0xb5
    "10110100", -- 1858 - 0x742  :  180 - 0xb4
    "10110101", -- 1859 - 0x743  :  181 - 0xb5
    "10110100", -- 1860 - 0x744  :  180 - 0xb4
    "10110101", -- 1861 - 0x745  :  181 - 0xb5
    "10110100", -- 1862 - 0x746  :  180 - 0xb4
    "10110101", -- 1863 - 0x747  :  181 - 0xb5
    "10110100", -- 1864 - 0x748  :  180 - 0xb4
    "10110101", -- 1865 - 0x749  :  181 - 0xb5
    "10110100", -- 1866 - 0x74a  :  180 - 0xb4
    "10110101", -- 1867 - 0x74b  :  181 - 0xb5
    "10110100", -- 1868 - 0x74c  :  180 - 0xb4
    "10110101", -- 1869 - 0x74d  :  181 - 0xb5
    "10110100", -- 1870 - 0x74e  :  180 - 0xb4
    "10110101", -- 1871 - 0x74f  :  181 - 0xb5
    "00100100", -- 1872 - 0x750  :   36 - 0x24
    "00100100", -- 1873 - 0x751  :   36 - 0x24
    "00100100", -- 1874 - 0x752  :   36 - 0x24
    "00100100", -- 1875 - 0x753  :   36 - 0x24
    "00100100", -- 1876 - 0x754  :   36 - 0x24
    "00100100", -- 1877 - 0x755  :   36 - 0x24
    "00100100", -- 1878 - 0x756  :   36 - 0x24
    "00100100", -- 1879 - 0x757  :   36 - 0x24
    "00100100", -- 1880 - 0x758  :   36 - 0x24
    "00100100", -- 1881 - 0x759  :   36 - 0x24
    "00100100", -- 1882 - 0x75a  :   36 - 0x24
    "00100100", -- 1883 - 0x75b  :   36 - 0x24
    "00100100", -- 1884 - 0x75c  :   36 - 0x24
    "00100100", -- 1885 - 0x75d  :   36 - 0x24
    "00100100", -- 1886 - 0x75e  :   36 - 0x24
    "00100100", -- 1887 - 0x75f  :   36 - 0x24
    "10110110", -- 1888 - 0x760  :  182 - 0xb6
    "10110111", -- 1889 - 0x761  :  183 - 0xb7
    "10110110", -- 1890 - 0x762  :  182 - 0xb6
    "10110111", -- 1891 - 0x763  :  183 - 0xb7
    "10110110", -- 1892 - 0x764  :  182 - 0xb6
    "10110111", -- 1893 - 0x765  :  183 - 0xb7
    "10110110", -- 1894 - 0x766  :  182 - 0xb6
    "10110111", -- 1895 - 0x767  :  183 - 0xb7
    "10110110", -- 1896 - 0x768  :  182 - 0xb6
    "10110111", -- 1897 - 0x769  :  183 - 0xb7
    "10110110", -- 1898 - 0x76a  :  182 - 0xb6
    "10110111", -- 1899 - 0x76b  :  183 - 0xb7
    "10110110", -- 1900 - 0x76c  :  182 - 0xb6
    "10110111", -- 1901 - 0x76d  :  183 - 0xb7
    "10110110", -- 1902 - 0x76e  :  182 - 0xb6
    "10110111", -- 1903 - 0x76f  :  183 - 0xb7
    "00100100", -- 1904 - 0x770  :   36 - 0x24
    "00100100", -- 1905 - 0x771  :   36 - 0x24
    "00100100", -- 1906 - 0x772  :   36 - 0x24
    "00100100", -- 1907 - 0x773  :   36 - 0x24
    "00100100", -- 1908 - 0x774  :   36 - 0x24
    "00100100", -- 1909 - 0x775  :   36 - 0x24
    "00100100", -- 1910 - 0x776  :   36 - 0x24
    "00100100", -- 1911 - 0x777  :   36 - 0x24
    "00100100", -- 1912 - 0x778  :   36 - 0x24
    "00100100", -- 1913 - 0x779  :   36 - 0x24
    "00100100", -- 1914 - 0x77a  :   36 - 0x24
    "00100100", -- 1915 - 0x77b  :   36 - 0x24
    "00100100", -- 1916 - 0x77c  :   36 - 0x24
    "00100100", -- 1917 - 0x77d  :   36 - 0x24
    "00100100", -- 1918 - 0x77e  :   36 - 0x24
    "00100100", -- 1919 - 0x77f  :   36 - 0x24
    "10110100", -- 1920 - 0x780  :  180 - 0xb4
    "10110101", -- 1921 - 0x781  :  181 - 0xb5
    "10110100", -- 1922 - 0x782  :  180 - 0xb4
    "10110101", -- 1923 - 0x783  :  181 - 0xb5
    "10110100", -- 1924 - 0x784  :  180 - 0xb4
    "10110101", -- 1925 - 0x785  :  181 - 0xb5
    "10110100", -- 1926 - 0x786  :  180 - 0xb4
    "10110101", -- 1927 - 0x787  :  181 - 0xb5
    "10110100", -- 1928 - 0x788  :  180 - 0xb4
    "10110101", -- 1929 - 0x789  :  181 - 0xb5
    "10110100", -- 1930 - 0x78a  :  180 - 0xb4
    "10110101", -- 1931 - 0x78b  :  181 - 0xb5
    "10110100", -- 1932 - 0x78c  :  180 - 0xb4
    "10110101", -- 1933 - 0x78d  :  181 - 0xb5
    "10110100", -- 1934 - 0x78e  :  180 - 0xb4
    "10110101", -- 1935 - 0x78f  :  181 - 0xb5
    "00100100", -- 1936 - 0x790  :   36 - 0x24
    "00100100", -- 1937 - 0x791  :   36 - 0x24
    "00100100", -- 1938 - 0x792  :   36 - 0x24
    "00100100", -- 1939 - 0x793  :   36 - 0x24
    "00100100", -- 1940 - 0x794  :   36 - 0x24
    "00100100", -- 1941 - 0x795  :   36 - 0x24
    "00100100", -- 1942 - 0x796  :   36 - 0x24
    "00100100", -- 1943 - 0x797  :   36 - 0x24
    "00100100", -- 1944 - 0x798  :   36 - 0x24
    "00100100", -- 1945 - 0x799  :   36 - 0x24
    "00100100", -- 1946 - 0x79a  :   36 - 0x24
    "00100100", -- 1947 - 0x79b  :   36 - 0x24
    "00100100", -- 1948 - 0x79c  :   36 - 0x24
    "00100100", -- 1949 - 0x79d  :   36 - 0x24
    "00100100", -- 1950 - 0x79e  :   36 - 0x24
    "00100100", -- 1951 - 0x79f  :   36 - 0x24
    "10110110", -- 1952 - 0x7a0  :  182 - 0xb6
    "10110111", -- 1953 - 0x7a1  :  183 - 0xb7
    "10110110", -- 1954 - 0x7a2  :  182 - 0xb6
    "10110111", -- 1955 - 0x7a3  :  183 - 0xb7
    "10110110", -- 1956 - 0x7a4  :  182 - 0xb6
    "10110111", -- 1957 - 0x7a5  :  183 - 0xb7
    "10110110", -- 1958 - 0x7a6  :  182 - 0xb6
    "10110111", -- 1959 - 0x7a7  :  183 - 0xb7
    "10110110", -- 1960 - 0x7a8  :  182 - 0xb6
    "10110111", -- 1961 - 0x7a9  :  183 - 0xb7
    "10110110", -- 1962 - 0x7aa  :  182 - 0xb6
    "10110111", -- 1963 - 0x7ab  :  183 - 0xb7
    "10110110", -- 1964 - 0x7ac  :  182 - 0xb6
    "10110111", -- 1965 - 0x7ad  :  183 - 0xb7
    "10110110", -- 1966 - 0x7ae  :  182 - 0xb6
    "10110111", -- 1967 - 0x7af  :  183 - 0xb7
    "00100100", -- 1968 - 0x7b0  :   36 - 0x24
    "00100100", -- 1969 - 0x7b1  :   36 - 0x24
    "00100100", -- 1970 - 0x7b2  :   36 - 0x24
    "00100100", -- 1971 - 0x7b3  :   36 - 0x24
    "00100100", -- 1972 - 0x7b4  :   36 - 0x24
    "00100100", -- 1973 - 0x7b5  :   36 - 0x24
    "00100100", -- 1974 - 0x7b6  :   36 - 0x24
    "00100100", -- 1975 - 0x7b7  :   36 - 0x24
    "00100100", -- 1976 - 0x7b8  :   36 - 0x24
    "00100100", -- 1977 - 0x7b9  :   36 - 0x24
    "00100100", -- 1978 - 0x7ba  :   36 - 0x24
    "00100100", -- 1979 - 0x7bb  :   36 - 0x24
    "00100100", -- 1980 - 0x7bc  :   36 - 0x24
    "00100100", -- 1981 - 0x7bd  :   36 - 0x24
    "00100100", -- 1982 - 0x7be  :   36 - 0x24
    "00100100", -- 1983 - 0x7bf  :   36 - 0x24
        ---- Attribute Table 1----
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0
    "10001000", -- 1993 - 0x7c9  :  136 - 0x88
    "10101010", -- 1994 - 0x7ca  :  170 - 0xaa
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00110000", -- 2003 - 0x7d3  :   48 - 0x30
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00110000", -- 2016 - 0x7e0  :   48 - 0x30
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "11010000", -- 2018 - 0x7e2  :  208 - 0xd0
    "11010000", -- 2019 - 0x7e3  :  208 - 0xd0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "01010000", -- 2032 - 0x7f0  :   80 - 0x50
    "01010000", -- 2033 - 0x7f1  :   80 - 0x50
    "01010000", -- 2034 - 0x7f2  :   80 - 0x50
    "01010000", -- 2035 - 0x7f3  :   80 - 0x50
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000101", -- 2040 - 0x7f8  :    5 - 0x5
    "00000101", -- 2041 - 0x7f9  :    5 - 0x5
    "00000101", -- 2042 - 0x7fa  :    5 - 0x5
    "00000101", -- 2043 - 0x7fb  :    5 - 0x5
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
