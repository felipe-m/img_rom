//- Autcmatically generated verilog ROM from a NES memory file----
//-   ATTRIBUTE TABLE SEPARATED FROM NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_attribute_tables


//-  Original memory dump file name: nova_ntable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_ATABLE_NOVA_00
  (
     //input     clk,   // clock
     input      [7-1:0] addr,  //128 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
      7'h0: dout  = 8'b00000000; //    0 :   0 - 0x0
      7'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      7'h2: dout  = 8'b00000000; //    2 :   0 - 0x0
      7'h3: dout  = 8'b00000000; //    3 :   0 - 0x0
      7'h4: dout  = 8'b00000000; //    4 :   0 - 0x0
      7'h5: dout  = 8'b00000000; //    5 :   0 - 0x0
      7'h6: dout  = 8'b00000000; //    6 :   0 - 0x0
      7'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      7'h8: dout  = 8'b00000000; //    8 :   0 - 0x0
      7'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      7'hA: dout  = 8'b00000000; //   10 :   0 - 0x0
      7'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      7'hC: dout  = 8'b00000000; //   12 :   0 - 0x0
      7'hD: dout  = 8'b00000000; //   13 :   0 - 0x0
      7'hE: dout  = 8'b00001000; //   14 :   8 - 0x8
      7'hF: dout  = 8'b00001000; //   15 :   8 - 0x8
      7'h10: dout  = 8'b00000000; //   16 :   0 - 0x0
      7'h11: dout  = 8'b00000000; //   17 :   0 - 0x0
      7'h12: dout  = 8'b00000000; //   18 :   0 - 0x0
      7'h13: dout  = 8'b00000000; //   19 :   0 - 0x0
      7'h14: dout  = 8'b00000000; //   20 :   0 - 0x0
      7'h15: dout  = 8'b01010001; //   21 :  81 - 0x51
      7'h16: dout  = 8'b01010000; //   22 :  80 - 0x50
      7'h17: dout  = 8'b01010000; //   23 :  80 - 0x50
      7'h18: dout  = 8'b00000000; //   24 :   0 - 0x0
      7'h19: dout  = 8'b00000000; //   25 :   0 - 0x0
      7'h1A: dout  = 8'b00000000; //   26 :   0 - 0x0
      7'h1B: dout  = 8'b00000000; //   27 :   0 - 0x0
      7'h1C: dout  = 8'b00000000; //   28 :   0 - 0x0
      7'h1D: dout  = 8'b00000000; //   29 :   0 - 0x0
      7'h1E: dout  = 8'b00000000; //   30 :   0 - 0x0
      7'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      7'h20: dout  = 8'b00000000; //   32 :   0 - 0x0
      7'h21: dout  = 8'b00000000; //   33 :   0 - 0x0
      7'h22: dout  = 8'b00000000; //   34 :   0 - 0x0
      7'h23: dout  = 8'b00000000; //   35 :   0 - 0x0
      7'h24: dout  = 8'b10100000; //   36 : 160 - 0xa0
      7'h25: dout  = 8'b10100000; //   37 : 160 - 0xa0
      7'h26: dout  = 8'b10100000; //   38 : 160 - 0xa0
      7'h27: dout  = 8'b10100000; //   39 : 160 - 0xa0
      7'h28: dout  = 8'b00000000; //   40 :   0 - 0x0
      7'h29: dout  = 8'b00000000; //   41 :   0 - 0x0
      7'h2A: dout  = 8'b00000000; //   42 :   0 - 0x0
      7'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      7'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      7'h2D: dout  = 8'b00000000; //   45 :   0 - 0x0
      7'h2E: dout  = 8'b00000000; //   46 :   0 - 0x0
      7'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      7'h30: dout  = 8'b00000000; //   48 :   0 - 0x0
      7'h31: dout  = 8'b00000010; //   49 :   2 - 0x2
      7'h32: dout  = 8'b00000000; //   50 :   0 - 0x0
      7'h33: dout  = 8'b00000000; //   51 :   0 - 0x0
      7'h34: dout  = 8'b00000000; //   52 :   0 - 0x0
      7'h35: dout  = 8'b00000000; //   53 :   0 - 0x0
      7'h36: dout  = 8'b00000000; //   54 :   0 - 0x0
      7'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      7'h38: dout  = 8'b00000000; //   56 :   0 - 0x0
      7'h39: dout  = 8'b00000000; //   57 :   0 - 0x0
      7'h3A: dout  = 8'b00000000; //   58 :   0 - 0x0
      7'h3B: dout  = 8'b00000000; //   59 :   0 - 0x0
      7'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      7'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      7'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      7'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      7'h40: dout  = 8'b00000000; //   64 :   0 - 0x0
      7'h41: dout  = 8'b00000000; //   65 :   0 - 0x0
      7'h42: dout  = 8'b10001000; //   66 : 136 - 0x88
      7'h43: dout  = 8'b00010001; //   67 :  17 - 0x11
      7'h44: dout  = 8'b00000000; //   68 :   0 - 0x0
      7'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      7'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      7'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      7'h48: dout  = 8'b00001010; //   72 :  10 - 0xa
      7'h49: dout  = 8'b00000010; //   73 :   2 - 0x2
      7'h4A: dout  = 8'b10001000; //   74 : 136 - 0x88
      7'h4B: dout  = 8'b00010001; //   75 :  17 - 0x11
      7'h4C: dout  = 8'b00000000; //   76 :   0 - 0x0
      7'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      7'h4E: dout  = 8'b00000000; //   78 :   0 - 0x0
      7'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      7'h50: dout  = 8'b01010100; //   80 :  84 - 0x54
      7'h51: dout  = 8'b00000101; //   81 :   5 - 0x5
      7'h52: dout  = 8'b00000101; //   82 :   5 - 0x5
      7'h53: dout  = 8'b00000001; //   83 :   1 - 0x1
      7'h54: dout  = 8'b00000000; //   84 :   0 - 0x0
      7'h55: dout  = 8'b00000000; //   85 :   0 - 0x0
      7'h56: dout  = 8'b10000000; //   86 : 128 - 0x80
      7'h57: dout  = 8'b10100000; //   87 : 160 - 0xa0
      7'h58: dout  = 8'b00000000; //   88 :   0 - 0x0
      7'h59: dout  = 8'b00000000; //   89 :   0 - 0x0
      7'h5A: dout  = 8'b00000000; //   90 :   0 - 0x0
      7'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      7'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      7'h5D: dout  = 8'b00000000; //   93 :   0 - 0x0
      7'h5E: dout  = 8'b01010000; //   94 :  80 - 0x50
      7'h5F: dout  = 8'b01010000; //   95 :  80 - 0x50
      7'h60: dout  = 8'b00000000; //   96 :   0 - 0x0
      7'h61: dout  = 8'b00000000; //   97 :   0 - 0x0
      7'h62: dout  = 8'b00000000; //   98 :   0 - 0x0
      7'h63: dout  = 8'b00000000; //   99 :   0 - 0x0
      7'h64: dout  = 8'b10000000; //  100 : 128 - 0x80
      7'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      7'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      7'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      7'h68: dout  = 8'b00000000; //  104 :   0 - 0x0
      7'h69: dout  = 8'b00000000; //  105 :   0 - 0x0
      7'h6A: dout  = 8'b00000000; //  106 :   0 - 0x0
      7'h6B: dout  = 8'b00000000; //  107 :   0 - 0x0
      7'h6C: dout  = 8'b00000000; //  108 :   0 - 0x0
      7'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      7'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      7'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      7'h70: dout  = 8'b00000000; //  112 :   0 - 0x0
      7'h71: dout  = 8'b00000000; //  113 :   0 - 0x0
      7'h72: dout  = 8'b00000010; //  114 :   2 - 0x2
      7'h73: dout  = 8'b00000000; //  115 :   0 - 0x0
      7'h74: dout  = 8'b00000000; //  116 :   0 - 0x0
      7'h75: dout  = 8'b00000000; //  117 :   0 - 0x0
      7'h76: dout  = 8'b00000000; //  118 :   0 - 0x0
      7'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      7'h78: dout  = 8'b00000000; //  120 :   0 - 0x0
      7'h79: dout  = 8'b00000000; //  121 :   0 - 0x0
      7'h7A: dout  = 8'b00000000; //  122 :   0 - 0x0
      7'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      7'h7C: dout  = 8'b00000000; //  124 :   0 - 0x0
      7'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      7'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      7'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
    endcase
  end

endmodule
