--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE WITH ONLY ONE COLOR PLANE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: donkeykong_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_DONKEYKONG_color0 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_DONKEYKONG_color0;

architecture BEHAVIORAL of ROM_PTABLE_DONKEYKONG_color0 is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000011", --    1 -  0x1  :    3 - 0x3
    "00000111", --    2 -  0x2  :    7 - 0x7
    "00000111", --    3 -  0x3  :    7 - 0x7
    "00001001", --    4 -  0x4  :    9 - 0x9
    "00001001", --    5 -  0x5  :    9 - 0x9
    "00011100", --    6 -  0x6  :   28 - 0x1c
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00001111", --    8 -  0x8  :   15 - 0xf -- Sprite 0x1
    "00001111", --    9 -  0x9  :   15 - 0xf
    "00001111", --   10 -  0xa  :   15 - 0xf
    "11111111", --   11 -  0xb  :  255 - 0xff
    "11111111", --   12 -  0xc  :  255 - 0xff
    "11111100", --   13 -  0xd  :  252 - 0xfc
    "10000001", --   14 -  0xe  :  129 - 0x81
    "00000001", --   15 -  0xf  :    1 - 0x1
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Sprite 0x2
    "11000000", --   17 - 0x11  :  192 - 0xc0
    "11111000", --   18 - 0x12  :  248 - 0xf8
    "10000000", --   19 - 0x13  :  128 - 0x80
    "00100000", --   20 - 0x14  :   32 - 0x20
    "10010000", --   21 - 0x15  :  144 - 0x90
    "00111100", --   22 - 0x16  :   60 - 0x3c
    "00000000", --   23 - 0x17  :    0 - 0x0
    "11000000", --   24 - 0x18  :  192 - 0xc0 -- Sprite 0x3
    "11000000", --   25 - 0x19  :  192 - 0xc0
    "11000000", --   26 - 0x1a  :  192 - 0xc0
    "11110000", --   27 - 0x1b  :  240 - 0xf0
    "11110000", --   28 - 0x1c  :  240 - 0xf0
    "11100000", --   29 - 0x1d  :  224 - 0xe0
    "11000000", --   30 - 0x1e  :  192 - 0xc0
    "11100000", --   31 - 0x1f  :  224 - 0xe0
    "00000111", --   32 - 0x20  :    7 - 0x7 -- Sprite 0x4
    "00001111", --   33 - 0x21  :   15 - 0xf
    "00001111", --   34 - 0x22  :   15 - 0xf
    "00010010", --   35 - 0x23  :   18 - 0x12
    "00010011", --   36 - 0x24  :   19 - 0x13
    "00111000", --   37 - 0x25  :   56 - 0x38
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00001111", --   39 - 0x27  :   15 - 0xf
    "00011111", --   40 - 0x28  :   31 - 0x1f -- Sprite 0x5
    "00011111", --   41 - 0x29  :   31 - 0x1f
    "00011111", --   42 - 0x2a  :   31 - 0x1f
    "00011000", --   43 - 0x2b  :   24 - 0x18
    "00011001", --   44 - 0x2c  :   25 - 0x19
    "00011110", --   45 - 0x2d  :   30 - 0x1e
    "00011100", --   46 - 0x2e  :   28 - 0x1c
    "00011110", --   47 - 0x2f  :   30 - 0x1e
    "10000000", --   48 - 0x30  :  128 - 0x80 -- Sprite 0x6
    "11110000", --   49 - 0x31  :  240 - 0xf0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "01000000", --   51 - 0x33  :   64 - 0x40
    "00100000", --   52 - 0x34  :   32 - 0x20
    "01111000", --   53 - 0x35  :  120 - 0x78
    "00000000", --   54 - 0x36  :    0 - 0x0
    "11000000", --   55 - 0x37  :  192 - 0xc0
    "11100000", --   56 - 0x38  :  224 - 0xe0 -- Sprite 0x7
    "01100000", --   57 - 0x39  :   96 - 0x60
    "11110000", --   58 - 0x3a  :  240 - 0xf0
    "11110000", --   59 - 0x3b  :  240 - 0xf0
    "11110000", --   60 - 0x3c  :  240 - 0xf0
    "11100000", --   61 - 0x3d  :  224 - 0xe0
    "11100000", --   62 - 0x3e  :  224 - 0xe0
    "11110000", --   63 - 0x3f  :  240 - 0xf0
    "00000111", --   64 - 0x40  :    7 - 0x7 -- Sprite 0x8
    "00001111", --   65 - 0x41  :   15 - 0xf
    "00001111", --   66 - 0x42  :   15 - 0xf
    "00010010", --   67 - 0x43  :   18 - 0x12
    "00010011", --   68 - 0x44  :   19 - 0x13
    "00111000", --   69 - 0x45  :   56 - 0x38
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00111111", --   71 - 0x47  :   63 - 0x3f
    "00111111", --   72 - 0x48  :   63 - 0x3f -- Sprite 0x9
    "00001110", --   73 - 0x49  :   14 - 0xe
    "00001111", --   74 - 0x4a  :   15 - 0xf
    "00011111", --   75 - 0x4b  :   31 - 0x1f
    "00111111", --   76 - 0x4c  :   63 - 0x3f
    "01111100", --   77 - 0x4d  :  124 - 0x7c
    "01110000", --   78 - 0x4e  :  112 - 0x70
    "00111000", --   79 - 0x4f  :   56 - 0x38
    "10000000", --   80 - 0x50  :  128 - 0x80 -- Sprite 0xa
    "11110000", --   81 - 0x51  :  240 - 0xf0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "01000000", --   83 - 0x53  :   64 - 0x40
    "00100000", --   84 - 0x54  :   32 - 0x20
    "01111000", --   85 - 0x55  :  120 - 0x78
    "00000000", --   86 - 0x56  :    0 - 0x0
    "11000000", --   87 - 0x57  :  192 - 0xc0
    "11110000", --   88 - 0x58  :  240 - 0xf0 -- Sprite 0xb
    "11111000", --   89 - 0x59  :  248 - 0xf8
    "11100100", --   90 - 0x5a  :  228 - 0xe4
    "11111100", --   91 - 0x5b  :  252 - 0xfc
    "11111100", --   92 - 0x5c  :  252 - 0xfc
    "01111100", --   93 - 0x5d  :  124 - 0x7c
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Sprite 0xc
    "00000010", --   97 - 0x61  :    2 - 0x2
    "00000110", --   98 - 0x62  :    6 - 0x6
    "00000111", --   99 - 0x63  :    7 - 0x7
    "00001001", --  100 - 0x64  :    9 - 0x9
    "00001001", --  101 - 0x65  :    9 - 0x9
    "00011101", --  102 - 0x66  :   29 - 0x1d
    "00000011", --  103 - 0x67  :    3 - 0x3
    "00001111", --  104 - 0x68  :   15 - 0xf -- Sprite 0xd
    "00001111", --  105 - 0x69  :   15 - 0xf
    "00001111", --  106 - 0x6a  :   15 - 0xf
    "11111111", --  107 - 0x6b  :  255 - 0xff
    "11111111", --  108 - 0x6c  :  255 - 0xff
    "11111100", --  109 - 0x6d  :  252 - 0xfc
    "10000001", --  110 - 0x6e  :  129 - 0x81
    "00000001", --  111 - 0x6f  :    1 - 0x1
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Sprite 0xe
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00111000", --  114 - 0x72  :   56 - 0x38
    "11000000", --  115 - 0x73  :  192 - 0xc0
    "11100000", --  116 - 0x74  :  224 - 0xe0
    "11010000", --  117 - 0x75  :  208 - 0xd0
    "11111100", --  118 - 0x76  :  252 - 0xfc
    "11000000", --  119 - 0x77  :  192 - 0xc0
    "11100000", --  120 - 0x78  :  224 - 0xe0 -- Sprite 0xf
    "11100000", --  121 - 0x79  :  224 - 0xe0
    "10110000", --  122 - 0x7a  :  176 - 0xb0
    "11110000", --  123 - 0x7b  :  240 - 0xf0
    "11110000", --  124 - 0x7c  :  240 - 0xf0
    "11100000", --  125 - 0x7d  :  224 - 0xe0
    "11000000", --  126 - 0x7e  :  192 - 0xc0
    "11100000", --  127 - 0x7f  :  224 - 0xe0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x10
    "00000011", --  129 - 0x81  :    3 - 0x3
    "00000111", --  130 - 0x82  :    7 - 0x7
    "00000111", --  131 - 0x83  :    7 - 0x7
    "00001001", --  132 - 0x84  :    9 - 0x9
    "00001001", --  133 - 0x85  :    9 - 0x9
    "00011100", --  134 - 0x86  :   28 - 0x1c
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00001111", --  136 - 0x88  :   15 - 0xf -- Sprite 0x11
    "00001111", --  137 - 0x89  :   15 - 0xf
    "00001111", --  138 - 0x8a  :   15 - 0xf
    "11111111", --  139 - 0x8b  :  255 - 0xff
    "11111111", --  140 - 0x8c  :  255 - 0xff
    "11111100", --  141 - 0x8d  :  252 - 0xfc
    "10000001", --  142 - 0x8e  :  129 - 0x81
    "00000001", --  143 - 0x8f  :    1 - 0x1
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Sprite 0x12
    "11000000", --  145 - 0x91  :  192 - 0xc0
    "11111000", --  146 - 0x92  :  248 - 0xf8
    "10000000", --  147 - 0x93  :  128 - 0x80
    "00100000", --  148 - 0x94  :   32 - 0x20
    "10010000", --  149 - 0x95  :  144 - 0x90
    "00111100", --  150 - 0x96  :   60 - 0x3c
    "00000000", --  151 - 0x97  :    0 - 0x0
    "11100000", --  152 - 0x98  :  224 - 0xe0 -- Sprite 0x13
    "11110000", --  153 - 0x99  :  240 - 0xf0
    "11110000", --  154 - 0x9a  :  240 - 0xf0
    "11110000", --  155 - 0x9b  :  240 - 0xf0
    "11110000", --  156 - 0x9c  :  240 - 0xf0
    "11100000", --  157 - 0x9d  :  224 - 0xe0
    "11000000", --  158 - 0x9e  :  192 - 0xc0
    "11100000", --  159 - 0x9f  :  224 - 0xe0
    "00000100", --  160 - 0xa0  :    4 - 0x4 -- Sprite 0x14
    "00001100", --  161 - 0xa1  :   12 - 0xc
    "00001100", --  162 - 0xa2  :   12 - 0xc
    "00010011", --  163 - 0xa3  :   19 - 0x13
    "00010011", --  164 - 0xa4  :   19 - 0x13
    "00111011", --  165 - 0xa5  :   59 - 0x3b
    "00000111", --  166 - 0xa6  :    7 - 0x7
    "00001111", --  167 - 0xa7  :   15 - 0xf
    "00001111", --  168 - 0xa8  :   15 - 0xf -- Sprite 0x15
    "00001111", --  169 - 0xa9  :   15 - 0xf
    "00001111", --  170 - 0xaa  :   15 - 0xf
    "00011111", --  171 - 0xab  :   31 - 0x1f
    "00011111", --  172 - 0xac  :   31 - 0x1f
    "00011110", --  173 - 0xad  :   30 - 0x1e
    "00011100", --  174 - 0xae  :   28 - 0x1c
    "00011110", --  175 - 0xaf  :   30 - 0x1e
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0x16
    "01110000", --  177 - 0xb1  :  112 - 0x70
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "11000000", --  179 - 0xb3  :  192 - 0xc0
    "10100000", --  180 - 0xb4  :  160 - 0xa0
    "11111000", --  181 - 0xb5  :  248 - 0xf8
    "10000000", --  182 - 0xb6  :  128 - 0x80
    "11000000", --  183 - 0xb7  :  192 - 0xc0
    "11100000", --  184 - 0xb8  :  224 - 0xe0 -- Sprite 0x17
    "01100000", --  185 - 0xb9  :   96 - 0x60
    "11110000", --  186 - 0xba  :  240 - 0xf0
    "11110000", --  187 - 0xbb  :  240 - 0xf0
    "11110000", --  188 - 0xbc  :  240 - 0xf0
    "11100000", --  189 - 0xbd  :  224 - 0xe0
    "11100000", --  190 - 0xbe  :  224 - 0xe0
    "11110000", --  191 - 0xbf  :  240 - 0xf0
    "00000111", --  192 - 0xc0  :    7 - 0x7 -- Sprite 0x18
    "00001111", --  193 - 0xc1  :   15 - 0xf
    "00001111", --  194 - 0xc2  :   15 - 0xf
    "00010010", --  195 - 0xc3  :   18 - 0x12
    "00010011", --  196 - 0xc4  :   19 - 0x13
    "00111000", --  197 - 0xc5  :   56 - 0x38
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00001111", --  199 - 0xc7  :   15 - 0xf
    "00011111", --  200 - 0xc8  :   31 - 0x1f -- Sprite 0x19
    "00011111", --  201 - 0xc9  :   31 - 0x1f
    "00011111", --  202 - 0xca  :   31 - 0x1f
    "00011111", --  203 - 0xcb  :   31 - 0x1f
    "00011111", --  204 - 0xcc  :   31 - 0x1f
    "00011110", --  205 - 0xcd  :   30 - 0x1e
    "00011100", --  206 - 0xce  :   28 - 0x1c
    "00011110", --  207 - 0xcf  :   30 - 0x1e
    "10000000", --  208 - 0xd0  :  128 - 0x80 -- Sprite 0x1a
    "11110000", --  209 - 0xd1  :  240 - 0xf0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "01000000", --  211 - 0xd3  :   64 - 0x40
    "00100000", --  212 - 0xd4  :   32 - 0x20
    "01111000", --  213 - 0xd5  :  120 - 0x78
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "11000000", --  215 - 0xd7  :  192 - 0xc0
    "11111000", --  216 - 0xd8  :  248 - 0xf8 -- Sprite 0x1b
    "11111000", --  217 - 0xd9  :  248 - 0xf8
    "11110000", --  218 - 0xda  :  240 - 0xf0
    "11110000", --  219 - 0xdb  :  240 - 0xf0
    "11110000", --  220 - 0xdc  :  240 - 0xf0
    "11100000", --  221 - 0xdd  :  224 - 0xe0
    "11100000", --  222 - 0xde  :  224 - 0xe0
    "11110000", --  223 - 0xdf  :  240 - 0xf0
    "00000100", --  224 - 0xe0  :    4 - 0x4 -- Sprite 0x1c
    "00001100", --  225 - 0xe1  :   12 - 0xc
    "00001100", --  226 - 0xe2  :   12 - 0xc
    "00010011", --  227 - 0xe3  :   19 - 0x13
    "00010011", --  228 - 0xe4  :   19 - 0x13
    "00111111", --  229 - 0xe5  :   63 - 0x3f
    "00000111", --  230 - 0xe6  :    7 - 0x7
    "00001111", --  231 - 0xe7  :   15 - 0xf
    "00001111", --  232 - 0xe8  :   15 - 0xf -- Sprite 0x1d
    "00001111", --  233 - 0xe9  :   15 - 0xf
    "00001111", --  234 - 0xea  :   15 - 0xf
    "00011111", --  235 - 0xeb  :   31 - 0x1f
    "00111111", --  236 - 0xec  :   63 - 0x3f
    "01111100", --  237 - 0xed  :  124 - 0x7c
    "01110000", --  238 - 0xee  :  112 - 0x70
    "00111000", --  239 - 0xef  :   56 - 0x38
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Sprite 0x1e
    "01110000", --  241 - 0xf1  :  112 - 0x70
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "11000000", --  243 - 0xf3  :  192 - 0xc0
    "10100000", --  244 - 0xf4  :  160 - 0xa0
    "11111000", --  245 - 0xf5  :  248 - 0xf8
    "10000000", --  246 - 0xf6  :  128 - 0x80
    "11000000", --  247 - 0xf7  :  192 - 0xc0
    "11000000", --  248 - 0xf8  :  192 - 0xc0 -- Sprite 0x1f
    "01100000", --  249 - 0xf9  :   96 - 0x60
    "11100100", --  250 - 0xfa  :  228 - 0xe4
    "11111100", --  251 - 0xfb  :  252 - 0xfc
    "11111100", --  252 - 0xfc  :  252 - 0xfc
    "01111100", --  253 - 0xfd  :  124 - 0x7c
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000111", --  256 - 0x100  :    7 - 0x7 -- Sprite 0x20
    "00001111", --  257 - 0x101  :   15 - 0xf
    "00001111", --  258 - 0x102  :   15 - 0xf
    "00010010", --  259 - 0x103  :   18 - 0x12
    "00010011", --  260 - 0x104  :   19 - 0x13
    "00111000", --  261 - 0x105  :   56 - 0x38
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000111", --  263 - 0x107  :    7 - 0x7
    "00001111", --  264 - 0x108  :   15 - 0xf -- Sprite 0x21
    "00001111", --  265 - 0x109  :   15 - 0xf
    "00001111", --  266 - 0x10a  :   15 - 0xf
    "00011111", --  267 - 0x10b  :   31 - 0x1f
    "00111111", --  268 - 0x10c  :   63 - 0x3f
    "01111100", --  269 - 0x10d  :  124 - 0x7c
    "01110000", --  270 - 0x10e  :  112 - 0x70
    "00111000", --  271 - 0x10f  :   56 - 0x38
    "10000000", --  272 - 0x110  :  128 - 0x80 -- Sprite 0x22
    "11110000", --  273 - 0x111  :  240 - 0xf0
    "00000000", --  274 - 0x112  :    0 - 0x0
    "01000000", --  275 - 0x113  :   64 - 0x40
    "00100000", --  276 - 0x114  :   32 - 0x20
    "01111000", --  277 - 0x115  :  120 - 0x78
    "00000000", --  278 - 0x116  :    0 - 0x0
    "11000000", --  279 - 0x117  :  192 - 0xc0
    "11111000", --  280 - 0x118  :  248 - 0xf8 -- Sprite 0x23
    "11111000", --  281 - 0x119  :  248 - 0xf8
    "11100000", --  282 - 0x11a  :  224 - 0xe0
    "11111100", --  283 - 0x11b  :  252 - 0xfc
    "11111100", --  284 - 0x11c  :  252 - 0xfc
    "01111100", --  285 - 0x11d  :  124 - 0x7c
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Sprite 0x24
    "00000111", --  289 - 0x121  :    7 - 0x7
    "00000111", --  290 - 0x122  :    7 - 0x7
    "00001111", --  291 - 0x123  :   15 - 0xf
    "00001111", --  292 - 0x124  :   15 - 0xf
    "00111000", --  293 - 0x125  :   56 - 0x38
    "01111111", --  294 - 0x126  :  127 - 0x7f
    "01111111", --  295 - 0x127  :  127 - 0x7f
    "00011111", --  296 - 0x128  :   31 - 0x1f -- Sprite 0x25
    "00011111", --  297 - 0x129  :   31 - 0x1f
    "00011111", --  298 - 0x12a  :   31 - 0x1f
    "00011111", --  299 - 0x12b  :   31 - 0x1f
    "00001111", --  300 - 0x12c  :   15 - 0xf
    "00001111", --  301 - 0x12d  :   15 - 0xf
    "00001111", --  302 - 0x12e  :   15 - 0xf
    "00000111", --  303 - 0x12f  :    7 - 0x7
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x26
    "11100000", --  305 - 0x131  :  224 - 0xe0
    "11111000", --  306 - 0x132  :  248 - 0xf8
    "11111100", --  307 - 0x133  :  252 - 0xfc
    "11111100", --  308 - 0x134  :  252 - 0xfc
    "00011100", --  309 - 0x135  :   28 - 0x1c
    "11111000", --  310 - 0x136  :  248 - 0xf8
    "11111000", --  311 - 0x137  :  248 - 0xf8
    "11111000", --  312 - 0x138  :  248 - 0xf8 -- Sprite 0x27
    "11111100", --  313 - 0x139  :  252 - 0xfc
    "11111100", --  314 - 0x13a  :  252 - 0xfc
    "11111000", --  315 - 0x13b  :  248 - 0xf8
    "01111000", --  316 - 0x13c  :  120 - 0x78
    "10000000", --  317 - 0x13d  :  128 - 0x80
    "11000000", --  318 - 0x13e  :  192 - 0xc0
    "11000000", --  319 - 0x13f  :  192 - 0xc0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Sprite 0x28
    "00000011", --  321 - 0x141  :    3 - 0x3
    "00000111", --  322 - 0x142  :    7 - 0x7
    "00000111", --  323 - 0x143  :    7 - 0x7
    "00001001", --  324 - 0x144  :    9 - 0x9
    "00001001", --  325 - 0x145  :    9 - 0x9
    "00011100", --  326 - 0x146  :   28 - 0x1c
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00011111", --  328 - 0x148  :   31 - 0x1f -- Sprite 0x29
    "00001111", --  329 - 0x149  :   15 - 0xf
    "00000111", --  330 - 0x14a  :    7 - 0x7
    "00110111", --  331 - 0x14b  :   55 - 0x37
    "01111111", --  332 - 0x14c  :  127 - 0x7f
    "11011111", --  333 - 0x14d  :  223 - 0xdf
    "00001111", --  334 - 0x14e  :   15 - 0xf
    "00000110", --  335 - 0x14f  :    6 - 0x6
    "00000000", --  336 - 0x150  :    0 - 0x0 -- Sprite 0x2a
    "11000000", --  337 - 0x151  :  192 - 0xc0
    "11111000", --  338 - 0x152  :  248 - 0xf8
    "10000000", --  339 - 0x153  :  128 - 0x80
    "00100000", --  340 - 0x154  :   32 - 0x20
    "10010000", --  341 - 0x155  :  144 - 0x90
    "00111100", --  342 - 0x156  :   60 - 0x3c
    "00000000", --  343 - 0x157  :    0 - 0x0
    "11100100", --  344 - 0x158  :  228 - 0xe4 -- Sprite 0x2b
    "11111110", --  345 - 0x159  :  254 - 0xfe
    "01110000", --  346 - 0x15a  :  112 - 0x70
    "11110001", --  347 - 0x15b  :  241 - 0xf1
    "11111111", --  348 - 0x15c  :  255 - 0xff
    "11111111", --  349 - 0x15d  :  255 - 0xff
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000111", --  352 - 0x160  :    7 - 0x7 -- Sprite 0x2c
    "00001111", --  353 - 0x161  :   15 - 0xf
    "00001111", --  354 - 0x162  :   15 - 0xf
    "00010010", --  355 - 0x163  :   18 - 0x12
    "00010011", --  356 - 0x164  :   19 - 0x13
    "00111000", --  357 - 0x165  :   56 - 0x38
    "01110000", --  358 - 0x166  :  112 - 0x70
    "11111111", --  359 - 0x167  :  255 - 0xff
    "11011111", --  360 - 0x168  :  223 - 0xdf -- Sprite 0x2d
    "00011110", --  361 - 0x169  :   30 - 0x1e
    "00011111", --  362 - 0x16a  :   31 - 0x1f
    "00011111", --  363 - 0x16b  :   31 - 0x1f
    "00011111", --  364 - 0x16c  :   31 - 0x1f
    "00001111", --  365 - 0x16d  :   15 - 0xf
    "00000111", --  366 - 0x16e  :    7 - 0x7
    "00000001", --  367 - 0x16f  :    1 - 0x1
    "10000000", --  368 - 0x170  :  128 - 0x80 -- Sprite 0x2e
    "11110000", --  369 - 0x171  :  240 - 0xf0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "01000000", --  371 - 0x173  :   64 - 0x40
    "00100000", --  372 - 0x174  :   32 - 0x20
    "01111000", --  373 - 0x175  :  120 - 0x78
    "00000000", --  374 - 0x176  :    0 - 0x0
    "11111100", --  375 - 0x177  :  252 - 0xfc
    "11110000", --  376 - 0x178  :  240 - 0xf0 -- Sprite 0x2f
    "11100000", --  377 - 0x179  :  224 - 0xe0
    "11100000", --  378 - 0x17a  :  224 - 0xe0
    "11110000", --  379 - 0x17b  :  240 - 0xf0
    "11111010", --  380 - 0x17c  :  250 - 0xfa
    "11111110", --  381 - 0x17d  :  254 - 0xfe
    "11111100", --  382 - 0x17e  :  252 - 0xfc
    "11011000", --  383 - 0x17f  :  216 - 0xd8
    "00000000", --  384 - 0x180  :    0 - 0x0 -- Sprite 0x30
    "00000000", --  385 - 0x181  :    0 - 0x0
    "00000111", --  386 - 0x182  :    7 - 0x7
    "00001000", --  387 - 0x183  :    8 - 0x8
    "00010000", --  388 - 0x184  :   16 - 0x10
    "00100000", --  389 - 0x185  :   32 - 0x20
    "01000000", --  390 - 0x186  :   64 - 0x40
    "01000000", --  391 - 0x187  :   64 - 0x40
    "01000000", --  392 - 0x188  :   64 - 0x40 -- Sprite 0x31
    "01000000", --  393 - 0x189  :   64 - 0x40
    "00100000", --  394 - 0x18a  :   32 - 0x20
    "00010000", --  395 - 0x18b  :   16 - 0x10
    "00001000", --  396 - 0x18c  :    8 - 0x8
    "00000111", --  397 - 0x18d  :    7 - 0x7
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Sprite 0x32
    "00000000", --  401 - 0x191  :    0 - 0x0
    "11100000", --  402 - 0x192  :  224 - 0xe0
    "00010000", --  403 - 0x193  :   16 - 0x10
    "00001000", --  404 - 0x194  :    8 - 0x8
    "00000100", --  405 - 0x195  :    4 - 0x4
    "00000010", --  406 - 0x196  :    2 - 0x2
    "00000010", --  407 - 0x197  :    2 - 0x2
    "00000010", --  408 - 0x198  :    2 - 0x2 -- Sprite 0x33
    "00000010", --  409 - 0x199  :    2 - 0x2
    "00000100", --  410 - 0x19a  :    4 - 0x4
    "00001000", --  411 - 0x19b  :    8 - 0x8
    "00010000", --  412 - 0x19c  :   16 - 0x10
    "11100000", --  413 - 0x19d  :  224 - 0xe0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- Sprite 0x34
    "00000000", --  417 - 0x1a1  :    0 - 0x0
    "00000000", --  418 - 0x1a2  :    0 - 0x0
    "00000000", --  419 - 0x1a3  :    0 - 0x0
    "00000011", --  420 - 0x1a4  :    3 - 0x3
    "00000100", --  421 - 0x1a5  :    4 - 0x4
    "00001000", --  422 - 0x1a6  :    8 - 0x8
    "00010000", --  423 - 0x1a7  :   16 - 0x10
    "00010000", --  424 - 0x1a8  :   16 - 0x10 -- Sprite 0x35
    "00001000", --  425 - 0x1a9  :    8 - 0x8
    "00000100", --  426 - 0x1aa  :    4 - 0x4
    "00000011", --  427 - 0x1ab  :    3 - 0x3
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x36
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00000000", --  434 - 0x1b2  :    0 - 0x0
    "00000000", --  435 - 0x1b3  :    0 - 0x0
    "11000000", --  436 - 0x1b4  :  192 - 0xc0
    "00100000", --  437 - 0x1b5  :   32 - 0x20
    "00010000", --  438 - 0x1b6  :   16 - 0x10
    "00001000", --  439 - 0x1b7  :    8 - 0x8
    "00001000", --  440 - 0x1b8  :    8 - 0x8 -- Sprite 0x37
    "00010000", --  441 - 0x1b9  :   16 - 0x10
    "00100000", --  442 - 0x1ba  :   32 - 0x20
    "11000000", --  443 - 0x1bb  :  192 - 0xc0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Sprite 0x38
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "00000000", --  453 - 0x1c5  :    0 - 0x0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000001", --  455 - 0x1c7  :    1 - 0x1
    "00000010", --  456 - 0x1c8  :    2 - 0x2 -- Sprite 0x39
    "00000001", --  457 - 0x1c9  :    1 - 0x1
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "00000000", --  467 - 0x1d3  :    0 - 0x0
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "00000000", --  469 - 0x1d5  :    0 - 0x0
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "10000000", --  472 - 0x1d8  :  128 - 0x80 -- Sprite 0x3b
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000001", --  483 - 0x1e3  :    1 - 0x1
    "00100001", --  484 - 0x1e4  :   33 - 0x21
    "00010000", --  485 - 0x1e5  :   16 - 0x10
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "01100000", --  488 - 0x1e8  :   96 - 0x60 -- Sprite 0x3d
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00010000", --  491 - 0x1eb  :   16 - 0x10
    "00100001", --  492 - 0x1ec  :   33 - 0x21
    "00000001", --  493 - 0x1ed  :    1 - 0x1
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Sprite 0x3e
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00001000", --  500 - 0x1f4  :    8 - 0x8
    "00010000", --  501 - 0x1f5  :   16 - 0x10
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "00001100", --  504 - 0x1f8  :   12 - 0xc -- Sprite 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00010000", --  507 - 0x1fb  :   16 - 0x10
    "00001000", --  508 - 0x1fc  :    8 - 0x8
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000100", --  512 - 0x200  :    4 - 0x4 -- Sprite 0x40
    "00000010", --  513 - 0x201  :    2 - 0x2
    "00000001", --  514 - 0x202  :    1 - 0x1
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0 -- Sprite 0x41
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000001", --  526 - 0x20e  :    1 - 0x1
    "00000011", --  527 - 0x20f  :    3 - 0x3
    "00000111", --  528 - 0x210  :    7 - 0x7 -- Sprite 0x42
    "00000111", --  529 - 0x211  :    7 - 0x7
    "00000111", --  530 - 0x212  :    7 - 0x7
    "00000011", --  531 - 0x213  :    3 - 0x3
    "00000001", --  532 - 0x214  :    1 - 0x1
    "00000000", --  533 - 0x215  :    0 - 0x0
    "00000000", --  534 - 0x216  :    0 - 0x0
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00000000", --  536 - 0x218  :    0 - 0x0 -- Sprite 0x43
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Sprite 0x44
    "01000010", --  545 - 0x221  :   66 - 0x42
    "00111001", --  546 - 0x222  :   57 - 0x39
    "11111111", --  547 - 0x223  :  255 - 0xff
    "11111111", --  548 - 0x224  :  255 - 0xff
    "11111111", --  549 - 0x225  :  255 - 0xff
    "11111111", --  550 - 0x226  :  255 - 0xff
    "11111111", --  551 - 0x227  :  255 - 0xff
    "01111111", --  552 - 0x228  :  127 - 0x7f -- Sprite 0x45
    "00111111", --  553 - 0x229  :   63 - 0x3f
    "00011111", --  554 - 0x22a  :   31 - 0x1f
    "00001111", --  555 - 0x22b  :   15 - 0xf
    "00011111", --  556 - 0x22c  :   31 - 0x1f
    "11111111", --  557 - 0x22d  :  255 - 0xff
    "11111111", --  558 - 0x22e  :  255 - 0xff
    "11111111", --  559 - 0x22f  :  255 - 0xff
    "11111000", --  560 - 0x230  :  248 - 0xf8 -- Sprite 0x46
    "11110111", --  561 - 0x231  :  247 - 0xf7
    "11101111", --  562 - 0x232  :  239 - 0xef
    "11111111", --  563 - 0x233  :  255 - 0xff
    "11111111", --  564 - 0x234  :  255 - 0xff
    "11111110", --  565 - 0x235  :  254 - 0xfe
    "01111110", --  566 - 0x236  :  126 - 0x7e
    "00111110", --  567 - 0x237  :   62 - 0x3e
    "00000111", --  568 - 0x238  :    7 - 0x7 -- Sprite 0x47
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Sprite 0x48
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "11000000", --  579 - 0x243  :  192 - 0xc0
    "11100000", --  580 - 0x244  :  224 - 0xe0
    "11110000", --  581 - 0x245  :  240 - 0xf0
    "11011011", --  582 - 0x246  :  219 - 0xdb
    "11110110", --  583 - 0x247  :  246 - 0xf6
    "11001011", --  584 - 0x248  :  203 - 0xcb -- Sprite 0x49
    "11100000", --  585 - 0x249  :  224 - 0xe0
    "11000100", --  586 - 0x24a  :  196 - 0xc4
    "00000010", --  587 - 0x24b  :    2 - 0x2
    "11010001", --  588 - 0x24c  :  209 - 0xd1
    "11100001", --  589 - 0x24d  :  225 - 0xe1
    "11010001", --  590 - 0x24e  :  209 - 0xd1
    "10000011", --  591 - 0x24f  :  131 - 0x83
    "00001111", --  592 - 0x250  :   15 - 0xf -- Sprite 0x4a
    "11111111", --  593 - 0x251  :  255 - 0xff
    "11100000", --  594 - 0x252  :  224 - 0xe0
    "10001111", --  595 - 0x253  :  143 - 0x8f
    "01101110", --  596 - 0x254  :  110 - 0x6e
    "01000100", --  597 - 0x255  :   68 - 0x44
    "11101110", --  598 - 0x256  :  238 - 0xee
    "01100000", --  599 - 0x257  :   96 - 0x60
    "10000011", --  600 - 0x258  :  131 - 0x83 -- Sprite 0x4b
    "11100000", --  601 - 0x259  :  224 - 0xe0
    "11100100", --  602 - 0x25a  :  228 - 0xe4
    "11000110", --  603 - 0x25b  :  198 - 0xc6
    "01100001", --  604 - 0x25c  :   97 - 0x61
    "00110011", --  605 - 0x25d  :   51 - 0x33
    "00011111", --  606 - 0x25e  :   31 - 0x1f
    "00001111", --  607 - 0x25f  :   15 - 0xf
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Sprite 0x4c
    "00000000", --  609 - 0x261  :    0 - 0x0
    "00000000", --  610 - 0x262  :    0 - 0x0
    "00000011", --  611 - 0x263  :    3 - 0x3
    "00000111", --  612 - 0x264  :    7 - 0x7
    "00001111", --  613 - 0x265  :   15 - 0xf
    "01011011", --  614 - 0x266  :   91 - 0x5b
    "10100111", --  615 - 0x267  :  167 - 0xa7
    "01110011", --  616 - 0x268  :  115 - 0x73 -- Sprite 0x4d
    "00000111", --  617 - 0x269  :    7 - 0x7
    "00100111", --  618 - 0x26a  :   39 - 0x27
    "01000000", --  619 - 0x26b  :   64 - 0x40
    "10001011", --  620 - 0x26c  :  139 - 0x8b
    "10000111", --  621 - 0x26d  :  135 - 0x87
    "10001011", --  622 - 0x26e  :  139 - 0x8b
    "11000001", --  623 - 0x26f  :  193 - 0xc1
    "11110000", --  624 - 0x270  :  240 - 0xf0 -- Sprite 0x4e
    "11111111", --  625 - 0x271  :  255 - 0xff
    "00001111", --  626 - 0x272  :   15 - 0xf
    "11100001", --  627 - 0x273  :  225 - 0xe1
    "11101100", --  628 - 0x274  :  236 - 0xec
    "01000100", --  629 - 0x275  :   68 - 0x44
    "11101110", --  630 - 0x276  :  238 - 0xee
    "00001100", --  631 - 0x277  :   12 - 0xc
    "10000000", --  632 - 0x278  :  128 - 0x80 -- Sprite 0x4f
    "00001110", --  633 - 0x279  :   14 - 0xe
    "01001110", --  634 - 0x27a  :   78 - 0x4e
    "11000110", --  635 - 0x27b  :  198 - 0xc6
    "00001100", --  636 - 0x27c  :   12 - 0xc
    "10011000", --  637 - 0x27d  :  152 - 0x98
    "11110000", --  638 - 0x27e  :  240 - 0xf0
    "11100000", --  639 - 0x27f  :  224 - 0xe0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x50
    "01000010", --  641 - 0x281  :   66 - 0x42
    "10011100", --  642 - 0x282  :  156 - 0x9c
    "11111111", --  643 - 0x283  :  255 - 0xff
    "11111111", --  644 - 0x284  :  255 - 0xff
    "11111111", --  645 - 0x285  :  255 - 0xff
    "11111111", --  646 - 0x286  :  255 - 0xff
    "11111111", --  647 - 0x287  :  255 - 0xff
    "11111110", --  648 - 0x288  :  254 - 0xfe -- Sprite 0x51
    "11111100", --  649 - 0x289  :  252 - 0xfc
    "11111000", --  650 - 0x28a  :  248 - 0xf8
    "11110000", --  651 - 0x28b  :  240 - 0xf0
    "11111000", --  652 - 0x28c  :  248 - 0xf8
    "11111111", --  653 - 0x28d  :  255 - 0xff
    "11111111", --  654 - 0x28e  :  255 - 0xff
    "11111111", --  655 - 0x28f  :  255 - 0xff
    "00011111", --  656 - 0x290  :   31 - 0x1f -- Sprite 0x52
    "11101111", --  657 - 0x291  :  239 - 0xef
    "11110111", --  658 - 0x292  :  247 - 0xf7
    "11111111", --  659 - 0x293  :  255 - 0xff
    "11111111", --  660 - 0x294  :  255 - 0xff
    "11111110", --  661 - 0x295  :  254 - 0xfe
    "01111100", --  662 - 0x296  :  124 - 0x7c
    "01110000", --  663 - 0x297  :  112 - 0x70
    "11100000", --  664 - 0x298  :  224 - 0xe0 -- Sprite 0x53
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00100000", --  672 - 0x2a0  :   32 - 0x20 -- Sprite 0x54
    "01000000", --  673 - 0x2a1  :   64 - 0x40
    "10000000", --  674 - 0x2a2  :  128 - 0x80
    "00000000", --  675 - 0x2a3  :    0 - 0x0
    "00000000", --  676 - 0x2a4  :    0 - 0x0
    "00000000", --  677 - 0x2a5  :    0 - 0x0
    "00000000", --  678 - 0x2a6  :    0 - 0x0
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- Sprite 0x55
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "10000000", --  686 - 0x2ae  :  128 - 0x80
    "11000000", --  687 - 0x2af  :  192 - 0xc0
    "11100000", --  688 - 0x2b0  :  224 - 0xe0 -- Sprite 0x56
    "11100000", --  689 - 0x2b1  :  224 - 0xe0
    "11100000", --  690 - 0x2b2  :  224 - 0xe0
    "11000000", --  691 - 0x2b3  :  192 - 0xc0
    "10000000", --  692 - 0x2b4  :  128 - 0x80
    "00000000", --  693 - 0x2b5  :    0 - 0x0
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "00000000", --  696 - 0x2b8  :    0 - 0x0 -- Sprite 0x57
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "11111111", --  704 - 0x2c0  :  255 - 0xff -- Sprite 0x58
    "11111111", --  705 - 0x2c1  :  255 - 0xff
    "11111111", --  706 - 0x2c2  :  255 - 0xff
    "11111111", --  707 - 0x2c3  :  255 - 0xff
    "11111111", --  708 - 0x2c4  :  255 - 0xff
    "11111111", --  709 - 0x2c5  :  255 - 0xff
    "11111111", --  710 - 0x2c6  :  255 - 0xff
    "11111111", --  711 - 0x2c7  :  255 - 0xff
    "11111111", --  712 - 0x2c8  :  255 - 0xff -- Sprite 0x59
    "11111111", --  713 - 0x2c9  :  255 - 0xff
    "11111111", --  714 - 0x2ca  :  255 - 0xff
    "11111111", --  715 - 0x2cb  :  255 - 0xff
    "11111111", --  716 - 0x2cc  :  255 - 0xff
    "11111111", --  717 - 0x2cd  :  255 - 0xff
    "11111111", --  718 - 0x2ce  :  255 - 0xff
    "11111111", --  719 - 0x2cf  :  255 - 0xff
    "11111111", --  720 - 0x2d0  :  255 - 0xff -- Sprite 0x5a
    "11111111", --  721 - 0x2d1  :  255 - 0xff
    "11111111", --  722 - 0x2d2  :  255 - 0xff
    "11111111", --  723 - 0x2d3  :  255 - 0xff
    "11111111", --  724 - 0x2d4  :  255 - 0xff
    "11111111", --  725 - 0x2d5  :  255 - 0xff
    "11111111", --  726 - 0x2d6  :  255 - 0xff
    "11111111", --  727 - 0x2d7  :  255 - 0xff
    "11111111", --  728 - 0x2d8  :  255 - 0xff -- Sprite 0x5b
    "11111111", --  729 - 0x2d9  :  255 - 0xff
    "11111111", --  730 - 0x2da  :  255 - 0xff
    "11111111", --  731 - 0x2db  :  255 - 0xff
    "11111111", --  732 - 0x2dc  :  255 - 0xff
    "11111111", --  733 - 0x2dd  :  255 - 0xff
    "11111111", --  734 - 0x2de  :  255 - 0xff
    "11111111", --  735 - 0x2df  :  255 - 0xff
    "11111111", --  736 - 0x2e0  :  255 - 0xff -- Sprite 0x5c
    "11111111", --  737 - 0x2e1  :  255 - 0xff
    "11111111", --  738 - 0x2e2  :  255 - 0xff
    "11111111", --  739 - 0x2e3  :  255 - 0xff
    "11111111", --  740 - 0x2e4  :  255 - 0xff
    "11111111", --  741 - 0x2e5  :  255 - 0xff
    "11111111", --  742 - 0x2e6  :  255 - 0xff
    "11111111", --  743 - 0x2e7  :  255 - 0xff
    "11111111", --  744 - 0x2e8  :  255 - 0xff -- Sprite 0x5d
    "11111111", --  745 - 0x2e9  :  255 - 0xff
    "11111111", --  746 - 0x2ea  :  255 - 0xff
    "11111111", --  747 - 0x2eb  :  255 - 0xff
    "11111111", --  748 - 0x2ec  :  255 - 0xff
    "11111111", --  749 - 0x2ed  :  255 - 0xff
    "11111111", --  750 - 0x2ee  :  255 - 0xff
    "11111111", --  751 - 0x2ef  :  255 - 0xff
    "11111111", --  752 - 0x2f0  :  255 - 0xff -- Sprite 0x5e
    "11111111", --  753 - 0x2f1  :  255 - 0xff
    "11111111", --  754 - 0x2f2  :  255 - 0xff
    "11111111", --  755 - 0x2f3  :  255 - 0xff
    "11111111", --  756 - 0x2f4  :  255 - 0xff
    "11111111", --  757 - 0x2f5  :  255 - 0xff
    "11111111", --  758 - 0x2f6  :  255 - 0xff
    "11111111", --  759 - 0x2f7  :  255 - 0xff
    "11111111", --  760 - 0x2f8  :  255 - 0xff -- Sprite 0x5f
    "11111111", --  761 - 0x2f9  :  255 - 0xff
    "11111111", --  762 - 0x2fa  :  255 - 0xff
    "11111111", --  763 - 0x2fb  :  255 - 0xff
    "11111111", --  764 - 0x2fc  :  255 - 0xff
    "11111111", --  765 - 0x2fd  :  255 - 0xff
    "11111111", --  766 - 0x2fe  :  255 - 0xff
    "11111111", --  767 - 0x2ff  :  255 - 0xff
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x60
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00011111", --  770 - 0x302  :   31 - 0x1f
    "00111111", --  771 - 0x303  :   63 - 0x3f
    "00111111", --  772 - 0x304  :   63 - 0x3f
    "01111111", --  773 - 0x305  :  127 - 0x7f
    "01111111", --  774 - 0x306  :  127 - 0x7f
    "01111111", --  775 - 0x307  :  127 - 0x7f
    "01111111", --  776 - 0x308  :  127 - 0x7f -- Sprite 0x61
    "00111110", --  777 - 0x309  :   62 - 0x3e
    "00011111", --  778 - 0x30a  :   31 - 0x1f
    "00011111", --  779 - 0x30b  :   31 - 0x1f
    "00001111", --  780 - 0x30c  :   15 - 0xf
    "00001111", --  781 - 0x30d  :   15 - 0xf
    "00001111", --  782 - 0x30e  :   15 - 0xf
    "00000111", --  783 - 0x30f  :    7 - 0x7
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Sprite 0x62
    "01100000", --  785 - 0x311  :   96 - 0x60
    "11110000", --  786 - 0x312  :  240 - 0xf0
    "11111000", --  787 - 0x313  :  248 - 0xf8
    "11111000", --  788 - 0x314  :  248 - 0xf8
    "11111000", --  789 - 0x315  :  248 - 0xf8
    "11111100", --  790 - 0x316  :  252 - 0xfc
    "11111100", --  791 - 0x317  :  252 - 0xfc
    "11111000", --  792 - 0x318  :  248 - 0xf8 -- Sprite 0x63
    "11110000", --  793 - 0x319  :  240 - 0xf0
    "11110000", --  794 - 0x31a  :  240 - 0xf0
    "11100000", --  795 - 0x31b  :  224 - 0xe0
    "10000000", --  796 - 0x31c  :  128 - 0x80
    "10000000", --  797 - 0x31d  :  128 - 0x80
    "11000000", --  798 - 0x31e  :  192 - 0xc0
    "11000000", --  799 - 0x31f  :  192 - 0xc0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Sprite 0x64
    "00011111", --  801 - 0x321  :   31 - 0x1f
    "00111111", --  802 - 0x322  :   63 - 0x3f
    "01111111", --  803 - 0x323  :  127 - 0x7f
    "11111111", --  804 - 0x324  :  255 - 0xff
    "11111111", --  805 - 0x325  :  255 - 0xff
    "00111110", --  806 - 0x326  :   62 - 0x3e
    "00001111", --  807 - 0x327  :   15 - 0xf
    "00000000", --  808 - 0x328  :    0 - 0x0 -- Sprite 0x65
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000001", --  811 - 0x32b  :    1 - 0x1
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "00000000", --  813 - 0x32d  :    0 - 0x0
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Sprite 0x66
    "11100000", --  817 - 0x331  :  224 - 0xe0
    "11110000", --  818 - 0x332  :  240 - 0xf0
    "11111100", --  819 - 0x333  :  252 - 0xfc
    "11111110", --  820 - 0x334  :  254 - 0xfe
    "11111110", --  821 - 0x335  :  254 - 0xfe
    "11111111", --  822 - 0x336  :  255 - 0xff
    "11111100", --  823 - 0x337  :  252 - 0xfc
    "01111100", --  824 - 0x338  :  124 - 0x7c -- Sprite 0x67
    "11111100", --  825 - 0x339  :  252 - 0xfc
    "11111000", --  826 - 0x33a  :  248 - 0xf8
    "11110000", --  827 - 0x33b  :  240 - 0xf0
    "11100000", --  828 - 0x33c  :  224 - 0xe0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x68
    "00000111", --  833 - 0x341  :    7 - 0x7
    "00000111", --  834 - 0x342  :    7 - 0x7
    "00001111", --  835 - 0x343  :   15 - 0xf
    "00001111", --  836 - 0x344  :   15 - 0xf
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00011111", --  838 - 0x346  :   31 - 0x1f
    "00111111", --  839 - 0x347  :   63 - 0x3f
    "01111111", --  840 - 0x348  :  127 - 0x7f -- Sprite 0x69
    "01111111", --  841 - 0x349  :  127 - 0x7f
    "00011111", --  842 - 0x34a  :   31 - 0x1f
    "00011111", --  843 - 0x34b  :   31 - 0x1f
    "00011111", --  844 - 0x34c  :   31 - 0x1f
    "00011110", --  845 - 0x34d  :   30 - 0x1e
    "00001111", --  846 - 0x34e  :   15 - 0xf
    "00011111", --  847 - 0x34f  :   31 - 0x1f
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Sprite 0x6a
    "11100000", --  849 - 0x351  :  224 - 0xe0
    "11100000", --  850 - 0x352  :  224 - 0xe0
    "11110000", --  851 - 0x353  :  240 - 0xf0
    "11110000", --  852 - 0x354  :  240 - 0xf0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "11111000", --  854 - 0x356  :  248 - 0xf8
    "11111100", --  855 - 0x357  :  252 - 0xfc
    "11111110", --  856 - 0x358  :  254 - 0xfe -- Sprite 0x6b
    "11111110", --  857 - 0x359  :  254 - 0xfe
    "11111000", --  858 - 0x35a  :  248 - 0xf8
    "11111000", --  859 - 0x35b  :  248 - 0xf8
    "11111000", --  860 - 0x35c  :  248 - 0xf8
    "01111000", --  861 - 0x35d  :  120 - 0x78
    "11110000", --  862 - 0x35e  :  240 - 0xf0
    "11111000", --  863 - 0x35f  :  248 - 0xf8
    "00000011", --  864 - 0x360  :    3 - 0x3 -- Sprite 0x6c
    "00000111", --  865 - 0x361  :    7 - 0x7
    "00000101", --  866 - 0x362  :    5 - 0x5
    "00001000", --  867 - 0x363  :    8 - 0x8
    "00011011", --  868 - 0x364  :   27 - 0x1b
    "00011001", --  869 - 0x365  :   25 - 0x19
    "00000101", --  870 - 0x366  :    5 - 0x5
    "00111111", --  871 - 0x367  :   63 - 0x3f
    "00111111", --  872 - 0x368  :   63 - 0x3f -- Sprite 0x6d
    "00001111", --  873 - 0x369  :   15 - 0xf
    "00000101", --  874 - 0x36a  :    5 - 0x5
    "00110111", --  875 - 0x36b  :   55 - 0x37
    "00111111", --  876 - 0x36c  :   63 - 0x3f
    "00111111", --  877 - 0x36d  :   63 - 0x3f
    "00111110", --  878 - 0x36e  :   62 - 0x3e
    "00011100", --  879 - 0x36f  :   28 - 0x1c
    "11100000", --  880 - 0x370  :  224 - 0xe0 -- Sprite 0x6e
    "11110000", --  881 - 0x371  :  240 - 0xf0
    "01010000", --  882 - 0x372  :   80 - 0x50
    "00001000", --  883 - 0x373  :    8 - 0x8
    "01101100", --  884 - 0x374  :  108 - 0x6c
    "11001100", --  885 - 0x375  :  204 - 0xcc
    "11010000", --  886 - 0x376  :  208 - 0xd0
    "11111110", --  887 - 0x377  :  254 - 0xfe
    "11111110", --  888 - 0x378  :  254 - 0xfe -- Sprite 0x6f
    "11111000", --  889 - 0x379  :  248 - 0xf8
    "11010000", --  890 - 0x37a  :  208 - 0xd0
    "11111011", --  891 - 0x37b  :  251 - 0xfb
    "11111111", --  892 - 0x37c  :  255 - 0xff
    "11111111", --  893 - 0x37d  :  255 - 0xff
    "00111110", --  894 - 0x37e  :   62 - 0x3e
    "00001100", --  895 - 0x37f  :   12 - 0xc
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Sprite 0x70
    "00000000", --  897 - 0x381  :    0 - 0x0
    "01111001", --  898 - 0x382  :  121 - 0x79
    "11111001", --  899 - 0x383  :  249 - 0xf9
    "11110011", --  900 - 0x384  :  243 - 0xf3
    "11111111", --  901 - 0x385  :  255 - 0xff
    "01111011", --  902 - 0x386  :  123 - 0x7b
    "00111111", --  903 - 0x387  :   63 - 0x3f
    "00111111", --  904 - 0x388  :   63 - 0x3f -- Sprite 0x71
    "00111111", --  905 - 0x389  :   63 - 0x3f
    "01111011", --  906 - 0x38a  :  123 - 0x7b
    "01111111", --  907 - 0x38b  :  127 - 0x7f
    "11111011", --  908 - 0x38c  :  251 - 0xfb
    "11110001", --  909 - 0x38d  :  241 - 0xf1
    "01111001", --  910 - 0x38e  :  121 - 0x79
    "00111000", --  911 - 0x38f  :   56 - 0x38
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Sprite 0x72
    "00000000", --  913 - 0x391  :    0 - 0x0
    "10000000", --  914 - 0x392  :  128 - 0x80
    "10110000", --  915 - 0x393  :  176 - 0xb0
    "10111000", --  916 - 0x394  :  184 - 0xb8
    "11000110", --  917 - 0x395  :  198 - 0xc6
    "10010011", --  918 - 0x396  :  147 - 0x93
    "11110111", --  919 - 0x397  :  247 - 0xf7
    "11100011", --  920 - 0x398  :  227 - 0xe3 -- Sprite 0x73
    "11110111", --  921 - 0x399  :  247 - 0xf7
    "10010011", --  922 - 0x39a  :  147 - 0x93
    "11000110", --  923 - 0x39b  :  198 - 0xc6
    "10111000", --  924 - 0x39c  :  184 - 0xb8
    "10110000", --  925 - 0x39d  :  176 - 0xb0
    "10000000", --  926 - 0x39e  :  128 - 0x80
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00110000", --  928 - 0x3a0  :   48 - 0x30 -- Sprite 0x74
    "01111100", --  929 - 0x3a1  :  124 - 0x7c
    "11111111", --  930 - 0x3a2  :  255 - 0xff
    "11111111", --  931 - 0x3a3  :  255 - 0xff
    "11011111", --  932 - 0x3a4  :  223 - 0xdf
    "00001011", --  933 - 0x3a5  :   11 - 0xb
    "00011111", --  934 - 0x3a6  :   31 - 0x1f
    "01111111", --  935 - 0x3a7  :  127 - 0x7f
    "01111111", --  936 - 0x3a8  :  127 - 0x7f -- Sprite 0x75
    "00001011", --  937 - 0x3a9  :   11 - 0xb
    "00110011", --  938 - 0x3aa  :   51 - 0x33
    "00110110", --  939 - 0x3ab  :   54 - 0x36
    "00010000", --  940 - 0x3ac  :   16 - 0x10
    "00001010", --  941 - 0x3ad  :   10 - 0xa
    "00001111", --  942 - 0x3ae  :   15 - 0xf
    "00000111", --  943 - 0x3af  :    7 - 0x7
    "00111000", --  944 - 0x3b0  :   56 - 0x38 -- Sprite 0x76
    "01111100", --  945 - 0x3b1  :  124 - 0x7c
    "11111100", --  946 - 0x3b2  :  252 - 0xfc
    "11111100", --  947 - 0x3b3  :  252 - 0xfc
    "11101100", --  948 - 0x3b4  :  236 - 0xec
    "10100000", --  949 - 0x3b5  :  160 - 0xa0
    "11110000", --  950 - 0x3b6  :  240 - 0xf0
    "11111100", --  951 - 0x3b7  :  252 - 0xfc
    "11111100", --  952 - 0x3b8  :  252 - 0xfc -- Sprite 0x77
    "10100000", --  953 - 0x3b9  :  160 - 0xa0
    "10011000", --  954 - 0x3ba  :  152 - 0x98
    "11011000", --  955 - 0x3bb  :  216 - 0xd8
    "00010000", --  956 - 0x3bc  :   16 - 0x10
    "10100000", --  957 - 0x3bd  :  160 - 0xa0
    "11100000", --  958 - 0x3be  :  224 - 0xe0
    "11000000", --  959 - 0x3bf  :  192 - 0xc0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x78
    "00000001", --  961 - 0x3c1  :    1 - 0x1
    "00001101", --  962 - 0x3c2  :   13 - 0xd
    "00011101", --  963 - 0x3c3  :   29 - 0x1d
    "01100011", --  964 - 0x3c4  :   99 - 0x63
    "11001001", --  965 - 0x3c5  :  201 - 0xc9
    "11101111", --  966 - 0x3c6  :  239 - 0xef
    "11000111", --  967 - 0x3c7  :  199 - 0xc7
    "11101111", --  968 - 0x3c8  :  239 - 0xef -- Sprite 0x79
    "11001001", --  969 - 0x3c9  :  201 - 0xc9
    "01100011", --  970 - 0x3ca  :   99 - 0x63
    "00011101", --  971 - 0x3cb  :   29 - 0x1d
    "00001101", --  972 - 0x3cc  :   13 - 0xd
    "00000001", --  973 - 0x3cd  :    1 - 0x1
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00011100", --  976 - 0x3d0  :   28 - 0x1c -- Sprite 0x7a
    "10011110", --  977 - 0x3d1  :  158 - 0x9e
    "10001111", --  978 - 0x3d2  :  143 - 0x8f
    "11011111", --  979 - 0x3d3  :  223 - 0xdf
    "11111110", --  980 - 0x3d4  :  254 - 0xfe
    "11011110", --  981 - 0x3d5  :  222 - 0xde
    "11111100", --  982 - 0x3d6  :  252 - 0xfc
    "11111100", --  983 - 0x3d7  :  252 - 0xfc
    "11111100", --  984 - 0x3d8  :  252 - 0xfc -- Sprite 0x7b
    "11011110", --  985 - 0x3d9  :  222 - 0xde
    "11111111", --  986 - 0x3da  :  255 - 0xff
    "11001111", --  987 - 0x3db  :  207 - 0xcf
    "10011111", --  988 - 0x3dc  :  159 - 0x9f
    "10011110", --  989 - 0x3dd  :  158 - 0x9e
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x7c
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00011110", --  996 - 0x3e4  :   30 - 0x1e
    "00111111", --  997 - 0x3e5  :   63 - 0x3f
    "01111101", --  998 - 0x3e6  :  125 - 0x7d
    "01111000", --  999 - 0x3e7  :  120 - 0x78
    "01111100", -- 1000 - 0x3e8  :  124 - 0x7c -- Sprite 0x7d
    "11111011", -- 1001 - 0x3e9  :  251 - 0xfb
    "11111111", -- 1002 - 0x3ea  :  255 - 0xff
    "11111111", -- 1003 - 0x3eb  :  255 - 0xff
    "01011111", -- 1004 - 0x3ec  :   95 - 0x5f
    "00011111", -- 1005 - 0x3ed  :   31 - 0x1f
    "00011111", -- 1006 - 0x3ee  :   31 - 0x1f
    "00011111", -- 1007 - 0x3ef  :   31 - 0x1f
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Sprite 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "10000000", -- 1013 - 0x3f5  :  128 - 0x80
    "10000000", -- 1014 - 0x3f6  :  128 - 0x80
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- Sprite 0x7f
    "00100001", -- 1017 - 0x3f9  :   33 - 0x21
    "10100010", -- 1018 - 0x3fa  :  162 - 0xa2
    "10100011", -- 1019 - 0x3fb  :  163 - 0xa3
    "10110011", -- 1020 - 0x3fc  :  179 - 0xb3
    "10001111", -- 1021 - 0x3fd  :  143 - 0x8f
    "00100111", -- 1022 - 0x3fe  :   39 - 0x27
    "11111110", -- 1023 - 0x3ff  :  254 - 0xfe
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Sprite 0x80
    "00000000", -- 1025 - 0x401  :    0 - 0x0
    "00000000", -- 1026 - 0x402  :    0 - 0x0
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000011", -- 1028 - 0x404  :    3 - 0x3
    "00001111", -- 1029 - 0x405  :   15 - 0xf
    "00011111", -- 1030 - 0x406  :   31 - 0x1f
    "00011111", -- 1031 - 0x407  :   31 - 0x1f
    "00011111", -- 1032 - 0x408  :   31 - 0x1f -- Sprite 0x81
    "00011111", -- 1033 - 0x409  :   31 - 0x1f
    "00001111", -- 1034 - 0x40a  :   15 - 0xf
    "00000011", -- 1035 - 0x40b  :    3 - 0x3
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Sprite 0x82
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "11000000", -- 1044 - 0x414  :  192 - 0xc0
    "11110000", -- 1045 - 0x415  :  240 - 0xf0
    "11111000", -- 1046 - 0x416  :  248 - 0xf8
    "11111000", -- 1047 - 0x417  :  248 - 0xf8
    "11111000", -- 1048 - 0x418  :  248 - 0xf8 -- Sprite 0x83
    "11111000", -- 1049 - 0x419  :  248 - 0xf8
    "11110000", -- 1050 - 0x41a  :  240 - 0xf0
    "11000000", -- 1051 - 0x41b  :  192 - 0xc0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- Sprite 0x84
    "00000000", -- 1057 - 0x421  :    0 - 0x0
    "00000000", -- 1058 - 0x422  :    0 - 0x0
    "00000000", -- 1059 - 0x423  :    0 - 0x0
    "00000011", -- 1060 - 0x424  :    3 - 0x3
    "00001111", -- 1061 - 0x425  :   15 - 0xf
    "00011111", -- 1062 - 0x426  :   31 - 0x1f
    "00011111", -- 1063 - 0x427  :   31 - 0x1f
    "00011111", -- 1064 - 0x428  :   31 - 0x1f -- Sprite 0x85
    "00011111", -- 1065 - 0x429  :   31 - 0x1f
    "00001111", -- 1066 - 0x42a  :   15 - 0xf
    "00000011", -- 1067 - 0x42b  :    3 - 0x3
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Sprite 0x86
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "11000000", -- 1076 - 0x434  :  192 - 0xc0
    "11110000", -- 1077 - 0x435  :  240 - 0xf0
    "11111000", -- 1078 - 0x436  :  248 - 0xf8
    "11111000", -- 1079 - 0x437  :  248 - 0xf8
    "11111000", -- 1080 - 0x438  :  248 - 0xf8 -- Sprite 0x87
    "11111000", -- 1081 - 0x439  :  248 - 0xf8
    "11110000", -- 1082 - 0x43a  :  240 - 0xf0
    "11000000", -- 1083 - 0x43b  :  192 - 0xc0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Sprite 0x88
    "00000000", -- 1089 - 0x441  :    0 - 0x0
    "00000000", -- 1090 - 0x442  :    0 - 0x0
    "00000000", -- 1091 - 0x443  :    0 - 0x0
    "00000011", -- 1092 - 0x444  :    3 - 0x3
    "00001111", -- 1093 - 0x445  :   15 - 0xf
    "00011111", -- 1094 - 0x446  :   31 - 0x1f
    "00011111", -- 1095 - 0x447  :   31 - 0x1f
    "00011111", -- 1096 - 0x448  :   31 - 0x1f -- Sprite 0x89
    "00011111", -- 1097 - 0x449  :   31 - 0x1f
    "00001111", -- 1098 - 0x44a  :   15 - 0xf
    "00000011", -- 1099 - 0x44b  :    3 - 0x3
    "00000000", -- 1100 - 0x44c  :    0 - 0x0
    "00000000", -- 1101 - 0x44d  :    0 - 0x0
    "00000000", -- 1102 - 0x44e  :    0 - 0x0
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Sprite 0x8a
    "00000000", -- 1105 - 0x451  :    0 - 0x0
    "00000000", -- 1106 - 0x452  :    0 - 0x0
    "00000000", -- 1107 - 0x453  :    0 - 0x0
    "11000000", -- 1108 - 0x454  :  192 - 0xc0
    "11110000", -- 1109 - 0x455  :  240 - 0xf0
    "11111000", -- 1110 - 0x456  :  248 - 0xf8
    "11111000", -- 1111 - 0x457  :  248 - 0xf8
    "11111000", -- 1112 - 0x458  :  248 - 0xf8 -- Sprite 0x8b
    "11111000", -- 1113 - 0x459  :  248 - 0xf8
    "11110000", -- 1114 - 0x45a  :  240 - 0xf0
    "11000000", -- 1115 - 0x45b  :  192 - 0xc0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00000000", -- 1117 - 0x45d  :    0 - 0x0
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Sprite 0x8c
    "00000000", -- 1121 - 0x461  :    0 - 0x0
    "00000000", -- 1122 - 0x462  :    0 - 0x0
    "00000000", -- 1123 - 0x463  :    0 - 0x0
    "00000011", -- 1124 - 0x464  :    3 - 0x3
    "00001111", -- 1125 - 0x465  :   15 - 0xf
    "00011111", -- 1126 - 0x466  :   31 - 0x1f
    "00011111", -- 1127 - 0x467  :   31 - 0x1f
    "00011111", -- 1128 - 0x468  :   31 - 0x1f -- Sprite 0x8d
    "00011111", -- 1129 - 0x469  :   31 - 0x1f
    "00001111", -- 1130 - 0x46a  :   15 - 0xf
    "00000011", -- 1131 - 0x46b  :    3 - 0x3
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0 -- Sprite 0x8e
    "00000000", -- 1137 - 0x471  :    0 - 0x0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "11000000", -- 1140 - 0x474  :  192 - 0xc0
    "11110000", -- 1141 - 0x475  :  240 - 0xf0
    "11111000", -- 1142 - 0x476  :  248 - 0xf8
    "11111000", -- 1143 - 0x477  :  248 - 0xf8
    "11111000", -- 1144 - 0x478  :  248 - 0xf8 -- Sprite 0x8f
    "11111000", -- 1145 - 0x479  :  248 - 0xf8
    "11110000", -- 1146 - 0x47a  :  240 - 0xf0
    "11000000", -- 1147 - 0x47b  :  192 - 0xc0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x90
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00001111", -- 1155 - 0x483  :   15 - 0xf
    "00110000", -- 1156 - 0x484  :   48 - 0x30
    "01100000", -- 1157 - 0x485  :   96 - 0x60
    "00111111", -- 1158 - 0x486  :   63 - 0x3f
    "01111111", -- 1159 - 0x487  :  127 - 0x7f
    "01111111", -- 1160 - 0x488  :  127 - 0x7f -- Sprite 0x91
    "00111111", -- 1161 - 0x489  :   63 - 0x3f
    "01100000", -- 1162 - 0x48a  :   96 - 0x60
    "00110000", -- 1163 - 0x48b  :   48 - 0x30
    "00001111", -- 1164 - 0x48c  :   15 - 0xf
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0 -- Sprite 0x92
    "00000000", -- 1169 - 0x491  :    0 - 0x0
    "00000000", -- 1170 - 0x492  :    0 - 0x0
    "11111000", -- 1171 - 0x493  :  248 - 0xf8
    "00000110", -- 1172 - 0x494  :    6 - 0x6
    "00000011", -- 1173 - 0x495  :    3 - 0x3
    "11111110", -- 1174 - 0x496  :  254 - 0xfe
    "11111111", -- 1175 - 0x497  :  255 - 0xff
    "11111111", -- 1176 - 0x498  :  255 - 0xff -- Sprite 0x93
    "11111110", -- 1177 - 0x499  :  254 - 0xfe
    "00000011", -- 1178 - 0x49a  :    3 - 0x3
    "00000110", -- 1179 - 0x49b  :    6 - 0x6
    "11111000", -- 1180 - 0x49c  :  248 - 0xf8
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- Sprite 0x94
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000000", -- 1186 - 0x4a2  :    0 - 0x0
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00101111", -- 1188 - 0x4a4  :   47 - 0x2f
    "00111111", -- 1189 - 0x4a5  :   63 - 0x3f
    "01100000", -- 1190 - 0x4a6  :   96 - 0x60
    "00100000", -- 1191 - 0x4a7  :   32 - 0x20
    "00100000", -- 1192 - 0x4a8  :   32 - 0x20 -- Sprite 0x95
    "01100000", -- 1193 - 0x4a9  :   96 - 0x60
    "00111111", -- 1194 - 0x4aa  :   63 - 0x3f
    "00101111", -- 1195 - 0x4ab  :   47 - 0x2f
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0 -- Sprite 0x96
    "00000000", -- 1201 - 0x4b1  :    0 - 0x0
    "00000000", -- 1202 - 0x4b2  :    0 - 0x0
    "00000000", -- 1203 - 0x4b3  :    0 - 0x0
    "11111010", -- 1204 - 0x4b4  :  250 - 0xfa
    "11111110", -- 1205 - 0x4b5  :  254 - 0xfe
    "00000011", -- 1206 - 0x4b6  :    3 - 0x3
    "00000010", -- 1207 - 0x4b7  :    2 - 0x2
    "00000010", -- 1208 - 0x4b8  :    2 - 0x2 -- Sprite 0x97
    "00000011", -- 1209 - 0x4b9  :    3 - 0x3
    "11111110", -- 1210 - 0x4ba  :  254 - 0xfe
    "11111010", -- 1211 - 0x4bb  :  250 - 0xfa
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- Sprite 0x98
    "01000100", -- 1217 - 0x4c1  :   68 - 0x44
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "01000001", -- 1219 - 0x4c3  :   65 - 0x41
    "00100000", -- 1220 - 0x4c4  :   32 - 0x20
    "01001011", -- 1221 - 0x4c5  :   75 - 0x4b
    "00100111", -- 1222 - 0x4c6  :   39 - 0x27
    "00011111", -- 1223 - 0x4c7  :   31 - 0x1f
    "00001111", -- 1224 - 0x4c8  :   15 - 0xf -- Sprite 0x99
    "00011110", -- 1225 - 0x4c9  :   30 - 0x1e
    "00011111", -- 1226 - 0x4ca  :   31 - 0x1f
    "00011111", -- 1227 - 0x4cb  :   31 - 0x1f
    "00011111", -- 1228 - 0x4cc  :   31 - 0x1f
    "00001111", -- 1229 - 0x4cd  :   15 - 0xf
    "00001111", -- 1230 - 0x4ce  :   15 - 0xf
    "00000011", -- 1231 - 0x4cf  :    3 - 0x3
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Sprite 0x9a
    "00100000", -- 1233 - 0x4d1  :   32 - 0x20
    "01010000", -- 1234 - 0x4d2  :   80 - 0x50
    "00100000", -- 1235 - 0x4d3  :   32 - 0x20
    "01100000", -- 1236 - 0x4d4  :   96 - 0x60
    "01001000", -- 1237 - 0x4d5  :   72 - 0x48
    "11100000", -- 1238 - 0x4d6  :  224 - 0xe0
    "11110000", -- 1239 - 0x4d7  :  240 - 0xf0
    "11111000", -- 1240 - 0x4d8  :  248 - 0xf8 -- Sprite 0x9b
    "01111000", -- 1241 - 0x4d9  :  120 - 0x78
    "00111100", -- 1242 - 0x4da  :   60 - 0x3c
    "00111100", -- 1243 - 0x4db  :   60 - 0x3c
    "00111100", -- 1244 - 0x4dc  :   60 - 0x3c
    "11111100", -- 1245 - 0x4dd  :  252 - 0xfc
    "11111000", -- 1246 - 0x4de  :  248 - 0xf8
    "11100000", -- 1247 - 0x4df  :  224 - 0xe0
    "00010000", -- 1248 - 0x4e0  :   16 - 0x10 -- Sprite 0x9c
    "00000001", -- 1249 - 0x4e1  :    1 - 0x1
    "00101010", -- 1250 - 0x4e2  :   42 - 0x2a
    "00001100", -- 1251 - 0x4e3  :   12 - 0xc
    "10100110", -- 1252 - 0x4e4  :  166 - 0xa6
    "00010111", -- 1253 - 0x4e5  :   23 - 0x17
    "00011111", -- 1254 - 0x4e6  :   31 - 0x1f
    "00011111", -- 1255 - 0x4e7  :   31 - 0x1f
    "01011110", -- 1256 - 0x4e8  :   94 - 0x5e -- Sprite 0x9d
    "00111100", -- 1257 - 0x4e9  :   60 - 0x3c
    "00111101", -- 1258 - 0x4ea  :   61 - 0x3d
    "00111101", -- 1259 - 0x4eb  :   61 - 0x3d
    "00111110", -- 1260 - 0x4ec  :   62 - 0x3e
    "00011111", -- 1261 - 0x4ed  :   31 - 0x1f
    "00001111", -- 1262 - 0x4ee  :   15 - 0xf
    "00000111", -- 1263 - 0x4ef  :    7 - 0x7
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0 -- Sprite 0x9e
    "00000000", -- 1265 - 0x4f1  :    0 - 0x0
    "10000000", -- 1266 - 0x4f2  :  128 - 0x80
    "11001000", -- 1267 - 0x4f3  :  200 - 0xc8
    "01100000", -- 1268 - 0x4f4  :   96 - 0x60
    "11100000", -- 1269 - 0x4f5  :  224 - 0xe0
    "11110100", -- 1270 - 0x4f6  :  244 - 0xf4
    "11111000", -- 1271 - 0x4f7  :  248 - 0xf8
    "01111100", -- 1272 - 0x4f8  :  124 - 0x7c -- Sprite 0x9f
    "00011100", -- 1273 - 0x4f9  :   28 - 0x1c
    "00101110", -- 1274 - 0x4fa  :   46 - 0x2e
    "00101110", -- 1275 - 0x4fb  :   46 - 0x2e
    "00011110", -- 1276 - 0x4fc  :   30 - 0x1e
    "11111100", -- 1277 - 0x4fd  :  252 - 0xfc
    "11111000", -- 1278 - 0x4fe  :  248 - 0xf8
    "11100000", -- 1279 - 0x4ff  :  224 - 0xe0
    "11111111", -- 1280 - 0x500  :  255 - 0xff -- Sprite 0xa0
    "11111111", -- 1281 - 0x501  :  255 - 0xff
    "00111000", -- 1282 - 0x502  :   56 - 0x38
    "01101100", -- 1283 - 0x503  :  108 - 0x6c
    "11000110", -- 1284 - 0x504  :  198 - 0xc6
    "10000011", -- 1285 - 0x505  :  131 - 0x83
    "11111111", -- 1286 - 0x506  :  255 - 0xff
    "11111111", -- 1287 - 0x507  :  255 - 0xff
    "11111111", -- 1288 - 0x508  :  255 - 0xff -- Sprite 0xa1
    "11111111", -- 1289 - 0x509  :  255 - 0xff
    "00111000", -- 1290 - 0x50a  :   56 - 0x38
    "01101100", -- 1291 - 0x50b  :  108 - 0x6c
    "11000110", -- 1292 - 0x50c  :  198 - 0xc6
    "10000011", -- 1293 - 0x50d  :  131 - 0x83
    "11111111", -- 1294 - 0x50e  :  255 - 0xff
    "11111111", -- 1295 - 0x50f  :  255 - 0xff
    "10010010", -- 1296 - 0x510  :  146 - 0x92 -- Sprite 0xa2
    "01010100", -- 1297 - 0x511  :   84 - 0x54
    "00111000", -- 1298 - 0x512  :   56 - 0x38
    "11111110", -- 1299 - 0x513  :  254 - 0xfe
    "00111000", -- 1300 - 0x514  :   56 - 0x38
    "01010100", -- 1301 - 0x515  :   84 - 0x54
    "10010010", -- 1302 - 0x516  :  146 - 0x92
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "11111111", -- 1304 - 0x518  :  255 - 0xff -- Sprite 0xa3
    "11111111", -- 1305 - 0x519  :  255 - 0xff
    "11111111", -- 1306 - 0x51a  :  255 - 0xff
    "11111111", -- 1307 - 0x51b  :  255 - 0xff
    "11111111", -- 1308 - 0x51c  :  255 - 0xff
    "11111111", -- 1309 - 0x51d  :  255 - 0xff
    "11111111", -- 1310 - 0x51e  :  255 - 0xff
    "11111111", -- 1311 - 0x51f  :  255 - 0xff
    "11111111", -- 1312 - 0x520  :  255 - 0xff -- Sprite 0xa4
    "11111111", -- 1313 - 0x521  :  255 - 0xff
    "11111111", -- 1314 - 0x522  :  255 - 0xff
    "11111111", -- 1315 - 0x523  :  255 - 0xff
    "11111111", -- 1316 - 0x524  :  255 - 0xff
    "11111111", -- 1317 - 0x525  :  255 - 0xff
    "11111111", -- 1318 - 0x526  :  255 - 0xff
    "11111111", -- 1319 - 0x527  :  255 - 0xff
    "11111111", -- 1320 - 0x528  :  255 - 0xff -- Sprite 0xa5
    "11111111", -- 1321 - 0x529  :  255 - 0xff
    "11111111", -- 1322 - 0x52a  :  255 - 0xff
    "11111111", -- 1323 - 0x52b  :  255 - 0xff
    "11111111", -- 1324 - 0x52c  :  255 - 0xff
    "11111111", -- 1325 - 0x52d  :  255 - 0xff
    "11111111", -- 1326 - 0x52e  :  255 - 0xff
    "11111111", -- 1327 - 0x52f  :  255 - 0xff
    "11111111", -- 1328 - 0x530  :  255 - 0xff -- Sprite 0xa6
    "11111111", -- 1329 - 0x531  :  255 - 0xff
    "11111111", -- 1330 - 0x532  :  255 - 0xff
    "11111111", -- 1331 - 0x533  :  255 - 0xff
    "11111111", -- 1332 - 0x534  :  255 - 0xff
    "11111111", -- 1333 - 0x535  :  255 - 0xff
    "11111111", -- 1334 - 0x536  :  255 - 0xff
    "11111111", -- 1335 - 0x537  :  255 - 0xff
    "11111111", -- 1336 - 0x538  :  255 - 0xff -- Sprite 0xa7
    "11111111", -- 1337 - 0x539  :  255 - 0xff
    "11111111", -- 1338 - 0x53a  :  255 - 0xff
    "11111111", -- 1339 - 0x53b  :  255 - 0xff
    "11111111", -- 1340 - 0x53c  :  255 - 0xff
    "11111111", -- 1341 - 0x53d  :  255 - 0xff
    "11111111", -- 1342 - 0x53e  :  255 - 0xff
    "11111111", -- 1343 - 0x53f  :  255 - 0xff
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Sprite 0xa8
    "00000000", -- 1345 - 0x541  :    0 - 0x0
    "00000000", -- 1346 - 0x542  :    0 - 0x0
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00100011", -- 1349 - 0x545  :   35 - 0x23
    "10010111", -- 1350 - 0x546  :  151 - 0x97
    "00101111", -- 1351 - 0x547  :   47 - 0x2f
    "01101110", -- 1352 - 0x548  :  110 - 0x6e -- Sprite 0xa9
    "11101111", -- 1353 - 0x549  :  239 - 0xef
    "11110111", -- 1354 - 0x54a  :  247 - 0xf7
    "11111111", -- 1355 - 0x54b  :  255 - 0xff
    "01111111", -- 1356 - 0x54c  :  127 - 0x7f
    "00111111", -- 1357 - 0x54d  :   63 - 0x3f
    "01011111", -- 1358 - 0x54e  :   95 - 0x5f
    "00001111", -- 1359 - 0x54f  :   15 - 0xf
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0xaa
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "11111000", -- 1364 - 0x554  :  248 - 0xf8
    "11111100", -- 1365 - 0x555  :  252 - 0xfc
    "11111110", -- 1366 - 0x556  :  254 - 0xfe
    "01011110", -- 1367 - 0x557  :   94 - 0x5e
    "01011110", -- 1368 - 0x558  :   94 - 0x5e -- Sprite 0xab
    "00001100", -- 1369 - 0x559  :   12 - 0xc
    "10011110", -- 1370 - 0x55a  :  158 - 0x9e
    "11111110", -- 1371 - 0x55b  :  254 - 0xfe
    "11111110", -- 1372 - 0x55c  :  254 - 0xfe
    "11111110", -- 1373 - 0x55d  :  254 - 0xfe
    "11111000", -- 1374 - 0x55e  :  248 - 0xf8
    "11000000", -- 1375 - 0x55f  :  192 - 0xc0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Sprite 0xac
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "00000000", -- 1380 - 0x564  :    0 - 0x0
    "00000011", -- 1381 - 0x565  :    3 - 0x3
    "00000111", -- 1382 - 0x566  :    7 - 0x7
    "00101111", -- 1383 - 0x567  :   47 - 0x2f
    "01001110", -- 1384 - 0x568  :   78 - 0x4e -- Sprite 0xad
    "01101110", -- 1385 - 0x569  :  110 - 0x6e
    "11111110", -- 1386 - 0x56a  :  254 - 0xfe
    "01111111", -- 1387 - 0x56b  :  127 - 0x7f
    "00111111", -- 1388 - 0x56c  :   63 - 0x3f
    "00011111", -- 1389 - 0x56d  :   31 - 0x1f
    "00001111", -- 1390 - 0x56e  :   15 - 0xf
    "00000011", -- 1391 - 0x56f  :    3 - 0x3
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0xae
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "11111000", -- 1396 - 0x574  :  248 - 0xf8
    "11111100", -- 1397 - 0x575  :  252 - 0xfc
    "11111110", -- 1398 - 0x576  :  254 - 0xfe
    "01010110", -- 1399 - 0x577  :   86 - 0x56
    "01010110", -- 1400 - 0x578  :   86 - 0x56 -- Sprite 0xaf
    "00001100", -- 1401 - 0x579  :   12 - 0xc
    "00001110", -- 1402 - 0x57a  :   14 - 0xe
    "00011111", -- 1403 - 0x57b  :   31 - 0x1f
    "11111111", -- 1404 - 0x57c  :  255 - 0xff
    "11111111", -- 1405 - 0x57d  :  255 - 0xff
    "11111110", -- 1406 - 0x57e  :  254 - 0xfe
    "11111000", -- 1407 - 0x57f  :  248 - 0xf8
    "11111111", -- 1408 - 0x580  :  255 - 0xff -- Sprite 0xb0
    "11111111", -- 1409 - 0x581  :  255 - 0xff
    "11111111", -- 1410 - 0x582  :  255 - 0xff
    "11111111", -- 1411 - 0x583  :  255 - 0xff
    "11111111", -- 1412 - 0x584  :  255 - 0xff
    "11111111", -- 1413 - 0x585  :  255 - 0xff
    "11111111", -- 1414 - 0x586  :  255 - 0xff
    "11111111", -- 1415 - 0x587  :  255 - 0xff
    "11111111", -- 1416 - 0x588  :  255 - 0xff -- Sprite 0xb1
    "11111111", -- 1417 - 0x589  :  255 - 0xff
    "11111111", -- 1418 - 0x58a  :  255 - 0xff
    "11111111", -- 1419 - 0x58b  :  255 - 0xff
    "11111111", -- 1420 - 0x58c  :  255 - 0xff
    "11111111", -- 1421 - 0x58d  :  255 - 0xff
    "11111111", -- 1422 - 0x58e  :  255 - 0xff
    "11111111", -- 1423 - 0x58f  :  255 - 0xff
    "11111111", -- 1424 - 0x590  :  255 - 0xff -- Sprite 0xb2
    "11111111", -- 1425 - 0x591  :  255 - 0xff
    "11111111", -- 1426 - 0x592  :  255 - 0xff
    "11111111", -- 1427 - 0x593  :  255 - 0xff
    "11111111", -- 1428 - 0x594  :  255 - 0xff
    "11111111", -- 1429 - 0x595  :  255 - 0xff
    "11111111", -- 1430 - 0x596  :  255 - 0xff
    "11111111", -- 1431 - 0x597  :  255 - 0xff
    "11111111", -- 1432 - 0x598  :  255 - 0xff -- Sprite 0xb3
    "11111111", -- 1433 - 0x599  :  255 - 0xff
    "11111111", -- 1434 - 0x59a  :  255 - 0xff
    "11111111", -- 1435 - 0x59b  :  255 - 0xff
    "11111111", -- 1436 - 0x59c  :  255 - 0xff
    "11111111", -- 1437 - 0x59d  :  255 - 0xff
    "11111111", -- 1438 - 0x59e  :  255 - 0xff
    "11111111", -- 1439 - 0x59f  :  255 - 0xff
    "11111111", -- 1440 - 0x5a0  :  255 - 0xff -- Sprite 0xb4
    "11111111", -- 1441 - 0x5a1  :  255 - 0xff
    "11111111", -- 1442 - 0x5a2  :  255 - 0xff
    "11111111", -- 1443 - 0x5a3  :  255 - 0xff
    "11111111", -- 1444 - 0x5a4  :  255 - 0xff
    "11111111", -- 1445 - 0x5a5  :  255 - 0xff
    "11111111", -- 1446 - 0x5a6  :  255 - 0xff
    "11111111", -- 1447 - 0x5a7  :  255 - 0xff
    "11111111", -- 1448 - 0x5a8  :  255 - 0xff -- Sprite 0xb5
    "11111111", -- 1449 - 0x5a9  :  255 - 0xff
    "11111111", -- 1450 - 0x5aa  :  255 - 0xff
    "11111111", -- 1451 - 0x5ab  :  255 - 0xff
    "11111111", -- 1452 - 0x5ac  :  255 - 0xff
    "11111111", -- 1453 - 0x5ad  :  255 - 0xff
    "11111111", -- 1454 - 0x5ae  :  255 - 0xff
    "11111111", -- 1455 - 0x5af  :  255 - 0xff
    "11111111", -- 1456 - 0x5b0  :  255 - 0xff -- Sprite 0xb6
    "11111111", -- 1457 - 0x5b1  :  255 - 0xff
    "11111111", -- 1458 - 0x5b2  :  255 - 0xff
    "11111111", -- 1459 - 0x5b3  :  255 - 0xff
    "11111111", -- 1460 - 0x5b4  :  255 - 0xff
    "11111111", -- 1461 - 0x5b5  :  255 - 0xff
    "11111111", -- 1462 - 0x5b6  :  255 - 0xff
    "11111111", -- 1463 - 0x5b7  :  255 - 0xff
    "11111111", -- 1464 - 0x5b8  :  255 - 0xff -- Sprite 0xb7
    "11111111", -- 1465 - 0x5b9  :  255 - 0xff
    "11111111", -- 1466 - 0x5ba  :  255 - 0xff
    "11111111", -- 1467 - 0x5bb  :  255 - 0xff
    "11111111", -- 1468 - 0x5bc  :  255 - 0xff
    "11111111", -- 1469 - 0x5bd  :  255 - 0xff
    "11111111", -- 1470 - 0x5be  :  255 - 0xff
    "11111111", -- 1471 - 0x5bf  :  255 - 0xff
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Sprite 0xb8
    "00000111", -- 1473 - 0x5c1  :    7 - 0x7
    "00001000", -- 1474 - 0x5c2  :    8 - 0x8
    "00010000", -- 1475 - 0x5c3  :   16 - 0x10
    "00010000", -- 1476 - 0x5c4  :   16 - 0x10
    "00100000", -- 1477 - 0x5c5  :   32 - 0x20
    "00100000", -- 1478 - 0x5c6  :   32 - 0x20
    "00100000", -- 1479 - 0x5c7  :   32 - 0x20
    "00011111", -- 1480 - 0x5c8  :   31 - 0x1f -- Sprite 0xb9
    "00101111", -- 1481 - 0x5c9  :   47 - 0x2f
    "00110111", -- 1482 - 0x5ca  :   55 - 0x37
    "00111010", -- 1483 - 0x5cb  :   58 - 0x3a
    "00111101", -- 1484 - 0x5cc  :   61 - 0x3d
    "00111110", -- 1485 - 0x5cd  :   62 - 0x3e
    "00111111", -- 1486 - 0x5ce  :   63 - 0x3f
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Sprite 0xba
    "00000101", -- 1489 - 0x5d1  :    5 - 0x5
    "00011001", -- 1490 - 0x5d2  :   25 - 0x19
    "00110011", -- 1491 - 0x5d3  :   51 - 0x33
    "01100011", -- 1492 - 0x5d4  :   99 - 0x63
    "11000111", -- 1493 - 0x5d5  :  199 - 0xc7
    "11000111", -- 1494 - 0x5d6  :  199 - 0xc7
    "11000100", -- 1495 - 0x5d7  :  196 - 0xc4
    "10000000", -- 1496 - 0x5d8  :  128 - 0x80 -- Sprite 0xbb
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000011", -- 1501 - 0x5dd  :    3 - 0x3
    "00000011", -- 1502 - 0x5de  :    3 - 0x3
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Sprite 0xbc
    "00000000", -- 1505 - 0x5e1  :    0 - 0x0
    "00000000", -- 1506 - 0x5e2  :    0 - 0x0
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "00000000", -- 1508 - 0x5e4  :    0 - 0x0
    "00000000", -- 1509 - 0x5e5  :    0 - 0x0
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- Sprite 0xbd
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00001111", -- 1514 - 0x5ea  :   15 - 0xf
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "10000000", -- 1516 - 0x5ec  :  128 - 0x80
    "01100011", -- 1517 - 0x5ed  :   99 - 0x63
    "00011110", -- 1518 - 0x5ee  :   30 - 0x1e
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000001", -- 1520 - 0x5f0  :    1 - 0x1 -- Sprite 0xbe
    "00000011", -- 1521 - 0x5f1  :    3 - 0x3
    "00011001", -- 1522 - 0x5f2  :   25 - 0x19
    "00111100", -- 1523 - 0x5f3  :   60 - 0x3c
    "00011001", -- 1524 - 0x5f4  :   25 - 0x19
    "00100011", -- 1525 - 0x5f5  :   35 - 0x23
    "01010001", -- 1526 - 0x5f6  :   81 - 0x51
    "00100000", -- 1527 - 0x5f7  :   32 - 0x20
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Sprite 0xbf
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0xc0
    "00111111", -- 1537 - 0x601  :   63 - 0x3f
    "00011111", -- 1538 - 0x602  :   31 - 0x1f
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000001", -- 1540 - 0x604  :    1 - 0x1
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000001", -- 1542 - 0x606  :    1 - 0x1
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00010001", -- 1544 - 0x608  :   17 - 0x11 -- Sprite 0xc1
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000001", -- 1546 - 0x60a  :    1 - 0x1
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000001", -- 1548 - 0x60c  :    1 - 0x1
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00011111", -- 1550 - 0x60e  :   31 - 0x1f
    "00111111", -- 1551 - 0x60f  :   63 - 0x3f
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0xc2
    "11111100", -- 1553 - 0x611  :  252 - 0xfc
    "11111000", -- 1554 - 0x612  :  248 - 0xf8
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "10000000", -- 1556 - 0x614  :  128 - 0x80
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "10000000", -- 1558 - 0x616  :  128 - 0x80
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "10001000", -- 1560 - 0x618  :  136 - 0x88 -- Sprite 0xc3
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "10000000", -- 1562 - 0x61a  :  128 - 0x80
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "10000000", -- 1564 - 0x61c  :  128 - 0x80
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "11111000", -- 1566 - 0x61e  :  248 - 0xf8
    "11111100", -- 1567 - 0x61f  :  252 - 0xfc
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00111111", -- 1573 - 0x625  :   63 - 0x3f
    "00011111", -- 1574 - 0x626  :   31 - 0x1f
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000001", -- 1576 - 0x628  :    1 - 0x1 -- Sprite 0xc5
    "00000001", -- 1577 - 0x629  :    1 - 0x1
    "01000001", -- 1578 - 0x62a  :   65 - 0x41
    "00000001", -- 1579 - 0x62b  :    1 - 0x1
    "00000001", -- 1580 - 0x62c  :    1 - 0x1
    "00000000", -- 1581 - 0x62d  :    0 - 0x0
    "00011111", -- 1582 - 0x62e  :   31 - 0x1f
    "00111111", -- 1583 - 0x62f  :   63 - 0x3f
    "00000000", -- 1584 - 0x630  :    0 - 0x0 -- Sprite 0xc6
    "00000000", -- 1585 - 0x631  :    0 - 0x0
    "00000000", -- 1586 - 0x632  :    0 - 0x0
    "00000000", -- 1587 - 0x633  :    0 - 0x0
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "11111100", -- 1589 - 0x635  :  252 - 0xfc
    "11111000", -- 1590 - 0x636  :  248 - 0xf8
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "10000000", -- 1592 - 0x638  :  128 - 0x80 -- Sprite 0xc7
    "10000000", -- 1593 - 0x639  :  128 - 0x80
    "10000010", -- 1594 - 0x63a  :  130 - 0x82
    "10000000", -- 1595 - 0x63b  :  128 - 0x80
    "10000000", -- 1596 - 0x63c  :  128 - 0x80
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "11111000", -- 1598 - 0x63e  :  248 - 0xf8
    "11111100", -- 1599 - 0x63f  :  252 - 0xfc
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0xc8
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00011110", -- 1603 - 0x643  :   30 - 0x1e
    "00111111", -- 1604 - 0x644  :   63 - 0x3f
    "00111111", -- 1605 - 0x645  :   63 - 0x3f
    "00111111", -- 1606 - 0x646  :   63 - 0x3f
    "00111111", -- 1607 - 0x647  :   63 - 0x3f
    "00011111", -- 1608 - 0x648  :   31 - 0x1f -- Sprite 0xc9
    "00001111", -- 1609 - 0x649  :   15 - 0xf
    "00000111", -- 1610 - 0x64a  :    7 - 0x7
    "00000011", -- 1611 - 0x64b  :    3 - 0x3
    "00000001", -- 1612 - 0x64c  :    1 - 0x1
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0xca
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00111100", -- 1619 - 0x653  :   60 - 0x3c
    "01111110", -- 1620 - 0x654  :  126 - 0x7e
    "11111110", -- 1621 - 0x655  :  254 - 0xfe
    "11111110", -- 1622 - 0x656  :  254 - 0xfe
    "11111110", -- 1623 - 0x657  :  254 - 0xfe
    "11111100", -- 1624 - 0x658  :  252 - 0xfc -- Sprite 0xcb
    "11111000", -- 1625 - 0x659  :  248 - 0xf8
    "11110000", -- 1626 - 0x65a  :  240 - 0xf0
    "11100000", -- 1627 - 0x65b  :  224 - 0xe0
    "11000000", -- 1628 - 0x65c  :  192 - 0xc0
    "10000000", -- 1629 - 0x65d  :  128 - 0x80
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "11111111", -- 1632 - 0x660  :  255 - 0xff -- Sprite 0xcc
    "11111111", -- 1633 - 0x661  :  255 - 0xff
    "11111111", -- 1634 - 0x662  :  255 - 0xff
    "11111111", -- 1635 - 0x663  :  255 - 0xff
    "11111111", -- 1636 - 0x664  :  255 - 0xff
    "11111111", -- 1637 - 0x665  :  255 - 0xff
    "11111111", -- 1638 - 0x666  :  255 - 0xff
    "11111111", -- 1639 - 0x667  :  255 - 0xff
    "11111111", -- 1640 - 0x668  :  255 - 0xff -- Sprite 0xcd
    "11111111", -- 1641 - 0x669  :  255 - 0xff
    "11111111", -- 1642 - 0x66a  :  255 - 0xff
    "11111111", -- 1643 - 0x66b  :  255 - 0xff
    "11111111", -- 1644 - 0x66c  :  255 - 0xff
    "11111111", -- 1645 - 0x66d  :  255 - 0xff
    "11111111", -- 1646 - 0x66e  :  255 - 0xff
    "11111111", -- 1647 - 0x66f  :  255 - 0xff
    "11111111", -- 1648 - 0x670  :  255 - 0xff -- Sprite 0xce
    "11111111", -- 1649 - 0x671  :  255 - 0xff
    "11111111", -- 1650 - 0x672  :  255 - 0xff
    "11111111", -- 1651 - 0x673  :  255 - 0xff
    "11111111", -- 1652 - 0x674  :  255 - 0xff
    "11111111", -- 1653 - 0x675  :  255 - 0xff
    "11111111", -- 1654 - 0x676  :  255 - 0xff
    "11111111", -- 1655 - 0x677  :  255 - 0xff
    "11111111", -- 1656 - 0x678  :  255 - 0xff -- Sprite 0xcf
    "11111111", -- 1657 - 0x679  :  255 - 0xff
    "11111111", -- 1658 - 0x67a  :  255 - 0xff
    "11111111", -- 1659 - 0x67b  :  255 - 0xff
    "11111111", -- 1660 - 0x67c  :  255 - 0xff
    "11111111", -- 1661 - 0x67d  :  255 - 0xff
    "11111111", -- 1662 - 0x67e  :  255 - 0xff
    "11111111", -- 1663 - 0x67f  :  255 - 0xff
    "00001000", -- 1664 - 0x680  :    8 - 0x8 -- Sprite 0xd0
    "00011001", -- 1665 - 0x681  :   25 - 0x19
    "00001001", -- 1666 - 0x682  :    9 - 0x9
    "00001001", -- 1667 - 0x683  :    9 - 0x9
    "00001001", -- 1668 - 0x684  :    9 - 0x9
    "00001001", -- 1669 - 0x685  :    9 - 0x9
    "00011100", -- 1670 - 0x686  :   28 - 0x1c
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00111000", -- 1672 - 0x688  :   56 - 0x38 -- Sprite 0xd1
    "00000101", -- 1673 - 0x689  :    5 - 0x5
    "00000101", -- 1674 - 0x68a  :    5 - 0x5
    "00011001", -- 1675 - 0x68b  :   25 - 0x19
    "00000101", -- 1676 - 0x68c  :    5 - 0x5
    "00000101", -- 1677 - 0x68d  :    5 - 0x5
    "00111000", -- 1678 - 0x68e  :   56 - 0x38
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00111100", -- 1680 - 0x690  :   60 - 0x3c -- Sprite 0xd2
    "00100001", -- 1681 - 0x691  :   33 - 0x21
    "00100001", -- 1682 - 0x692  :   33 - 0x21
    "00111101", -- 1683 - 0x693  :   61 - 0x3d
    "00000101", -- 1684 - 0x694  :    5 - 0x5
    "00000101", -- 1685 - 0x695  :    5 - 0x5
    "00111000", -- 1686 - 0x696  :   56 - 0x38
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00011000", -- 1688 - 0x698  :   24 - 0x18 -- Sprite 0xd3
    "00100101", -- 1689 - 0x699  :   37 - 0x25
    "00100101", -- 1690 - 0x69a  :   37 - 0x25
    "00011001", -- 1691 - 0x69b  :   25 - 0x19
    "00100101", -- 1692 - 0x69c  :   37 - 0x25
    "00100101", -- 1693 - 0x69d  :   37 - 0x25
    "00011000", -- 1694 - 0x69e  :   24 - 0x18
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "11000110", -- 1696 - 0x6a0  :  198 - 0xc6 -- Sprite 0xd4
    "00101001", -- 1697 - 0x6a1  :   41 - 0x29
    "00101001", -- 1698 - 0x6a2  :   41 - 0x29
    "00101001", -- 1699 - 0x6a3  :   41 - 0x29
    "00101001", -- 1700 - 0x6a4  :   41 - 0x29
    "00101001", -- 1701 - 0x6a5  :   41 - 0x29
    "11000110", -- 1702 - 0x6a6  :  198 - 0xc6
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0 -- Sprite 0xd5
    "00000000", -- 1705 - 0x6a9  :    0 - 0x0
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "00000000", -- 1715 - 0x6b3  :    0 - 0x0
    "00111100", -- 1716 - 0x6b4  :   60 - 0x3c
    "10110110", -- 1717 - 0x6b5  :  182 - 0xb6
    "01111100", -- 1718 - 0x6b6  :  124 - 0x7c
    "11111000", -- 1719 - 0x6b7  :  248 - 0xf8
    "00000011", -- 1720 - 0x6b8  :    3 - 0x3 -- Sprite 0xd7
    "00000011", -- 1721 - 0x6b9  :    3 - 0x3
    "00000011", -- 1722 - 0x6ba  :    3 - 0x3
    "00000111", -- 1723 - 0x6bb  :    7 - 0x7
    "00001100", -- 1724 - 0x6bc  :   12 - 0xc
    "00011011", -- 1725 - 0x6bd  :   27 - 0x1b
    "01110111", -- 1726 - 0x6be  :  119 - 0x77
    "00000111", -- 1727 - 0x6bf  :    7 - 0x7
    "00001111", -- 1728 - 0x6c0  :   15 - 0xf -- Sprite 0xd8
    "00001111", -- 1729 - 0x6c1  :   15 - 0xf
    "00011111", -- 1730 - 0x6c2  :   31 - 0x1f
    "00111111", -- 1731 - 0x6c3  :   63 - 0x3f
    "01111111", -- 1732 - 0x6c4  :  127 - 0x7f
    "00111111", -- 1733 - 0x6c5  :   63 - 0x3f
    "00000000", -- 1734 - 0x6c6  :    0 - 0x0
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "11100000", -- 1736 - 0x6c8  :  224 - 0xe0 -- Sprite 0xd9
    "11110000", -- 1737 - 0x6c9  :  240 - 0xf0
    "11110000", -- 1738 - 0x6ca  :  240 - 0xf0
    "11110000", -- 1739 - 0x6cb  :  240 - 0xf0
    "00011000", -- 1740 - 0x6cc  :   24 - 0x18
    "11111100", -- 1741 - 0x6cd  :  252 - 0xfc
    "11111100", -- 1742 - 0x6ce  :  252 - 0xfc
    "11111100", -- 1743 - 0x6cf  :  252 - 0xfc
    "11111000", -- 1744 - 0x6d0  :  248 - 0xf8 -- Sprite 0xda
    "11111100", -- 1745 - 0x6d1  :  252 - 0xfc
    "11111111", -- 1746 - 0x6d2  :  255 - 0xff
    "11111111", -- 1747 - 0x6d3  :  255 - 0xff
    "11111110", -- 1748 - 0x6d4  :  254 - 0xfe
    "11110000", -- 1749 - 0x6d5  :  240 - 0xf0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000011", -- 1752 - 0x6d8  :    3 - 0x3 -- Sprite 0xdb
    "00000011", -- 1753 - 0x6d9  :    3 - 0x3
    "00000011", -- 1754 - 0x6da  :    3 - 0x3
    "00000011", -- 1755 - 0x6db  :    3 - 0x3
    "00000001", -- 1756 - 0x6dc  :    1 - 0x1
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000111", -- 1758 - 0x6de  :    7 - 0x7
    "00011111", -- 1759 - 0x6df  :   31 - 0x1f
    "11111111", -- 1760 - 0x6e0  :  255 - 0xff -- Sprite 0xdc
    "11111111", -- 1761 - 0x6e1  :  255 - 0xff
    "01111111", -- 1762 - 0x6e2  :  127 - 0x7f
    "00111111", -- 1763 - 0x6e3  :   63 - 0x3f
    "00001111", -- 1764 - 0x6e4  :   15 - 0xf
    "00000011", -- 1765 - 0x6e5  :    3 - 0x3
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "11100000", -- 1768 - 0x6e8  :  224 - 0xe0 -- Sprite 0xdd
    "11110000", -- 1769 - 0x6e9  :  240 - 0xf0
    "11110000", -- 1770 - 0x6ea  :  240 - 0xf0
    "11100000", -- 1771 - 0x6eb  :  224 - 0xe0
    "11111110", -- 1772 - 0x6ec  :  254 - 0xfe
    "00111100", -- 1773 - 0x6ed  :   60 - 0x3c
    "11110000", -- 1774 - 0x6ee  :  240 - 0xf0
    "11111100", -- 1775 - 0x6ef  :  252 - 0xfc
    "11111100", -- 1776 - 0x6f0  :  252 - 0xfc -- Sprite 0xde
    "11111000", -- 1777 - 0x6f1  :  248 - 0xf8
    "11111000", -- 1778 - 0x6f2  :  248 - 0xf8
    "11111000", -- 1779 - 0x6f3  :  248 - 0xf8
    "11111000", -- 1780 - 0x6f4  :  248 - 0xf8
    "11111000", -- 1781 - 0x6f5  :  248 - 0xf8
    "11111000", -- 1782 - 0x6f6  :  248 - 0xf8
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "11111111", -- 1784 - 0x6f8  :  255 - 0xff -- Sprite 0xdf
    "11111111", -- 1785 - 0x6f9  :  255 - 0xff
    "11111111", -- 1786 - 0x6fa  :  255 - 0xff
    "11111111", -- 1787 - 0x6fb  :  255 - 0xff
    "11111111", -- 1788 - 0x6fc  :  255 - 0xff
    "11111111", -- 1789 - 0x6fd  :  255 - 0xff
    "11111111", -- 1790 - 0x6fe  :  255 - 0xff
    "11111111", -- 1791 - 0x6ff  :  255 - 0xff
    "11111111", -- 1792 - 0x700  :  255 - 0xff -- Sprite 0xe0
    "11111111", -- 1793 - 0x701  :  255 - 0xff
    "11111111", -- 1794 - 0x702  :  255 - 0xff
    "11111111", -- 1795 - 0x703  :  255 - 0xff
    "11111111", -- 1796 - 0x704  :  255 - 0xff
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "11111111", -- 1798 - 0x706  :  255 - 0xff
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "11111111", -- 1800 - 0x708  :  255 - 0xff -- Sprite 0xe1
    "11111111", -- 1801 - 0x709  :  255 - 0xff
    "11111111", -- 1802 - 0x70a  :  255 - 0xff
    "11111111", -- 1803 - 0x70b  :  255 - 0xff
    "11111111", -- 1804 - 0x70c  :  255 - 0xff
    "11111111", -- 1805 - 0x70d  :  255 - 0xff
    "11111111", -- 1806 - 0x70e  :  255 - 0xff
    "11111111", -- 1807 - 0x70f  :  255 - 0xff
    "11111111", -- 1808 - 0x710  :  255 - 0xff -- Sprite 0xe2
    "11111111", -- 1809 - 0x711  :  255 - 0xff
    "11111111", -- 1810 - 0x712  :  255 - 0xff
    "11111111", -- 1811 - 0x713  :  255 - 0xff
    "11111111", -- 1812 - 0x714  :  255 - 0xff
    "11111111", -- 1813 - 0x715  :  255 - 0xff
    "11111111", -- 1814 - 0x716  :  255 - 0xff
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "11111111", -- 1816 - 0x718  :  255 - 0xff -- Sprite 0xe3
    "11111111", -- 1817 - 0x719  :  255 - 0xff
    "11111111", -- 1818 - 0x71a  :  255 - 0xff
    "11111111", -- 1819 - 0x71b  :  255 - 0xff
    "11111111", -- 1820 - 0x71c  :  255 - 0xff
    "11111111", -- 1821 - 0x71d  :  255 - 0xff
    "11111111", -- 1822 - 0x71e  :  255 - 0xff
    "11111111", -- 1823 - 0x71f  :  255 - 0xff
    "11111111", -- 1824 - 0x720  :  255 - 0xff -- Sprite 0xe4
    "11111111", -- 1825 - 0x721  :  255 - 0xff
    "11111111", -- 1826 - 0x722  :  255 - 0xff
    "11111111", -- 1827 - 0x723  :  255 - 0xff
    "11111111", -- 1828 - 0x724  :  255 - 0xff
    "11111111", -- 1829 - 0x725  :  255 - 0xff
    "11111111", -- 1830 - 0x726  :  255 - 0xff
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "11111111", -- 1832 - 0x728  :  255 - 0xff -- Sprite 0xe5
    "11111111", -- 1833 - 0x729  :  255 - 0xff
    "11111111", -- 1834 - 0x72a  :  255 - 0xff
    "11111111", -- 1835 - 0x72b  :  255 - 0xff
    "11111111", -- 1836 - 0x72c  :  255 - 0xff
    "11111111", -- 1837 - 0x72d  :  255 - 0xff
    "11111111", -- 1838 - 0x72e  :  255 - 0xff
    "11111111", -- 1839 - 0x72f  :  255 - 0xff
    "11111111", -- 1840 - 0x730  :  255 - 0xff -- Sprite 0xe6
    "11111111", -- 1841 - 0x731  :  255 - 0xff
    "11111111", -- 1842 - 0x732  :  255 - 0xff
    "11111111", -- 1843 - 0x733  :  255 - 0xff
    "11111111", -- 1844 - 0x734  :  255 - 0xff
    "11111111", -- 1845 - 0x735  :  255 - 0xff
    "11111111", -- 1846 - 0x736  :  255 - 0xff
    "11111111", -- 1847 - 0x737  :  255 - 0xff
    "11111111", -- 1848 - 0x738  :  255 - 0xff -- Sprite 0xe7
    "11111111", -- 1849 - 0x739  :  255 - 0xff
    "11111111", -- 1850 - 0x73a  :  255 - 0xff
    "11111111", -- 1851 - 0x73b  :  255 - 0xff
    "11111111", -- 1852 - 0x73c  :  255 - 0xff
    "11111111", -- 1853 - 0x73d  :  255 - 0xff
    "11111111", -- 1854 - 0x73e  :  255 - 0xff
    "11111111", -- 1855 - 0x73f  :  255 - 0xff
    "11111111", -- 1856 - 0x740  :  255 - 0xff -- Sprite 0xe8
    "11111111", -- 1857 - 0x741  :  255 - 0xff
    "11111111", -- 1858 - 0x742  :  255 - 0xff
    "11111111", -- 1859 - 0x743  :  255 - 0xff
    "11111111", -- 1860 - 0x744  :  255 - 0xff
    "11111111", -- 1861 - 0x745  :  255 - 0xff
    "11111111", -- 1862 - 0x746  :  255 - 0xff
    "11111111", -- 1863 - 0x747  :  255 - 0xff
    "11111111", -- 1864 - 0x748  :  255 - 0xff -- Sprite 0xe9
    "11111111", -- 1865 - 0x749  :  255 - 0xff
    "11111111", -- 1866 - 0x74a  :  255 - 0xff
    "11111111", -- 1867 - 0x74b  :  255 - 0xff
    "11111111", -- 1868 - 0x74c  :  255 - 0xff
    "11111111", -- 1869 - 0x74d  :  255 - 0xff
    "11111111", -- 1870 - 0x74e  :  255 - 0xff
    "11111111", -- 1871 - 0x74f  :  255 - 0xff
    "11111111", -- 1872 - 0x750  :  255 - 0xff -- Sprite 0xea
    "11111111", -- 1873 - 0x751  :  255 - 0xff
    "11111111", -- 1874 - 0x752  :  255 - 0xff
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "11111111", -- 1876 - 0x754  :  255 - 0xff
    "11111111", -- 1877 - 0x755  :  255 - 0xff
    "11111111", -- 1878 - 0x756  :  255 - 0xff
    "11111111", -- 1879 - 0x757  :  255 - 0xff
    "11111111", -- 1880 - 0x758  :  255 - 0xff -- Sprite 0xeb
    "11111111", -- 1881 - 0x759  :  255 - 0xff
    "11111111", -- 1882 - 0x75a  :  255 - 0xff
    "11111111", -- 1883 - 0x75b  :  255 - 0xff
    "11111111", -- 1884 - 0x75c  :  255 - 0xff
    "11111111", -- 1885 - 0x75d  :  255 - 0xff
    "11111111", -- 1886 - 0x75e  :  255 - 0xff
    "11111111", -- 1887 - 0x75f  :  255 - 0xff
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0xec
    "00000001", -- 1889 - 0x761  :    1 - 0x1
    "00000011", -- 1890 - 0x762  :    3 - 0x3
    "00110011", -- 1891 - 0x763  :   51 - 0x33
    "00011001", -- 1892 - 0x764  :   25 - 0x19
    "00001111", -- 1893 - 0x765  :   15 - 0xf
    "00111111", -- 1894 - 0x766  :   63 - 0x3f
    "00011111", -- 1895 - 0x767  :   31 - 0x1f
    "00101011", -- 1896 - 0x768  :   43 - 0x2b -- Sprite 0xed
    "00000111", -- 1897 - 0x769  :    7 - 0x7
    "00000101", -- 1898 - 0x76a  :    5 - 0x5
    "00001101", -- 1899 - 0x76b  :   13 - 0xd
    "00001011", -- 1900 - 0x76c  :   11 - 0xb
    "00011011", -- 1901 - 0x76d  :   27 - 0x1b
    "00011011", -- 1902 - 0x76e  :   27 - 0x1b
    "00111011", -- 1903 - 0x76f  :   59 - 0x3b
    "00001001", -- 1904 - 0x770  :    9 - 0x9 -- Sprite 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000111", -- 1906 - 0x772  :    7 - 0x7
    "00000111", -- 1907 - 0x773  :    7 - 0x7
    "00001111", -- 1908 - 0x774  :   15 - 0xf
    "00001101", -- 1909 - 0x775  :   13 - 0xd
    "00000001", -- 1910 - 0x776  :    1 - 0x1
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "11111000", -- 1912 - 0x778  :  248 - 0xf8 -- Sprite 0xef
    "11111100", -- 1913 - 0x779  :  252 - 0xfc
    "11111000", -- 1914 - 0x77a  :  248 - 0xf8
    "11101100", -- 1915 - 0x77b  :  236 - 0xec
    "11111000", -- 1916 - 0x77c  :  248 - 0xf8
    "11110000", -- 1917 - 0x77d  :  240 - 0xf0
    "11000000", -- 1918 - 0x77e  :  192 - 0xc0
    "11000000", -- 1919 - 0x77f  :  192 - 0xc0
    "11110000", -- 1920 - 0x780  :  240 - 0xf0 -- Sprite 0xf0
    "11111000", -- 1921 - 0x781  :  248 - 0xf8
    "11111000", -- 1922 - 0x782  :  248 - 0xf8
    "11101000", -- 1923 - 0x783  :  232 - 0xe8
    "11001100", -- 1924 - 0x784  :  204 - 0xcc
    "11100110", -- 1925 - 0x785  :  230 - 0xe6
    "11111011", -- 1926 - 0x786  :  251 - 0xfb
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11111111", -- 1928 - 0x788  :  255 - 0xff -- Sprite 0xf1
    "11111110", -- 1929 - 0x789  :  254 - 0xfe
    "11111110", -- 1930 - 0x78a  :  254 - 0xfe
    "11111110", -- 1931 - 0x78b  :  254 - 0xfe
    "11111110", -- 1932 - 0x78c  :  254 - 0xfe
    "10001111", -- 1933 - 0x78d  :  143 - 0x8f
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000001", -- 1936 - 0x790  :    1 - 0x1 -- Sprite 0xf2
    "00001111", -- 1937 - 0x791  :   15 - 0xf
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000100", -- 1940 - 0x794  :    4 - 0x4
    "00011110", -- 1941 - 0x795  :   30 - 0x1e
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000011", -- 1943 - 0x797  :    3 - 0x3
    "00000111", -- 1944 - 0x798  :    7 - 0x7 -- Sprite 0xf3
    "00001111", -- 1945 - 0x799  :   15 - 0xf
    "00011111", -- 1946 - 0x79a  :   31 - 0x1f
    "00001111", -- 1947 - 0x79b  :   15 - 0xf
    "00000111", -- 1948 - 0x79c  :    7 - 0x7
    "00001111", -- 1949 - 0x79d  :   15 - 0xf
    "00001111", -- 1950 - 0x79e  :   15 - 0xf
    "00000011", -- 1951 - 0x79f  :    3 - 0x3
    "11100000", -- 1952 - 0x7a0  :  224 - 0xe0 -- Sprite 0xf4
    "11110000", -- 1953 - 0x7a1  :  240 - 0xf0
    "11110000", -- 1954 - 0x7a2  :  240 - 0xf0
    "01001000", -- 1955 - 0x7a3  :   72 - 0x48
    "11001000", -- 1956 - 0x7a4  :  200 - 0xc8
    "10011100", -- 1957 - 0x7a5  :  156 - 0x9c
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "11110000", -- 1959 - 0x7a7  :  240 - 0xf0
    "11111000", -- 1960 - 0x7a8  :  248 - 0xf8 -- Sprite 0xf5
    "11111100", -- 1961 - 0x7a9  :  252 - 0xfc
    "11111100", -- 1962 - 0x7aa  :  252 - 0xfc
    "11111000", -- 1963 - 0x7ab  :  248 - 0xf8
    "11111000", -- 1964 - 0x7ac  :  248 - 0xf8
    "01111000", -- 1965 - 0x7ad  :  120 - 0x78
    "01110000", -- 1966 - 0x7ae  :  112 - 0x70
    "01100000", -- 1967 - 0x7af  :   96 - 0x60
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0xf6
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "01111100", -- 1970 - 0x7b2  :  124 - 0x7c
    "10001010", -- 1971 - 0x7b3  :  138 - 0x8a
    "11111110", -- 1972 - 0x7b4  :  254 - 0xfe
    "11111110", -- 1973 - 0x7b5  :  254 - 0xfe
    "11111110", -- 1974 - 0x7b6  :  254 - 0xfe
    "11111110", -- 1975 - 0x7b7  :  254 - 0xfe
    "11111110", -- 1976 - 0x7b8  :  254 - 0xfe -- Sprite 0xf7
    "01111100", -- 1977 - 0x7b9  :  124 - 0x7c
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000111", -- 1984 - 0x7c0  :    7 - 0x7 -- Sprite 0xf8
    "00001011", -- 1985 - 0x7c1  :   11 - 0xb
    "00001111", -- 1986 - 0x7c2  :   15 - 0xf
    "00001011", -- 1987 - 0x7c3  :   11 - 0xb
    "00001011", -- 1988 - 0x7c4  :   11 - 0xb
    "00001011", -- 1989 - 0x7c5  :   11 - 0xb
    "00001011", -- 1990 - 0x7c6  :   11 - 0xb
    "00000111", -- 1991 - 0x7c7  :    7 - 0x7
    "11000000", -- 1992 - 0x7c8  :  192 - 0xc0 -- Sprite 0xf9
    "11100000", -- 1993 - 0x7c9  :  224 - 0xe0
    "11100000", -- 1994 - 0x7ca  :  224 - 0xe0
    "11100000", -- 1995 - 0x7cb  :  224 - 0xe0
    "11100000", -- 1996 - 0x7cc  :  224 - 0xe0
    "11100000", -- 1997 - 0x7cd  :  224 - 0xe0
    "11100000", -- 1998 - 0x7ce  :  224 - 0xe0
    "11000000", -- 1999 - 0x7cf  :  192 - 0xc0
    "00000011", -- 2000 - 0x7d0  :    3 - 0x3 -- Sprite 0xfa
    "00000111", -- 2001 - 0x7d1  :    7 - 0x7
    "00000111", -- 2002 - 0x7d2  :    7 - 0x7
    "00000111", -- 2003 - 0x7d3  :    7 - 0x7
    "00000111", -- 2004 - 0x7d4  :    7 - 0x7
    "00000111", -- 2005 - 0x7d5  :    7 - 0x7
    "00000111", -- 2006 - 0x7d6  :    7 - 0x7
    "00000011", -- 2007 - 0x7d7  :    3 - 0x3
    "11100000", -- 2008 - 0x7d8  :  224 - 0xe0 -- Sprite 0xfb
    "11010000", -- 2009 - 0x7d9  :  208 - 0xd0
    "11010000", -- 2010 - 0x7da  :  208 - 0xd0
    "11010000", -- 2011 - 0x7db  :  208 - 0xd0
    "11010000", -- 2012 - 0x7dc  :  208 - 0xd0
    "11110000", -- 2013 - 0x7dd  :  240 - 0xf0
    "11010000", -- 2014 - 0x7de  :  208 - 0xd0
    "11100000", -- 2015 - 0x7df  :  224 - 0xe0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0xfc
    "00000001", -- 2017 - 0x7e1  :    1 - 0x1
    "00010011", -- 2018 - 0x7e2  :   19 - 0x13
    "00110111", -- 2019 - 0x7e3  :   55 - 0x37
    "00111011", -- 2020 - 0x7e4  :   59 - 0x3b
    "01110100", -- 2021 - 0x7e5  :  116 - 0x74
    "01111010", -- 2022 - 0x7e6  :  122 - 0x7a
    "00111110", -- 2023 - 0x7e7  :   62 - 0x3e
    "11011000", -- 2024 - 0x7e8  :  216 - 0xd8 -- Sprite 0xfd
    "10011000", -- 2025 - 0x7e9  :  152 - 0x98
    "10101000", -- 2026 - 0x7ea  :  168 - 0xa8
    "11011000", -- 2027 - 0x7eb  :  216 - 0xd8
    "11011010", -- 2028 - 0x7ec  :  218 - 0xda
    "01110100", -- 2029 - 0x7ed  :  116 - 0x74
    "00101000", -- 2030 - 0x7ee  :   40 - 0x28
    "11001000", -- 2031 - 0x7ef  :  200 - 0xc8
    "00001000", -- 2032 - 0x7f0  :    8 - 0x8 -- Sprite 0xfe
    "01011001", -- 2033 - 0x7f1  :   89 - 0x59
    "00110000", -- 2034 - 0x7f2  :   48 - 0x30
    "01110001", -- 2035 - 0x7f3  :  113 - 0x71
    "01111001", -- 2036 - 0x7f4  :  121 - 0x79
    "00101011", -- 2037 - 0x7f5  :   43 - 0x2b
    "00110110", -- 2038 - 0x7f6  :   54 - 0x36
    "00010110", -- 2039 - 0x7f7  :   22 - 0x16
    "11000110", -- 2040 - 0x7f8  :  198 - 0xc6 -- Sprite 0xff
    "11000100", -- 2041 - 0x7f9  :  196 - 0xc4
    "11001100", -- 2042 - 0x7fa  :  204 - 0xcc
    "11001100", -- 2043 - 0x7fb  :  204 - 0xcc
    "10111000", -- 2044 - 0x7fc  :  184 - 0xb8
    "01111100", -- 2045 - 0x7fd  :  124 - 0x7c
    "11101100", -- 2046 - 0x7fe  :  236 - 0xec
    "11001000", -- 2047 - 0x7ff  :  200 - 0xc8
          -- Background pattern Table
    "00111000", -- 2048 - 0x800  :   56 - 0x38 -- Background 0x0
    "01001100", -- 2049 - 0x801  :   76 - 0x4c
    "11000110", -- 2050 - 0x802  :  198 - 0xc6
    "11000110", -- 2051 - 0x803  :  198 - 0xc6
    "11000110", -- 2052 - 0x804  :  198 - 0xc6
    "01100100", -- 2053 - 0x805  :  100 - 0x64
    "00111000", -- 2054 - 0x806  :   56 - 0x38
    "00000000", -- 2055 - 0x807  :    0 - 0x0
    "00011000", -- 2056 - 0x808  :   24 - 0x18 -- Background 0x1
    "00111000", -- 2057 - 0x809  :   56 - 0x38
    "00011000", -- 2058 - 0x80a  :   24 - 0x18
    "00011000", -- 2059 - 0x80b  :   24 - 0x18
    "00011000", -- 2060 - 0x80c  :   24 - 0x18
    "00011000", -- 2061 - 0x80d  :   24 - 0x18
    "01111110", -- 2062 - 0x80e  :  126 - 0x7e
    "00000000", -- 2063 - 0x80f  :    0 - 0x0
    "01111100", -- 2064 - 0x810  :  124 - 0x7c -- Background 0x2
    "11000110", -- 2065 - 0x811  :  198 - 0xc6
    "00001110", -- 2066 - 0x812  :   14 - 0xe
    "00111100", -- 2067 - 0x813  :   60 - 0x3c
    "01111000", -- 2068 - 0x814  :  120 - 0x78
    "11100000", -- 2069 - 0x815  :  224 - 0xe0
    "11111110", -- 2070 - 0x816  :  254 - 0xfe
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "01111110", -- 2072 - 0x818  :  126 - 0x7e -- Background 0x3
    "00001100", -- 2073 - 0x819  :   12 - 0xc
    "00011000", -- 2074 - 0x81a  :   24 - 0x18
    "00111100", -- 2075 - 0x81b  :   60 - 0x3c
    "00000110", -- 2076 - 0x81c  :    6 - 0x6
    "11000110", -- 2077 - 0x81d  :  198 - 0xc6
    "01111100", -- 2078 - 0x81e  :  124 - 0x7c
    "00000000", -- 2079 - 0x81f  :    0 - 0x0
    "00011100", -- 2080 - 0x820  :   28 - 0x1c -- Background 0x4
    "00111100", -- 2081 - 0x821  :   60 - 0x3c
    "01101100", -- 2082 - 0x822  :  108 - 0x6c
    "11001100", -- 2083 - 0x823  :  204 - 0xcc
    "11111110", -- 2084 - 0x824  :  254 - 0xfe
    "00001100", -- 2085 - 0x825  :   12 - 0xc
    "00001100", -- 2086 - 0x826  :   12 - 0xc
    "00000000", -- 2087 - 0x827  :    0 - 0x0
    "11111100", -- 2088 - 0x828  :  252 - 0xfc -- Background 0x5
    "11000000", -- 2089 - 0x829  :  192 - 0xc0
    "11111100", -- 2090 - 0x82a  :  252 - 0xfc
    "00000110", -- 2091 - 0x82b  :    6 - 0x6
    "00000110", -- 2092 - 0x82c  :    6 - 0x6
    "11000110", -- 2093 - 0x82d  :  198 - 0xc6
    "01111100", -- 2094 - 0x82e  :  124 - 0x7c
    "00000000", -- 2095 - 0x82f  :    0 - 0x0
    "00111100", -- 2096 - 0x830  :   60 - 0x3c -- Background 0x6
    "01100000", -- 2097 - 0x831  :   96 - 0x60
    "11000000", -- 2098 - 0x832  :  192 - 0xc0
    "11111100", -- 2099 - 0x833  :  252 - 0xfc
    "11000110", -- 2100 - 0x834  :  198 - 0xc6
    "11000110", -- 2101 - 0x835  :  198 - 0xc6
    "01111100", -- 2102 - 0x836  :  124 - 0x7c
    "00000000", -- 2103 - 0x837  :    0 - 0x0
    "11111110", -- 2104 - 0x838  :  254 - 0xfe -- Background 0x7
    "11000110", -- 2105 - 0x839  :  198 - 0xc6
    "00001100", -- 2106 - 0x83a  :   12 - 0xc
    "00011000", -- 2107 - 0x83b  :   24 - 0x18
    "00110000", -- 2108 - 0x83c  :   48 - 0x30
    "00110000", -- 2109 - 0x83d  :   48 - 0x30
    "00110000", -- 2110 - 0x83e  :   48 - 0x30
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "01111000", -- 2112 - 0x840  :  120 - 0x78 -- Background 0x8
    "11000100", -- 2113 - 0x841  :  196 - 0xc4
    "11100100", -- 2114 - 0x842  :  228 - 0xe4
    "01111000", -- 2115 - 0x843  :  120 - 0x78
    "10000110", -- 2116 - 0x844  :  134 - 0x86
    "10000110", -- 2117 - 0x845  :  134 - 0x86
    "01111100", -- 2118 - 0x846  :  124 - 0x7c
    "00000000", -- 2119 - 0x847  :    0 - 0x0
    "01111100", -- 2120 - 0x848  :  124 - 0x7c -- Background 0x9
    "11000110", -- 2121 - 0x849  :  198 - 0xc6
    "11000110", -- 2122 - 0x84a  :  198 - 0xc6
    "01111110", -- 2123 - 0x84b  :  126 - 0x7e
    "00000110", -- 2124 - 0x84c  :    6 - 0x6
    "00001100", -- 2125 - 0x84d  :   12 - 0xc
    "01111000", -- 2126 - 0x84e  :  120 - 0x78
    "00000000", -- 2127 - 0x84f  :    0 - 0x0
    "00111000", -- 2128 - 0x850  :   56 - 0x38 -- Background 0xa
    "01101100", -- 2129 - 0x851  :  108 - 0x6c
    "11000110", -- 2130 - 0x852  :  198 - 0xc6
    "11000110", -- 2131 - 0x853  :  198 - 0xc6
    "11111110", -- 2132 - 0x854  :  254 - 0xfe
    "11000110", -- 2133 - 0x855  :  198 - 0xc6
    "11000110", -- 2134 - 0x856  :  198 - 0xc6
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "11111100", -- 2136 - 0x858  :  252 - 0xfc -- Background 0xb
    "11000110", -- 2137 - 0x859  :  198 - 0xc6
    "11000110", -- 2138 - 0x85a  :  198 - 0xc6
    "11111100", -- 2139 - 0x85b  :  252 - 0xfc
    "11000110", -- 2140 - 0x85c  :  198 - 0xc6
    "11000110", -- 2141 - 0x85d  :  198 - 0xc6
    "11111100", -- 2142 - 0x85e  :  252 - 0xfc
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "00111100", -- 2144 - 0x860  :   60 - 0x3c -- Background 0xc
    "01100110", -- 2145 - 0x861  :  102 - 0x66
    "11000000", -- 2146 - 0x862  :  192 - 0xc0
    "11000000", -- 2147 - 0x863  :  192 - 0xc0
    "11000000", -- 2148 - 0x864  :  192 - 0xc0
    "01100110", -- 2149 - 0x865  :  102 - 0x66
    "00111100", -- 2150 - 0x866  :   60 - 0x3c
    "00000000", -- 2151 - 0x867  :    0 - 0x0
    "11111000", -- 2152 - 0x868  :  248 - 0xf8 -- Background 0xd
    "11001100", -- 2153 - 0x869  :  204 - 0xcc
    "11000110", -- 2154 - 0x86a  :  198 - 0xc6
    "11000110", -- 2155 - 0x86b  :  198 - 0xc6
    "11000110", -- 2156 - 0x86c  :  198 - 0xc6
    "11001100", -- 2157 - 0x86d  :  204 - 0xcc
    "11111000", -- 2158 - 0x86e  :  248 - 0xf8
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "11111110", -- 2160 - 0x870  :  254 - 0xfe -- Background 0xe
    "11000000", -- 2161 - 0x871  :  192 - 0xc0
    "11000000", -- 2162 - 0x872  :  192 - 0xc0
    "11111100", -- 2163 - 0x873  :  252 - 0xfc
    "11000000", -- 2164 - 0x874  :  192 - 0xc0
    "11000000", -- 2165 - 0x875  :  192 - 0xc0
    "11111110", -- 2166 - 0x876  :  254 - 0xfe
    "00000000", -- 2167 - 0x877  :    0 - 0x0
    "11111110", -- 2168 - 0x878  :  254 - 0xfe -- Background 0xf
    "11000000", -- 2169 - 0x879  :  192 - 0xc0
    "11000000", -- 2170 - 0x87a  :  192 - 0xc0
    "11111100", -- 2171 - 0x87b  :  252 - 0xfc
    "11000000", -- 2172 - 0x87c  :  192 - 0xc0
    "11000000", -- 2173 - 0x87d  :  192 - 0xc0
    "11000000", -- 2174 - 0x87e  :  192 - 0xc0
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "00111110", -- 2176 - 0x880  :   62 - 0x3e -- Background 0x10
    "01100000", -- 2177 - 0x881  :   96 - 0x60
    "11000000", -- 2178 - 0x882  :  192 - 0xc0
    "11011110", -- 2179 - 0x883  :  222 - 0xde
    "11000110", -- 2180 - 0x884  :  198 - 0xc6
    "01100110", -- 2181 - 0x885  :  102 - 0x66
    "01111110", -- 2182 - 0x886  :  126 - 0x7e
    "00000000", -- 2183 - 0x887  :    0 - 0x0
    "11000110", -- 2184 - 0x888  :  198 - 0xc6 -- Background 0x11
    "11000110", -- 2185 - 0x889  :  198 - 0xc6
    "11000110", -- 2186 - 0x88a  :  198 - 0xc6
    "11111110", -- 2187 - 0x88b  :  254 - 0xfe
    "11000110", -- 2188 - 0x88c  :  198 - 0xc6
    "11000110", -- 2189 - 0x88d  :  198 - 0xc6
    "11000110", -- 2190 - 0x88e  :  198 - 0xc6
    "00000000", -- 2191 - 0x88f  :    0 - 0x0
    "01111110", -- 2192 - 0x890  :  126 - 0x7e -- Background 0x12
    "00011000", -- 2193 - 0x891  :   24 - 0x18
    "00011000", -- 2194 - 0x892  :   24 - 0x18
    "00011000", -- 2195 - 0x893  :   24 - 0x18
    "00011000", -- 2196 - 0x894  :   24 - 0x18
    "00011000", -- 2197 - 0x895  :   24 - 0x18
    "01111110", -- 2198 - 0x896  :  126 - 0x7e
    "00000000", -- 2199 - 0x897  :    0 - 0x0
    "00011110", -- 2200 - 0x898  :   30 - 0x1e -- Background 0x13
    "00000110", -- 2201 - 0x899  :    6 - 0x6
    "00000110", -- 2202 - 0x89a  :    6 - 0x6
    "00000110", -- 2203 - 0x89b  :    6 - 0x6
    "11000110", -- 2204 - 0x89c  :  198 - 0xc6
    "11000110", -- 2205 - 0x89d  :  198 - 0xc6
    "01111100", -- 2206 - 0x89e  :  124 - 0x7c
    "00000000", -- 2207 - 0x89f  :    0 - 0x0
    "11000110", -- 2208 - 0x8a0  :  198 - 0xc6 -- Background 0x14
    "11001100", -- 2209 - 0x8a1  :  204 - 0xcc
    "11011000", -- 2210 - 0x8a2  :  216 - 0xd8
    "11110000", -- 2211 - 0x8a3  :  240 - 0xf0
    "11111000", -- 2212 - 0x8a4  :  248 - 0xf8
    "11011100", -- 2213 - 0x8a5  :  220 - 0xdc
    "11001110", -- 2214 - 0x8a6  :  206 - 0xce
    "00000000", -- 2215 - 0x8a7  :    0 - 0x0
    "01100000", -- 2216 - 0x8a8  :   96 - 0x60 -- Background 0x15
    "01100000", -- 2217 - 0x8a9  :   96 - 0x60
    "01100000", -- 2218 - 0x8aa  :   96 - 0x60
    "01100000", -- 2219 - 0x8ab  :   96 - 0x60
    "01100000", -- 2220 - 0x8ac  :   96 - 0x60
    "01100000", -- 2221 - 0x8ad  :   96 - 0x60
    "01111110", -- 2222 - 0x8ae  :  126 - 0x7e
    "00000000", -- 2223 - 0x8af  :    0 - 0x0
    "11000110", -- 2224 - 0x8b0  :  198 - 0xc6 -- Background 0x16
    "11101110", -- 2225 - 0x8b1  :  238 - 0xee
    "11111110", -- 2226 - 0x8b2  :  254 - 0xfe
    "11111110", -- 2227 - 0x8b3  :  254 - 0xfe
    "11010110", -- 2228 - 0x8b4  :  214 - 0xd6
    "11000110", -- 2229 - 0x8b5  :  198 - 0xc6
    "11000110", -- 2230 - 0x8b6  :  198 - 0xc6
    "00000000", -- 2231 - 0x8b7  :    0 - 0x0
    "11000110", -- 2232 - 0x8b8  :  198 - 0xc6 -- Background 0x17
    "11100110", -- 2233 - 0x8b9  :  230 - 0xe6
    "11110110", -- 2234 - 0x8ba  :  246 - 0xf6
    "11111110", -- 2235 - 0x8bb  :  254 - 0xfe
    "11011110", -- 2236 - 0x8bc  :  222 - 0xde
    "11001110", -- 2237 - 0x8bd  :  206 - 0xce
    "11000110", -- 2238 - 0x8be  :  198 - 0xc6
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "01111100", -- 2240 - 0x8c0  :  124 - 0x7c -- Background 0x18
    "11000110", -- 2241 - 0x8c1  :  198 - 0xc6
    "11000110", -- 2242 - 0x8c2  :  198 - 0xc6
    "11000110", -- 2243 - 0x8c3  :  198 - 0xc6
    "11000110", -- 2244 - 0x8c4  :  198 - 0xc6
    "11000110", -- 2245 - 0x8c5  :  198 - 0xc6
    "01111100", -- 2246 - 0x8c6  :  124 - 0x7c
    "00000000", -- 2247 - 0x8c7  :    0 - 0x0
    "11111100", -- 2248 - 0x8c8  :  252 - 0xfc -- Background 0x19
    "11000110", -- 2249 - 0x8c9  :  198 - 0xc6
    "11000110", -- 2250 - 0x8ca  :  198 - 0xc6
    "11000110", -- 2251 - 0x8cb  :  198 - 0xc6
    "11111100", -- 2252 - 0x8cc  :  252 - 0xfc
    "11000000", -- 2253 - 0x8cd  :  192 - 0xc0
    "11000000", -- 2254 - 0x8ce  :  192 - 0xc0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "01111100", -- 2256 - 0x8d0  :  124 - 0x7c -- Background 0x1a
    "11000110", -- 2257 - 0x8d1  :  198 - 0xc6
    "11000110", -- 2258 - 0x8d2  :  198 - 0xc6
    "11000110", -- 2259 - 0x8d3  :  198 - 0xc6
    "11011110", -- 2260 - 0x8d4  :  222 - 0xde
    "11001100", -- 2261 - 0x8d5  :  204 - 0xcc
    "01111010", -- 2262 - 0x8d6  :  122 - 0x7a
    "00000000", -- 2263 - 0x8d7  :    0 - 0x0
    "11111100", -- 2264 - 0x8d8  :  252 - 0xfc -- Background 0x1b
    "11000110", -- 2265 - 0x8d9  :  198 - 0xc6
    "11000110", -- 2266 - 0x8da  :  198 - 0xc6
    "11001110", -- 2267 - 0x8db  :  206 - 0xce
    "11111000", -- 2268 - 0x8dc  :  248 - 0xf8
    "11011100", -- 2269 - 0x8dd  :  220 - 0xdc
    "11001110", -- 2270 - 0x8de  :  206 - 0xce
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "01111000", -- 2272 - 0x8e0  :  120 - 0x78 -- Background 0x1c
    "11001100", -- 2273 - 0x8e1  :  204 - 0xcc
    "11000000", -- 2274 - 0x8e2  :  192 - 0xc0
    "01111100", -- 2275 - 0x8e3  :  124 - 0x7c
    "00000110", -- 2276 - 0x8e4  :    6 - 0x6
    "11000110", -- 2277 - 0x8e5  :  198 - 0xc6
    "01111100", -- 2278 - 0x8e6  :  124 - 0x7c
    "00000000", -- 2279 - 0x8e7  :    0 - 0x0
    "01111110", -- 2280 - 0x8e8  :  126 - 0x7e -- Background 0x1d
    "00011000", -- 2281 - 0x8e9  :   24 - 0x18
    "00011000", -- 2282 - 0x8ea  :   24 - 0x18
    "00011000", -- 2283 - 0x8eb  :   24 - 0x18
    "00011000", -- 2284 - 0x8ec  :   24 - 0x18
    "00011000", -- 2285 - 0x8ed  :   24 - 0x18
    "00011000", -- 2286 - 0x8ee  :   24 - 0x18
    "00000000", -- 2287 - 0x8ef  :    0 - 0x0
    "11000110", -- 2288 - 0x8f0  :  198 - 0xc6 -- Background 0x1e
    "11000110", -- 2289 - 0x8f1  :  198 - 0xc6
    "11000110", -- 2290 - 0x8f2  :  198 - 0xc6
    "11000110", -- 2291 - 0x8f3  :  198 - 0xc6
    "11000110", -- 2292 - 0x8f4  :  198 - 0xc6
    "11000110", -- 2293 - 0x8f5  :  198 - 0xc6
    "01111100", -- 2294 - 0x8f6  :  124 - 0x7c
    "00000000", -- 2295 - 0x8f7  :    0 - 0x0
    "11000110", -- 2296 - 0x8f8  :  198 - 0xc6 -- Background 0x1f
    "11000110", -- 2297 - 0x8f9  :  198 - 0xc6
    "11000110", -- 2298 - 0x8fa  :  198 - 0xc6
    "11101110", -- 2299 - 0x8fb  :  238 - 0xee
    "01111100", -- 2300 - 0x8fc  :  124 - 0x7c
    "00111000", -- 2301 - 0x8fd  :   56 - 0x38
    "00010000", -- 2302 - 0x8fe  :   16 - 0x10
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "11000110", -- 2304 - 0x900  :  198 - 0xc6 -- Background 0x20
    "11000110", -- 2305 - 0x901  :  198 - 0xc6
    "11010110", -- 2306 - 0x902  :  214 - 0xd6
    "11111110", -- 2307 - 0x903  :  254 - 0xfe
    "11111110", -- 2308 - 0x904  :  254 - 0xfe
    "11101110", -- 2309 - 0x905  :  238 - 0xee
    "11000110", -- 2310 - 0x906  :  198 - 0xc6
    "00000000", -- 2311 - 0x907  :    0 - 0x0
    "11000110", -- 2312 - 0x908  :  198 - 0xc6 -- Background 0x21
    "11101110", -- 2313 - 0x909  :  238 - 0xee
    "01111100", -- 2314 - 0x90a  :  124 - 0x7c
    "00111000", -- 2315 - 0x90b  :   56 - 0x38
    "01111100", -- 2316 - 0x90c  :  124 - 0x7c
    "11101110", -- 2317 - 0x90d  :  238 - 0xee
    "11000110", -- 2318 - 0x90e  :  198 - 0xc6
    "00000000", -- 2319 - 0x90f  :    0 - 0x0
    "01100110", -- 2320 - 0x910  :  102 - 0x66 -- Background 0x22
    "01100110", -- 2321 - 0x911  :  102 - 0x66
    "01100110", -- 2322 - 0x912  :  102 - 0x66
    "00111100", -- 2323 - 0x913  :   60 - 0x3c
    "00011000", -- 2324 - 0x914  :   24 - 0x18
    "00011000", -- 2325 - 0x915  :   24 - 0x18
    "00011000", -- 2326 - 0x916  :   24 - 0x18
    "00000000", -- 2327 - 0x917  :    0 - 0x0
    "11111110", -- 2328 - 0x918  :  254 - 0xfe -- Background 0x23
    "00001110", -- 2329 - 0x919  :   14 - 0xe
    "00011100", -- 2330 - 0x91a  :   28 - 0x1c
    "00111000", -- 2331 - 0x91b  :   56 - 0x38
    "01110000", -- 2332 - 0x91c  :  112 - 0x70
    "11100000", -- 2333 - 0x91d  :  224 - 0xe0
    "11111110", -- 2334 - 0x91e  :  254 - 0xfe
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "00000000", -- 2336 - 0x920  :    0 - 0x0 -- Background 0x24
    "00000000", -- 2337 - 0x921  :    0 - 0x0
    "00000000", -- 2338 - 0x922  :    0 - 0x0
    "00000000", -- 2339 - 0x923  :    0 - 0x0
    "00000000", -- 2340 - 0x924  :    0 - 0x0
    "00000000", -- 2341 - 0x925  :    0 - 0x0
    "00000000", -- 2342 - 0x926  :    0 - 0x0
    "00000000", -- 2343 - 0x927  :    0 - 0x0
    "00000000", -- 2344 - 0x928  :    0 - 0x0 -- Background 0x25
    "00000000", -- 2345 - 0x929  :    0 - 0x0
    "00000110", -- 2346 - 0x92a  :    6 - 0x6
    "00001110", -- 2347 - 0x92b  :   14 - 0xe
    "00001000", -- 2348 - 0x92c  :    8 - 0x8
    "00001000", -- 2349 - 0x92d  :    8 - 0x8
    "00001000", -- 2350 - 0x92e  :    8 - 0x8
    "00001000", -- 2351 - 0x92f  :    8 - 0x8
    "00000000", -- 2352 - 0x930  :    0 - 0x0 -- Background 0x26
    "01111000", -- 2353 - 0x931  :  120 - 0x78
    "01100101", -- 2354 - 0x932  :  101 - 0x65
    "01111001", -- 2355 - 0x933  :  121 - 0x79
    "01100101", -- 2356 - 0x934  :  101 - 0x65
    "01100101", -- 2357 - 0x935  :  101 - 0x65
    "01111000", -- 2358 - 0x936  :  120 - 0x78
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "00000000", -- 2360 - 0x938  :    0 - 0x0 -- Background 0x27
    "11100100", -- 2361 - 0x939  :  228 - 0xe4
    "10010110", -- 2362 - 0x93a  :  150 - 0x96
    "10010110", -- 2363 - 0x93b  :  150 - 0x96
    "10010111", -- 2364 - 0x93c  :  151 - 0x97
    "10010110", -- 2365 - 0x93d  :  150 - 0x96
    "11100110", -- 2366 - 0x93e  :  230 - 0xe6
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Background 0x28
    "01011001", -- 2369 - 0x941  :   89 - 0x59
    "01011001", -- 2370 - 0x942  :   89 - 0x59
    "01011001", -- 2371 - 0x943  :   89 - 0x59
    "01011001", -- 2372 - 0x944  :   89 - 0x59
    "11011001", -- 2373 - 0x945  :  217 - 0xd9
    "01001110", -- 2374 - 0x946  :   78 - 0x4e
    "00000000", -- 2375 - 0x947  :    0 - 0x0
    "00000000", -- 2376 - 0x948  :    0 - 0x0 -- Background 0x29
    "00111100", -- 2377 - 0x949  :   60 - 0x3c
    "01110000", -- 2378 - 0x94a  :  112 - 0x70
    "01110000", -- 2379 - 0x94b  :  112 - 0x70
    "00111100", -- 2380 - 0x94c  :   60 - 0x3c
    "00001100", -- 2381 - 0x94d  :   12 - 0xc
    "01111000", -- 2382 - 0x94e  :  120 - 0x78
    "00000000", -- 2383 - 0x94f  :    0 - 0x0
    "00000000", -- 2384 - 0x950  :    0 - 0x0 -- Background 0x2a
    "00000000", -- 2385 - 0x951  :    0 - 0x0
    "11000110", -- 2386 - 0x952  :  198 - 0xc6
    "11101110", -- 2387 - 0x953  :  238 - 0xee
    "00101000", -- 2388 - 0x954  :   40 - 0x28
    "00101000", -- 2389 - 0x955  :   40 - 0x28
    "00101000", -- 2390 - 0x956  :   40 - 0x28
    "00101000", -- 2391 - 0x957  :   40 - 0x28
    "00001000", -- 2392 - 0x958  :    8 - 0x8 -- Background 0x2b
    "00001000", -- 2393 - 0x959  :    8 - 0x8
    "00001000", -- 2394 - 0x95a  :    8 - 0x8
    "00001000", -- 2395 - 0x95b  :    8 - 0x8
    "00001110", -- 2396 - 0x95c  :   14 - 0xe
    "00000110", -- 2397 - 0x95d  :    6 - 0x6
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "00101000", -- 2400 - 0x960  :   40 - 0x28 -- Background 0x2c
    "00101000", -- 2401 - 0x961  :   40 - 0x28
    "00101000", -- 2402 - 0x962  :   40 - 0x28
    "00101000", -- 2403 - 0x963  :   40 - 0x28
    "11101110", -- 2404 - 0x964  :  238 - 0xee
    "11000110", -- 2405 - 0x965  :  198 - 0xc6
    "00000000", -- 2406 - 0x966  :    0 - 0x0
    "00000000", -- 2407 - 0x967  :    0 - 0x0
    "00000000", -- 2408 - 0x968  :    0 - 0x0 -- Background 0x2d
    "00000000", -- 2409 - 0x969  :    0 - 0x0
    "01100000", -- 2410 - 0x96a  :   96 - 0x60
    "01110000", -- 2411 - 0x96b  :  112 - 0x70
    "00010000", -- 2412 - 0x96c  :   16 - 0x10
    "00010000", -- 2413 - 0x96d  :   16 - 0x10
    "00010000", -- 2414 - 0x96e  :   16 - 0x10
    "00010000", -- 2415 - 0x96f  :   16 - 0x10
    "00011100", -- 2416 - 0x970  :   28 - 0x1c -- Background 0x2e
    "00111110", -- 2417 - 0x971  :   62 - 0x3e
    "00111100", -- 2418 - 0x972  :   60 - 0x3c
    "00111000", -- 2419 - 0x973  :   56 - 0x38
    "00110000", -- 2420 - 0x974  :   48 - 0x30
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "01100000", -- 2422 - 0x976  :   96 - 0x60
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "00010000", -- 2424 - 0x978  :   16 - 0x10 -- Background 0x2f
    "00010000", -- 2425 - 0x979  :   16 - 0x10
    "00010000", -- 2426 - 0x97a  :   16 - 0x10
    "00010000", -- 2427 - 0x97b  :   16 - 0x10
    "01110000", -- 2428 - 0x97c  :  112 - 0x70
    "01100000", -- 2429 - 0x97d  :   96 - 0x60
    "00000000", -- 2430 - 0x97e  :    0 - 0x0
    "00000000", -- 2431 - 0x97f  :    0 - 0x0
    "11111111", -- 2432 - 0x980  :  255 - 0xff -- Background 0x30
    "11111111", -- 2433 - 0x981  :  255 - 0xff
    "00111000", -- 2434 - 0x982  :   56 - 0x38
    "01101100", -- 2435 - 0x983  :  108 - 0x6c
    "11000110", -- 2436 - 0x984  :  198 - 0xc6
    "10000011", -- 2437 - 0x985  :  131 - 0x83
    "11111111", -- 2438 - 0x986  :  255 - 0xff
    "11111111", -- 2439 - 0x987  :  255 - 0xff
    "11111111", -- 2440 - 0x988  :  255 - 0xff -- Background 0x31
    "00111000", -- 2441 - 0x989  :   56 - 0x38
    "01101100", -- 2442 - 0x98a  :  108 - 0x6c
    "11000110", -- 2443 - 0x98b  :  198 - 0xc6
    "10000011", -- 2444 - 0x98c  :  131 - 0x83
    "11111111", -- 2445 - 0x98d  :  255 - 0xff
    "11111111", -- 2446 - 0x98e  :  255 - 0xff
    "00000000", -- 2447 - 0x98f  :    0 - 0x0
    "00111000", -- 2448 - 0x990  :   56 - 0x38 -- Background 0x32
    "01101100", -- 2449 - 0x991  :  108 - 0x6c
    "11000110", -- 2450 - 0x992  :  198 - 0xc6
    "10000011", -- 2451 - 0x993  :  131 - 0x83
    "11111111", -- 2452 - 0x994  :  255 - 0xff
    "11111111", -- 2453 - 0x995  :  255 - 0xff
    "00000000", -- 2454 - 0x996  :    0 - 0x0
    "00000000", -- 2455 - 0x997  :    0 - 0x0
    "01101100", -- 2456 - 0x998  :  108 - 0x6c -- Background 0x33
    "11000110", -- 2457 - 0x999  :  198 - 0xc6
    "10000011", -- 2458 - 0x99a  :  131 - 0x83
    "11111111", -- 2459 - 0x99b  :  255 - 0xff
    "11111111", -- 2460 - 0x99c  :  255 - 0xff
    "00000000", -- 2461 - 0x99d  :    0 - 0x0
    "00000000", -- 2462 - 0x99e  :    0 - 0x0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "11000110", -- 2464 - 0x9a0  :  198 - 0xc6 -- Background 0x34
    "10000011", -- 2465 - 0x9a1  :  131 - 0x83
    "11111111", -- 2466 - 0x9a2  :  255 - 0xff
    "11111111", -- 2467 - 0x9a3  :  255 - 0xff
    "00000000", -- 2468 - 0x9a4  :    0 - 0x0
    "00000000", -- 2469 - 0x9a5  :    0 - 0x0
    "00000000", -- 2470 - 0x9a6  :    0 - 0x0
    "00000000", -- 2471 - 0x9a7  :    0 - 0x0
    "10000011", -- 2472 - 0x9a8  :  131 - 0x83 -- Background 0x35
    "11111111", -- 2473 - 0x9a9  :  255 - 0xff
    "11111111", -- 2474 - 0x9aa  :  255 - 0xff
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00000000", -- 2476 - 0x9ac  :    0 - 0x0
    "00000000", -- 2477 - 0x9ad  :    0 - 0x0
    "00000000", -- 2478 - 0x9ae  :    0 - 0x0
    "00000000", -- 2479 - 0x9af  :    0 - 0x0
    "11111111", -- 2480 - 0x9b0  :  255 - 0xff -- Background 0x36
    "11111111", -- 2481 - 0x9b1  :  255 - 0xff
    "00000000", -- 2482 - 0x9b2  :    0 - 0x0
    "00000000", -- 2483 - 0x9b3  :    0 - 0x0
    "00000000", -- 2484 - 0x9b4  :    0 - 0x0
    "00000000", -- 2485 - 0x9b5  :    0 - 0x0
    "00000000", -- 2486 - 0x9b6  :    0 - 0x0
    "00000000", -- 2487 - 0x9b7  :    0 - 0x0
    "11111111", -- 2488 - 0x9b8  :  255 - 0xff -- Background 0x37
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "00000000", -- 2490 - 0x9ba  :    0 - 0x0
    "00000000", -- 2491 - 0x9bb  :    0 - 0x0
    "00000000", -- 2492 - 0x9bc  :    0 - 0x0
    "00000000", -- 2493 - 0x9bd  :    0 - 0x0
    "00000000", -- 2494 - 0x9be  :    0 - 0x0
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0 -- Background 0x38
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000000", -- 2498 - 0x9c2  :    0 - 0x0
    "00000000", -- 2499 - 0x9c3  :    0 - 0x0
    "00000000", -- 2500 - 0x9c4  :    0 - 0x0
    "00000000", -- 2501 - 0x9c5  :    0 - 0x0
    "00000000", -- 2502 - 0x9c6  :    0 - 0x0
    "11111111", -- 2503 - 0x9c7  :  255 - 0xff
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0 -- Background 0x39
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "11111111", -- 2510 - 0x9ce  :  255 - 0xff
    "11111111", -- 2511 - 0x9cf  :  255 - 0xff
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0 -- Background 0x3a
    "00000000", -- 2513 - 0x9d1  :    0 - 0x0
    "00000000", -- 2514 - 0x9d2  :    0 - 0x0
    "00000000", -- 2515 - 0x9d3  :    0 - 0x0
    "00000000", -- 2516 - 0x9d4  :    0 - 0x0
    "11111111", -- 2517 - 0x9d5  :  255 - 0xff
    "11111111", -- 2518 - 0x9d6  :  255 - 0xff
    "00111000", -- 2519 - 0x9d7  :   56 - 0x38
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0 -- Background 0x3b
    "00000000", -- 2521 - 0x9d9  :    0 - 0x0
    "00000000", -- 2522 - 0x9da  :    0 - 0x0
    "00000000", -- 2523 - 0x9db  :    0 - 0x0
    "11111111", -- 2524 - 0x9dc  :  255 - 0xff
    "11111111", -- 2525 - 0x9dd  :  255 - 0xff
    "00111000", -- 2526 - 0x9de  :   56 - 0x38
    "01101100", -- 2527 - 0x9df  :  108 - 0x6c
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0 -- Background 0x3c
    "00000000", -- 2529 - 0x9e1  :    0 - 0x0
    "00000000", -- 2530 - 0x9e2  :    0 - 0x0
    "11111111", -- 2531 - 0x9e3  :  255 - 0xff
    "11111111", -- 2532 - 0x9e4  :  255 - 0xff
    "00111000", -- 2533 - 0x9e5  :   56 - 0x38
    "01101100", -- 2534 - 0x9e6  :  108 - 0x6c
    "11000110", -- 2535 - 0x9e7  :  198 - 0xc6
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0 -- Background 0x3d
    "00000000", -- 2537 - 0x9e9  :    0 - 0x0
    "11111111", -- 2538 - 0x9ea  :  255 - 0xff
    "11111111", -- 2539 - 0x9eb  :  255 - 0xff
    "00111000", -- 2540 - 0x9ec  :   56 - 0x38
    "01101100", -- 2541 - 0x9ed  :  108 - 0x6c
    "11000110", -- 2542 - 0x9ee  :  198 - 0xc6
    "10000011", -- 2543 - 0x9ef  :  131 - 0x83
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0 -- Background 0x3e
    "11111111", -- 2545 - 0x9f1  :  255 - 0xff
    "11111111", -- 2546 - 0x9f2  :  255 - 0xff
    "00111000", -- 2547 - 0x9f3  :   56 - 0x38
    "01101100", -- 2548 - 0x9f4  :  108 - 0x6c
    "11000110", -- 2549 - 0x9f5  :  198 - 0xc6
    "10000011", -- 2550 - 0x9f6  :  131 - 0x83
    "11111111", -- 2551 - 0x9f7  :  255 - 0xff
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00000000", -- 2560 - 0xa00  :    0 - 0x0 -- Background 0x40
    "00000000", -- 2561 - 0xa01  :    0 - 0x0
    "00000000", -- 2562 - 0xa02  :    0 - 0x0
    "00000000", -- 2563 - 0xa03  :    0 - 0x0
    "00000000", -- 2564 - 0xa04  :    0 - 0x0
    "00000000", -- 2565 - 0xa05  :    0 - 0x0
    "00000000", -- 2566 - 0xa06  :    0 - 0x0
    "11111111", -- 2567 - 0xa07  :  255 - 0xff
    "00000000", -- 2568 - 0xa08  :    0 - 0x0 -- Background 0x41
    "00000000", -- 2569 - 0xa09  :    0 - 0x0
    "00000000", -- 2570 - 0xa0a  :    0 - 0x0
    "00000000", -- 2571 - 0xa0b  :    0 - 0x0
    "00000000", -- 2572 - 0xa0c  :    0 - 0x0
    "11111111", -- 2573 - 0xa0d  :  255 - 0xff
    "11111111", -- 2574 - 0xa0e  :  255 - 0xff
    "00111000", -- 2575 - 0xa0f  :   56 - 0x38
    "00000000", -- 2576 - 0xa10  :    0 - 0x0 -- Background 0x42
    "00000000", -- 2577 - 0xa11  :    0 - 0x0
    "00000000", -- 2578 - 0xa12  :    0 - 0x0
    "00000000", -- 2579 - 0xa13  :    0 - 0x0
    "11111111", -- 2580 - 0xa14  :  255 - 0xff
    "11111111", -- 2581 - 0xa15  :  255 - 0xff
    "00111000", -- 2582 - 0xa16  :   56 - 0x38
    "01101100", -- 2583 - 0xa17  :  108 - 0x6c
    "00000000", -- 2584 - 0xa18  :    0 - 0x0 -- Background 0x43
    "00000000", -- 2585 - 0xa19  :    0 - 0x0
    "00000000", -- 2586 - 0xa1a  :    0 - 0x0
    "11111111", -- 2587 - 0xa1b  :  255 - 0xff
    "11111111", -- 2588 - 0xa1c  :  255 - 0xff
    "00111000", -- 2589 - 0xa1d  :   56 - 0x38
    "01101100", -- 2590 - 0xa1e  :  108 - 0x6c
    "11000110", -- 2591 - 0xa1f  :  198 - 0xc6
    "00000000", -- 2592 - 0xa20  :    0 - 0x0 -- Background 0x44
    "00000000", -- 2593 - 0xa21  :    0 - 0x0
    "11111111", -- 2594 - 0xa22  :  255 - 0xff
    "11111111", -- 2595 - 0xa23  :  255 - 0xff
    "00111000", -- 2596 - 0xa24  :   56 - 0x38
    "01101100", -- 2597 - 0xa25  :  108 - 0x6c
    "11000110", -- 2598 - 0xa26  :  198 - 0xc6
    "10000011", -- 2599 - 0xa27  :  131 - 0x83
    "00000000", -- 2600 - 0xa28  :    0 - 0x0 -- Background 0x45
    "11111111", -- 2601 - 0xa29  :  255 - 0xff
    "11111111", -- 2602 - 0xa2a  :  255 - 0xff
    "00111000", -- 2603 - 0xa2b  :   56 - 0x38
    "01101100", -- 2604 - 0xa2c  :  108 - 0x6c
    "11000110", -- 2605 - 0xa2d  :  198 - 0xc6
    "10000011", -- 2606 - 0xa2e  :  131 - 0x83
    "11111111", -- 2607 - 0xa2f  :  255 - 0xff
    "11111111", -- 2608 - 0xa30  :  255 - 0xff -- Background 0x46
    "00111000", -- 2609 - 0xa31  :   56 - 0x38
    "01101100", -- 2610 - 0xa32  :  108 - 0x6c
    "11000110", -- 2611 - 0xa33  :  198 - 0xc6
    "10000011", -- 2612 - 0xa34  :  131 - 0x83
    "11111111", -- 2613 - 0xa35  :  255 - 0xff
    "11111111", -- 2614 - 0xa36  :  255 - 0xff
    "00000000", -- 2615 - 0xa37  :    0 - 0x0
    "00111000", -- 2616 - 0xa38  :   56 - 0x38 -- Background 0x47
    "01101100", -- 2617 - 0xa39  :  108 - 0x6c
    "11000110", -- 2618 - 0xa3a  :  198 - 0xc6
    "10000011", -- 2619 - 0xa3b  :  131 - 0x83
    "11111111", -- 2620 - 0xa3c  :  255 - 0xff
    "11111111", -- 2621 - 0xa3d  :  255 - 0xff
    "00000000", -- 2622 - 0xa3e  :    0 - 0x0
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "01101100", -- 2624 - 0xa40  :  108 - 0x6c -- Background 0x48
    "11000110", -- 2625 - 0xa41  :  198 - 0xc6
    "10000011", -- 2626 - 0xa42  :  131 - 0x83
    "11111111", -- 2627 - 0xa43  :  255 - 0xff
    "11111111", -- 2628 - 0xa44  :  255 - 0xff
    "00000000", -- 2629 - 0xa45  :    0 - 0x0
    "00000000", -- 2630 - 0xa46  :    0 - 0x0
    "00000000", -- 2631 - 0xa47  :    0 - 0x0
    "11000110", -- 2632 - 0xa48  :  198 - 0xc6 -- Background 0x49
    "10000011", -- 2633 - 0xa49  :  131 - 0x83
    "11111111", -- 2634 - 0xa4a  :  255 - 0xff
    "11111111", -- 2635 - 0xa4b  :  255 - 0xff
    "00000000", -- 2636 - 0xa4c  :    0 - 0x0
    "00000000", -- 2637 - 0xa4d  :    0 - 0x0
    "00000000", -- 2638 - 0xa4e  :    0 - 0x0
    "00000000", -- 2639 - 0xa4f  :    0 - 0x0
    "10000011", -- 2640 - 0xa50  :  131 - 0x83 -- Background 0x4a
    "11111111", -- 2641 - 0xa51  :  255 - 0xff
    "11111111", -- 2642 - 0xa52  :  255 - 0xff
    "00000000", -- 2643 - 0xa53  :    0 - 0x0
    "00000000", -- 2644 - 0xa54  :    0 - 0x0
    "00000000", -- 2645 - 0xa55  :    0 - 0x0
    "00000000", -- 2646 - 0xa56  :    0 - 0x0
    "00000000", -- 2647 - 0xa57  :    0 - 0x0
    "11111111", -- 2648 - 0xa58  :  255 - 0xff -- Background 0x4b
    "11111111", -- 2649 - 0xa59  :  255 - 0xff
    "00000000", -- 2650 - 0xa5a  :    0 - 0x0
    "00000000", -- 2651 - 0xa5b  :    0 - 0x0
    "00000000", -- 2652 - 0xa5c  :    0 - 0x0
    "00000000", -- 2653 - 0xa5d  :    0 - 0x0
    "00000000", -- 2654 - 0xa5e  :    0 - 0x0
    "00000000", -- 2655 - 0xa5f  :    0 - 0x0
    "10111111", -- 2656 - 0xa60  :  191 - 0xbf -- Background 0x4c
    "01011111", -- 2657 - 0xa61  :   95 - 0x5f
    "01011111", -- 2658 - 0xa62  :   95 - 0x5f
    "01011111", -- 2659 - 0xa63  :   95 - 0x5f
    "00000000", -- 2660 - 0xa64  :    0 - 0x0
    "01011111", -- 2661 - 0xa65  :   95 - 0x5f
    "01010001", -- 2662 - 0xa66  :   81 - 0x51
    "01010101", -- 2663 - 0xa67  :   85 - 0x55
    "01010001", -- 2664 - 0xa68  :   81 - 0x51 -- Background 0x4d
    "01011111", -- 2665 - 0xa69  :   95 - 0x5f
    "00000000", -- 2666 - 0xa6a  :    0 - 0x0
    "01011111", -- 2667 - 0xa6b  :   95 - 0x5f
    "01011111", -- 2668 - 0xa6c  :   95 - 0x5f
    "01011111", -- 2669 - 0xa6d  :   95 - 0x5f
    "01011111", -- 2670 - 0xa6e  :   95 - 0x5f
    "10111111", -- 2671 - 0xa6f  :  191 - 0xbf
    "11111111", -- 2672 - 0xa70  :  255 - 0xff -- Background 0x4e
    "11111110", -- 2673 - 0xa71  :  254 - 0xfe
    "11111110", -- 2674 - 0xa72  :  254 - 0xfe
    "11111110", -- 2675 - 0xa73  :  254 - 0xfe
    "00000000", -- 2676 - 0xa74  :    0 - 0x0
    "11111110", -- 2677 - 0xa75  :  254 - 0xfe
    "00100110", -- 2678 - 0xa76  :   38 - 0x26
    "00100110", -- 2679 - 0xa77  :   38 - 0x26
    "00100010", -- 2680 - 0xa78  :   34 - 0x22 -- Background 0x4f
    "11111110", -- 2681 - 0xa79  :  254 - 0xfe
    "00000000", -- 2682 - 0xa7a  :    0 - 0x0
    "11111110", -- 2683 - 0xa7b  :  254 - 0xfe
    "11111110", -- 2684 - 0xa7c  :  254 - 0xfe
    "11111110", -- 2685 - 0xa7d  :  254 - 0xfe
    "11111110", -- 2686 - 0xa7e  :  254 - 0xfe
    "11111111", -- 2687 - 0xa7f  :  255 - 0xff
    "00000111", -- 2688 - 0xa80  :    7 - 0x7 -- Background 0x50
    "00000000", -- 2689 - 0xa81  :    0 - 0x0
    "00001111", -- 2690 - 0xa82  :   15 - 0xf
    "00011111", -- 2691 - 0xa83  :   31 - 0x1f
    "00011111", -- 2692 - 0xa84  :   31 - 0x1f
    "00011111", -- 2693 - 0xa85  :   31 - 0x1f
    "00011111", -- 2694 - 0xa86  :   31 - 0x1f
    "00011111", -- 2695 - 0xa87  :   31 - 0x1f
    "00011111", -- 2696 - 0xa88  :   31 - 0x1f -- Background 0x51
    "00011111", -- 2697 - 0xa89  :   31 - 0x1f
    "00011111", -- 2698 - 0xa8a  :   31 - 0x1f
    "00011111", -- 2699 - 0xa8b  :   31 - 0x1f
    "00011111", -- 2700 - 0xa8c  :   31 - 0x1f
    "00001111", -- 2701 - 0xa8d  :   15 - 0xf
    "00000000", -- 2702 - 0xa8e  :    0 - 0x0
    "00000111", -- 2703 - 0xa8f  :    7 - 0x7
    "00000111", -- 2704 - 0xa90  :    7 - 0x7 -- Background 0x52
    "00000000", -- 2705 - 0xa91  :    0 - 0x0
    "00001111", -- 2706 - 0xa92  :   15 - 0xf
    "00011111", -- 2707 - 0xa93  :   31 - 0x1f
    "00011111", -- 2708 - 0xa94  :   31 - 0x1f
    "00011111", -- 2709 - 0xa95  :   31 - 0x1f
    "00011111", -- 2710 - 0xa96  :   31 - 0x1f
    "00011111", -- 2711 - 0xa97  :   31 - 0x1f
    "00011111", -- 2712 - 0xa98  :   31 - 0x1f -- Background 0x53
    "00011111", -- 2713 - 0xa99  :   31 - 0x1f
    "00011111", -- 2714 - 0xa9a  :   31 - 0x1f
    "00011111", -- 2715 - 0xa9b  :   31 - 0x1f
    "00011111", -- 2716 - 0xa9c  :   31 - 0x1f
    "00001111", -- 2717 - 0xa9d  :   15 - 0xf
    "00000000", -- 2718 - 0xa9e  :    0 - 0x0
    "00000111", -- 2719 - 0xa9f  :    7 - 0x7
    "11100000", -- 2720 - 0xaa0  :  224 - 0xe0 -- Background 0x54
    "00000000", -- 2721 - 0xaa1  :    0 - 0x0
    "11110001", -- 2722 - 0xaa2  :  241 - 0xf1
    "11111011", -- 2723 - 0xaa3  :  251 - 0xfb
    "11111011", -- 2724 - 0xaa4  :  251 - 0xfb
    "11111011", -- 2725 - 0xaa5  :  251 - 0xfb
    "11111011", -- 2726 - 0xaa6  :  251 - 0xfb
    "11111011", -- 2727 - 0xaa7  :  251 - 0xfb
    "11111011", -- 2728 - 0xaa8  :  251 - 0xfb -- Background 0x55
    "11111011", -- 2729 - 0xaa9  :  251 - 0xfb
    "11111011", -- 2730 - 0xaaa  :  251 - 0xfb
    "11111011", -- 2731 - 0xaab  :  251 - 0xfb
    "11111011", -- 2732 - 0xaac  :  251 - 0xfb
    "11110001", -- 2733 - 0xaad  :  241 - 0xf1
    "00000000", -- 2734 - 0xaae  :    0 - 0x0
    "11100000", -- 2735 - 0xaaf  :  224 - 0xe0
    "11100000", -- 2736 - 0xab0  :  224 - 0xe0 -- Background 0x56
    "00000000", -- 2737 - 0xab1  :    0 - 0x0
    "11110001", -- 2738 - 0xab2  :  241 - 0xf1
    "11111011", -- 2739 - 0xab3  :  251 - 0xfb
    "11111011", -- 2740 - 0xab4  :  251 - 0xfb
    "11111011", -- 2741 - 0xab5  :  251 - 0xfb
    "11111011", -- 2742 - 0xab6  :  251 - 0xfb
    "11111011", -- 2743 - 0xab7  :  251 - 0xfb
    "11111011", -- 2744 - 0xab8  :  251 - 0xfb -- Background 0x57
    "11111011", -- 2745 - 0xab9  :  251 - 0xfb
    "11111011", -- 2746 - 0xaba  :  251 - 0xfb
    "11111011", -- 2747 - 0xabb  :  251 - 0xfb
    "11111011", -- 2748 - 0xabc  :  251 - 0xfb
    "11110001", -- 2749 - 0xabd  :  241 - 0xf1
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "11100000", -- 2751 - 0xabf  :  224 - 0xe0
    "11111100", -- 2752 - 0xac0  :  252 - 0xfc -- Background 0x58
    "00000000", -- 2753 - 0xac1  :    0 - 0x0
    "11111110", -- 2754 - 0xac2  :  254 - 0xfe
    "11111111", -- 2755 - 0xac3  :  255 - 0xff
    "11111111", -- 2756 - 0xac4  :  255 - 0xff
    "11111111", -- 2757 - 0xac5  :  255 - 0xff
    "11111111", -- 2758 - 0xac6  :  255 - 0xff
    "11111111", -- 2759 - 0xac7  :  255 - 0xff
    "11111111", -- 2760 - 0xac8  :  255 - 0xff -- Background 0x59
    "11111111", -- 2761 - 0xac9  :  255 - 0xff
    "11111111", -- 2762 - 0xaca  :  255 - 0xff
    "11111111", -- 2763 - 0xacb  :  255 - 0xff
    "11111111", -- 2764 - 0xacc  :  255 - 0xff
    "11111110", -- 2765 - 0xacd  :  254 - 0xfe
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "11111100", -- 2767 - 0xacf  :  252 - 0xfc
    "11111100", -- 2768 - 0xad0  :  252 - 0xfc -- Background 0x5a
    "00000000", -- 2769 - 0xad1  :    0 - 0x0
    "11111110", -- 2770 - 0xad2  :  254 - 0xfe
    "11111111", -- 2771 - 0xad3  :  255 - 0xff
    "11111111", -- 2772 - 0xad4  :  255 - 0xff
    "11111111", -- 2773 - 0xad5  :  255 - 0xff
    "11111111", -- 2774 - 0xad6  :  255 - 0xff
    "11111111", -- 2775 - 0xad7  :  255 - 0xff
    "11111111", -- 2776 - 0xad8  :  255 - 0xff -- Background 0x5b
    "11111111", -- 2777 - 0xad9  :  255 - 0xff
    "11111111", -- 2778 - 0xada  :  255 - 0xff
    "11111111", -- 2779 - 0xadb  :  255 - 0xff
    "11111111", -- 2780 - 0xadc  :  255 - 0xff
    "11111110", -- 2781 - 0xadd  :  254 - 0xfe
    "00000000", -- 2782 - 0xade  :    0 - 0x0
    "11111100", -- 2783 - 0xadf  :  252 - 0xfc
    "00000000", -- 2784 - 0xae0  :    0 - 0x0 -- Background 0x5c
    "00000000", -- 2785 - 0xae1  :    0 - 0x0
    "00011111", -- 2786 - 0xae2  :   31 - 0x1f
    "00010000", -- 2787 - 0xae3  :   16 - 0x10
    "00010000", -- 2788 - 0xae4  :   16 - 0x10
    "00011111", -- 2789 - 0xae5  :   31 - 0x1f
    "00000000", -- 2790 - 0xae6  :    0 - 0x0
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "00000000", -- 2792 - 0xae8  :    0 - 0x0 -- Background 0x5d
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "11111000", -- 2794 - 0xaea  :  248 - 0xf8
    "00001000", -- 2795 - 0xaeb  :    8 - 0x8
    "00001000", -- 2796 - 0xaec  :    8 - 0x8
    "11111000", -- 2797 - 0xaed  :  248 - 0xf8
    "00000000", -- 2798 - 0xaee  :    0 - 0x0
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "00000000", -- 2800 - 0xaf0  :    0 - 0x0 -- Background 0x5e
    "00000001", -- 2801 - 0xaf1  :    1 - 0x1
    "00000010", -- 2802 - 0xaf2  :    2 - 0x2
    "00000010", -- 2803 - 0xaf3  :    2 - 0x2
    "11110001", -- 2804 - 0xaf4  :  241 - 0xf1
    "00001000", -- 2805 - 0xaf5  :    8 - 0x8
    "00000100", -- 2806 - 0xaf6  :    4 - 0x4
    "00000011", -- 2807 - 0xaf7  :    3 - 0x3
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0 -- Background 0x5f
    "10000000", -- 2809 - 0xaf9  :  128 - 0x80
    "01000000", -- 2810 - 0xafa  :   64 - 0x40
    "01000000", -- 2811 - 0xafb  :   64 - 0x40
    "10001111", -- 2812 - 0xafc  :  143 - 0x8f
    "00010000", -- 2813 - 0xafd  :   16 - 0x10
    "00100000", -- 2814 - 0xafe  :   32 - 0x20
    "11000000", -- 2815 - 0xaff  :  192 - 0xc0
    "00000011", -- 2816 - 0xb00  :    3 - 0x3 -- Background 0x60
    "00000100", -- 2817 - 0xb01  :    4 - 0x4
    "00001000", -- 2818 - 0xb02  :    8 - 0x8
    "11110001", -- 2819 - 0xb03  :  241 - 0xf1
    "00000010", -- 2820 - 0xb04  :    2 - 0x2
    "00000010", -- 2821 - 0xb05  :    2 - 0x2
    "00000001", -- 2822 - 0xb06  :    1 - 0x1
    "00000000", -- 2823 - 0xb07  :    0 - 0x0
    "11000000", -- 2824 - 0xb08  :  192 - 0xc0 -- Background 0x61
    "00100000", -- 2825 - 0xb09  :   32 - 0x20
    "00010000", -- 2826 - 0xb0a  :   16 - 0x10
    "10001111", -- 2827 - 0xb0b  :  143 - 0x8f
    "01000000", -- 2828 - 0xb0c  :   64 - 0x40
    "01000000", -- 2829 - 0xb0d  :   64 - 0x40
    "10000000", -- 2830 - 0xb0e  :  128 - 0x80
    "00000000", -- 2831 - 0xb0f  :    0 - 0x0
    "11111111", -- 2832 - 0xb10  :  255 - 0xff -- Background 0x62
    "11111111", -- 2833 - 0xb11  :  255 - 0xff
    "11000011", -- 2834 - 0xb12  :  195 - 0xc3
    "10000001", -- 2835 - 0xb13  :  129 - 0x81
    "10000001", -- 2836 - 0xb14  :  129 - 0x81
    "11000011", -- 2837 - 0xb15  :  195 - 0xc3
    "11111111", -- 2838 - 0xb16  :  255 - 0xff
    "11111111", -- 2839 - 0xb17  :  255 - 0xff
    "11111111", -- 2840 - 0xb18  :  255 - 0xff -- Background 0x63
    "10011001", -- 2841 - 0xb19  :  153 - 0x99
    "00000000", -- 2842 - 0xb1a  :    0 - 0x0
    "00000000", -- 2843 - 0xb1b  :    0 - 0x0
    "00000000", -- 2844 - 0xb1c  :    0 - 0x0
    "10000001", -- 2845 - 0xb1d  :  129 - 0x81
    "10000001", -- 2846 - 0xb1e  :  129 - 0x81
    "10000001", -- 2847 - 0xb1f  :  129 - 0x81
    "00000000", -- 2848 - 0xb20  :    0 - 0x0 -- Background 0x64
    "00000000", -- 2849 - 0xb21  :    0 - 0x0
    "00000000", -- 2850 - 0xb22  :    0 - 0x0
    "00000000", -- 2851 - 0xb23  :    0 - 0x0
    "01100000", -- 2852 - 0xb24  :   96 - 0x60
    "01100000", -- 2853 - 0xb25  :   96 - 0x60
    "00000000", -- 2854 - 0xb26  :    0 - 0x0
    "00000000", -- 2855 - 0xb27  :    0 - 0x0
    "00000000", -- 2856 - 0xb28  :    0 - 0x0 -- Background 0x65
    "00000000", -- 2857 - 0xb29  :    0 - 0x0
    "00000000", -- 2858 - 0xb2a  :    0 - 0x0
    "00000000", -- 2859 - 0xb2b  :    0 - 0x0
    "01101100", -- 2860 - 0xb2c  :  108 - 0x6c
    "01101100", -- 2861 - 0xb2d  :  108 - 0x6c
    "00001000", -- 2862 - 0xb2e  :    8 - 0x8
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "00111100", -- 2864 - 0xb30  :   60 - 0x3c -- Background 0x66
    "00011000", -- 2865 - 0xb31  :   24 - 0x18
    "00011000", -- 2866 - 0xb32  :   24 - 0x18
    "00011000", -- 2867 - 0xb33  :   24 - 0x18
    "00011000", -- 2868 - 0xb34  :   24 - 0x18
    "00011000", -- 2869 - 0xb35  :   24 - 0x18
    "00111100", -- 2870 - 0xb36  :   60 - 0x3c
    "00000000", -- 2871 - 0xb37  :    0 - 0x0
    "11111111", -- 2872 - 0xb38  :  255 - 0xff -- Background 0x67
    "01100110", -- 2873 - 0xb39  :  102 - 0x66
    "01100110", -- 2874 - 0xb3a  :  102 - 0x66
    "01100110", -- 2875 - 0xb3b  :  102 - 0x66
    "01100110", -- 2876 - 0xb3c  :  102 - 0x66
    "01100110", -- 2877 - 0xb3d  :  102 - 0x66
    "01100110", -- 2878 - 0xb3e  :  102 - 0x66
    "11111111", -- 2879 - 0xb3f  :  255 - 0xff
    "00000011", -- 2880 - 0xb40  :    3 - 0x3 -- Background 0x68
    "00000001", -- 2881 - 0xb41  :    1 - 0x1
    "00000000", -- 2882 - 0xb42  :    0 - 0x0
    "00000000", -- 2883 - 0xb43  :    0 - 0x0
    "00000000", -- 2884 - 0xb44  :    0 - 0x0
    "00000000", -- 2885 - 0xb45  :    0 - 0x0
    "00000000", -- 2886 - 0xb46  :    0 - 0x0
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "10000011", -- 2888 - 0xb48  :  131 - 0x83 -- Background 0x69
    "11010001", -- 2889 - 0xb49  :  209 - 0xd1
    "11100001", -- 2890 - 0xb4a  :  225 - 0xe1
    "11010001", -- 2891 - 0xb4b  :  209 - 0xd1
    "00000010", -- 2892 - 0xb4c  :    2 - 0x2
    "10000100", -- 2893 - 0xb4d  :  132 - 0x84
    "11110000", -- 2894 - 0xb4e  :  240 - 0xf0
    "11001110", -- 2895 - 0xb4f  :  206 - 0xce
    "11000000", -- 2896 - 0xb50  :  192 - 0xc0 -- Background 0x6a
    "10000000", -- 2897 - 0xb51  :  128 - 0x80
    "00000000", -- 2898 - 0xb52  :    0 - 0x0
    "00000000", -- 2899 - 0xb53  :    0 - 0x0
    "00000000", -- 2900 - 0xb54  :    0 - 0x0
    "00000000", -- 2901 - 0xb55  :    0 - 0x0
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "11000001", -- 2904 - 0xb58  :  193 - 0xc1 -- Background 0x6b
    "10001011", -- 2905 - 0xb59  :  139 - 0x8b
    "10000111", -- 2906 - 0xb5a  :  135 - 0x87
    "10001011", -- 2907 - 0xb5b  :  139 - 0x8b
    "01000000", -- 2908 - 0xb5c  :   64 - 0x40
    "00100001", -- 2909 - 0xb5d  :   33 - 0x21
    "00001111", -- 2910 - 0xb5e  :   15 - 0xf
    "11010011", -- 2911 - 0xb5f  :  211 - 0xd3
    "11111111", -- 2912 - 0xb60  :  255 - 0xff -- Background 0x6c
    "11111111", -- 2913 - 0xb61  :  255 - 0xff
    "11111111", -- 2914 - 0xb62  :  255 - 0xff
    "00011111", -- 2915 - 0xb63  :   31 - 0x1f
    "00001111", -- 2916 - 0xb64  :   15 - 0xf
    "00011110", -- 2917 - 0xb65  :   30 - 0x1e
    "00111111", -- 2918 - 0xb66  :   63 - 0x3f
    "01111111", -- 2919 - 0xb67  :  127 - 0x7f
    "11111111", -- 2920 - 0xb68  :  255 - 0xff -- Background 0x6d
    "11111111", -- 2921 - 0xb69  :  255 - 0xff
    "11111111", -- 2922 - 0xb6a  :  255 - 0xff
    "11111000", -- 2923 - 0xb6b  :  248 - 0xf8
    "11110000", -- 2924 - 0xb6c  :  240 - 0xf0
    "01111000", -- 2925 - 0xb6d  :  120 - 0x78
    "11111100", -- 2926 - 0xb6e  :  252 - 0xfc
    "11111110", -- 2927 - 0xb6f  :  254 - 0xfe
    "00000000", -- 2928 - 0xb70  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 2929 - 0xb71  :    0 - 0x0
    "00000000", -- 2930 - 0xb72  :    0 - 0x0
    "00000000", -- 2931 - 0xb73  :    0 - 0x0
    "00000000", -- 2932 - 0xb74  :    0 - 0x0
    "00111100", -- 2933 - 0xb75  :   60 - 0x3c
    "01000010", -- 2934 - 0xb76  :   66 - 0x42
    "10000001", -- 2935 - 0xb77  :  129 - 0x81
    "10000001", -- 2936 - 0xb78  :  129 - 0x81 -- Background 0x6f
    "10111101", -- 2937 - 0xb79  :  189 - 0xbd
    "01111110", -- 2938 - 0xb7a  :  126 - 0x7e
    "11111111", -- 2939 - 0xb7b  :  255 - 0xff
    "11100111", -- 2940 - 0xb7c  :  231 - 0xe7
    "11111111", -- 2941 - 0xb7d  :  255 - 0xff
    "11111111", -- 2942 - 0xb7e  :  255 - 0xff
    "11111111", -- 2943 - 0xb7f  :  255 - 0xff
    "00000001", -- 2944 - 0xb80  :    1 - 0x1 -- Background 0x70
    "00000111", -- 2945 - 0xb81  :    7 - 0x7
    "00011111", -- 2946 - 0xb82  :   31 - 0x1f
    "00111111", -- 2947 - 0xb83  :   63 - 0x3f
    "01111111", -- 2948 - 0xb84  :  127 - 0x7f
    "11111111", -- 2949 - 0xb85  :  255 - 0xff
    "11111111", -- 2950 - 0xb86  :  255 - 0xff
    "11011101", -- 2951 - 0xb87  :  221 - 0xdd
    "10001001", -- 2952 - 0xb88  :  137 - 0x89 -- Background 0x71
    "00000001", -- 2953 - 0xb89  :    1 - 0x1
    "00000001", -- 2954 - 0xb8a  :    1 - 0x1
    "00000001", -- 2955 - 0xb8b  :    1 - 0x1
    "00000001", -- 2956 - 0xb8c  :    1 - 0x1
    "00000001", -- 2957 - 0xb8d  :    1 - 0x1
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "10000000", -- 2960 - 0xb90  :  128 - 0x80 -- Background 0x72
    "11100000", -- 2961 - 0xb91  :  224 - 0xe0
    "11111000", -- 2962 - 0xb92  :  248 - 0xf8
    "11111100", -- 2963 - 0xb93  :  252 - 0xfc
    "11111110", -- 2964 - 0xb94  :  254 - 0xfe
    "11111111", -- 2965 - 0xb95  :  255 - 0xff
    "11111111", -- 2966 - 0xb96  :  255 - 0xff
    "00111011", -- 2967 - 0xb97  :   59 - 0x3b
    "00010001", -- 2968 - 0xb98  :   17 - 0x11 -- Background 0x73
    "00000000", -- 2969 - 0xb99  :    0 - 0x0
    "00000000", -- 2970 - 0xb9a  :    0 - 0x0
    "00000000", -- 2971 - 0xb9b  :    0 - 0x0
    "00000000", -- 2972 - 0xb9c  :    0 - 0x0
    "01000000", -- 2973 - 0xb9d  :   64 - 0x40
    "10000000", -- 2974 - 0xb9e  :  128 - 0x80
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "00000001", -- 2976 - 0xba0  :    1 - 0x1 -- Background 0x74
    "00000001", -- 2977 - 0xba1  :    1 - 0x1
    "00000001", -- 2978 - 0xba2  :    1 - 0x1
    "00000001", -- 2979 - 0xba3  :    1 - 0x1
    "00000001", -- 2980 - 0xba4  :    1 - 0x1
    "00000001", -- 2981 - 0xba5  :    1 - 0x1
    "00000001", -- 2982 - 0xba6  :    1 - 0x1
    "00000001", -- 2983 - 0xba7  :    1 - 0x1
    "10000000", -- 2984 - 0xba8  :  128 - 0x80 -- Background 0x75
    "10000000", -- 2985 - 0xba9  :  128 - 0x80
    "10000000", -- 2986 - 0xbaa  :  128 - 0x80
    "10000000", -- 2987 - 0xbab  :  128 - 0x80
    "10000000", -- 2988 - 0xbac  :  128 - 0x80
    "10000000", -- 2989 - 0xbad  :  128 - 0x80
    "10000000", -- 2990 - 0xbae  :  128 - 0x80
    "10000000", -- 2991 - 0xbaf  :  128 - 0x80
    "00000001", -- 2992 - 0xbb0  :    1 - 0x1 -- Background 0x76
    "00000011", -- 2993 - 0xbb1  :    3 - 0x3
    "00000000", -- 2994 - 0xbb2  :    0 - 0x0
    "00000000", -- 2995 - 0xbb3  :    0 - 0x0
    "00000011", -- 2996 - 0xbb4  :    3 - 0x3
    "00011001", -- 2997 - 0xbb5  :   25 - 0x19
    "00000000", -- 2998 - 0xbb6  :    0 - 0x0
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "00000000", -- 3000 - 0xbb8  :    0 - 0x0 -- Background 0x77
    "00000000", -- 3001 - 0xbb9  :    0 - 0x0
    "01111100", -- 3002 - 0xbba  :  124 - 0x7c
    "00000010", -- 3003 - 0xbbb  :    2 - 0x2
    "00000001", -- 3004 - 0xbbc  :    1 - 0x1
    "00000000", -- 3005 - 0xbbd  :    0 - 0x0
    "00000000", -- 3006 - 0xbbe  :    0 - 0x0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Background 0x78
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000001", -- 3010 - 0xbc2  :    1 - 0x1
    "00000001", -- 3011 - 0xbc3  :    1 - 0x1
    "00000011", -- 3012 - 0xbc4  :    3 - 0x3
    "00000111", -- 3013 - 0xbc5  :    7 - 0x7
    "00000111", -- 3014 - 0xbc6  :    7 - 0x7
    "00001111", -- 3015 - 0xbc7  :   15 - 0xf
    "00001111", -- 3016 - 0xbc8  :   15 - 0xf -- Background 0x79
    "00000111", -- 3017 - 0xbc9  :    7 - 0x7
    "00001111", -- 3018 - 0xbca  :   15 - 0xf
    "00000111", -- 3019 - 0xbcb  :    7 - 0x7
    "00000001", -- 3020 - 0xbcc  :    1 - 0x1
    "00010000", -- 3021 - 0xbcd  :   16 - 0x10
    "00100000", -- 3022 - 0xbce  :   32 - 0x20
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "11111000", -- 3024 - 0xbd0  :  248 - 0xf8 -- Background 0x7a
    "11111110", -- 3025 - 0xbd1  :  254 - 0xfe
    "01111111", -- 3026 - 0xbd2  :  127 - 0x7f
    "00011111", -- 3027 - 0xbd3  :   31 - 0x1f
    "00001111", -- 3028 - 0xbd4  :   15 - 0xf
    "00011001", -- 3029 - 0xbd5  :   25 - 0x19
    "00110000", -- 3030 - 0xbd6  :   48 - 0x30
    "01110000", -- 3031 - 0xbd7  :  112 - 0x70
    "11111011", -- 3032 - 0xbd8  :  251 - 0xfb -- Background 0x7b
    "01110011", -- 3033 - 0xbd9  :  115 - 0x73
    "00100111", -- 3034 - 0xbda  :   39 - 0x27
    "00001111", -- 3035 - 0xbdb  :   15 - 0xf
    "00011111", -- 3036 - 0xbdc  :   31 - 0x1f
    "00011111", -- 3037 - 0xbdd  :   31 - 0x1f
    "00111111", -- 3038 - 0xbde  :   63 - 0x3f
    "01111111", -- 3039 - 0xbdf  :  127 - 0x7f
    "11111111", -- 3040 - 0xbe0  :  255 - 0xff -- Background 0x7c
    "11111111", -- 3041 - 0xbe1  :  255 - 0xff
    "11111111", -- 3042 - 0xbe2  :  255 - 0xff
    "11111111", -- 3043 - 0xbe3  :  255 - 0xff
    "11111110", -- 3044 - 0xbe4  :  254 - 0xfe
    "11111101", -- 3045 - 0xbe5  :  253 - 0xfd
    "11111000", -- 3046 - 0xbe6  :  248 - 0xf8
    "11110110", -- 3047 - 0xbe7  :  246 - 0xf6
    "11101111", -- 3048 - 0xbe8  :  239 - 0xef -- Background 0x7d
    "11001111", -- 3049 - 0xbe9  :  207 - 0xcf
    "10011111", -- 3050 - 0xbea  :  159 - 0x9f
    "00011111", -- 3051 - 0xbeb  :   31 - 0x1f
    "00001111", -- 3052 - 0xbec  :   15 - 0xf
    "00101101", -- 3053 - 0xbed  :   45 - 0x2d
    "01010000", -- 3054 - 0xbee  :   80 - 0x50
    "01000000", -- 3055 - 0xbef  :   64 - 0x40
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00000000", -- 3058 - 0xbf2  :    0 - 0x0
    "00000000", -- 3059 - 0xbf3  :    0 - 0x0
    "11100000", -- 3060 - 0xbf4  :  224 - 0xe0
    "11111110", -- 3061 - 0xbf5  :  254 - 0xfe
    "11111111", -- 3062 - 0xbf6  :  255 - 0xff
    "11110011", -- 3063 - 0xbf7  :  243 - 0xf3
    "11111011", -- 3064 - 0xbf8  :  251 - 0xfb -- Background 0x7f
    "11111011", -- 3065 - 0xbf9  :  251 - 0xfb
    "11111011", -- 3066 - 0xbfa  :  251 - 0xfb
    "11111011", -- 3067 - 0xbfb  :  251 - 0xfb
    "11111011", -- 3068 - 0xbfc  :  251 - 0xfb
    "11110011", -- 3069 - 0xbfd  :  243 - 0xf3
    "11110111", -- 3070 - 0xbfe  :  247 - 0xf7
    "11100111", -- 3071 - 0xbff  :  231 - 0xe7
    "11001111", -- 3072 - 0xc00  :  207 - 0xcf -- Background 0x80
    "10011111", -- 3073 - 0xc01  :  159 - 0x9f
    "00111111", -- 3074 - 0xc02  :   63 - 0x3f
    "00111111", -- 3075 - 0xc03  :   63 - 0x3f
    "00111111", -- 3076 - 0xc04  :   63 - 0x3f
    "00001111", -- 3077 - 0xc05  :   15 - 0xf
    "00000011", -- 3078 - 0xc06  :    3 - 0x3
    "00000000", -- 3079 - 0xc07  :    0 - 0x0
    "11000000", -- 3080 - 0xc08  :  192 - 0xc0 -- Background 0x81
    "11110000", -- 3081 - 0xc09  :  240 - 0xf0
    "11111100", -- 3082 - 0xc0a  :  252 - 0xfc
    "11110000", -- 3083 - 0xc0b  :  240 - 0xf0
    "11110000", -- 3084 - 0xc0c  :  240 - 0xf0
    "10011000", -- 3085 - 0xc0d  :  152 - 0x98
    "00001000", -- 3086 - 0xc0e  :    8 - 0x8
    "00000000", -- 3087 - 0xc0f  :    0 - 0x0
    "00000000", -- 3088 - 0xc10  :    0 - 0x0 -- Background 0x82
    "00000000", -- 3089 - 0xc11  :    0 - 0x0
    "00000000", -- 3090 - 0xc12  :    0 - 0x0
    "00000000", -- 3091 - 0xc13  :    0 - 0x0
    "00000000", -- 3092 - 0xc14  :    0 - 0x0
    "00000000", -- 3093 - 0xc15  :    0 - 0x0
    "10000000", -- 3094 - 0xc16  :  128 - 0x80
    "11000000", -- 3095 - 0xc17  :  192 - 0xc0
    "11100000", -- 3096 - 0xc18  :  224 - 0xe0 -- Background 0x83
    "11100000", -- 3097 - 0xc19  :  224 - 0xe0
    "11110000", -- 3098 - 0xc1a  :  240 - 0xf0
    "11110000", -- 3099 - 0xc1b  :  240 - 0xf0
    "11110000", -- 3100 - 0xc1c  :  240 - 0xf0
    "11110000", -- 3101 - 0xc1d  :  240 - 0xf0
    "11111000", -- 3102 - 0xc1e  :  248 - 0xf8
    "11111000", -- 3103 - 0xc1f  :  248 - 0xf8
    "11111110", -- 3104 - 0xc20  :  254 - 0xfe -- Background 0x84
    "11111111", -- 3105 - 0xc21  :  255 - 0xff
    "11111111", -- 3106 - 0xc22  :  255 - 0xff
    "11111111", -- 3107 - 0xc23  :  255 - 0xff
    "11111111", -- 3108 - 0xc24  :  255 - 0xff
    "11111111", -- 3109 - 0xc25  :  255 - 0xff
    "11111111", -- 3110 - 0xc26  :  255 - 0xff
    "11111111", -- 3111 - 0xc27  :  255 - 0xff
    "00111111", -- 3112 - 0xc28  :   63 - 0x3f -- Background 0x85
    "00011111", -- 3113 - 0xc29  :   31 - 0x1f
    "00011111", -- 3114 - 0xc2a  :   31 - 0x1f
    "00001111", -- 3115 - 0xc2b  :   15 - 0xf
    "00000111", -- 3116 - 0xc2c  :    7 - 0x7
    "00000000", -- 3117 - 0xc2d  :    0 - 0x0
    "00000000", -- 3118 - 0xc2e  :    0 - 0x0
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "00000000", -- 3120 - 0xc30  :    0 - 0x0 -- Background 0x86
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "11000000", -- 3122 - 0xc32  :  192 - 0xc0
    "11100000", -- 3123 - 0xc33  :  224 - 0xe0
    "11110000", -- 3124 - 0xc34  :  240 - 0xf0
    "11110000", -- 3125 - 0xc35  :  240 - 0xf0
    "11110000", -- 3126 - 0xc36  :  240 - 0xf0
    "11111000", -- 3127 - 0xc37  :  248 - 0xf8
    "11111001", -- 3128 - 0xc38  :  249 - 0xf9 -- Background 0x87
    "11111111", -- 3129 - 0xc39  :  255 - 0xff
    "11111111", -- 3130 - 0xc3a  :  255 - 0xff
    "11111111", -- 3131 - 0xc3b  :  255 - 0xff
    "11111111", -- 3132 - 0xc3c  :  255 - 0xff
    "00001110", -- 3133 - 0xc3d  :   14 - 0xe
    "00000010", -- 3134 - 0xc3e  :    2 - 0x2
    "00010100", -- 3135 - 0xc3f  :   20 - 0x14
    "10000000", -- 3136 - 0xc40  :  128 - 0x80 -- Background 0x88
    "10100000", -- 3137 - 0xc41  :  160 - 0xa0
    "00100000", -- 3138 - 0xc42  :   32 - 0x20
    "00100000", -- 3139 - 0xc43  :   32 - 0x20
    "10100000", -- 3140 - 0xc44  :  160 - 0xa0
    "10000000", -- 3141 - 0xc45  :  128 - 0x80
    "00000000", -- 3142 - 0xc46  :    0 - 0x0
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00000001", -- 3144 - 0xc48  :    1 - 0x1 -- Background 0x89
    "00000101", -- 3145 - 0xc49  :    5 - 0x5
    "00000100", -- 3146 - 0xc4a  :    4 - 0x4
    "00000100", -- 3147 - 0xc4b  :    4 - 0x4
    "00000101", -- 3148 - 0xc4c  :    5 - 0x5
    "00000001", -- 3149 - 0xc4d  :    1 - 0x1
    "00000000", -- 3150 - 0xc4e  :    0 - 0x0
    "00000000", -- 3151 - 0xc4f  :    0 - 0x0
    "00000000", -- 3152 - 0xc50  :    0 - 0x0 -- Background 0x8a
    "00000000", -- 3153 - 0xc51  :    0 - 0x0
    "00000011", -- 3154 - 0xc52  :    3 - 0x3
    "00000111", -- 3155 - 0xc53  :    7 - 0x7
    "00001111", -- 3156 - 0xc54  :   15 - 0xf
    "00001111", -- 3157 - 0xc55  :   15 - 0xf
    "00001111", -- 3158 - 0xc56  :   15 - 0xf
    "00001111", -- 3159 - 0xc57  :   15 - 0xf
    "10011111", -- 3160 - 0xc58  :  159 - 0x9f -- Background 0x8b
    "11111111", -- 3161 - 0xc59  :  255 - 0xff
    "11111111", -- 3162 - 0xc5a  :  255 - 0xff
    "11111111", -- 3163 - 0xc5b  :  255 - 0xff
    "11111111", -- 3164 - 0xc5c  :  255 - 0xff
    "01110000", -- 3165 - 0xc5d  :  112 - 0x70
    "01000000", -- 3166 - 0xc5e  :   64 - 0x40
    "00101000", -- 3167 - 0xc5f  :   40 - 0x28
    "00000000", -- 3168 - 0xc60  :    0 - 0x0 -- Background 0x8c
    "00000000", -- 3169 - 0xc61  :    0 - 0x0
    "00000000", -- 3170 - 0xc62  :    0 - 0x0
    "00000000", -- 3171 - 0xc63  :    0 - 0x0
    "00000000", -- 3172 - 0xc64  :    0 - 0x0
    "00000000", -- 3173 - 0xc65  :    0 - 0x0
    "00000001", -- 3174 - 0xc66  :    1 - 0x1
    "00000011", -- 3175 - 0xc67  :    3 - 0x3
    "00000111", -- 3176 - 0xc68  :    7 - 0x7 -- Background 0x8d
    "00000111", -- 3177 - 0xc69  :    7 - 0x7
    "00001111", -- 3178 - 0xc6a  :   15 - 0xf
    "00001111", -- 3179 - 0xc6b  :   15 - 0xf
    "00001111", -- 3180 - 0xc6c  :   15 - 0xf
    "00001111", -- 3181 - 0xc6d  :   15 - 0xf
    "00011111", -- 3182 - 0xc6e  :   31 - 0x1f
    "00011111", -- 3183 - 0xc6f  :   31 - 0x1f
    "01111111", -- 3184 - 0xc70  :  127 - 0x7f -- Background 0x8e
    "11111111", -- 3185 - 0xc71  :  255 - 0xff
    "11111111", -- 3186 - 0xc72  :  255 - 0xff
    "11111111", -- 3187 - 0xc73  :  255 - 0xff
    "11111111", -- 3188 - 0xc74  :  255 - 0xff
    "11111111", -- 3189 - 0xc75  :  255 - 0xff
    "11111111", -- 3190 - 0xc76  :  255 - 0xff
    "11111111", -- 3191 - 0xc77  :  255 - 0xff
    "11111100", -- 3192 - 0xc78  :  252 - 0xfc -- Background 0x8f
    "11111000", -- 3193 - 0xc79  :  248 - 0xf8
    "11111000", -- 3194 - 0xc7a  :  248 - 0xf8
    "11110000", -- 3195 - 0xc7b  :  240 - 0xf0
    "11100000", -- 3196 - 0xc7c  :  224 - 0xe0
    "00000000", -- 3197 - 0xc7d  :    0 - 0x0
    "00000000", -- 3198 - 0xc7e  :    0 - 0x0
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Background 0x90
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000111", -- 3204 - 0xc84  :    7 - 0x7
    "01111111", -- 3205 - 0xc85  :  127 - 0x7f
    "11111111", -- 3206 - 0xc86  :  255 - 0xff
    "11001111", -- 3207 - 0xc87  :  207 - 0xcf
    "11011111", -- 3208 - 0xc88  :  223 - 0xdf -- Background 0x91
    "11011111", -- 3209 - 0xc89  :  223 - 0xdf
    "11011111", -- 3210 - 0xc8a  :  223 - 0xdf
    "11011111", -- 3211 - 0xc8b  :  223 - 0xdf
    "11011111", -- 3212 - 0xc8c  :  223 - 0xdf
    "11001111", -- 3213 - 0xc8d  :  207 - 0xcf
    "11101111", -- 3214 - 0xc8e  :  239 - 0xef
    "11100111", -- 3215 - 0xc8f  :  231 - 0xe7
    "11110011", -- 3216 - 0xc90  :  243 - 0xf3 -- Background 0x92
    "11111001", -- 3217 - 0xc91  :  249 - 0xf9
    "11111100", -- 3218 - 0xc92  :  252 - 0xfc
    "11111100", -- 3219 - 0xc93  :  252 - 0xfc
    "11111100", -- 3220 - 0xc94  :  252 - 0xfc
    "11110000", -- 3221 - 0xc95  :  240 - 0xf0
    "11000000", -- 3222 - 0xc96  :  192 - 0xc0
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "00000011", -- 3224 - 0xc98  :    3 - 0x3 -- Background 0x93
    "00001111", -- 3225 - 0xc99  :   15 - 0xf
    "00111111", -- 3226 - 0xc9a  :   63 - 0x3f
    "00001111", -- 3227 - 0xc9b  :   15 - 0xf
    "00001111", -- 3228 - 0xc9c  :   15 - 0xf
    "00011001", -- 3229 - 0xc9d  :   25 - 0x19
    "00010000", -- 3230 - 0xc9e  :   16 - 0x10
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00011111", -- 3232 - 0xca0  :   31 - 0x1f -- Background 0x94
    "01111111", -- 3233 - 0xca1  :  127 - 0x7f
    "11111110", -- 3234 - 0xca2  :  254 - 0xfe
    "11111000", -- 3235 - 0xca3  :  248 - 0xf8
    "11110000", -- 3236 - 0xca4  :  240 - 0xf0
    "10011000", -- 3237 - 0xca5  :  152 - 0x98
    "00001100", -- 3238 - 0xca6  :   12 - 0xc
    "00001110", -- 3239 - 0xca7  :   14 - 0xe
    "11011111", -- 3240 - 0xca8  :  223 - 0xdf -- Background 0x95
    "11001110", -- 3241 - 0xca9  :  206 - 0xce
    "11100100", -- 3242 - 0xcaa  :  228 - 0xe4
    "11110000", -- 3243 - 0xcab  :  240 - 0xf0
    "11111000", -- 3244 - 0xcac  :  248 - 0xf8
    "11111000", -- 3245 - 0xcad  :  248 - 0xf8
    "11111100", -- 3246 - 0xcae  :  252 - 0xfc
    "11111110", -- 3247 - 0xcaf  :  254 - 0xfe
    "11111111", -- 3248 - 0xcb0  :  255 - 0xff -- Background 0x96
    "11111111", -- 3249 - 0xcb1  :  255 - 0xff
    "11111111", -- 3250 - 0xcb2  :  255 - 0xff
    "11111111", -- 3251 - 0xcb3  :  255 - 0xff
    "01111111", -- 3252 - 0xcb4  :  127 - 0x7f
    "10111111", -- 3253 - 0xcb5  :  191 - 0xbf
    "00011111", -- 3254 - 0xcb6  :   31 - 0x1f
    "01101111", -- 3255 - 0xcb7  :  111 - 0x6f
    "11110111", -- 3256 - 0xcb8  :  247 - 0xf7 -- Background 0x97
    "11110011", -- 3257 - 0xcb9  :  243 - 0xf3
    "11111001", -- 3258 - 0xcba  :  249 - 0xf9
    "11111000", -- 3259 - 0xcbb  :  248 - 0xf8
    "11110000", -- 3260 - 0xcbc  :  240 - 0xf0
    "10110100", -- 3261 - 0xcbd  :  180 - 0xb4
    "00001010", -- 3262 - 0xcbe  :   10 - 0xa
    "00000010", -- 3263 - 0xcbf  :    2 - 0x2
    "10000000", -- 3264 - 0xcc0  :  128 - 0x80 -- Background 0x98
    "11000000", -- 3265 - 0xcc1  :  192 - 0xc0
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "00000000", -- 3267 - 0xcc3  :    0 - 0x0
    "11000000", -- 3268 - 0xcc4  :  192 - 0xc0
    "10011000", -- 3269 - 0xcc5  :  152 - 0x98
    "00000000", -- 3270 - 0xcc6  :    0 - 0x0
    "00000000", -- 3271 - 0xcc7  :    0 - 0x0
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0 -- Background 0x99
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00111110", -- 3274 - 0xcca  :   62 - 0x3e
    "01000000", -- 3275 - 0xccb  :   64 - 0x40
    "10000000", -- 3276 - 0xccc  :  128 - 0x80
    "00000000", -- 3277 - 0xccd  :    0 - 0x0
    "00000000", -- 3278 - 0xcce  :    0 - 0x0
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0 -- Background 0x9a
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "10000000", -- 3282 - 0xcd2  :  128 - 0x80
    "10000000", -- 3283 - 0xcd3  :  128 - 0x80
    "11000000", -- 3284 - 0xcd4  :  192 - 0xc0
    "11100000", -- 3285 - 0xcd5  :  224 - 0xe0
    "11100000", -- 3286 - 0xcd6  :  224 - 0xe0
    "11110000", -- 3287 - 0xcd7  :  240 - 0xf0
    "11110000", -- 3288 - 0xcd8  :  240 - 0xf0 -- Background 0x9b
    "11100000", -- 3289 - 0xcd9  :  224 - 0xe0
    "11110000", -- 3290 - 0xcda  :  240 - 0xf0
    "11100000", -- 3291 - 0xcdb  :  224 - 0xe0
    "10000000", -- 3292 - 0xcdc  :  128 - 0x80
    "00001000", -- 3293 - 0xcdd  :    8 - 0x8
    "00000100", -- 3294 - 0xcde  :    4 - 0x4
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Background 0x9c
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000001", -- 3298 - 0xce2  :    1 - 0x1
    "00000011", -- 3299 - 0xce3  :    3 - 0x3
    "00000011", -- 3300 - 0xce4  :    3 - 0x3
    "00000011", -- 3301 - 0xce5  :    3 - 0x3
    "00000111", -- 3302 - 0xce6  :    7 - 0x7
    "00000111", -- 3303 - 0xce7  :    7 - 0x7
    "00000111", -- 3304 - 0xce8  :    7 - 0x7 -- Background 0x9d
    "00000011", -- 3305 - 0xce9  :    3 - 0x3
    "00000011", -- 3306 - 0xcea  :    3 - 0x3
    "00000011", -- 3307 - 0xceb  :    3 - 0x3
    "00000011", -- 3308 - 0xcec  :    3 - 0x3
    "00000011", -- 3309 - 0xced  :    3 - 0x3
    "00000011", -- 3310 - 0xcee  :    3 - 0x3
    "00000001", -- 3311 - 0xcef  :    1 - 0x1
    "00000000", -- 3312 - 0xcf0  :    0 - 0x0 -- Background 0x9e
    "00000000", -- 3313 - 0xcf1  :    0 - 0x0
    "00000000", -- 3314 - 0xcf2  :    0 - 0x0
    "00000000", -- 3315 - 0xcf3  :    0 - 0x0
    "00000000", -- 3316 - 0xcf4  :    0 - 0x0
    "00000001", -- 3317 - 0xcf5  :    1 - 0x1
    "00000010", -- 3318 - 0xcf6  :    2 - 0x2
    "00000100", -- 3319 - 0xcf7  :    4 - 0x4
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0 -- Background 0x9f
    "00000000", -- 3321 - 0xcf9  :    0 - 0x0
    "00000000", -- 3322 - 0xcfa  :    0 - 0x0
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00011100", -- 3326 - 0xcfe  :   28 - 0x1c
    "00111011", -- 3327 - 0xcff  :   59 - 0x3b
    "01111110", -- 3328 - 0xd00  :  126 - 0x7e -- Background 0xa0
    "11111110", -- 3329 - 0xd01  :  254 - 0xfe
    "11111111", -- 3330 - 0xd02  :  255 - 0xff
    "11111111", -- 3331 - 0xd03  :  255 - 0xff
    "11111111", -- 3332 - 0xd04  :  255 - 0xff
    "11111111", -- 3333 - 0xd05  :  255 - 0xff
    "11111101", -- 3334 - 0xd06  :  253 - 0xfd
    "11111001", -- 3335 - 0xd07  :  249 - 0xf9
    "11110011", -- 3336 - 0xd08  :  243 - 0xf3 -- Background 0xa1
    "11110111", -- 3337 - 0xd09  :  247 - 0xf7
    "11110110", -- 3338 - 0xd0a  :  246 - 0xf6
    "11101110", -- 3339 - 0xd0b  :  238 - 0xee
    "11111101", -- 3340 - 0xd0c  :  253 - 0xfd
    "11111100", -- 3341 - 0xd0d  :  252 - 0xfc
    "11111000", -- 3342 - 0xd0e  :  248 - 0xf8
    "11100001", -- 3343 - 0xd0f  :  225 - 0xe1
    "11010011", -- 3344 - 0xd10  :  211 - 0xd3 -- Background 0xa2
    "11001011", -- 3345 - 0xd11  :  203 - 0xcb
    "11000011", -- 3346 - 0xd12  :  195 - 0xc3
    "11100001", -- 3347 - 0xd13  :  225 - 0xe1
    "11111001", -- 3348 - 0xd14  :  249 - 0xf9
    "00111001", -- 3349 - 0xd15  :   57 - 0x39
    "01000010", -- 3350 - 0xd16  :   66 - 0x42
    "00000000", -- 3351 - 0xd17  :    0 - 0x0
    "00000111", -- 3352 - 0xd18  :    7 - 0x7 -- Background 0xa3
    "00001111", -- 3353 - 0xd19  :   15 - 0xf
    "00011001", -- 3354 - 0xd1a  :   25 - 0x19
    "00110000", -- 3355 - 0xd1b  :   48 - 0x30
    "01100011", -- 3356 - 0xd1c  :   99 - 0x63
    "01110010", -- 3357 - 0xd1d  :  114 - 0x72
    "01110000", -- 3358 - 0xd1e  :  112 - 0x70
    "00000001", -- 3359 - 0xd1f  :    1 - 0x1
    "00000000", -- 3360 - 0xd20  :    0 - 0x0 -- Background 0xa4
    "00011111", -- 3361 - 0xd21  :   31 - 0x1f
    "00100000", -- 3362 - 0xd22  :   32 - 0x20
    "11000000", -- 3363 - 0xd23  :  192 - 0xc0
    "11000000", -- 3364 - 0xd24  :  192 - 0xc0
    "11110000", -- 3365 - 0xd25  :  240 - 0xf0
    "11111111", -- 3366 - 0xd26  :  255 - 0xff
    "11111111", -- 3367 - 0xd27  :  255 - 0xff
    "10101011", -- 3368 - 0xd28  :  171 - 0xab -- Background 0xa5
    "11000001", -- 3369 - 0xd29  :  193 - 0xc1
    "10000001", -- 3370 - 0xd2a  :  129 - 0x81
    "10010001", -- 3371 - 0xd2b  :  145 - 0x91
    "10000010", -- 3372 - 0xd2c  :  130 - 0x82
    "11111100", -- 3373 - 0xd2d  :  252 - 0xfc
    "11100000", -- 3374 - 0xd2e  :  224 - 0xe0
    "11001110", -- 3375 - 0xd2f  :  206 - 0xce
    "11100101", -- 3376 - 0xd30  :  229 - 0xe5 -- Background 0xa6
    "11011010", -- 3377 - 0xd31  :  218 - 0xda
    "11110000", -- 3378 - 0xd32  :  240 - 0xf0
    "11100000", -- 3379 - 0xd33  :  224 - 0xe0
    "11000000", -- 3380 - 0xd34  :  192 - 0xc0
    "00000000", -- 3381 - 0xd35  :    0 - 0x0
    "00000000", -- 3382 - 0xd36  :    0 - 0x0
    "00000000", -- 3383 - 0xd37  :    0 - 0x0
    "11110000", -- 3384 - 0xd38  :  240 - 0xf0 -- Background 0xa7
    "11111000", -- 3385 - 0xd39  :  248 - 0xf8
    "11001100", -- 3386 - 0xd3a  :  204 - 0xcc
    "10000110", -- 3387 - 0xd3b  :  134 - 0x86
    "01100010", -- 3388 - 0xd3c  :   98 - 0x62
    "00100110", -- 3389 - 0xd3d  :   38 - 0x26
    "00000110", -- 3390 - 0xd3e  :    6 - 0x6
    "11000000", -- 3391 - 0xd3f  :  192 - 0xc0
    "00000000", -- 3392 - 0xd40  :    0 - 0x0 -- Background 0xa8
    "11111100", -- 3393 - 0xd41  :  252 - 0xfc
    "00000110", -- 3394 - 0xd42  :    6 - 0x6
    "00000011", -- 3395 - 0xd43  :    3 - 0x3
    "00000001", -- 3396 - 0xd44  :    1 - 0x1
    "00000111", -- 3397 - 0xd45  :    7 - 0x7
    "11111111", -- 3398 - 0xd46  :  255 - 0xff
    "11111111", -- 3399 - 0xd47  :  255 - 0xff
    "11010101", -- 3400 - 0xd48  :  213 - 0xd5 -- Background 0xa9
    "10000011", -- 3401 - 0xd49  :  131 - 0x83
    "10000001", -- 3402 - 0xd4a  :  129 - 0x81
    "10001001", -- 3403 - 0xd4b  :  137 - 0x89
    "01000001", -- 3404 - 0xd4c  :   65 - 0x41
    "00111111", -- 3405 - 0xd4d  :   63 - 0x3f
    "00000111", -- 3406 - 0xd4e  :    7 - 0x7
    "11010011", -- 3407 - 0xd4f  :  211 - 0xd3
    "01101111", -- 3408 - 0xd50  :  111 - 0x6f -- Background 0xaa
    "11011011", -- 3409 - 0xd51  :  219 - 0xdb
    "00001111", -- 3410 - 0xd52  :   15 - 0xf
    "00000111", -- 3411 - 0xd53  :    7 - 0x7
    "00000011", -- 3412 - 0xd54  :    3 - 0x3
    "00000000", -- 3413 - 0xd55  :    0 - 0x0
    "00000000", -- 3414 - 0xd56  :    0 - 0x0
    "00000000", -- 3415 - 0xd57  :    0 - 0x0
    "00000000", -- 3416 - 0xd58  :    0 - 0x0 -- Background 0xab
    "00000000", -- 3417 - 0xd59  :    0 - 0x0
    "00000000", -- 3418 - 0xd5a  :    0 - 0x0
    "00000000", -- 3419 - 0xd5b  :    0 - 0x0
    "00000000", -- 3420 - 0xd5c  :    0 - 0x0
    "00000000", -- 3421 - 0xd5d  :    0 - 0x0
    "00111000", -- 3422 - 0xd5e  :   56 - 0x38
    "11011100", -- 3423 - 0xd5f  :  220 - 0xdc
    "01111110", -- 3424 - 0xd60  :  126 - 0x7e -- Background 0xac
    "01111111", -- 3425 - 0xd61  :  127 - 0x7f
    "01111111", -- 3426 - 0xd62  :  127 - 0x7f
    "11111111", -- 3427 - 0xd63  :  255 - 0xff
    "11111111", -- 3428 - 0xd64  :  255 - 0xff
    "11111111", -- 3429 - 0xd65  :  255 - 0xff
    "10111111", -- 3430 - 0xd66  :  191 - 0xbf
    "10011111", -- 3431 - 0xd67  :  159 - 0x9f
    "11001111", -- 3432 - 0xd68  :  207 - 0xcf -- Background 0xad
    "11101111", -- 3433 - 0xd69  :  239 - 0xef
    "01101111", -- 3434 - 0xd6a  :  111 - 0x6f
    "01110111", -- 3435 - 0xd6b  :  119 - 0x77
    "10111111", -- 3436 - 0xd6c  :  191 - 0xbf
    "00111111", -- 3437 - 0xd6d  :   63 - 0x3f
    "00011111", -- 3438 - 0xd6e  :   31 - 0x1f
    "10000111", -- 3439 - 0xd6f  :  135 - 0x87
    "11001011", -- 3440 - 0xd70  :  203 - 0xcb -- Background 0xae
    "11010011", -- 3441 - 0xd71  :  211 - 0xd3
    "11000011", -- 3442 - 0xd72  :  195 - 0xc3
    "10000111", -- 3443 - 0xd73  :  135 - 0x87
    "10011111", -- 3444 - 0xd74  :  159 - 0x9f
    "10011100", -- 3445 - 0xd75  :  156 - 0x9c
    "01000010", -- 3446 - 0xd76  :   66 - 0x42
    "00000000", -- 3447 - 0xd77  :    0 - 0x0
    "00000000", -- 3448 - 0xd78  :    0 - 0x0 -- Background 0xaf
    "00000000", -- 3449 - 0xd79  :    0 - 0x0
    "10000000", -- 3450 - 0xd7a  :  128 - 0x80
    "11000000", -- 3451 - 0xd7b  :  192 - 0xc0
    "11000000", -- 3452 - 0xd7c  :  192 - 0xc0
    "11000000", -- 3453 - 0xd7d  :  192 - 0xc0
    "11100000", -- 3454 - 0xd7e  :  224 - 0xe0
    "11100000", -- 3455 - 0xd7f  :  224 - 0xe0
    "11100000", -- 3456 - 0xd80  :  224 - 0xe0 -- Background 0xb0
    "11000000", -- 3457 - 0xd81  :  192 - 0xc0
    "11000000", -- 3458 - 0xd82  :  192 - 0xc0
    "11000000", -- 3459 - 0xd83  :  192 - 0xc0
    "11000000", -- 3460 - 0xd84  :  192 - 0xc0
    "11000000", -- 3461 - 0xd85  :  192 - 0xc0
    "11000000", -- 3462 - 0xd86  :  192 - 0xc0
    "10000000", -- 3463 - 0xd87  :  128 - 0x80
    "00000000", -- 3464 - 0xd88  :    0 - 0x0 -- Background 0xb1
    "00000000", -- 3465 - 0xd89  :    0 - 0x0
    "00000000", -- 3466 - 0xd8a  :    0 - 0x0
    "00000000", -- 3467 - 0xd8b  :    0 - 0x0
    "00000000", -- 3468 - 0xd8c  :    0 - 0x0
    "10000000", -- 3469 - 0xd8d  :  128 - 0x80
    "01000000", -- 3470 - 0xd8e  :   64 - 0x40
    "00100000", -- 3471 - 0xd8f  :   32 - 0x20
    "00000000", -- 3472 - 0xd90  :    0 - 0x0 -- Background 0xb2
    "00000000", -- 3473 - 0xd91  :    0 - 0x0
    "00000000", -- 3474 - 0xd92  :    0 - 0x0
    "00000001", -- 3475 - 0xd93  :    1 - 0x1
    "00000011", -- 3476 - 0xd94  :    3 - 0x3
    "00000111", -- 3477 - 0xd95  :    7 - 0x7
    "00000111", -- 3478 - 0xd96  :    7 - 0x7
    "00000111", -- 3479 - 0xd97  :    7 - 0x7
    "00000011", -- 3480 - 0xd98  :    3 - 0x3 -- Background 0xb3
    "00000001", -- 3481 - 0xd99  :    1 - 0x1
    "00000000", -- 3482 - 0xd9a  :    0 - 0x0
    "00000000", -- 3483 - 0xd9b  :    0 - 0x0
    "00000000", -- 3484 - 0xd9c  :    0 - 0x0
    "00000000", -- 3485 - 0xd9d  :    0 - 0x0
    "00000001", -- 3486 - 0xd9e  :    1 - 0x1
    "00000001", -- 3487 - 0xd9f  :    1 - 0x1
    "00000001", -- 3488 - 0xda0  :    1 - 0x1 -- Background 0xb4
    "00000001", -- 3489 - 0xda1  :    1 - 0x1
    "00000111", -- 3490 - 0xda2  :    7 - 0x7
    "00000011", -- 3491 - 0xda3  :    3 - 0x3
    "00000100", -- 3492 - 0xda4  :    4 - 0x4
    "00000000", -- 3493 - 0xda5  :    0 - 0x0
    "00000000", -- 3494 - 0xda6  :    0 - 0x0
    "00000000", -- 3495 - 0xda7  :    0 - 0x0
    "00000000", -- 3496 - 0xda8  :    0 - 0x0 -- Background 0xb5
    "00000000", -- 3497 - 0xda9  :    0 - 0x0
    "00000000", -- 3498 - 0xdaa  :    0 - 0x0
    "00000000", -- 3499 - 0xdab  :    0 - 0x0
    "00000000", -- 3500 - 0xdac  :    0 - 0x0
    "00000000", -- 3501 - 0xdad  :    0 - 0x0
    "00000000", -- 3502 - 0xdae  :    0 - 0x0
    "00000111", -- 3503 - 0xdaf  :    7 - 0x7
    "00001110", -- 3504 - 0xdb0  :   14 - 0xe -- Background 0xb6
    "00111110", -- 3505 - 0xdb1  :   62 - 0x3e
    "01111111", -- 3506 - 0xdb2  :  127 - 0x7f
    "11111111", -- 3507 - 0xdb3  :  255 - 0xff
    "11111111", -- 3508 - 0xdb4  :  255 - 0xff
    "11101111", -- 3509 - 0xdb5  :  239 - 0xef
    "11110111", -- 3510 - 0xdb6  :  247 - 0xf7
    "11111000", -- 3511 - 0xdb7  :  248 - 0xf8
    "11111111", -- 3512 - 0xdb8  :  255 - 0xff -- Background 0xb7
    "11111111", -- 3513 - 0xdb9  :  255 - 0xff
    "11111111", -- 3514 - 0xdba  :  255 - 0xff
    "00011111", -- 3515 - 0xdbb  :   31 - 0x1f
    "00011111", -- 3516 - 0xdbc  :   31 - 0x1f
    "01111111", -- 3517 - 0xdbd  :  127 - 0x7f
    "11111111", -- 3518 - 0xdbe  :  255 - 0xff
    "11111110", -- 3519 - 0xdbf  :  254 - 0xfe
    "11111111", -- 3520 - 0xdc0  :  255 - 0xff -- Background 0xb8
    "11111111", -- 3521 - 0xdc1  :  255 - 0xff
    "11111111", -- 3522 - 0xdc2  :  255 - 0xff
    "11111100", -- 3523 - 0xdc3  :  252 - 0xfc
    "11111000", -- 3524 - 0xdc4  :  248 - 0xf8
    "10000000", -- 3525 - 0xdc5  :  128 - 0x80
    "00000000", -- 3526 - 0xdc6  :    0 - 0x0
    "00000000", -- 3527 - 0xdc7  :    0 - 0x0
    "00110000", -- 3528 - 0xdc8  :   48 - 0x30 -- Background 0xb9
    "01111111", -- 3529 - 0xdc9  :  127 - 0x7f
    "01111111", -- 3530 - 0xdca  :  127 - 0x7f
    "00111111", -- 3531 - 0xdcb  :   63 - 0x3f
    "10000111", -- 3532 - 0xdcc  :  135 - 0x87
    "11110000", -- 3533 - 0xdcd  :  240 - 0xf0
    "11111111", -- 3534 - 0xdce  :  255 - 0xff
    "11111111", -- 3535 - 0xdcf  :  255 - 0xff
    "11100101", -- 3536 - 0xdd0  :  229 - 0xe5 -- Background 0xba
    "11011010", -- 3537 - 0xdd1  :  218 - 0xda
    "11000000", -- 3538 - 0xdd2  :  192 - 0xc0
    "00000000", -- 3539 - 0xdd3  :    0 - 0x0
    "00000000", -- 3540 - 0xdd4  :    0 - 0x0
    "00000000", -- 3541 - 0xdd5  :    0 - 0x0
    "00000000", -- 3542 - 0xdd6  :    0 - 0x0
    "00000000", -- 3543 - 0xdd7  :    0 - 0x0
    "00000110", -- 3544 - 0xdd8  :    6 - 0x6 -- Background 0xbb
    "11111111", -- 3545 - 0xdd9  :  255 - 0xff
    "11111111", -- 3546 - 0xdda  :  255 - 0xff
    "11111110", -- 3547 - 0xddb  :  254 - 0xfe
    "11110001", -- 3548 - 0xddc  :  241 - 0xf1
    "00000111", -- 3549 - 0xddd  :    7 - 0x7
    "11111111", -- 3550 - 0xdde  :  255 - 0xff
    "11111111", -- 3551 - 0xddf  :  255 - 0xff
    "00000000", -- 3552 - 0xde0  :    0 - 0x0 -- Background 0xbc
    "00000001", -- 3553 - 0xde1  :    1 - 0x1
    "00000010", -- 3554 - 0xde2  :    2 - 0x2
    "00000111", -- 3555 - 0xde3  :    7 - 0x7
    "00000000", -- 3556 - 0xde4  :    0 - 0x0
    "00000000", -- 3557 - 0xde5  :    0 - 0x0
    "00100000", -- 3558 - 0xde6  :   32 - 0x20
    "11111111", -- 3559 - 0xde7  :  255 - 0xff
    "01111111", -- 3560 - 0xde8  :  127 - 0x7f -- Background 0xbd
    "01111111", -- 3561 - 0xde9  :  127 - 0x7f
    "01111111", -- 3562 - 0xdea  :  127 - 0x7f
    "11111111", -- 3563 - 0xdeb  :  255 - 0xff
    "11111111", -- 3564 - 0xdec  :  255 - 0xff
    "11111111", -- 3565 - 0xded  :  255 - 0xff
    "11111111", -- 3566 - 0xdee  :  255 - 0xff
    "11111110", -- 3567 - 0xdef  :  254 - 0xfe
    "11111100", -- 3568 - 0xdf0  :  252 - 0xfc -- Background 0xbe
    "10111000", -- 3569 - 0xdf1  :  184 - 0xb8
    "01111000", -- 3570 - 0xdf2  :  120 - 0x78
    "01111000", -- 3571 - 0xdf3  :  120 - 0x78
    "10110000", -- 3572 - 0xdf4  :  176 - 0xb0
    "01111000", -- 3573 - 0xdf5  :  120 - 0x78
    "11111100", -- 3574 - 0xdf6  :  252 - 0xfc
    "11111110", -- 3575 - 0xdf7  :  254 - 0xfe
    "11111111", -- 3576 - 0xdf8  :  255 - 0xff -- Background 0xbf
    "11111111", -- 3577 - 0xdf9  :  255 - 0xff
    "11111111", -- 3578 - 0xdfa  :  255 - 0xff
    "11111111", -- 3579 - 0xdfb  :  255 - 0xff
    "11111111", -- 3580 - 0xdfc  :  255 - 0xff
    "10011100", -- 3581 - 0xdfd  :  156 - 0x9c
    "01000010", -- 3582 - 0xdfe  :   66 - 0x42
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "00000000", -- 3584 - 0xe00  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 3585 - 0xe01  :    0 - 0x0
    "00100000", -- 3586 - 0xe02  :   32 - 0x20
    "01000000", -- 3587 - 0xe03  :   64 - 0x40
    "10001010", -- 3588 - 0xe04  :  138 - 0x8a
    "00011110", -- 3589 - 0xe05  :   30 - 0x1e
    "01111110", -- 3590 - 0xe06  :  126 - 0x7e
    "10111110", -- 3591 - 0xe07  :  190 - 0xbe
    "11011111", -- 3592 - 0xe08  :  223 - 0xdf -- Background 0xc1
    "11111111", -- 3593 - 0xe09  :  255 - 0xff
    "11111110", -- 3594 - 0xe0a  :  254 - 0xfe
    "11111100", -- 3595 - 0xe0b  :  252 - 0xfc
    "11110000", -- 3596 - 0xe0c  :  240 - 0xf0
    "11100000", -- 3597 - 0xe0d  :  224 - 0xe0
    "10000000", -- 3598 - 0xe0e  :  128 - 0x80
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "00000000", -- 3600 - 0xe10  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 3601 - 0xe11  :    0 - 0x0
    "00000100", -- 3602 - 0xe12  :    4 - 0x4
    "00000010", -- 3603 - 0xe13  :    2 - 0x2
    "01010001", -- 3604 - 0xe14  :   81 - 0x51
    "01111000", -- 3605 - 0xe15  :  120 - 0x78
    "01111110", -- 3606 - 0xe16  :  126 - 0x7e
    "11111101", -- 3607 - 0xe17  :  253 - 0xfd
    "11111011", -- 3608 - 0xe18  :  251 - 0xfb -- Background 0xc3
    "11111111", -- 3609 - 0xe19  :  255 - 0xff
    "01111111", -- 3610 - 0xe1a  :  127 - 0x7f
    "00111111", -- 3611 - 0xe1b  :   63 - 0x3f
    "00001111", -- 3612 - 0xe1c  :   15 - 0xf
    "00000111", -- 3613 - 0xe1d  :    7 - 0x7
    "00000001", -- 3614 - 0xe1e  :    1 - 0x1
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "00000000", -- 3616 - 0xe20  :    0 - 0x0 -- Background 0xc4
    "10000000", -- 3617 - 0xe21  :  128 - 0x80
    "01000000", -- 3618 - 0xe22  :   64 - 0x40
    "11100000", -- 3619 - 0xe23  :  224 - 0xe0
    "00000000", -- 3620 - 0xe24  :    0 - 0x0
    "00000000", -- 3621 - 0xe25  :    0 - 0x0
    "00000100", -- 3622 - 0xe26  :    4 - 0x4
    "11111111", -- 3623 - 0xe27  :  255 - 0xff
    "11111110", -- 3624 - 0xe28  :  254 - 0xfe -- Background 0xc5
    "11111110", -- 3625 - 0xe29  :  254 - 0xfe
    "11111110", -- 3626 - 0xe2a  :  254 - 0xfe
    "11111111", -- 3627 - 0xe2b  :  255 - 0xff
    "11111111", -- 3628 - 0xe2c  :  255 - 0xff
    "11111111", -- 3629 - 0xe2d  :  255 - 0xff
    "11111111", -- 3630 - 0xe2e  :  255 - 0xff
    "01111111", -- 3631 - 0xe2f  :  127 - 0x7f
    "00111111", -- 3632 - 0xe30  :   63 - 0x3f -- Background 0xc6
    "00011101", -- 3633 - 0xe31  :   29 - 0x1d
    "00011110", -- 3634 - 0xe32  :   30 - 0x1e
    "00011110", -- 3635 - 0xe33  :   30 - 0x1e
    "00001101", -- 3636 - 0xe34  :   13 - 0xd
    "00011110", -- 3637 - 0xe35  :   30 - 0x1e
    "00111111", -- 3638 - 0xe36  :   63 - 0x3f
    "01111111", -- 3639 - 0xe37  :  127 - 0x7f
    "11111111", -- 3640 - 0xe38  :  255 - 0xff -- Background 0xc7
    "11111111", -- 3641 - 0xe39  :  255 - 0xff
    "11111111", -- 3642 - 0xe3a  :  255 - 0xff
    "11111111", -- 3643 - 0xe3b  :  255 - 0xff
    "11111111", -- 3644 - 0xe3c  :  255 - 0xff
    "00111001", -- 3645 - 0xe3d  :   57 - 0x39
    "01000010", -- 3646 - 0xe3e  :   66 - 0x42
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "01101111", -- 3648 - 0xe40  :  111 - 0x6f -- Background 0xc8
    "11011011", -- 3649 - 0xe41  :  219 - 0xdb
    "00000011", -- 3650 - 0xe42  :    3 - 0x3
    "00000000", -- 3651 - 0xe43  :    0 - 0x0
    "00000000", -- 3652 - 0xe44  :    0 - 0x0
    "00000000", -- 3653 - 0xe45  :    0 - 0x0
    "00000000", -- 3654 - 0xe46  :    0 - 0x0
    "00000000", -- 3655 - 0xe47  :    0 - 0x0
    "00000000", -- 3656 - 0xe48  :    0 - 0x0 -- Background 0xc9
    "00000000", -- 3657 - 0xe49  :    0 - 0x0
    "00000000", -- 3658 - 0xe4a  :    0 - 0x0
    "00000000", -- 3659 - 0xe4b  :    0 - 0x0
    "00000000", -- 3660 - 0xe4c  :    0 - 0x0
    "00000000", -- 3661 - 0xe4d  :    0 - 0x0
    "00000000", -- 3662 - 0xe4e  :    0 - 0x0
    "11100000", -- 3663 - 0xe4f  :  224 - 0xe0
    "01110000", -- 3664 - 0xe50  :  112 - 0x70 -- Background 0xca
    "01111100", -- 3665 - 0xe51  :  124 - 0x7c
    "01111110", -- 3666 - 0xe52  :  126 - 0x7e
    "11111111", -- 3667 - 0xe53  :  255 - 0xff
    "11111111", -- 3668 - 0xe54  :  255 - 0xff
    "11110111", -- 3669 - 0xe55  :  247 - 0xf7
    "11101111", -- 3670 - 0xe56  :  239 - 0xef
    "00011111", -- 3671 - 0xe57  :   31 - 0x1f
    "11111111", -- 3672 - 0xe58  :  255 - 0xff -- Background 0xcb
    "11111111", -- 3673 - 0xe59  :  255 - 0xff
    "11111111", -- 3674 - 0xe5a  :  255 - 0xff
    "11111000", -- 3675 - 0xe5b  :  248 - 0xf8
    "11111000", -- 3676 - 0xe5c  :  248 - 0xf8
    "11111110", -- 3677 - 0xe5d  :  254 - 0xfe
    "11111111", -- 3678 - 0xe5e  :  255 - 0xff
    "11111111", -- 3679 - 0xe5f  :  255 - 0xff
    "11111111", -- 3680 - 0xe60  :  255 - 0xff -- Background 0xcc
    "11111111", -- 3681 - 0xe61  :  255 - 0xff
    "11111111", -- 3682 - 0xe62  :  255 - 0xff
    "00111111", -- 3683 - 0xe63  :   63 - 0x3f
    "00011110", -- 3684 - 0xe64  :   30 - 0x1e
    "00000001", -- 3685 - 0xe65  :    1 - 0x1
    "00000000", -- 3686 - 0xe66  :    0 - 0x0
    "00000000", -- 3687 - 0xe67  :    0 - 0x0
    "00000000", -- 3688 - 0xe68  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 3689 - 0xe69  :    0 - 0x0
    "00000000", -- 3690 - 0xe6a  :    0 - 0x0
    "10000000", -- 3691 - 0xe6b  :  128 - 0x80
    "11000000", -- 3692 - 0xe6c  :  192 - 0xc0
    "11100000", -- 3693 - 0xe6d  :  224 - 0xe0
    "11100000", -- 3694 - 0xe6e  :  224 - 0xe0
    "11100000", -- 3695 - 0xe6f  :  224 - 0xe0
    "11000000", -- 3696 - 0xe70  :  192 - 0xc0 -- Background 0xce
    "10000000", -- 3697 - 0xe71  :  128 - 0x80
    "00000000", -- 3698 - 0xe72  :    0 - 0x0
    "00000000", -- 3699 - 0xe73  :    0 - 0x0
    "00000000", -- 3700 - 0xe74  :    0 - 0x0
    "00000000", -- 3701 - 0xe75  :    0 - 0x0
    "10000000", -- 3702 - 0xe76  :  128 - 0x80
    "10000000", -- 3703 - 0xe77  :  128 - 0x80
    "10000000", -- 3704 - 0xe78  :  128 - 0x80 -- Background 0xcf
    "10000000", -- 3705 - 0xe79  :  128 - 0x80
    "11100000", -- 3706 - 0xe7a  :  224 - 0xe0
    "11000000", -- 3707 - 0xe7b  :  192 - 0xc0
    "00100000", -- 3708 - 0xe7c  :   32 - 0x20
    "00000000", -- 3709 - 0xe7d  :    0 - 0x0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "00011111", -- 3712 - 0xe80  :   31 - 0x1f -- Background 0xd0
    "00000110", -- 3713 - 0xe81  :    6 - 0x6
    "00000110", -- 3714 - 0xe82  :    6 - 0x6
    "00000110", -- 3715 - 0xe83  :    6 - 0x6
    "00000110", -- 3716 - 0xe84  :    6 - 0x6
    "00000110", -- 3717 - 0xe85  :    6 - 0x6
    "00000110", -- 3718 - 0xe86  :    6 - 0x6
    "00000000", -- 3719 - 0xe87  :    0 - 0x0
    "00111001", -- 3720 - 0xe88  :   57 - 0x39 -- Background 0xd1
    "01100101", -- 3721 - 0xe89  :  101 - 0x65
    "01100101", -- 3722 - 0xe8a  :  101 - 0x65
    "01100101", -- 3723 - 0xe8b  :  101 - 0x65
    "01100101", -- 3724 - 0xe8c  :  101 - 0x65
    "01100101", -- 3725 - 0xe8d  :  101 - 0x65
    "00111001", -- 3726 - 0xe8e  :   57 - 0x39
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "11100000", -- 3728 - 0xe90  :  224 - 0xe0 -- Background 0xd2
    "10110000", -- 3729 - 0xe91  :  176 - 0xb0
    "10110000", -- 3730 - 0xe92  :  176 - 0xb0
    "10110110", -- 3731 - 0xe93  :  182 - 0xb6
    "11100110", -- 3732 - 0xe94  :  230 - 0xe6
    "10000000", -- 3733 - 0xe95  :  128 - 0x80
    "10000000", -- 3734 - 0xe96  :  128 - 0x80
    "00000000", -- 3735 - 0xe97  :    0 - 0x0
    "00111100", -- 3736 - 0xe98  :   60 - 0x3c -- Background 0xd3
    "01000010", -- 3737 - 0xe99  :   66 - 0x42
    "10011001", -- 3738 - 0xe9a  :  153 - 0x99
    "10100001", -- 3739 - 0xe9b  :  161 - 0xa1
    "10100001", -- 3740 - 0xe9c  :  161 - 0xa1
    "10011001", -- 3741 - 0xe9d  :  153 - 0x99
    "01000010", -- 3742 - 0xe9e  :   66 - 0x42
    "00111100", -- 3743 - 0xe9f  :   60 - 0x3c
    "00000000", -- 3744 - 0xea0  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 3745 - 0xea1  :    0 - 0x0
    "00000000", -- 3746 - 0xea2  :    0 - 0x0
    "00000011", -- 3747 - 0xea3  :    3 - 0x3
    "00000110", -- 3748 - 0xea4  :    6 - 0x6
    "00000000", -- 3749 - 0xea5  :    0 - 0x0
    "00000001", -- 3750 - 0xea6  :    1 - 0x1
    "00000111", -- 3751 - 0xea7  :    7 - 0x7
    "00001111", -- 3752 - 0xea8  :   15 - 0xf -- Background 0xd5
    "00011111", -- 3753 - 0xea9  :   31 - 0x1f
    "00111111", -- 3754 - 0xeaa  :   63 - 0x3f
    "01111111", -- 3755 - 0xeab  :  127 - 0x7f
    "01111111", -- 3756 - 0xeac  :  127 - 0x7f
    "01111111", -- 3757 - 0xead  :  127 - 0x7f
    "11111111", -- 3758 - 0xeae  :  255 - 0xff
    "01111111", -- 3759 - 0xeaf  :  127 - 0x7f
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 3761 - 0xeb1  :    0 - 0x0
    "00000000", -- 3762 - 0xeb2  :    0 - 0x0
    "10000000", -- 3763 - 0xeb3  :  128 - 0x80
    "00000000", -- 3764 - 0xeb4  :    0 - 0x0
    "00000000", -- 3765 - 0xeb5  :    0 - 0x0
    "00000000", -- 3766 - 0xeb6  :    0 - 0x0
    "10100000", -- 3767 - 0xeb7  :  160 - 0xa0
    "11100000", -- 3768 - 0xeb8  :  224 - 0xe0 -- Background 0xd7
    "11110000", -- 3769 - 0xeb9  :  240 - 0xf0
    "11100000", -- 3770 - 0xeba  :  224 - 0xe0
    "11011101", -- 3771 - 0xebb  :  221 - 0xdd
    "11111010", -- 3772 - 0xebc  :  250 - 0xfa
    "11101011", -- 3773 - 0xebd  :  235 - 0xeb
    "10000000", -- 3774 - 0xebe  :  128 - 0x80
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Background 0xd8
    "00000000", -- 3777 - 0xec1  :    0 - 0x0
    "00000000", -- 3778 - 0xec2  :    0 - 0x0
    "00000011", -- 3779 - 0xec3  :    3 - 0x3
    "00000110", -- 3780 - 0xec4  :    6 - 0x6
    "00000000", -- 3781 - 0xec5  :    0 - 0x0
    "00000001", -- 3782 - 0xec6  :    1 - 0x1
    "00000001", -- 3783 - 0xec7  :    1 - 0x1
    "00001011", -- 3784 - 0xec8  :   11 - 0xb -- Background 0xd9
    "00000111", -- 3785 - 0xec9  :    7 - 0x7
    "00000011", -- 3786 - 0xeca  :    3 - 0x3
    "01011101", -- 3787 - 0xecb  :   93 - 0x5d
    "10101111", -- 3788 - 0xecc  :  175 - 0xaf
    "01010011", -- 3789 - 0xecd  :   83 - 0x53
    "00000000", -- 3790 - 0xece  :    0 - 0x0
    "00000000", -- 3791 - 0xecf  :    0 - 0x0
    "00000000", -- 3792 - 0xed0  :    0 - 0x0 -- Background 0xda
    "00000000", -- 3793 - 0xed1  :    0 - 0x0
    "00000000", -- 3794 - 0xed2  :    0 - 0x0
    "10000000", -- 3795 - 0xed3  :  128 - 0x80
    "00000000", -- 3796 - 0xed4  :    0 - 0x0
    "00000000", -- 3797 - 0xed5  :    0 - 0x0
    "01100000", -- 3798 - 0xed6  :   96 - 0x60
    "11110000", -- 3799 - 0xed7  :  240 - 0xf0
    "11111000", -- 3800 - 0xed8  :  248 - 0xf8 -- Background 0xdb
    "11111100", -- 3801 - 0xed9  :  252 - 0xfc
    "11111100", -- 3802 - 0xeda  :  252 - 0xfc
    "11111110", -- 3803 - 0xedb  :  254 - 0xfe
    "11111110", -- 3804 - 0xedc  :  254 - 0xfe
    "11111111", -- 3805 - 0xedd  :  255 - 0xff
    "11111111", -- 3806 - 0xede  :  255 - 0xff
    "01111110", -- 3807 - 0xedf  :  126 - 0x7e
    "00000000", -- 3808 - 0xee0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000000", -- 3811 - 0xee3  :    0 - 0x0
    "00000000", -- 3812 - 0xee4  :    0 - 0x0
    "00000000", -- 3813 - 0xee5  :    0 - 0x0
    "00100001", -- 3814 - 0xee6  :   33 - 0x21
    "00111111", -- 3815 - 0xee7  :   63 - 0x3f
    "00111111", -- 3816 - 0xee8  :   63 - 0x3f -- Background 0xdd
    "00011111", -- 3817 - 0xee9  :   31 - 0x1f
    "00011111", -- 3818 - 0xeea  :   31 - 0x1f
    "00001111", -- 3819 - 0xeeb  :   15 - 0xf
    "00000111", -- 3820 - 0xeec  :    7 - 0x7
    "00000011", -- 3821 - 0xeed  :    3 - 0x3
    "00000000", -- 3822 - 0xeee  :    0 - 0x0
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "00111110", -- 3824 - 0xef0  :   62 - 0x3e -- Background 0xde
    "00011110", -- 3825 - 0xef1  :   30 - 0x1e
    "00011110", -- 3826 - 0xef2  :   30 - 0x1e
    "00001110", -- 3827 - 0xef3  :   14 - 0xe
    "00001111", -- 3828 - 0xef4  :   15 - 0xf
    "00011111", -- 3829 - 0xef5  :   31 - 0x1f
    "10011111", -- 3830 - 0xef6  :  159 - 0x9f
    "10011111", -- 3831 - 0xef7  :  159 - 0x9f
    "11011111", -- 3832 - 0xef8  :  223 - 0xdf -- Background 0xdf
    "11111111", -- 3833 - 0xef9  :  255 - 0xff
    "11111111", -- 3834 - 0xefa  :  255 - 0xff
    "11111111", -- 3835 - 0xefb  :  255 - 0xff
    "11111111", -- 3836 - 0xefc  :  255 - 0xff
    "11011111", -- 3837 - 0xefd  :  223 - 0xdf
    "11100111", -- 3838 - 0xefe  :  231 - 0xe7
    "00000000", -- 3839 - 0xeff  :    0 - 0x0
    "00100000", -- 3840 - 0xf00  :   32 - 0x20 -- Background 0xe0
    "00001111", -- 3841 - 0xf01  :   15 - 0xf
    "00110000", -- 3842 - 0xf02  :   48 - 0x30
    "01000000", -- 3843 - 0xf03  :   64 - 0x40
    "10011000", -- 3844 - 0xf04  :  152 - 0x98
    "00111110", -- 3845 - 0xf05  :   62 - 0x3e
    "00011111", -- 3846 - 0xf06  :   31 - 0x1f
    "00000000", -- 3847 - 0xf07  :    0 - 0x0
    "10000001", -- 3848 - 0xf08  :  129 - 0x81 -- Background 0xe1
    "00110110", -- 3849 - 0xf09  :   54 - 0x36
    "00101110", -- 3850 - 0xf0a  :   46 - 0x2e
    "10101111", -- 3851 - 0xf0b  :  175 - 0xaf
    "10101110", -- 3852 - 0xf0c  :  174 - 0xae
    "11010001", -- 3853 - 0xf0d  :  209 - 0xd1
    "11101111", -- 3854 - 0xf0e  :  239 - 0xef
    "10000111", -- 3855 - 0xf0f  :  135 - 0x87
    "00000010", -- 3856 - 0xf10  :    2 - 0x2 -- Background 0xe2
    "11111000", -- 3857 - 0xf11  :  248 - 0xf8
    "00000110", -- 3858 - 0xf12  :    6 - 0x6
    "00000001", -- 3859 - 0xf13  :    1 - 0x1
    "00001100", -- 3860 - 0xf14  :   12 - 0xc
    "00111110", -- 3861 - 0xf15  :   62 - 0x3e
    "11111100", -- 3862 - 0xf16  :  252 - 0xfc
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "11000000", -- 3864 - 0xf18  :  192 - 0xc0 -- Background 0xe3
    "00110110", -- 3865 - 0xf19  :   54 - 0x36
    "00111110", -- 3866 - 0xf1a  :   62 - 0x3e
    "01111010", -- 3867 - 0xf1b  :  122 - 0x7a
    "10110110", -- 3868 - 0xf1c  :  182 - 0xb6
    "11001101", -- 3869 - 0xf1d  :  205 - 0xcd
    "11111011", -- 3870 - 0xf1e  :  251 - 0xfb
    "11110000", -- 3871 - 0xf1f  :  240 - 0xf0
    "00111110", -- 3872 - 0xf20  :   62 - 0x3e -- Background 0xe4
    "00111100", -- 3873 - 0xf21  :   60 - 0x3c
    "00111100", -- 3874 - 0xf22  :   60 - 0x3c
    "00111000", -- 3875 - 0xf23  :   56 - 0x38
    "11111000", -- 3876 - 0xf24  :  248 - 0xf8
    "01111100", -- 3877 - 0xf25  :  124 - 0x7c
    "01111110", -- 3878 - 0xf26  :  126 - 0x7e
    "01111000", -- 3879 - 0xf27  :  120 - 0x78
    "11111000", -- 3880 - 0xf28  :  248 - 0xf8 -- Background 0xe5
    "01111111", -- 3881 - 0xf29  :  127 - 0x7f
    "01111111", -- 3882 - 0xf2a  :  127 - 0x7f
    "11111110", -- 3883 - 0xf2b  :  254 - 0xfe
    "11111111", -- 3884 - 0xf2c  :  255 - 0xff
    "11111111", -- 3885 - 0xf2d  :  255 - 0xff
    "11110011", -- 3886 - 0xf2e  :  243 - 0xf3
    "10000001", -- 3887 - 0xf2f  :  129 - 0x81
    "00000000", -- 3888 - 0xf30  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 3889 - 0xf31  :    0 - 0x0
    "00000000", -- 3890 - 0xf32  :    0 - 0x0
    "00010000", -- 3891 - 0xf33  :   16 - 0x10
    "01000000", -- 3892 - 0xf34  :   64 - 0x40
    "00100000", -- 3893 - 0xf35  :   32 - 0x20
    "00000000", -- 3894 - 0xf36  :    0 - 0x0
    "00000000", -- 3895 - 0xf37  :    0 - 0x0
    "00000110", -- 3896 - 0xf38  :    6 - 0x6 -- Background 0xe7
    "00001110", -- 3897 - 0xf39  :   14 - 0xe
    "01111110", -- 3898 - 0xf3a  :  126 - 0x7e
    "11111110", -- 3899 - 0xf3b  :  254 - 0xfe
    "11111110", -- 3900 - 0xf3c  :  254 - 0xfe
    "11111100", -- 3901 - 0xf3d  :  252 - 0xfc
    "11111000", -- 3902 - 0xf3e  :  248 - 0xf8
    "11110000", -- 3903 - 0xf3f  :  240 - 0xf0
    "00000000", -- 3904 - 0xf40  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 3905 - 0xf41  :    0 - 0x0
    "00000000", -- 3906 - 0xf42  :    0 - 0x0
    "00000000", -- 3907 - 0xf43  :    0 - 0x0
    "00000000", -- 3908 - 0xf44  :    0 - 0x0
    "00000000", -- 3909 - 0xf45  :    0 - 0x0
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "00000001", -- 3911 - 0xf47  :    1 - 0x1
    "00000010", -- 3912 - 0xf48  :    2 - 0x2 -- Background 0xe9
    "00000000", -- 3913 - 0xf49  :    0 - 0x0
    "00001000", -- 3914 - 0xf4a  :    8 - 0x8
    "00000001", -- 3915 - 0xf4b  :    1 - 0x1
    "00010011", -- 3916 - 0xf4c  :   19 - 0x13
    "00000001", -- 3917 - 0xf4d  :    1 - 0x1
    "00000000", -- 3918 - 0xf4e  :    0 - 0x0
    "00000000", -- 3919 - 0xf4f  :    0 - 0x0
    "00000000", -- 3920 - 0xf50  :    0 - 0x0 -- Background 0xea
    "00000000", -- 3921 - 0xf51  :    0 - 0x0
    "00000000", -- 3922 - 0xf52  :    0 - 0x0
    "00000000", -- 3923 - 0xf53  :    0 - 0x0
    "00000000", -- 3924 - 0xf54  :    0 - 0x0
    "00000000", -- 3925 - 0xf55  :    0 - 0x0
    "00000000", -- 3926 - 0xf56  :    0 - 0x0
    "00000000", -- 3927 - 0xf57  :    0 - 0x0
    "00000000", -- 3928 - 0xf58  :    0 - 0x0 -- Background 0xeb
    "01000011", -- 3929 - 0xf59  :   67 - 0x43
    "01111111", -- 3930 - 0xf5a  :  127 - 0x7f
    "01111111", -- 3931 - 0xf5b  :  127 - 0x7f
    "01111111", -- 3932 - 0xf5c  :  127 - 0x7f
    "00111111", -- 3933 - 0xf5d  :   63 - 0x3f
    "00011111", -- 3934 - 0xf5e  :   31 - 0x1f
    "00000111", -- 3935 - 0xf5f  :    7 - 0x7
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Background 0xec
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00000000", -- 3941 - 0xf65  :    0 - 0x0
    "11000000", -- 3942 - 0xf66  :  192 - 0xc0
    "00000000", -- 3943 - 0xf67  :    0 - 0x0
    "00010000", -- 3944 - 0xf68  :   16 - 0x10 -- Background 0xed
    "00111000", -- 3945 - 0xf69  :   56 - 0x38
    "10111111", -- 3946 - 0xf6a  :  191 - 0xbf
    "11111111", -- 3947 - 0xf6b  :  255 - 0xff
    "11111111", -- 3948 - 0xf6c  :  255 - 0xff
    "11111111", -- 3949 - 0xf6d  :  255 - 0xff
    "11111111", -- 3950 - 0xf6e  :  255 - 0xff
    "11111111", -- 3951 - 0xf6f  :  255 - 0xff
    "01111110", -- 3952 - 0xf70  :  126 - 0x7e -- Background 0xee
    "00011110", -- 3953 - 0xf71  :   30 - 0x1e
    "00011110", -- 3954 - 0xf72  :   30 - 0x1e
    "00001110", -- 3955 - 0xf73  :   14 - 0xe
    "00001111", -- 3956 - 0xf74  :   15 - 0xf
    "00011110", -- 3957 - 0xf75  :   30 - 0x1e
    "00011110", -- 3958 - 0xf76  :   30 - 0x1e
    "00111110", -- 3959 - 0xf77  :   62 - 0x3e
    "01111111", -- 3960 - 0xf78  :  127 - 0x7f -- Background 0xef
    "01111111", -- 3961 - 0xf79  :  127 - 0x7f
    "10111111", -- 3962 - 0xf7a  :  191 - 0xbf
    "11111111", -- 3963 - 0xf7b  :  255 - 0xff
    "11111111", -- 3964 - 0xf7c  :  255 - 0xff
    "11111111", -- 3965 - 0xf7d  :  255 - 0xff
    "11100111", -- 3966 - 0xf7e  :  231 - 0xe7
    "11000000", -- 3967 - 0xf7f  :  192 - 0xc0
    "00000000", -- 3968 - 0xf80  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 3969 - 0xf81  :    0 - 0x0
    "00010000", -- 3970 - 0xf82  :   16 - 0x10
    "11111101", -- 3971 - 0xf83  :  253 - 0xfd
    "11111010", -- 3972 - 0xf84  :  250 - 0xfa
    "11101011", -- 3973 - 0xf85  :  235 - 0xeb
    "10000000", -- 3974 - 0xf86  :  128 - 0x80
    "00000000", -- 3975 - 0xf87  :    0 - 0x0
    "00100000", -- 3976 - 0xf88  :   32 - 0x20 -- Background 0xf1
    "00011111", -- 3977 - 0xf89  :   31 - 0x1f
    "01100000", -- 3978 - 0xf8a  :   96 - 0x60
    "10001110", -- 3979 - 0xf8b  :  142 - 0x8e
    "00111111", -- 3980 - 0xf8c  :   63 - 0x3f
    "01111111", -- 3981 - 0xf8d  :  127 - 0x7f
    "01111111", -- 3982 - 0xf8e  :  127 - 0x7f
    "01111100", -- 3983 - 0xf8f  :  124 - 0x7c
    "00111001", -- 3984 - 0xf90  :   57 - 0x39 -- Background 0xf2
    "00110110", -- 3985 - 0xf91  :   54 - 0x36
    "00101110", -- 3986 - 0xf92  :   46 - 0x2e
    "10101111", -- 3987 - 0xf93  :  175 - 0xaf
    "10101110", -- 3988 - 0xf94  :  174 - 0xae
    "11010001", -- 3989 - 0xf95  :  209 - 0xd1
    "11101111", -- 3990 - 0xf96  :  239 - 0xef
    "10000111", -- 3991 - 0xf97  :  135 - 0x87
    "00000000", -- 3992 - 0xf98  :    0 - 0x0 -- Background 0xf3
    "00000000", -- 3993 - 0xf99  :    0 - 0x0
    "00000100", -- 3994 - 0xf9a  :    4 - 0x4
    "01011111", -- 3995 - 0xf9b  :   95 - 0x5f
    "10101111", -- 3996 - 0xf9c  :  175 - 0xaf
    "01010011", -- 3997 - 0xf9d  :   83 - 0x53
    "00000000", -- 3998 - 0xf9e  :    0 - 0x0
    "00000000", -- 3999 - 0xf9f  :    0 - 0x0
    "00000010", -- 4000 - 0xfa0  :    2 - 0x2 -- Background 0xf4
    "11111100", -- 4001 - 0xfa1  :  252 - 0xfc
    "00000011", -- 4002 - 0xfa2  :    3 - 0x3
    "00111000", -- 4003 - 0xfa3  :   56 - 0x38
    "11111110", -- 4004 - 0xfa4  :  254 - 0xfe
    "11111111", -- 4005 - 0xfa5  :  255 - 0xff
    "11111111", -- 4006 - 0xfa6  :  255 - 0xff
    "00011110", -- 4007 - 0xfa7  :   30 - 0x1e
    "11000000", -- 4008 - 0xfa8  :  192 - 0xc0 -- Background 0xf5
    "00110110", -- 4009 - 0xfa9  :   54 - 0x36
    "00111110", -- 4010 - 0xfaa  :   62 - 0x3e
    "01111010", -- 4011 - 0xfab  :  122 - 0x7a
    "10110110", -- 4012 - 0xfac  :  182 - 0xb6
    "11001101", -- 4013 - 0xfad  :  205 - 0xcd
    "11111011", -- 4014 - 0xfae  :  251 - 0xfb
    "11110000", -- 4015 - 0xfaf  :  240 - 0xf0
    "00000000", -- 4016 - 0xfb0  :    0 - 0x0 -- Background 0xf6
    "00000000", -- 4017 - 0xfb1  :    0 - 0x0
    "00000000", -- 4018 - 0xfb2  :    0 - 0x0
    "00000000", -- 4019 - 0xfb3  :    0 - 0x0
    "00000000", -- 4020 - 0xfb4  :    0 - 0x0
    "00001110", -- 4021 - 0xfb5  :   14 - 0xe
    "00001000", -- 4022 - 0xfb6  :    8 - 0x8
    "00001000", -- 4023 - 0xfb7  :    8 - 0x8
    "00011111", -- 4024 - 0xfb8  :   31 - 0x1f -- Background 0xf7
    "00111111", -- 4025 - 0xfb9  :   63 - 0x3f
    "11111111", -- 4026 - 0xfba  :  255 - 0xff
    "11111111", -- 4027 - 0xfbb  :  255 - 0xff
    "11111111", -- 4028 - 0xfbc  :  255 - 0xff
    "11111111", -- 4029 - 0xfbd  :  255 - 0xff
    "11111111", -- 4030 - 0xfbe  :  255 - 0xff
    "01111111", -- 4031 - 0xfbf  :  127 - 0x7f
    "00111111", -- 4032 - 0xfc0  :   63 - 0x3f -- Background 0xf8
    "00111110", -- 4033 - 0xfc1  :   62 - 0x3e
    "00111100", -- 4034 - 0xfc2  :   60 - 0x3c
    "10111000", -- 4035 - 0xfc3  :  184 - 0xb8
    "01111000", -- 4036 - 0xfc4  :  120 - 0x78
    "01111000", -- 4037 - 0xfc5  :  120 - 0x78
    "01111110", -- 4038 - 0xfc6  :  126 - 0x7e
    "01111110", -- 4039 - 0xfc7  :  126 - 0x7e
    "11111101", -- 4040 - 0xfc8  :  253 - 0xfd -- Background 0xf9
    "01111001", -- 4041 - 0xfc9  :  121 - 0x79
    "01111011", -- 4042 - 0xfca  :  123 - 0x7b
    "11111111", -- 4043 - 0xfcb  :  255 - 0xff
    "11111111", -- 4044 - 0xfcc  :  255 - 0xff
    "11111111", -- 4045 - 0xfcd  :  255 - 0xff
    "11110011", -- 4046 - 0xfce  :  243 - 0xf3
    "10000000", -- 4047 - 0xfcf  :  128 - 0x80
    "00000000", -- 4048 - 0xfd0  :    0 - 0x0 -- Background 0xfa
    "00000000", -- 4049 - 0xfd1  :    0 - 0x0
    "00000000", -- 4050 - 0xfd2  :    0 - 0x0
    "00000000", -- 4051 - 0xfd3  :    0 - 0x0
    "00000000", -- 4052 - 0xfd4  :    0 - 0x0
    "00000000", -- 4053 - 0xfd5  :    0 - 0x0
    "00000000", -- 4054 - 0xfd6  :    0 - 0x0
    "00000000", -- 4055 - 0xfd7  :    0 - 0x0
    "00010000", -- 4056 - 0xfd8  :   16 - 0x10 -- Background 0xfb
    "10000100", -- 4057 - 0xfd9  :  132 - 0x84
    "11100000", -- 4058 - 0xfda  :  224 - 0xe0
    "11000000", -- 4059 - 0xfdb  :  192 - 0xc0
    "10000000", -- 4060 - 0xfdc  :  128 - 0x80
    "10000000", -- 4061 - 0xfdd  :  128 - 0x80
    "00000000", -- 4062 - 0xfde  :    0 - 0x0
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00000000", -- 4064 - 0xfe0  :    0 - 0x0 -- Background 0xfc
    "01001000", -- 4065 - 0xfe1  :   72 - 0x48
    "00100000", -- 4066 - 0xfe2  :   32 - 0x20
    "00000000", -- 4067 - 0xfe3  :    0 - 0x0
    "00000000", -- 4068 - 0xfe4  :    0 - 0x0
    "00000100", -- 4069 - 0xfe5  :    4 - 0x4
    "00001110", -- 4070 - 0xfe6  :   14 - 0xe
    "11111110", -- 4071 - 0xfe7  :  254 - 0xfe
    "11111110", -- 4072 - 0xfe8  :  254 - 0xfe -- Background 0xfd
    "11111100", -- 4073 - 0xfe9  :  252 - 0xfc
    "11111100", -- 4074 - 0xfea  :  252 - 0xfc
    "11111000", -- 4075 - 0xfeb  :  248 - 0xf8
    "11110000", -- 4076 - 0xfec  :  240 - 0xf0
    "11100000", -- 4077 - 0xfed  :  224 - 0xe0
    "10000000", -- 4078 - 0xfee  :  128 - 0x80
    "00000000", -- 4079 - 0xfef  :    0 - 0x0
    "00001111", -- 4080 - 0xff0  :   15 - 0xf -- Background 0xfe
    "00000110", -- 4081 - 0xff1  :    6 - 0x6
    "00000110", -- 4082 - 0xff2  :    6 - 0x6
    "00000110", -- 4083 - 0xff3  :    6 - 0x6
    "00000110", -- 4084 - 0xff4  :    6 - 0x6
    "00000110", -- 4085 - 0xff5  :    6 - 0x6
    "00001111", -- 4086 - 0xff6  :   15 - 0xf
    "00000000", -- 4087 - 0xff7  :    0 - 0x0
    "11110000", -- 4088 - 0xff8  :  240 - 0xf0 -- Background 0xff
    "01100000", -- 4089 - 0xff9  :   96 - 0x60
    "01100000", -- 4090 - 0xffa  :   96 - 0x60
    "01100110", -- 4091 - 0xffb  :  102 - 0x66
    "01100110", -- 4092 - 0xffc  :  102 - 0x66
    "01100000", -- 4093 - 0xffd  :   96 - 0x60
    "11110000", -- 4094 - 0xffe  :  240 - 0xf0
    "00000000"  -- 4095 - 0xfff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
