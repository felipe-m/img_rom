--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: lawnmower_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_LAWN is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(13-1 downto 0);  --8192 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_LAWN;

architecture BEHAVIORAL of ROM_PTABLE_LAWN is
  signal addr_int  : natural range 0 to 2**13-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Pattern Table 0---------
    "11111111", --    0 -  0x0  :  255 - 0xff -- Sprite 0x0
    "11111111", --    1 -  0x1  :  255 - 0xff
    "11111111", --    2 -  0x2  :  255 - 0xff
    "11111111", --    3 -  0x3  :  255 - 0xff
    "11111111", --    4 -  0x4  :  255 - 0xff
    "11111111", --    5 -  0x5  :  255 - 0xff
    "11111111", --    6 -  0x6  :  255 - 0xff
    "11111111", --    7 -  0x7  :  255 - 0xff
    "00000000", --    8 -  0x8  :    0 - 0x0
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "11111111", --   16 - 0x10  :  255 - 0xff -- Sprite 0x1
    "11111111", --   17 - 0x11  :  255 - 0xff
    "11111111", --   18 - 0x12  :  255 - 0xff
    "11111111", --   19 - 0x13  :  255 - 0xff
    "11111111", --   20 - 0x14  :  255 - 0xff
    "11111111", --   21 - 0x15  :  255 - 0xff
    "11111100", --   22 - 0x16  :  252 - 0xfc
    "11111100", --   23 - 0x17  :  252 - 0xfc
    "00000000", --   24 - 0x18  :    0 - 0x0
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000111", --   29 - 0x1d  :    7 - 0x7
    "00000111", --   30 - 0x1e  :    7 - 0x7
    "00000110", --   31 - 0x1f  :    6 - 0x6
    "11111111", --   32 - 0x20  :  255 - 0xff -- Sprite 0x2
    "11111111", --   33 - 0x21  :  255 - 0xff
    "11111111", --   34 - 0x22  :  255 - 0xff
    "11111111", --   35 - 0x23  :  255 - 0xff
    "11111111", --   36 - 0x24  :  255 - 0xff
    "11111111", --   37 - 0x25  :  255 - 0xff
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "11111111", --   45 - 0x2d  :  255 - 0xff
    "11111111", --   46 - 0x2e  :  255 - 0xff
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "11111111", --   48 - 0x30  :  255 - 0xff -- Sprite 0x3
    "11111111", --   49 - 0x31  :  255 - 0xff
    "11111111", --   50 - 0x32  :  255 - 0xff
    "11111111", --   51 - 0x33  :  255 - 0xff
    "11111111", --   52 - 0x34  :  255 - 0xff
    "11111111", --   53 - 0x35  :  255 - 0xff
    "00011111", --   54 - 0x36  :   31 - 0x1f
    "01000111", --   55 - 0x37  :   71 - 0x47
    "00000000", --   56 - 0x38  :    0 - 0x0
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "11100000", --   61 - 0x3d  :  224 - 0xe0
    "11100000", --   62 - 0x3e  :  224 - 0xe0
    "01100000", --   63 - 0x3f  :   96 - 0x60
    "11111111", --   64 - 0x40  :  255 - 0xff -- Sprite 0x4
    "11111111", --   65 - 0x41  :  255 - 0xff
    "11111111", --   66 - 0x42  :  255 - 0xff
    "11111111", --   67 - 0x43  :  255 - 0xff
    "11111111", --   68 - 0x44  :  255 - 0xff
    "11111111", --   69 - 0x45  :  255 - 0xff
    "11100000", --   70 - 0x46  :  224 - 0xe0
    "10000000", --   71 - 0x47  :  128 - 0x80
    "00000000", --   72 - 0x48  :    0 - 0x0
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00011111", --   77 - 0x4d  :   31 - 0x1f
    "01111111", --   78 - 0x4e  :  127 - 0x7f
    "11110000", --   79 - 0x4f  :  240 - 0xf0
    "11111111", --   80 - 0x50  :  255 - 0xff -- Sprite 0x5
    "11111111", --   81 - 0x51  :  255 - 0xff
    "11111111", --   82 - 0x52  :  255 - 0xff
    "11111111", --   83 - 0x53  :  255 - 0xff
    "11111111", --   84 - 0x54  :  255 - 0xff
    "11110111", --   85 - 0x55  :  247 - 0xf7
    "00000001", --   86 - 0x56  :    1 - 0x1
    "00000100", --   87 - 0x57  :    4 - 0x4
    "00000000", --   88 - 0x58  :    0 - 0x0
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "11111000", --   93 - 0x5d  :  248 - 0xf8
    "11111110", --   94 - 0x5e  :  254 - 0xfe
    "00001111", --   95 - 0x5f  :   15 - 0xf
    "11111111", --   96 - 0x60  :  255 - 0xff -- Sprite 0x6
    "11111111", --   97 - 0x61  :  255 - 0xff
    "11111111", --   98 - 0x62  :  255 - 0xff
    "11111111", --   99 - 0x63  :  255 - 0xff
    "11111111", --  100 - 0x64  :  255 - 0xff
    "11011111", --  101 - 0x65  :  223 - 0xdf
    "00011100", --  102 - 0x66  :   28 - 0x1c
    "01000100", --  103 - 0x67  :   68 - 0x44
    "00000000", --  104 - 0x68  :    0 - 0x0
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "11100111", --  109 - 0x6d  :  231 - 0xe7
    "11100111", --  110 - 0x6e  :  231 - 0xe7
    "01100110", --  111 - 0x6f  :  102 - 0x66
    "11111111", --  112 - 0x70  :  255 - 0xff -- Sprite 0x7
    "11111111", --  113 - 0x71  :  255 - 0xff
    "11111111", --  114 - 0x72  :  255 - 0xff
    "11111111", --  115 - 0x73  :  255 - 0xff
    "11111111", --  116 - 0x74  :  255 - 0xff
    "10111111", --  117 - 0x75  :  191 - 0xbf
    "00111100", --  118 - 0x76  :   60 - 0x3c
    "01001100", --  119 - 0x77  :   76 - 0x4c
    "00000000", --  120 - 0x78  :    0 - 0x0
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "11000111", --  125 - 0x7d  :  199 - 0xc7
    "11000111", --  126 - 0x7e  :  199 - 0xc7
    "01100110", --  127 - 0x7f  :  102 - 0x66
    "11111100", --  128 - 0x80  :  252 - 0xfc -- Sprite 0x8
    "11111100", --  129 - 0x81  :  252 - 0xfc
    "11111100", --  130 - 0x82  :  252 - 0xfc
    "11111100", --  131 - 0x83  :  252 - 0xfc
    "11111100", --  132 - 0x84  :  252 - 0xfc
    "11111100", --  133 - 0x85  :  252 - 0xfc
    "11111100", --  134 - 0x86  :  252 - 0xfc
    "11111100", --  135 - 0x87  :  252 - 0xfc
    "00000110", --  136 - 0x88  :    6 - 0x6
    "00000110", --  137 - 0x89  :    6 - 0x6
    "00000110", --  138 - 0x8a  :    6 - 0x6
    "00000110", --  139 - 0x8b  :    6 - 0x6
    "00000110", --  140 - 0x8c  :    6 - 0x6
    "00000110", --  141 - 0x8d  :    6 - 0x6
    "00000110", --  142 - 0x8e  :    6 - 0x6
    "00000110", --  143 - 0x8f  :    6 - 0x6
    "00010000", --  144 - 0x90  :   16 - 0x10 -- Sprite 0x9
    "00111000", --  145 - 0x91  :   56 - 0x38
    "01111100", --  146 - 0x92  :  124 - 0x7c
    "11111000", --  147 - 0x93  :  248 - 0xf8
    "01110000", --  148 - 0x94  :  112 - 0x70
    "00100010", --  149 - 0x95  :   34 - 0x22
    "00000101", --  150 - 0x96  :    5 - 0x5
    "00000010", --  151 - 0x97  :    2 - 0x2
    "11111111", --  152 - 0x98  :  255 - 0xff
    "11111111", --  153 - 0x99  :  255 - 0xff
    "11111111", --  154 - 0x9a  :  255 - 0xff
    "11111111", --  155 - 0x9b  :  255 - 0xff
    "11111111", --  156 - 0x9c  :  255 - 0xff
    "11111111", --  157 - 0x9d  :  255 - 0xff
    "11111111", --  158 - 0x9e  :  255 - 0xff
    "11111111", --  159 - 0x9f  :  255 - 0xff
    "01000111", --  160 - 0xa0  :   71 - 0x47 -- Sprite 0xa
    "01000111", --  161 - 0xa1  :   71 - 0x47
    "01000111", --  162 - 0xa2  :   71 - 0x47
    "01000111", --  163 - 0xa3  :   71 - 0x47
    "01000111", --  164 - 0xa4  :   71 - 0x47
    "01000111", --  165 - 0xa5  :   71 - 0x47
    "01000111", --  166 - 0xa6  :   71 - 0x47
    "01000111", --  167 - 0xa7  :   71 - 0x47
    "01100000", --  168 - 0xa8  :   96 - 0x60
    "01100000", --  169 - 0xa9  :   96 - 0x60
    "01100000", --  170 - 0xaa  :   96 - 0x60
    "01100000", --  171 - 0xab  :   96 - 0x60
    "01100000", --  172 - 0xac  :   96 - 0x60
    "01100000", --  173 - 0xad  :   96 - 0x60
    "01100000", --  174 - 0xae  :   96 - 0x60
    "01100000", --  175 - 0xaf  :   96 - 0x60
    "11111111", --  176 - 0xb0  :  255 - 0xff -- Sprite 0xb
    "11111110", --  177 - 0xb1  :  254 - 0xfe
    "11111110", --  178 - 0xb2  :  254 - 0xfe
    "11111100", --  179 - 0xb3  :  252 - 0xfc
    "11111100", --  180 - 0xb4  :  252 - 0xfc
    "11111100", --  181 - 0xb5  :  252 - 0xfc
    "11111100", --  182 - 0xb6  :  252 - 0xfc
    "11111100", --  183 - 0xb7  :  252 - 0xfc
    "00000001", --  184 - 0xb8  :    1 - 0x1
    "00000011", --  185 - 0xb9  :    3 - 0x3
    "00000011", --  186 - 0xba  :    3 - 0x3
    "00000111", --  187 - 0xbb  :    7 - 0x7
    "00000110", --  188 - 0xbc  :    6 - 0x6
    "00000110", --  189 - 0xbd  :    6 - 0x6
    "00000110", --  190 - 0xbe  :    6 - 0x6
    "00000110", --  191 - 0xbf  :    6 - 0x6
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0xc
    "00001000", --  193 - 0xc1  :    8 - 0x8
    "00011100", --  194 - 0xc2  :   28 - 0x1c
    "00111000", --  195 - 0xc3  :   56 - 0x38
    "01110000", --  196 - 0xc4  :  112 - 0x70
    "00100010", --  197 - 0xc5  :   34 - 0x22
    "00000101", --  198 - 0xc6  :    5 - 0x5
    "00000010", --  199 - 0xc7  :    2 - 0x2
    "11000111", --  200 - 0xc8  :  199 - 0xc7
    "10011111", --  201 - 0xc9  :  159 - 0x9f
    "00111111", --  202 - 0xca  :   63 - 0x3f
    "01111111", --  203 - 0xcb  :  127 - 0x7f
    "01111111", --  204 - 0xcc  :  127 - 0x7f
    "11111111", --  205 - 0xcd  :  255 - 0xff
    "11111111", --  206 - 0xce  :  255 - 0xff
    "11111111", --  207 - 0xcf  :  255 - 0xff
    "00000010", --  208 - 0xd0  :    2 - 0x2 -- Sprite 0xd
    "00110001", --  209 - 0xd1  :   49 - 0x31
    "01111000", --  210 - 0xd2  :  120 - 0x78
    "11111000", --  211 - 0xd3  :  248 - 0xf8
    "01110000", --  212 - 0xd4  :  112 - 0x70
    "00100010", --  213 - 0xd5  :   34 - 0x22
    "00000101", --  214 - 0xd6  :    5 - 0x5
    "00000010", --  215 - 0xd7  :    2 - 0x2
    "11100011", --  216 - 0xd8  :  227 - 0xe3
    "11111001", --  217 - 0xd9  :  249 - 0xf9
    "11111100", --  218 - 0xda  :  252 - 0xfc
    "11111110", --  219 - 0xdb  :  254 - 0xfe
    "11111110", --  220 - 0xdc  :  254 - 0xfe
    "11111111", --  221 - 0xdd  :  255 - 0xff
    "11111111", --  222 - 0xde  :  255 - 0xff
    "11111111", --  223 - 0xdf  :  255 - 0xff
    "01111100", --  224 - 0xe0  :  124 - 0x7c -- Sprite 0xe
    "00111100", --  225 - 0xe1  :   60 - 0x3c
    "10011100", --  226 - 0xe2  :  156 - 0x9c
    "10001100", --  227 - 0xe3  :  140 - 0x8c
    "01001100", --  228 - 0xe4  :   76 - 0x4c
    "01000100", --  229 - 0xe5  :   68 - 0x44
    "01000100", --  230 - 0xe6  :   68 - 0x44
    "01000100", --  231 - 0xe7  :   68 - 0x44
    "10000110", --  232 - 0xe8  :  134 - 0x86
    "11000110", --  233 - 0xe9  :  198 - 0xc6
    "11000110", --  234 - 0xea  :  198 - 0xc6
    "11100110", --  235 - 0xeb  :  230 - 0xe6
    "01100110", --  236 - 0xec  :  102 - 0x66
    "01100110", --  237 - 0xed  :  102 - 0x66
    "01100110", --  238 - 0xee  :  102 - 0x66
    "01100110", --  239 - 0xef  :  102 - 0x66
    "01000100", --  240 - 0xf0  :   68 - 0x44 -- Sprite 0xf
    "01000100", --  241 - 0xf1  :   68 - 0x44
    "01000100", --  242 - 0xf2  :   68 - 0x44
    "01000100", --  243 - 0xf3  :   68 - 0x44
    "01000100", --  244 - 0xf4  :   68 - 0x44
    "01000100", --  245 - 0xf5  :   68 - 0x44
    "01000100", --  246 - 0xf6  :   68 - 0x44
    "01000100", --  247 - 0xf7  :   68 - 0x44
    "01100110", --  248 - 0xf8  :  102 - 0x66
    "01100110", --  249 - 0xf9  :  102 - 0x66
    "01100110", --  250 - 0xfa  :  102 - 0x66
    "01100110", --  251 - 0xfb  :  102 - 0x66
    "01100110", --  252 - 0xfc  :  102 - 0x66
    "01100110", --  253 - 0xfd  :  102 - 0x66
    "01100110", --  254 - 0xfe  :  102 - 0x66
    "01100110", --  255 - 0xff  :  102 - 0x66
    "01001100", --  256 - 0x100  :   76 - 0x4c -- Sprite 0x10
    "00100100", --  257 - 0x101  :   36 - 0x24
    "00100100", --  258 - 0x102  :   36 - 0x24
    "10010100", --  259 - 0x103  :  148 - 0x94
    "00010000", --  260 - 0x104  :   16 - 0x10
    "00001000", --  261 - 0x105  :    8 - 0x8
    "00001000", --  262 - 0x106  :    8 - 0x8
    "00000100", --  263 - 0x107  :    4 - 0x4
    "01100110", --  264 - 0x108  :  102 - 0x66
    "00110110", --  265 - 0x109  :   54 - 0x36
    "10110110", --  266 - 0x10a  :  182 - 0xb6
    "10011110", --  267 - 0x10b  :  158 - 0x9e
    "11011110", --  268 - 0x10c  :  222 - 0xde
    "11001110", --  269 - 0x10d  :  206 - 0xce
    "11101110", --  270 - 0x10e  :  238 - 0xee
    "11100110", --  271 - 0x10f  :  230 - 0xe6
    "00000000", --  272 - 0x110  :    0 - 0x0 -- Sprite 0x11
    "00111100", --  273 - 0x111  :   60 - 0x3c
    "01000000", --  274 - 0x112  :   64 - 0x40
    "01000100", --  275 - 0x113  :   68 - 0x44
    "01000100", --  276 - 0x114  :   68 - 0x44
    "01000100", --  277 - 0x115  :   68 - 0x44
    "01000100", --  278 - 0x116  :   68 - 0x44
    "01000100", --  279 - 0x117  :   68 - 0x44
    "10000001", --  280 - 0x118  :  129 - 0x81
    "00111100", --  281 - 0x119  :   60 - 0x3c
    "01111110", --  282 - 0x11a  :  126 - 0x7e
    "01100110", --  283 - 0x11b  :  102 - 0x66
    "01100110", --  284 - 0x11c  :  102 - 0x66
    "01100110", --  285 - 0x11d  :  102 - 0x66
    "01100110", --  286 - 0x11e  :  102 - 0x66
    "01100110", --  287 - 0x11f  :  102 - 0x66
    "00000100", --  288 - 0x120  :    4 - 0x4 -- Sprite 0x12
    "00010010", --  289 - 0x121  :   18 - 0x12
    "00110010", --  290 - 0x122  :   50 - 0x32
    "01111000", --  291 - 0x123  :  120 - 0x78
    "11111000", --  292 - 0x124  :  248 - 0xf8
    "01110000", --  293 - 0x125  :  112 - 0x70
    "00100100", --  294 - 0x126  :   36 - 0x24
    "00000000", --  295 - 0x127  :    0 - 0x0
    "11110110", --  296 - 0x128  :  246 - 0xf6
    "11110010", --  297 - 0x129  :  242 - 0xf2
    "11111010", --  298 - 0x12a  :  250 - 0xfa
    "11111000", --  299 - 0x12b  :  248 - 0xf8
    "11111100", --  300 - 0x12c  :  252 - 0xfc
    "11111100", --  301 - 0x12d  :  252 - 0xfc
    "11111110", --  302 - 0x12e  :  254 - 0xfe
    "11111110", --  303 - 0x12f  :  254 - 0xfe
    "01000100", --  304 - 0x130  :   68 - 0x44 -- Sprite 0x13
    "01000100", --  305 - 0x131  :   68 - 0x44
    "01000100", --  306 - 0x132  :   68 - 0x44
    "01000100", --  307 - 0x133  :   68 - 0x44
    "01000100", --  308 - 0x134  :   68 - 0x44
    "01000100", --  309 - 0x135  :   68 - 0x44
    "01000100", --  310 - 0x136  :   68 - 0x44
    "01011100", --  311 - 0x137  :   92 - 0x5c
    "01100110", --  312 - 0x138  :  102 - 0x66
    "01100110", --  313 - 0x139  :  102 - 0x66
    "01100110", --  314 - 0x13a  :  102 - 0x66
    "01100110", --  315 - 0x13b  :  102 - 0x66
    "01100110", --  316 - 0x13c  :  102 - 0x66
    "01100110", --  317 - 0x13d  :  102 - 0x66
    "01100110", --  318 - 0x13e  :  102 - 0x66
    "01111110", --  319 - 0x13f  :  126 - 0x7e
    "00010000", --  320 - 0x140  :   16 - 0x10 -- Sprite 0x14
    "00111000", --  321 - 0x141  :   56 - 0x38
    "00111100", --  322 - 0x142  :   60 - 0x3c
    "00111000", --  323 - 0x143  :   56 - 0x38
    "00010000", --  324 - 0x144  :   16 - 0x10
    "00000010", --  325 - 0x145  :    2 - 0x2
    "01000101", --  326 - 0x146  :   69 - 0x45
    "01000010", --  327 - 0x147  :   66 - 0x42
    "11111111", --  328 - 0x148  :  255 - 0xff
    "01111111", --  329 - 0x149  :  127 - 0x7f
    "01111111", --  330 - 0x14a  :  127 - 0x7f
    "00111111", --  331 - 0x14b  :   63 - 0x3f
    "00111111", --  332 - 0x14c  :   63 - 0x3f
    "00011111", --  333 - 0x14d  :   31 - 0x1f
    "01011111", --  334 - 0x14e  :   95 - 0x5f
    "01001111", --  335 - 0x14f  :   79 - 0x4f
    "01000100", --  336 - 0x150  :   68 - 0x44 -- Sprite 0x15
    "01000100", --  337 - 0x151  :   68 - 0x44
    "01000100", --  338 - 0x152  :   68 - 0x44
    "01000100", --  339 - 0x153  :   68 - 0x44
    "01000100", --  340 - 0x154  :   68 - 0x44
    "01011100", --  341 - 0x155  :   92 - 0x5c
    "01000000", --  342 - 0x156  :   64 - 0x40
    "00000000", --  343 - 0x157  :    0 - 0x0
    "01100110", --  344 - 0x158  :  102 - 0x66
    "01100110", --  345 - 0x159  :  102 - 0x66
    "01100110", --  346 - 0x15a  :  102 - 0x66
    "01100110", --  347 - 0x15b  :  102 - 0x66
    "01100110", --  348 - 0x15c  :  102 - 0x66
    "01111110", --  349 - 0x15d  :  126 - 0x7e
    "01111110", --  350 - 0x15e  :  126 - 0x7e
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "01000000", --  352 - 0x160  :   64 - 0x40 -- Sprite 0x16
    "01000000", --  353 - 0x161  :   64 - 0x40
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00011000", --  356 - 0x164  :   24 - 0x18
    "00111000", --  357 - 0x165  :   56 - 0x38
    "00010000", --  358 - 0x166  :   16 - 0x10
    "00000000", --  359 - 0x167  :    0 - 0x0
    "01111110", --  360 - 0x168  :  126 - 0x7e
    "01100110", --  361 - 0x169  :  102 - 0x66
    "01000010", --  362 - 0x16a  :   66 - 0x42
    "00011000", --  363 - 0x16b  :   24 - 0x18
    "00111100", --  364 - 0x16c  :   60 - 0x3c
    "01111110", --  365 - 0x16d  :  126 - 0x7e
    "11111111", --  366 - 0x16e  :  255 - 0xff
    "11111111", --  367 - 0x16f  :  255 - 0xff
    "01000000", --  368 - 0x170  :   64 - 0x40 -- Sprite 0x17
    "01000000", --  369 - 0x171  :   64 - 0x40
    "01000000", --  370 - 0x172  :   64 - 0x40
    "01000000", --  371 - 0x173  :   64 - 0x40
    "01010000", --  372 - 0x174  :   80 - 0x50
    "01010000", --  373 - 0x175  :   80 - 0x50
    "01001000", --  374 - 0x176  :   72 - 0x48
    "01001000", --  375 - 0x177  :   72 - 0x48
    "01101111", --  376 - 0x178  :  111 - 0x6f
    "01100111", --  377 - 0x179  :  103 - 0x67
    "01110111", --  378 - 0x17a  :  119 - 0x77
    "01110011", --  379 - 0x17b  :  115 - 0x73
    "01111011", --  380 - 0x17c  :  123 - 0x7b
    "01111001", --  381 - 0x17d  :  121 - 0x79
    "01101101", --  382 - 0x17e  :  109 - 0x6d
    "01101100", --  383 - 0x17f  :  108 - 0x6c
    "01000111", --  384 - 0x180  :   71 - 0x47 -- Sprite 0x18
    "01000111", --  385 - 0x181  :   71 - 0x47
    "01000111", --  386 - 0x182  :   71 - 0x47
    "01000111", --  387 - 0x183  :   71 - 0x47
    "01000111", --  388 - 0x184  :   71 - 0x47
    "01011111", --  389 - 0x185  :   95 - 0x5f
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00000000", --  391 - 0x187  :    0 - 0x0
    "01100000", --  392 - 0x188  :   96 - 0x60
    "01100000", --  393 - 0x189  :   96 - 0x60
    "01100000", --  394 - 0x18a  :   96 - 0x60
    "01100000", --  395 - 0x18b  :   96 - 0x60
    "01100000", --  396 - 0x18c  :   96 - 0x60
    "01111111", --  397 - 0x18d  :  127 - 0x7f
    "01111111", --  398 - 0x18e  :  127 - 0x7f
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "11111100", --  400 - 0x190  :  252 - 0xfc -- Sprite 0x19
    "11111100", --  401 - 0x191  :  252 - 0xfc
    "11111100", --  402 - 0x192  :  252 - 0xfc
    "11111100", --  403 - 0x193  :  252 - 0xfc
    "11111100", --  404 - 0x194  :  252 - 0xfc
    "11011100", --  405 - 0x195  :  220 - 0xdc
    "00011100", --  406 - 0x196  :   28 - 0x1c
    "01000100", --  407 - 0x197  :   68 - 0x44
    "00000110", --  408 - 0x198  :    6 - 0x6
    "00000110", --  409 - 0x199  :    6 - 0x6
    "00000110", --  410 - 0x19a  :    6 - 0x6
    "00000110", --  411 - 0x19b  :    6 - 0x6
    "00000110", --  412 - 0x19c  :    6 - 0x6
    "11100110", --  413 - 0x19d  :  230 - 0xe6
    "11100110", --  414 - 0x19e  :  230 - 0xe6
    "01100110", --  415 - 0x19f  :  102 - 0x66
    "00010000", --  416 - 0x1a0  :   16 - 0x10 -- Sprite 0x1a
    "00111000", --  417 - 0x1a1  :   56 - 0x38
    "01111100", --  418 - 0x1a2  :  124 - 0x7c
    "11100000", --  419 - 0x1a3  :  224 - 0xe0
    "01000000", --  420 - 0x1a4  :   64 - 0x40
    "00000000", --  421 - 0x1a5  :    0 - 0x0
    "00010000", --  422 - 0x1a6  :   16 - 0x10
    "00100000", --  423 - 0x1a7  :   32 - 0x20
    "11111111", --  424 - 0x1a8  :  255 - 0xff
    "11111111", --  425 - 0x1a9  :  255 - 0xff
    "11111111", --  426 - 0x1aa  :  255 - 0xff
    "11111111", --  427 - 0x1ab  :  255 - 0xff
    "11100111", --  428 - 0x1ac  :  231 - 0xe7
    "11000011", --  429 - 0x1ad  :  195 - 0xc3
    "10011001", --  430 - 0x1ae  :  153 - 0x99
    "00111100", --  431 - 0x1af  :   60 - 0x3c
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x1b
    "01111100", --  433 - 0x1b1  :  124 - 0x7c
    "01000000", --  434 - 0x1b2  :   64 - 0x40
    "01000100", --  435 - 0x1b3  :   68 - 0x44
    "01000100", --  436 - 0x1b4  :   68 - 0x44
    "01000100", --  437 - 0x1b5  :   68 - 0x44
    "01000100", --  438 - 0x1b6  :   68 - 0x44
    "01000100", --  439 - 0x1b7  :   68 - 0x44
    "00000000", --  440 - 0x1b8  :    0 - 0x0
    "01111110", --  441 - 0x1b9  :  126 - 0x7e
    "01111110", --  442 - 0x1ba  :  126 - 0x7e
    "01100110", --  443 - 0x1bb  :  102 - 0x66
    "01100110", --  444 - 0x1bc  :  102 - 0x66
    "01100110", --  445 - 0x1bd  :  102 - 0x66
    "01100110", --  446 - 0x1be  :  102 - 0x66
    "01100110", --  447 - 0x1bf  :  102 - 0x66
    "00010000", --  448 - 0x1c0  :   16 - 0x10 -- Sprite 0x1c
    "00111000", --  449 - 0x1c1  :   56 - 0x38
    "01110001", --  450 - 0x1c2  :  113 - 0x71
    "11100010", --  451 - 0x1c3  :  226 - 0xe2
    "01000100", --  452 - 0x1c4  :   68 - 0x44
    "00001000", --  453 - 0x1c5  :    8 - 0x8
    "00010000", --  454 - 0x1c6  :   16 - 0x10
    "00100000", --  455 - 0x1c7  :   32 - 0x20
    "11111110", --  456 - 0x1c8  :  254 - 0xfe
    "11111100", --  457 - 0x1c9  :  252 - 0xfc
    "11111001", --  458 - 0x1ca  :  249 - 0xf9
    "11110011", --  459 - 0x1cb  :  243 - 0xf3
    "11100111", --  460 - 0x1cc  :  231 - 0xe7
    "11001110", --  461 - 0x1cd  :  206 - 0xce
    "10011100", --  462 - 0x1ce  :  156 - 0x9c
    "00111000", --  463 - 0x1cf  :   56 - 0x38
    "01000000", --  464 - 0x1d0  :   64 - 0x40 -- Sprite 0x1d
    "10000100", --  465 - 0x1d1  :  132 - 0x84
    "00000010", --  466 - 0x1d2  :    2 - 0x2
    "00000111", --  467 - 0x1d3  :    7 - 0x7
    "00001111", --  468 - 0x1d4  :   15 - 0xf
    "00011111", --  469 - 0x1d5  :   31 - 0x1f
    "00111111", --  470 - 0x1d6  :   63 - 0x3f
    "01111111", --  471 - 0x1d7  :  127 - 0x7f
    "01111110", --  472 - 0x1d8  :  126 - 0x7e
    "11100111", --  473 - 0x1d9  :  231 - 0xe7
    "11000011", --  474 - 0x1da  :  195 - 0xc3
    "10000001", --  475 - 0x1db  :  129 - 0x81
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00010000", --  480 - 0x1e0  :   16 - 0x10 -- Sprite 0x1e
    "00011000", --  481 - 0x1e1  :   24 - 0x18
    "00001100", --  482 - 0x1e2  :   12 - 0xc
    "00000110", --  483 - 0x1e3  :    6 - 0x6
    "10000000", --  484 - 0x1e4  :  128 - 0x80
    "11000000", --  485 - 0x1e5  :  192 - 0xc0
    "11100000", --  486 - 0x1e6  :  224 - 0xe0
    "11110000", --  487 - 0x1e7  :  240 - 0xf0
    "01111111", --  488 - 0x1e8  :  127 - 0x7f
    "00111111", --  489 - 0x1e9  :   63 - 0x3f
    "10011111", --  490 - 0x1ea  :  159 - 0x9f
    "11001111", --  491 - 0x1eb  :  207 - 0xcf
    "11100111", --  492 - 0x1ec  :  231 - 0xe7
    "01110011", --  493 - 0x1ed  :  115 - 0x73
    "00111001", --  494 - 0x1ee  :   57 - 0x39
    "00011100", --  495 - 0x1ef  :   28 - 0x1c
    "11111100", --  496 - 0x1f0  :  252 - 0xfc -- Sprite 0x1f
    "11111101", --  497 - 0x1f1  :  253 - 0xfd
    "11111100", --  498 - 0x1f2  :  252 - 0xfc
    "11111110", --  499 - 0x1f3  :  254 - 0xfe
    "11111110", --  500 - 0x1f4  :  254 - 0xfe
    "11111111", --  501 - 0x1f5  :  255 - 0xff
    "11111111", --  502 - 0x1f6  :  255 - 0xff
    "11111111", --  503 - 0x1f7  :  255 - 0xff
    "00000110", --  504 - 0x1f8  :    6 - 0x6
    "00000111", --  505 - 0x1f9  :    7 - 0x7
    "00000111", --  506 - 0x1fa  :    7 - 0x7
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Sprite 0x20
    "11111111", --  513 - 0x201  :  255 - 0xff
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "11111111", --  517 - 0x205  :  255 - 0xff
    "11111111", --  518 - 0x206  :  255 - 0xff
    "11111111", --  519 - 0x207  :  255 - 0xff
    "00000000", --  520 - 0x208  :    0 - 0x0
    "11111111", --  521 - 0x209  :  255 - 0xff
    "11111111", --  522 - 0x20a  :  255 - 0xff
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "01000100", --  528 - 0x210  :   68 - 0x44 -- Sprite 0x21
    "11000101", --  529 - 0x211  :  197 - 0xc5
    "00000000", --  530 - 0x212  :    0 - 0x0
    "00000110", --  531 - 0x213  :    6 - 0x6
    "00000110", --  532 - 0x214  :    6 - 0x6
    "11111111", --  533 - 0x215  :  255 - 0xff
    "11111111", --  534 - 0x216  :  255 - 0xff
    "11111111", --  535 - 0x217  :  255 - 0xff
    "01100110", --  536 - 0x218  :  102 - 0x66
    "11100111", --  537 - 0x219  :  231 - 0xe7
    "11100111", --  538 - 0x21a  :  231 - 0xe7
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "01000000", --  544 - 0x220  :   64 - 0x40 -- Sprite 0x22
    "10000001", --  545 - 0x221  :  129 - 0x81
    "00000011", --  546 - 0x222  :    3 - 0x3
    "00000111", --  547 - 0x223  :    7 - 0x7
    "00001111", --  548 - 0x224  :   15 - 0xf
    "11111111", --  549 - 0x225  :  255 - 0xff
    "11111111", --  550 - 0x226  :  255 - 0xff
    "11111111", --  551 - 0x227  :  255 - 0xff
    "01110000", --  552 - 0x228  :  112 - 0x70
    "11100000", --  553 - 0x229  :  224 - 0xe0
    "11000000", --  554 - 0x22a  :  192 - 0xc0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "11111000", --  560 - 0x230  :  248 - 0xf8 -- Sprite 0x23
    "11111100", --  561 - 0x231  :  252 - 0xfc
    "11111110", --  562 - 0x232  :  254 - 0xfe
    "11111110", --  563 - 0x233  :  254 - 0xfe
    "11111111", --  564 - 0x234  :  255 - 0xff
    "11111111", --  565 - 0x235  :  255 - 0xff
    "11111111", --  566 - 0x236  :  255 - 0xff
    "11111111", --  567 - 0x237  :  255 - 0xff
    "00001110", --  568 - 0x238  :   14 - 0xe
    "00000111", --  569 - 0x239  :    7 - 0x7
    "00000011", --  570 - 0x23a  :    3 - 0x3
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "01000111", --  576 - 0x240  :   71 - 0x47 -- Sprite 0x24
    "11000111", --  577 - 0x241  :  199 - 0xc7
    "00000111", --  578 - 0x242  :    7 - 0x7
    "00000111", --  579 - 0x243  :    7 - 0x7
    "00000111", --  580 - 0x244  :    7 - 0x7
    "11111111", --  581 - 0x245  :  255 - 0xff
    "11111111", --  582 - 0x246  :  255 - 0xff
    "11111111", --  583 - 0x247  :  255 - 0xff
    "01100000", --  584 - 0x248  :   96 - 0x60
    "11100000", --  585 - 0x249  :  224 - 0xe0
    "11100000", --  586 - 0x24a  :  224 - 0xe0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "11111111", --  592 - 0x250  :  255 - 0xff -- Sprite 0x25
    "11111111", --  593 - 0x251  :  255 - 0xff
    "11111111", --  594 - 0x252  :  255 - 0xff
    "11111111", --  595 - 0x253  :  255 - 0xff
    "11111111", --  596 - 0x254  :  255 - 0xff
    "11111111", --  597 - 0x255  :  255 - 0xff
    "00011111", --  598 - 0x256  :   31 - 0x1f
    "00001111", --  599 - 0x257  :   15 - 0xf
    "00000000", --  600 - 0x258  :    0 - 0x0
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "11000000", --  605 - 0x25d  :  192 - 0xc0
    "11100000", --  606 - 0x25e  :  224 - 0xe0
    "01110000", --  607 - 0x25f  :  112 - 0x70
    "11111111", --  608 - 0x260  :  255 - 0xff -- Sprite 0x26
    "11111111", --  609 - 0x261  :  255 - 0xff
    "11111111", --  610 - 0x262  :  255 - 0xff
    "11111111", --  611 - 0x263  :  255 - 0xff
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111111", --  613 - 0x265  :  255 - 0xff
    "11111100", --  614 - 0x266  :  252 - 0xfc
    "11111000", --  615 - 0x267  :  248 - 0xf8
    "00000000", --  616 - 0x268  :    0 - 0x0
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000011", --  621 - 0x26d  :    3 - 0x3
    "00000111", --  622 - 0x26e  :    7 - 0x7
    "00001110", --  623 - 0x26f  :   14 - 0xe
    "00100111", --  624 - 0x270  :   39 - 0x27 -- Sprite 0x27
    "00010011", --  625 - 0x271  :   19 - 0x13
    "00001001", --  626 - 0x272  :    9 - 0x9
    "11000100", --  627 - 0x273  :  196 - 0xc4
    "01100010", --  628 - 0x274  :   98 - 0x62
    "00100001", --  629 - 0x275  :   33 - 0x21
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00111000", --  632 - 0x278  :   56 - 0x38
    "10011100", --  633 - 0x279  :  156 - 0x9c
    "11001110", --  634 - 0x27a  :  206 - 0xce
    "11100111", --  635 - 0x27b  :  231 - 0xe7
    "11110011", --  636 - 0x27c  :  243 - 0xf3
    "11111001", --  637 - 0x27d  :  249 - 0xf9
    "11111100", --  638 - 0x27e  :  252 - 0xfc
    "11111110", --  639 - 0x27f  :  254 - 0xfe
    "11111111", --  640 - 0x280  :  255 - 0xff -- Sprite 0x28
    "11111111", --  641 - 0x281  :  255 - 0xff
    "11111111", --  642 - 0x282  :  255 - 0xff
    "11111111", --  643 - 0x283  :  255 - 0xff
    "01111111", --  644 - 0x284  :  127 - 0x7f
    "00111110", --  645 - 0x285  :   62 - 0x3e
    "10011100", --  646 - 0x286  :  156 - 0x9c
    "01001000", --  647 - 0x287  :   72 - 0x48
    "00000000", --  648 - 0x288  :    0 - 0x0
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "10000001", --  652 - 0x28c  :  129 - 0x81
    "11000011", --  653 - 0x28d  :  195 - 0xc3
    "11100111", --  654 - 0x28e  :  231 - 0xe7
    "01111110", --  655 - 0x28f  :  126 - 0x7e
    "11110000", --  656 - 0x290  :  240 - 0xf0 -- Sprite 0x29
    "11100000", --  657 - 0x291  :  224 - 0xe0
    "11000000", --  658 - 0x292  :  192 - 0xc0
    "10000000", --  659 - 0x293  :  128 - 0x80
    "00000000", --  660 - 0x294  :    0 - 0x0
    "00000010", --  661 - 0x295  :    2 - 0x2
    "00000101", --  662 - 0x296  :    5 - 0x5
    "00000010", --  663 - 0x297  :    2 - 0x2
    "00011100", --  664 - 0x298  :   28 - 0x1c
    "00111001", --  665 - 0x299  :   57 - 0x39
    "01110011", --  666 - 0x29a  :  115 - 0x73
    "11100111", --  667 - 0x29b  :  231 - 0xe7
    "11001111", --  668 - 0x29c  :  207 - 0xcf
    "10011111", --  669 - 0x29d  :  159 - 0x9f
    "00111111", --  670 - 0x29e  :   63 - 0x3f
    "01111111", --  671 - 0x29f  :  127 - 0x7f
    "01000111", --  672 - 0x2a0  :   71 - 0x47 -- Sprite 0x2a
    "01000110", --  673 - 0x2a1  :   70 - 0x46
    "01000110", --  674 - 0x2a2  :   70 - 0x46
    "01000100", --  675 - 0x2a3  :   68 - 0x44
    "01000100", --  676 - 0x2a4  :   68 - 0x44
    "01000100", --  677 - 0x2a5  :   68 - 0x44
    "01000100", --  678 - 0x2a6  :   68 - 0x44
    "01000100", --  679 - 0x2a7  :   68 - 0x44
    "01100001", --  680 - 0x2a8  :   97 - 0x61
    "01100011", --  681 - 0x2a9  :   99 - 0x63
    "01100011", --  682 - 0x2aa  :   99 - 0x63
    "01100111", --  683 - 0x2ab  :  103 - 0x67
    "01100110", --  684 - 0x2ac  :  102 - 0x66
    "01100110", --  685 - 0x2ad  :  102 - 0x66
    "01100110", --  686 - 0x2ae  :  102 - 0x66
    "01100110", --  687 - 0x2af  :  102 - 0x66
    "01111111", --  688 - 0x2b0  :  127 - 0x7f -- Sprite 0x2b
    "00111111", --  689 - 0x2b1  :   63 - 0x3f
    "10011111", --  690 - 0x2b2  :  159 - 0x9f
    "10001111", --  691 - 0x2b3  :  143 - 0x8f
    "01001111", --  692 - 0x2b4  :   79 - 0x4f
    "01000111", --  693 - 0x2b5  :   71 - 0x47
    "01000111", --  694 - 0x2b6  :   71 - 0x47
    "01000111", --  695 - 0x2b7  :   71 - 0x47
    "10000000", --  696 - 0x2b8  :  128 - 0x80
    "11000000", --  697 - 0x2b9  :  192 - 0xc0
    "11000000", --  698 - 0x2ba  :  192 - 0xc0
    "11100000", --  699 - 0x2bb  :  224 - 0xe0
    "01100000", --  700 - 0x2bc  :   96 - 0x60
    "01100000", --  701 - 0x2bd  :   96 - 0x60
    "01100000", --  702 - 0x2be  :   96 - 0x60
    "01100000", --  703 - 0x2bf  :   96 - 0x60
    "00100000", --  704 - 0x2c0  :   32 - 0x20 -- Sprite 0x2c
    "00010000", --  705 - 0x2c1  :   16 - 0x10
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "11000000", --  707 - 0x2c3  :  192 - 0xc0
    "01100000", --  708 - 0x2c4  :   96 - 0x60
    "00100010", --  709 - 0x2c5  :   34 - 0x22
    "00000101", --  710 - 0x2c6  :    5 - 0x5
    "00000010", --  711 - 0x2c7  :    2 - 0x2
    "00111100", --  712 - 0x2c8  :   60 - 0x3c
    "10011001", --  713 - 0x2c9  :  153 - 0x99
    "11000011", --  714 - 0x2ca  :  195 - 0xc3
    "11100111", --  715 - 0x2cb  :  231 - 0xe7
    "11111111", --  716 - 0x2cc  :  255 - 0xff
    "11111111", --  717 - 0x2cd  :  255 - 0xff
    "11111111", --  718 - 0x2ce  :  255 - 0xff
    "11111111", --  719 - 0x2cf  :  255 - 0xff
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x2d
    "01111111", --  721 - 0x2d1  :  127 - 0x7f
    "01000000", --  722 - 0x2d2  :   64 - 0x40
    "01000000", --  723 - 0x2d3  :   64 - 0x40
    "01000000", --  724 - 0x2d4  :   64 - 0x40
    "01000111", --  725 - 0x2d5  :   71 - 0x47
    "01000111", --  726 - 0x2d6  :   71 - 0x47
    "01000111", --  727 - 0x2d7  :   71 - 0x47
    "00000000", --  728 - 0x2d8  :    0 - 0x0
    "01111111", --  729 - 0x2d9  :  127 - 0x7f
    "01111111", --  730 - 0x2da  :  127 - 0x7f
    "01100000", --  731 - 0x2db  :   96 - 0x60
    "01100000", --  732 - 0x2dc  :   96 - 0x60
    "01100000", --  733 - 0x2dd  :   96 - 0x60
    "01100000", --  734 - 0x2de  :   96 - 0x60
    "01100000", --  735 - 0x2df  :   96 - 0x60
    "01000100", --  736 - 0x2e0  :   68 - 0x44 -- Sprite 0x2e
    "11000100", --  737 - 0x2e1  :  196 - 0xc4
    "00000100", --  738 - 0x2e2  :    4 - 0x4
    "00000100", --  739 - 0x2e3  :    4 - 0x4
    "00000100", --  740 - 0x2e4  :    4 - 0x4
    "11111100", --  741 - 0x2e5  :  252 - 0xfc
    "11111100", --  742 - 0x2e6  :  252 - 0xfc
    "11111100", --  743 - 0x2e7  :  252 - 0xfc
    "01100110", --  744 - 0x2e8  :  102 - 0x66
    "11100110", --  745 - 0x2e9  :  230 - 0xe6
    "11100110", --  746 - 0x2ea  :  230 - 0xe6
    "00000110", --  747 - 0x2eb  :    6 - 0x6
    "00000110", --  748 - 0x2ec  :    6 - 0x6
    "00000110", --  749 - 0x2ed  :    6 - 0x6
    "00000110", --  750 - 0x2ee  :    6 - 0x6
    "00000110", --  751 - 0x2ef  :    6 - 0x6
    "00000001", --  752 - 0x2f0  :    1 - 0x1 -- Sprite 0x2f
    "01111100", --  753 - 0x2f1  :  124 - 0x7c
    "01000000", --  754 - 0x2f2  :   64 - 0x40
    "01000100", --  755 - 0x2f3  :   68 - 0x44
    "01000100", --  756 - 0x2f4  :   68 - 0x44
    "01000100", --  757 - 0x2f5  :   68 - 0x44
    "01000100", --  758 - 0x2f6  :   68 - 0x44
    "01000100", --  759 - 0x2f7  :   68 - 0x44
    "00000001", --  760 - 0x2f8  :    1 - 0x1
    "01111100", --  761 - 0x2f9  :  124 - 0x7c
    "01111110", --  762 - 0x2fa  :  126 - 0x7e
    "01100110", --  763 - 0x2fb  :  102 - 0x66
    "01100110", --  764 - 0x2fc  :  102 - 0x66
    "01100110", --  765 - 0x2fd  :  102 - 0x66
    "01100110", --  766 - 0x2fe  :  102 - 0x66
    "01100110", --  767 - 0x2ff  :  102 - 0x66
    "00010000", --  768 - 0x300  :   16 - 0x10 -- Sprite 0x30
    "00111000", --  769 - 0x301  :   56 - 0x38
    "00111100", --  770 - 0x302  :   60 - 0x3c
    "00011000", --  771 - 0x303  :   24 - 0x18
    "00000000", --  772 - 0x304  :    0 - 0x0
    "01000010", --  773 - 0x305  :   66 - 0x42
    "01000100", --  774 - 0x306  :   68 - 0x44
    "01001000", --  775 - 0x307  :   72 - 0x48
    "11111111", --  776 - 0x308  :  255 - 0xff
    "11111111", --  777 - 0x309  :  255 - 0xff
    "01111110", --  778 - 0x30a  :  126 - 0x7e
    "00111100", --  779 - 0x30b  :   60 - 0x3c
    "00011000", --  780 - 0x30c  :   24 - 0x18
    "01000010", --  781 - 0x30d  :   66 - 0x42
    "01100110", --  782 - 0x30e  :  102 - 0x66
    "01111110", --  783 - 0x30f  :  126 - 0x7e
    "01000111", --  784 - 0x310  :   71 - 0x47 -- Sprite 0x31
    "01011111", --  785 - 0x311  :   95 - 0x5f
    "00000000", --  786 - 0x312  :    0 - 0x0
    "00000000", --  787 - 0x313  :    0 - 0x0
    "01110000", --  788 - 0x314  :  112 - 0x70
    "00100010", --  789 - 0x315  :   34 - 0x22
    "00000101", --  790 - 0x316  :    5 - 0x5
    "00000010", --  791 - 0x317  :    2 - 0x2
    "01100000", --  792 - 0x318  :   96 - 0x60
    "01111111", --  793 - 0x319  :  127 - 0x7f
    "01111111", --  794 - 0x31a  :  127 - 0x7f
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "11111111", --  796 - 0x31c  :  255 - 0xff
    "11111111", --  797 - 0x31d  :  255 - 0xff
    "11111111", --  798 - 0x31e  :  255 - 0xff
    "11111111", --  799 - 0x31f  :  255 - 0xff
    "11111111", --  800 - 0x320  :  255 - 0xff -- Sprite 0x32
    "11111111", --  801 - 0x321  :  255 - 0xff
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "01110000", --  804 - 0x324  :  112 - 0x70
    "00100010", --  805 - 0x325  :   34 - 0x22
    "00000101", --  806 - 0x326  :    5 - 0x5
    "00000010", --  807 - 0x327  :    2 - 0x2
    "00000000", --  808 - 0x328  :    0 - 0x0
    "11111111", --  809 - 0x329  :  255 - 0xff
    "11111111", --  810 - 0x32a  :  255 - 0xff
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "11111111", --  812 - 0x32c  :  255 - 0xff
    "11111111", --  813 - 0x32d  :  255 - 0xff
    "11111111", --  814 - 0x32e  :  255 - 0xff
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "11111111", --  816 - 0x330  :  255 - 0xff -- Sprite 0x33
    "11011111", --  817 - 0x331  :  223 - 0xdf
    "00011111", --  818 - 0x332  :   31 - 0x1f
    "01000111", --  819 - 0x333  :   71 - 0x47
    "01000111", --  820 - 0x334  :   71 - 0x47
    "01000111", --  821 - 0x335  :   71 - 0x47
    "01000111", --  822 - 0x336  :   71 - 0x47
    "01000111", --  823 - 0x337  :   71 - 0x47
    "00000000", --  824 - 0x338  :    0 - 0x0
    "11100000", --  825 - 0x339  :  224 - 0xe0
    "11100000", --  826 - 0x33a  :  224 - 0xe0
    "01100000", --  827 - 0x33b  :   96 - 0x60
    "01100000", --  828 - 0x33c  :   96 - 0x60
    "01100000", --  829 - 0x33d  :   96 - 0x60
    "01100000", --  830 - 0x33e  :   96 - 0x60
    "01100000", --  831 - 0x33f  :   96 - 0x60
    "01000100", --  832 - 0x340  :   68 - 0x44 -- Sprite 0x34
    "01000100", --  833 - 0x341  :   68 - 0x44
    "01000100", --  834 - 0x342  :   68 - 0x44
    "01000100", --  835 - 0x343  :   68 - 0x44
    "01000100", --  836 - 0x344  :   68 - 0x44
    "01000100", --  837 - 0x345  :   68 - 0x44
    "01000100", --  838 - 0x346  :   68 - 0x44
    "01000100", --  839 - 0x347  :   68 - 0x44
    "01111110", --  840 - 0x348  :  126 - 0x7e
    "01100110", --  841 - 0x349  :  102 - 0x66
    "01100110", --  842 - 0x34a  :  102 - 0x66
    "01100110", --  843 - 0x34b  :  102 - 0x66
    "01100110", --  844 - 0x34c  :  102 - 0x66
    "01100110", --  845 - 0x34d  :  102 - 0x66
    "01100110", --  846 - 0x34e  :  102 - 0x66
    "01100110", --  847 - 0x34f  :  102 - 0x66
    "00010000", --  848 - 0x350  :   16 - 0x10 -- Sprite 0x35
    "00111000", --  849 - 0x351  :   56 - 0x38
    "01111100", --  850 - 0x352  :  124 - 0x7c
    "11111000", --  851 - 0x353  :  248 - 0xf8
    "00000000", --  852 - 0x354  :    0 - 0x0
    "01111111", --  853 - 0x355  :  127 - 0x7f
    "01000000", --  854 - 0x356  :   64 - 0x40
    "01000000", --  855 - 0x357  :   64 - 0x40
    "11111111", --  856 - 0x358  :  255 - 0xff
    "11111111", --  857 - 0x359  :  255 - 0xff
    "11111111", --  858 - 0x35a  :  255 - 0xff
    "11111111", --  859 - 0x35b  :  255 - 0xff
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "01111111", --  861 - 0x35d  :  127 - 0x7f
    "01111111", --  862 - 0x35e  :  127 - 0x7f
    "01100000", --  863 - 0x35f  :   96 - 0x60
    "00010000", --  864 - 0x360  :   16 - 0x10 -- Sprite 0x36
    "00111000", --  865 - 0x361  :   56 - 0x38
    "01111100", --  866 - 0x362  :  124 - 0x7c
    "11111000", --  867 - 0x363  :  248 - 0xf8
    "00000000", --  868 - 0x364  :    0 - 0x0
    "11111111", --  869 - 0x365  :  255 - 0xff
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "11111111", --  872 - 0x368  :  255 - 0xff
    "11111111", --  873 - 0x369  :  255 - 0xff
    "11111111", --  874 - 0x36a  :  255 - 0xff
    "11111111", --  875 - 0x36b  :  255 - 0xff
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "11111111", --  877 - 0x36d  :  255 - 0xff
    "11111111", --  878 - 0x36e  :  255 - 0xff
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "01000111", --  880 - 0x370  :   71 - 0x47 -- Sprite 0x37
    "01000111", --  881 - 0x371  :   71 - 0x47
    "01000111", --  882 - 0x372  :   71 - 0x47
    "01000111", --  883 - 0x373  :   71 - 0x47
    "01000111", --  884 - 0x374  :   71 - 0x47
    "11000111", --  885 - 0x375  :  199 - 0xc7
    "00000111", --  886 - 0x376  :    7 - 0x7
    "00000111", --  887 - 0x377  :    7 - 0x7
    "01100000", --  888 - 0x378  :   96 - 0x60
    "01100000", --  889 - 0x379  :   96 - 0x60
    "01100000", --  890 - 0x37a  :   96 - 0x60
    "01100000", --  891 - 0x37b  :   96 - 0x60
    "01100000", --  892 - 0x37c  :   96 - 0x60
    "11100000", --  893 - 0x37d  :  224 - 0xe0
    "11100000", --  894 - 0x37e  :  224 - 0xe0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "01000100", --  896 - 0x380  :   68 - 0x44 -- Sprite 0x38
    "01000100", --  897 - 0x381  :   68 - 0x44
    "01000100", --  898 - 0x382  :   68 - 0x44
    "01000100", --  899 - 0x383  :   68 - 0x44
    "01000100", --  900 - 0x384  :   68 - 0x44
    "01011000", --  901 - 0x385  :   88 - 0x58
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "01100110", --  904 - 0x388  :  102 - 0x66
    "01100110", --  905 - 0x389  :  102 - 0x66
    "01100110", --  906 - 0x38a  :  102 - 0x66
    "01100110", --  907 - 0x38b  :  102 - 0x66
    "01100110", --  908 - 0x38c  :  102 - 0x66
    "01111110", --  909 - 0x38d  :  126 - 0x7e
    "01111100", --  910 - 0x38e  :  124 - 0x7c
    "00000001", --  911 - 0x38f  :    1 - 0x1
    "00010000", --  912 - 0x390  :   16 - 0x10 -- Sprite 0x39
    "00111000", --  913 - 0x391  :   56 - 0x38
    "01111100", --  914 - 0x392  :  124 - 0x7c
    "11111000", --  915 - 0x393  :  248 - 0xf8
    "01110000", --  916 - 0x394  :  112 - 0x70
    "00100010", --  917 - 0x395  :   34 - 0x22
    "00000100", --  918 - 0x396  :    4 - 0x4
    "00000000", --  919 - 0x397  :    0 - 0x0
    "11111111", --  920 - 0x398  :  255 - 0xff
    "11111111", --  921 - 0x399  :  255 - 0xff
    "11111111", --  922 - 0x39a  :  255 - 0xff
    "11111111", --  923 - 0x39b  :  255 - 0xff
    "11111111", --  924 - 0x39c  :  255 - 0xff
    "11111111", --  925 - 0x39d  :  255 - 0xff
    "11111111", --  926 - 0x39e  :  255 - 0xff
    "11111110", --  927 - 0x39f  :  254 - 0xfe
    "01000100", --  928 - 0x3a0  :   68 - 0x44 -- Sprite 0x3a
    "01000100", --  929 - 0x3a1  :   68 - 0x44
    "01000100", --  930 - 0x3a2  :   68 - 0x44
    "01000100", --  931 - 0x3a3  :   68 - 0x44
    "01000100", --  932 - 0x3a4  :   68 - 0x44
    "01011000", --  933 - 0x3a5  :   88 - 0x58
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "01100110", --  936 - 0x3a8  :  102 - 0x66
    "01100110", --  937 - 0x3a9  :  102 - 0x66
    "01100110", --  938 - 0x3aa  :  102 - 0x66
    "01100110", --  939 - 0x3ab  :  102 - 0x66
    "01100110", --  940 - 0x3ac  :  102 - 0x66
    "01111110", --  941 - 0x3ad  :  126 - 0x7e
    "00111100", --  942 - 0x3ae  :   60 - 0x3c
    "10000001", --  943 - 0x3af  :  129 - 0x81
    "01000000", --  944 - 0x3b0  :   64 - 0x40 -- Sprite 0x3b
    "01000111", --  945 - 0x3b1  :   71 - 0x47
    "01000111", --  946 - 0x3b2  :   71 - 0x47
    "01000111", --  947 - 0x3b3  :   71 - 0x47
    "01000111", --  948 - 0x3b4  :   71 - 0x47
    "01011111", --  949 - 0x3b5  :   95 - 0x5f
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "01100000", --  952 - 0x3b8  :   96 - 0x60
    "01100000", --  953 - 0x3b9  :   96 - 0x60
    "01100000", --  954 - 0x3ba  :   96 - 0x60
    "01100000", --  955 - 0x3bb  :   96 - 0x60
    "01100000", --  956 - 0x3bc  :   96 - 0x60
    "01111111", --  957 - 0x3bd  :  127 - 0x7f
    "01111111", --  958 - 0x3be  :  127 - 0x7f
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x3c
    "11111111", --  961 - 0x3c1  :  255 - 0xff
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "11111111", --  963 - 0x3c3  :  255 - 0xff
    "11111111", --  964 - 0x3c4  :  255 - 0xff
    "11111111", --  965 - 0x3c5  :  255 - 0xff
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "11111111", --  973 - 0x3cd  :  255 - 0xff
    "11111111", --  974 - 0x3ce  :  255 - 0xff
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000111", --  976 - 0x3d0  :    7 - 0x7 -- Sprite 0x3d
    "11111111", --  977 - 0x3d1  :  255 - 0xff
    "11111111", --  978 - 0x3d2  :  255 - 0xff
    "11111111", --  979 - 0x3d3  :  255 - 0xff
    "11111111", --  980 - 0x3d4  :  255 - 0xff
    "11111111", --  981 - 0x3d5  :  255 - 0xff
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "11111111", --  989 - 0x3dd  :  255 - 0xff
    "11111111", --  990 - 0x3de  :  255 - 0xff
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00010000", --  992 - 0x3e0  :   16 - 0x10 -- Sprite 0x3e
    "00111000", --  993 - 0x3e1  :   56 - 0x38
    "01110001", --  994 - 0x3e2  :  113 - 0x71
    "11100010", --  995 - 0x3e3  :  226 - 0xe2
    "01100010", --  996 - 0x3e4  :   98 - 0x62
    "00100001", --  997 - 0x3e5  :   33 - 0x21
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "11111110", -- 1000 - 0x3e8  :  254 - 0xfe
    "11111100", -- 1001 - 0x3e9  :  252 - 0xfc
    "11111001", -- 1002 - 0x3ea  :  249 - 0xf9
    "11110011", -- 1003 - 0x3eb  :  243 - 0xf3
    "11110011", -- 1004 - 0x3ec  :  243 - 0xf3
    "11111001", -- 1005 - 0x3ed  :  249 - 0xf9
    "11111100", -- 1006 - 0x3ee  :  252 - 0xfc
    "11111110", -- 1007 - 0x3ef  :  254 - 0xfe
    "10000111", -- 1008 - 0x3f0  :  135 - 0x87 -- Sprite 0x3f
    "10000111", -- 1009 - 0x3f1  :  135 - 0x87
    "00000111", -- 1010 - 0x3f2  :    7 - 0x7
    "00001111", -- 1011 - 0x3f3  :   15 - 0xf
    "00001111", -- 1012 - 0x3f4  :   15 - 0xf
    "00011111", -- 1013 - 0x3f5  :   31 - 0x1f
    "10011111", -- 1014 - 0x3f6  :  159 - 0x9f
    "10001111", -- 1015 - 0x3f7  :  143 - 0x8f
    "11100000", -- 1016 - 0x3f8  :  224 - 0xe0
    "11000000", -- 1017 - 0x3f9  :  192 - 0xc0
    "11000000", -- 1018 - 0x3fa  :  192 - 0xc0
    "10000000", -- 1019 - 0x3fb  :  128 - 0x80
    "10000000", -- 1020 - 0x3fc  :  128 - 0x80
    "11000000", -- 1021 - 0x3fd  :  192 - 0xc0
    "11000000", -- 1022 - 0x3fe  :  192 - 0xc0
    "11100000", -- 1023 - 0x3ff  :  224 - 0xe0
    "01000100", -- 1024 - 0x400  :   68 - 0x44 -- Sprite 0x40
    "01000100", -- 1025 - 0x401  :   68 - 0x44
    "01000100", -- 1026 - 0x402  :   68 - 0x44
    "01000100", -- 1027 - 0x403  :   68 - 0x44
    "01000100", -- 1028 - 0x404  :   68 - 0x44
    "01000110", -- 1029 - 0x405  :   70 - 0x46
    "01000110", -- 1030 - 0x406  :   70 - 0x46
    "01000111", -- 1031 - 0x407  :   71 - 0x47
    "01100110", -- 1032 - 0x408  :  102 - 0x66
    "01100110", -- 1033 - 0x409  :  102 - 0x66
    "01100110", -- 1034 - 0x40a  :  102 - 0x66
    "01100110", -- 1035 - 0x40b  :  102 - 0x66
    "01100111", -- 1036 - 0x40c  :  103 - 0x67
    "01100011", -- 1037 - 0x40d  :   99 - 0x63
    "01100011", -- 1038 - 0x40e  :   99 - 0x63
    "01100001", -- 1039 - 0x40f  :   97 - 0x61
    "00010000", -- 1040 - 0x410  :   16 - 0x10 -- Sprite 0x41
    "00111000", -- 1041 - 0x411  :   56 - 0x38
    "01111100", -- 1042 - 0x412  :  124 - 0x7c
    "01111000", -- 1043 - 0x413  :  120 - 0x78
    "00110000", -- 1044 - 0x414  :   48 - 0x30
    "00000010", -- 1045 - 0x415  :    2 - 0x2
    "00000101", -- 1046 - 0x416  :    5 - 0x5
    "00000010", -- 1047 - 0x417  :    2 - 0x2
    "11111111", -- 1048 - 0x418  :  255 - 0xff
    "11111111", -- 1049 - 0x419  :  255 - 0xff
    "11111111", -- 1050 - 0x41a  :  255 - 0xff
    "01111111", -- 1051 - 0x41b  :  127 - 0x7f
    "01111111", -- 1052 - 0x41c  :  127 - 0x7f
    "00111111", -- 1053 - 0x41d  :   63 - 0x3f
    "10011111", -- 1054 - 0x41e  :  159 - 0x9f
    "11000111", -- 1055 - 0x41f  :  199 - 0xc7
    "00010000", -- 1056 - 0x420  :   16 - 0x10 -- Sprite 0x42
    "00111000", -- 1057 - 0x421  :   56 - 0x38
    "01111100", -- 1058 - 0x422  :  124 - 0x7c
    "11111000", -- 1059 - 0x423  :  248 - 0xf8
    "01110000", -- 1060 - 0x424  :  112 - 0x70
    "00100000", -- 1061 - 0x425  :   32 - 0x20
    "00000001", -- 1062 - 0x426  :    1 - 0x1
    "00000010", -- 1063 - 0x427  :    2 - 0x2
    "11111111", -- 1064 - 0x428  :  255 - 0xff
    "11111111", -- 1065 - 0x429  :  255 - 0xff
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "11111110", -- 1067 - 0x42b  :  254 - 0xfe
    "11111110", -- 1068 - 0x42c  :  254 - 0xfe
    "11111100", -- 1069 - 0x42d  :  252 - 0xfc
    "11111001", -- 1070 - 0x42e  :  249 - 0xf9
    "11100011", -- 1071 - 0x42f  :  227 - 0xe3
    "01000100", -- 1072 - 0x430  :   68 - 0x44 -- Sprite 0x43
    "01000100", -- 1073 - 0x431  :   68 - 0x44
    "01000100", -- 1074 - 0x432  :   68 - 0x44
    "01000100", -- 1075 - 0x433  :   68 - 0x44
    "10000100", -- 1076 - 0x434  :  132 - 0x84
    "10000100", -- 1077 - 0x435  :  132 - 0x84
    "00000100", -- 1078 - 0x436  :    4 - 0x4
    "00001100", -- 1079 - 0x437  :   12 - 0xc
    "01100110", -- 1080 - 0x438  :  102 - 0x66
    "01100110", -- 1081 - 0x439  :  102 - 0x66
    "01100110", -- 1082 - 0x43a  :  102 - 0x66
    "01100110", -- 1083 - 0x43b  :  102 - 0x66
    "11100110", -- 1084 - 0x43c  :  230 - 0xe6
    "11000110", -- 1085 - 0x43d  :  198 - 0xc6
    "11000110", -- 1086 - 0x43e  :  198 - 0xc6
    "10000110", -- 1087 - 0x43f  :  134 - 0x86
    "00010000", -- 1088 - 0x440  :   16 - 0x10 -- Sprite 0x44
    "00111000", -- 1089 - 0x441  :   56 - 0x38
    "01111100", -- 1090 - 0x442  :  124 - 0x7c
    "11111000", -- 1091 - 0x443  :  248 - 0xf8
    "01110000", -- 1092 - 0x444  :  112 - 0x70
    "00100010", -- 1093 - 0x445  :   34 - 0x22
    "00000101", -- 1094 - 0x446  :    5 - 0x5
    "00000010", -- 1095 - 0x447  :    2 - 0x2
    "11111110", -- 1096 - 0x448  :  254 - 0xfe
    "11111111", -- 1097 - 0x449  :  255 - 0xff
    "11111111", -- 1098 - 0x44a  :  255 - 0xff
    "11111111", -- 1099 - 0x44b  :  255 - 0xff
    "11111111", -- 1100 - 0x44c  :  255 - 0xff
    "11111111", -- 1101 - 0x44d  :  255 - 0xff
    "11111111", -- 1102 - 0x44e  :  255 - 0xff
    "11111111", -- 1103 - 0x44f  :  255 - 0xff
    "01001111", -- 1104 - 0x450  :   79 - 0x4f -- Sprite 0x45
    "01000111", -- 1105 - 0x451  :   71 - 0x47
    "01000111", -- 1106 - 0x452  :   71 - 0x47
    "01000111", -- 1107 - 0x453  :   71 - 0x47
    "01000111", -- 1108 - 0x454  :   71 - 0x47
    "01000111", -- 1109 - 0x455  :   71 - 0x47
    "01000111", -- 1110 - 0x456  :   71 - 0x47
    "01000111", -- 1111 - 0x457  :   71 - 0x47
    "01100000", -- 1112 - 0x458  :   96 - 0x60
    "01100000", -- 1113 - 0x459  :   96 - 0x60
    "01100000", -- 1114 - 0x45a  :   96 - 0x60
    "01100000", -- 1115 - 0x45b  :   96 - 0x60
    "01100000", -- 1116 - 0x45c  :   96 - 0x60
    "01100000", -- 1117 - 0x45d  :   96 - 0x60
    "01100000", -- 1118 - 0x45e  :   96 - 0x60
    "01100000", -- 1119 - 0x45f  :   96 - 0x60
    "10100000", -- 1120 - 0x460  :  160 - 0xa0 -- Sprite 0x46
    "10011111", -- 1121 - 0x461  :  159 - 0x9f
    "11000000", -- 1122 - 0x462  :  192 - 0xc0
    "11100000", -- 1123 - 0x463  :  224 - 0xe0
    "11111000", -- 1124 - 0x464  :  248 - 0xf8
    "11111111", -- 1125 - 0x465  :  255 - 0xff
    "11111111", -- 1126 - 0x466  :  255 - 0xff
    "11111111", -- 1127 - 0x467  :  255 - 0xff
    "11110000", -- 1128 - 0x468  :  240 - 0xf0
    "01111111", -- 1129 - 0x469  :  127 - 0x7f
    "00011111", -- 1130 - 0x46a  :   31 - 0x1f
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00001100", -- 1136 - 0x470  :   12 - 0xc -- Sprite 0x47
    "11110000", -- 1137 - 0x471  :  240 - 0xf0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "00000001", -- 1140 - 0x474  :    1 - 0x1
    "11111111", -- 1141 - 0x475  :  255 - 0xff
    "11111111", -- 1142 - 0x476  :  255 - 0xff
    "11111111", -- 1143 - 0x477  :  255 - 0xff
    "00001111", -- 1144 - 0x478  :   15 - 0xf
    "11111110", -- 1145 - 0x479  :  254 - 0xfe
    "11111000", -- 1146 - 0x47a  :  248 - 0xf8
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00001100", -- 1152 - 0x480  :   12 - 0xc -- Sprite 0x48
    "00011101", -- 1153 - 0x481  :   29 - 0x1d
    "00111000", -- 1154 - 0x482  :   56 - 0x38
    "01111110", -- 1155 - 0x483  :  126 - 0x7e
    "11111110", -- 1156 - 0x484  :  254 - 0xfe
    "11111111", -- 1157 - 0x485  :  255 - 0xff
    "11111111", -- 1158 - 0x486  :  255 - 0xff
    "11111111", -- 1159 - 0x487  :  255 - 0xff
    "00000110", -- 1160 - 0x488  :    6 - 0x6
    "00000111", -- 1161 - 0x489  :    7 - 0x7
    "00000111", -- 1162 - 0x48a  :    7 - 0x7
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "11111111", -- 1168 - 0x490  :  255 - 0xff -- Sprite 0x49
    "11111111", -- 1169 - 0x491  :  255 - 0xff
    "11111111", -- 1170 - 0x492  :  255 - 0xff
    "11111111", -- 1171 - 0x493  :  255 - 0xff
    "11111111", -- 1172 - 0x494  :  255 - 0xff
    "11111111", -- 1173 - 0x495  :  255 - 0xff
    "11111111", -- 1174 - 0x496  :  255 - 0xff
    "11111111", -- 1175 - 0x497  :  255 - 0xff
    "00000000", -- 1176 - 0x498  :    0 - 0x0
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "11111111", -- 1184 - 0x4a0  :  255 - 0xff -- Sprite 0x4a
    "11101111", -- 1185 - 0x4a1  :  239 - 0xef
    "11111101", -- 1186 - 0x4a2  :  253 - 0xfd
    "11111111", -- 1187 - 0x4a3  :  255 - 0xff
    "11111111", -- 1188 - 0x4a4  :  255 - 0xff
    "11101111", -- 1189 - 0x4a5  :  239 - 0xef
    "11111110", -- 1190 - 0x4a6  :  254 - 0xfe
    "11111111", -- 1191 - 0x4a7  :  255 - 0xff
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0
    "01110110", -- 1193 - 0x4a9  :  118 - 0x76
    "01010111", -- 1194 - 0x4aa  :   87 - 0x57
    "01010101", -- 1195 - 0x4ab  :   85 - 0x55
    "01010101", -- 1196 - 0x4ac  :   85 - 0x55
    "01110101", -- 1197 - 0x4ad  :  117 - 0x75
    "01000111", -- 1198 - 0x4ae  :   71 - 0x47
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "11111111", -- 1200 - 0x4b0  :  255 - 0xff -- Sprite 0x4b
    "11101010", -- 1201 - 0x4b1  :  234 - 0xea
    "11111111", -- 1202 - 0x4b2  :  255 - 0xff
    "10101111", -- 1203 - 0x4b3  :  175 - 0xaf
    "11111111", -- 1204 - 0x4b4  :  255 - 0xff
    "11111111", -- 1205 - 0x4b5  :  255 - 0xff
    "11111010", -- 1206 - 0x4b6  :  250 - 0xfa
    "11111111", -- 1207 - 0x4b7  :  255 - 0xff
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0
    "01110111", -- 1209 - 0x4b9  :  119 - 0x77
    "00010101", -- 1210 - 0x4ba  :   21 - 0x15
    "01110101", -- 1211 - 0x4bb  :  117 - 0x75
    "01000101", -- 1212 - 0x4bc  :   69 - 0x45
    "01000101", -- 1213 - 0x4bd  :   69 - 0x45
    "01110111", -- 1214 - 0x4be  :  119 - 0x77
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Sprite 0x4c
    "11111111", -- 1217 - 0x4c1  :  255 - 0xff
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111111", -- 1219 - 0x4c3  :  255 - 0xff
    "11111111", -- 1220 - 0x4c4  :  255 - 0xff
    "11111111", -- 1221 - 0x4c5  :  255 - 0xff
    "11111110", -- 1222 - 0x4c6  :  254 - 0xfe
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0
    "00100100", -- 1225 - 0x4c9  :   36 - 0x24
    "01101100", -- 1226 - 0x4ca  :  108 - 0x6c
    "00100100", -- 1227 - 0x4cb  :   36 - 0x24
    "00100100", -- 1228 - 0x4cc  :   36 - 0x24
    "00100100", -- 1229 - 0x4cd  :   36 - 0x24
    "00100101", -- 1230 - 0x4ce  :   37 - 0x25
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "11111111", -- 1232 - 0x4d0  :  255 - 0xff -- Sprite 0x4d
    "10111111", -- 1233 - 0x4d1  :  191 - 0xbf
    "11111110", -- 1234 - 0x4d2  :  254 - 0xfe
    "10101111", -- 1235 - 0x4d3  :  175 - 0xaf
    "11111111", -- 1236 - 0x4d4  :  255 - 0xff
    "11111111", -- 1237 - 0x4d5  :  255 - 0xff
    "11101111", -- 1238 - 0x4d6  :  239 - 0xef
    "11111111", -- 1239 - 0x4d7  :  255 - 0xff
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0
    "01110100", -- 1241 - 0x4d9  :  116 - 0x74
    "01000111", -- 1242 - 0x4da  :   71 - 0x47
    "01110101", -- 1243 - 0x4db  :  117 - 0x75
    "00010101", -- 1244 - 0x4dc  :   21 - 0x15
    "00010101", -- 1245 - 0x4dd  :   21 - 0x15
    "01110101", -- 1246 - 0x4de  :  117 - 0x75
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "11111111", -- 1248 - 0x4e0  :  255 - 0xff -- Sprite 0x4e
    "11111111", -- 1249 - 0x4e1  :  255 - 0xff
    "11111011", -- 1250 - 0x4e2  :  251 - 0xfb
    "11111111", -- 1251 - 0x4e3  :  255 - 0xff
    "11111111", -- 1252 - 0x4e4  :  255 - 0xff
    "11111111", -- 1253 - 0x4e5  :  255 - 0xff
    "11111110", -- 1254 - 0x4e6  :  254 - 0xfe
    "11111111", -- 1255 - 0x4e7  :  255 - 0xff
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0
    "01000000", -- 1257 - 0x4e9  :   64 - 0x40
    "00011101", -- 1258 - 0x4ea  :   29 - 0x1d
    "01010101", -- 1259 - 0x4eb  :   85 - 0x55
    "01010001", -- 1260 - 0x4ec  :   81 - 0x51
    "01010001", -- 1261 - 0x4ed  :   81 - 0x51
    "01010001", -- 1262 - 0x4ee  :   81 - 0x51
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "11111111", -- 1264 - 0x4f0  :  255 - 0xff -- Sprite 0x4f
    "11111111", -- 1265 - 0x4f1  :  255 - 0xff
    "11110111", -- 1266 - 0x4f2  :  247 - 0xf7
    "11111110", -- 1267 - 0x4f3  :  254 - 0xfe
    "11111011", -- 1268 - 0x4f4  :  251 - 0xfb
    "11111111", -- 1269 - 0x4f5  :  255 - 0xff
    "11101111", -- 1270 - 0x4f6  :  239 - 0xef
    "11111101", -- 1271 - 0x4f7  :  253 - 0xfd
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "01001000", -- 1274 - 0x4fa  :   72 - 0x48
    "01000001", -- 1275 - 0x4fb  :   65 - 0x41
    "01000100", -- 1276 - 0x4fc  :   68 - 0x44
    "01000000", -- 1277 - 0x4fd  :   64 - 0x40
    "11010000", -- 1278 - 0x4fe  :  208 - 0xd0
    "00000010", -- 1279 - 0x4ff  :    2 - 0x2
    "11111111", -- 1280 - 0x500  :  255 - 0xff -- Sprite 0x50
    "11111111", -- 1281 - 0x501  :  255 - 0xff
    "00000011", -- 1282 - 0x502  :    3 - 0x3
    "00000001", -- 1283 - 0x503  :    1 - 0x1
    "11101110", -- 1284 - 0x504  :  238 - 0xee
    "00000000", -- 1285 - 0x505  :    0 - 0x0
    "11101110", -- 1286 - 0x506  :  238 - 0xee
    "11101110", -- 1287 - 0x507  :  238 - 0xee
    "00000000", -- 1288 - 0x508  :    0 - 0x0
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "11111100", -- 1290 - 0x50a  :  252 - 0xfc
    "11111110", -- 1291 - 0x50b  :  254 - 0xfe
    "11101110", -- 1292 - 0x50c  :  238 - 0xee
    "11101110", -- 1293 - 0x50d  :  238 - 0xee
    "11101110", -- 1294 - 0x50e  :  238 - 0xee
    "11101110", -- 1295 - 0x50f  :  238 - 0xee
    "11111111", -- 1296 - 0x510  :  255 - 0xff -- Sprite 0x51
    "11111111", -- 1297 - 0x511  :  255 - 0xff
    "00000011", -- 1298 - 0x512  :    3 - 0x3
    "00000001", -- 1299 - 0x513  :    1 - 0x1
    "11101110", -- 1300 - 0x514  :  238 - 0xee
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "11101110", -- 1302 - 0x516  :  238 - 0xee
    "11101110", -- 1303 - 0x517  :  238 - 0xee
    "00000000", -- 1304 - 0x518  :    0 - 0x0
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "11111100", -- 1306 - 0x51a  :  252 - 0xfc
    "11111110", -- 1307 - 0x51b  :  254 - 0xfe
    "11101110", -- 1308 - 0x51c  :  238 - 0xee
    "11101110", -- 1309 - 0x51d  :  238 - 0xee
    "11101110", -- 1310 - 0x51e  :  238 - 0xee
    "11101110", -- 1311 - 0x51f  :  238 - 0xee
    "11111111", -- 1312 - 0x520  :  255 - 0xff -- Sprite 0x52
    "11111111", -- 1313 - 0x521  :  255 - 0xff
    "00000001", -- 1314 - 0x522  :    1 - 0x1
    "00000000", -- 1315 - 0x523  :    0 - 0x0
    "11100000", -- 1316 - 0x524  :  224 - 0xe0
    "00001111", -- 1317 - 0x525  :   15 - 0xf
    "11111111", -- 1318 - 0x526  :  255 - 0xff
    "11111011", -- 1319 - 0x527  :  251 - 0xfb
    "00000000", -- 1320 - 0x528  :    0 - 0x0
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "11111110", -- 1322 - 0x52a  :  254 - 0xfe
    "11111110", -- 1323 - 0x52b  :  254 - 0xfe
    "11100000", -- 1324 - 0x52c  :  224 - 0xe0
    "11100000", -- 1325 - 0x52d  :  224 - 0xe0
    "11111000", -- 1326 - 0x52e  :  248 - 0xf8
    "11111000", -- 1327 - 0x52f  :  248 - 0xf8
    "11111111", -- 1328 - 0x530  :  255 - 0xff -- Sprite 0x53
    "11111111", -- 1329 - 0x531  :  255 - 0xff
    "10000011", -- 1330 - 0x532  :  131 - 0x83
    "00000001", -- 1331 - 0x533  :    1 - 0x1
    "11101110", -- 1332 - 0x534  :  238 - 0xee
    "00000000", -- 1333 - 0x535  :    0 - 0x0
    "11111111", -- 1334 - 0x536  :  255 - 0xff
    "11111111", -- 1335 - 0x537  :  255 - 0xff
    "00000000", -- 1336 - 0x538  :    0 - 0x0
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "01111100", -- 1338 - 0x53a  :  124 - 0x7c
    "11111110", -- 1339 - 0x53b  :  254 - 0xfe
    "11101110", -- 1340 - 0x53c  :  238 - 0xee
    "11100000", -- 1341 - 0x53d  :  224 - 0xe0
    "11111100", -- 1342 - 0x53e  :  252 - 0xfc
    "01111110", -- 1343 - 0x53f  :  126 - 0x7e
    "11111111", -- 1344 - 0x540  :  255 - 0xff -- Sprite 0x54
    "11111111", -- 1345 - 0x541  :  255 - 0xff
    "00000001", -- 1346 - 0x542  :    1 - 0x1
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "10111000", -- 1348 - 0x544  :  184 - 0xb8
    "11000011", -- 1349 - 0x545  :  195 - 0xc3
    "11111011", -- 1350 - 0x546  :  251 - 0xfb
    "11111011", -- 1351 - 0x547  :  251 - 0xfb
    "00000000", -- 1352 - 0x548  :    0 - 0x0
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "11111110", -- 1354 - 0x54a  :  254 - 0xfe
    "11111110", -- 1355 - 0x54b  :  254 - 0xfe
    "00111000", -- 1356 - 0x54c  :   56 - 0x38
    "00111000", -- 1357 - 0x54d  :   56 - 0x38
    "00111000", -- 1358 - 0x54e  :   56 - 0x38
    "00111000", -- 1359 - 0x54f  :   56 - 0x38
    "11111111", -- 1360 - 0x550  :  255 - 0xff -- Sprite 0x55
    "11111111", -- 1361 - 0x551  :  255 - 0xff
    "10000011", -- 1362 - 0x552  :  131 - 0x83
    "00000001", -- 1363 - 0x553  :    1 - 0x1
    "11101110", -- 1364 - 0x554  :  238 - 0xee
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "11101110", -- 1366 - 0x556  :  238 - 0xee
    "11101110", -- 1367 - 0x557  :  238 - 0xee
    "00000000", -- 1368 - 0x558  :    0 - 0x0
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "01111100", -- 1370 - 0x55a  :  124 - 0x7c
    "11111110", -- 1371 - 0x55b  :  254 - 0xfe
    "11101110", -- 1372 - 0x55c  :  238 - 0xee
    "11101110", -- 1373 - 0x55d  :  238 - 0xee
    "11101110", -- 1374 - 0x55e  :  238 - 0xee
    "11101110", -- 1375 - 0x55f  :  238 - 0xee
    "11111111", -- 1376 - 0x560  :  255 - 0xff -- Sprite 0x56
    "11111111", -- 1377 - 0x561  :  255 - 0xff
    "00011111", -- 1378 - 0x562  :   31 - 0x1f
    "00001111", -- 1379 - 0x563  :   15 - 0xf
    "11101111", -- 1380 - 0x564  :  239 - 0xef
    "00001111", -- 1381 - 0x565  :   15 - 0xf
    "11101111", -- 1382 - 0x566  :  239 - 0xef
    "11101111", -- 1383 - 0x567  :  239 - 0xef
    "00000000", -- 1384 - 0x568  :    0 - 0x0
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "11100000", -- 1386 - 0x56a  :  224 - 0xe0
    "11100000", -- 1387 - 0x56b  :  224 - 0xe0
    "11100000", -- 1388 - 0x56c  :  224 - 0xe0
    "11100000", -- 1389 - 0x56d  :  224 - 0xe0
    "11100000", -- 1390 - 0x56e  :  224 - 0xe0
    "11100000", -- 1391 - 0x56f  :  224 - 0xe0
    "11111111", -- 1392 - 0x570  :  255 - 0xff -- Sprite 0x57
    "11111111", -- 1393 - 0x571  :  255 - 0xff
    "00010001", -- 1394 - 0x572  :   17 - 0x11
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "11101110", -- 1396 - 0x574  :  238 - 0xee
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "11101110", -- 1398 - 0x576  :  238 - 0xee
    "11101110", -- 1399 - 0x577  :  238 - 0xee
    "00000000", -- 1400 - 0x578  :    0 - 0x0
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "11101110", -- 1402 - 0x57a  :  238 - 0xee
    "11101110", -- 1403 - 0x57b  :  238 - 0xee
    "11101110", -- 1404 - 0x57c  :  238 - 0xee
    "11101110", -- 1405 - 0x57d  :  238 - 0xee
    "11101110", -- 1406 - 0x57e  :  238 - 0xee
    "11101110", -- 1407 - 0x57f  :  238 - 0xee
    "11111111", -- 1408 - 0x580  :  255 - 0xff -- Sprite 0x58
    "11111111", -- 1409 - 0x581  :  255 - 0xff
    "01110001", -- 1410 - 0x582  :  113 - 0x71
    "00110000", -- 1411 - 0x583  :   48 - 0x30
    "11111110", -- 1412 - 0x584  :  254 - 0xfe
    "00000000", -- 1413 - 0x585  :    0 - 0x0
    "11111110", -- 1414 - 0x586  :  254 - 0xfe
    "11101110", -- 1415 - 0x587  :  238 - 0xee
    "00000000", -- 1416 - 0x588  :    0 - 0x0
    "00000000", -- 1417 - 0x589  :    0 - 0x0
    "10001110", -- 1418 - 0x58a  :  142 - 0x8e
    "11001110", -- 1419 - 0x58b  :  206 - 0xce
    "11101110", -- 1420 - 0x58c  :  238 - 0xee
    "11111110", -- 1421 - 0x58d  :  254 - 0xfe
    "11111110", -- 1422 - 0x58e  :  254 - 0xfe
    "11101110", -- 1423 - 0x58f  :  238 - 0xee
    "11111111", -- 1424 - 0x590  :  255 - 0xff -- Sprite 0x59
    "11111111", -- 1425 - 0x591  :  255 - 0xff
    "00000011", -- 1426 - 0x592  :    3 - 0x3
    "00000001", -- 1427 - 0x593  :    1 - 0x1
    "11101110", -- 1428 - 0x594  :  238 - 0xee
    "00000000", -- 1429 - 0x595  :    0 - 0x0
    "11101110", -- 1430 - 0x596  :  238 - 0xee
    "11101110", -- 1431 - 0x597  :  238 - 0xee
    "00000000", -- 1432 - 0x598  :    0 - 0x0
    "00000000", -- 1433 - 0x599  :    0 - 0x0
    "11111100", -- 1434 - 0x59a  :  252 - 0xfc
    "11111110", -- 1435 - 0x59b  :  254 - 0xfe
    "11101110", -- 1436 - 0x59c  :  238 - 0xee
    "11101110", -- 1437 - 0x59d  :  238 - 0xee
    "11101110", -- 1438 - 0x59e  :  238 - 0xee
    "11101110", -- 1439 - 0x59f  :  238 - 0xee
    "11111111", -- 1440 - 0x5a0  :  255 - 0xff -- Sprite 0x5a
    "11111111", -- 1441 - 0x5a1  :  255 - 0xff
    "10000011", -- 1442 - 0x5a2  :  131 - 0x83
    "00000001", -- 1443 - 0x5a3  :    1 - 0x1
    "11101110", -- 1444 - 0x5a4  :  238 - 0xee
    "00000000", -- 1445 - 0x5a5  :    0 - 0x0
    "11101110", -- 1446 - 0x5a6  :  238 - 0xee
    "11101110", -- 1447 - 0x5a7  :  238 - 0xee
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "01111100", -- 1450 - 0x5aa  :  124 - 0x7c
    "11111110", -- 1451 - 0x5ab  :  254 - 0xfe
    "11101110", -- 1452 - 0x5ac  :  238 - 0xee
    "11101110", -- 1453 - 0x5ad  :  238 - 0xee
    "11101110", -- 1454 - 0x5ae  :  238 - 0xee
    "11101110", -- 1455 - 0x5af  :  238 - 0xee
    "11111111", -- 1456 - 0x5b0  :  255 - 0xff -- Sprite 0x5b
    "11111111", -- 1457 - 0x5b1  :  255 - 0xff
    "00000001", -- 1458 - 0x5b2  :    1 - 0x1
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "11100000", -- 1460 - 0x5b4  :  224 - 0xe0
    "00001111", -- 1461 - 0x5b5  :   15 - 0xf
    "11111111", -- 1462 - 0x5b6  :  255 - 0xff
    "11111011", -- 1463 - 0x5b7  :  251 - 0xfb
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "11111110", -- 1466 - 0x5ba  :  254 - 0xfe
    "11111110", -- 1467 - 0x5bb  :  254 - 0xfe
    "11100000", -- 1468 - 0x5bc  :  224 - 0xe0
    "11100000", -- 1469 - 0x5bd  :  224 - 0xe0
    "11111000", -- 1470 - 0x5be  :  248 - 0xf8
    "11111000", -- 1471 - 0x5bf  :  248 - 0xf8
    "11111111", -- 1472 - 0x5c0  :  255 - 0xff -- Sprite 0x5c
    "11111111", -- 1473 - 0x5c1  :  255 - 0xff
    "11111111", -- 1474 - 0x5c2  :  255 - 0xff
    "11111111", -- 1475 - 0x5c3  :  255 - 0xff
    "11111111", -- 1476 - 0x5c4  :  255 - 0xff
    "11111111", -- 1477 - 0x5c5  :  255 - 0xff
    "11111111", -- 1478 - 0x5c6  :  255 - 0xff
    "11011101", -- 1479 - 0x5c7  :  221 - 0xdd
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "00000000", -- 1482 - 0x5ca  :    0 - 0x0
    "00000000", -- 1483 - 0x5cb  :    0 - 0x0
    "00000000", -- 1484 - 0x5cc  :    0 - 0x0
    "00000000", -- 1485 - 0x5cd  :    0 - 0x0
    "11001100", -- 1486 - 0x5ce  :  204 - 0xcc
    "11001100", -- 1487 - 0x5cf  :  204 - 0xcc
    "11111111", -- 1488 - 0x5d0  :  255 - 0xff -- Sprite 0x5d
    "11111111", -- 1489 - 0x5d1  :  255 - 0xff
    "00000001", -- 1490 - 0x5d2  :    1 - 0x1
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "11100000", -- 1492 - 0x5d4  :  224 - 0xe0
    "00001111", -- 1493 - 0x5d5  :   15 - 0xf
    "11111111", -- 1494 - 0x5d6  :  255 - 0xff
    "11111011", -- 1495 - 0x5d7  :  251 - 0xfb
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "11111110", -- 1498 - 0x5da  :  254 - 0xfe
    "11111110", -- 1499 - 0x5db  :  254 - 0xfe
    "11100000", -- 1500 - 0x5dc  :  224 - 0xe0
    "11100000", -- 1501 - 0x5dd  :  224 - 0xe0
    "11111000", -- 1502 - 0x5de  :  248 - 0xf8
    "11111000", -- 1503 - 0x5df  :  248 - 0xf8
    "11111111", -- 1504 - 0x5e0  :  255 - 0xff -- Sprite 0x5e
    "11111111", -- 1505 - 0x5e1  :  255 - 0xff
    "00010001", -- 1506 - 0x5e2  :   17 - 0x11
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "11101110", -- 1508 - 0x5e4  :  238 - 0xee
    "00000000", -- 1509 - 0x5e5  :    0 - 0x0
    "11101110", -- 1510 - 0x5e6  :  238 - 0xee
    "11101110", -- 1511 - 0x5e7  :  238 - 0xee
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "11101110", -- 1514 - 0x5ea  :  238 - 0xee
    "11101110", -- 1515 - 0x5eb  :  238 - 0xee
    "11101110", -- 1516 - 0x5ec  :  238 - 0xee
    "11101110", -- 1517 - 0x5ed  :  238 - 0xee
    "11101110", -- 1518 - 0x5ee  :  238 - 0xee
    "11101110", -- 1519 - 0x5ef  :  238 - 0xee
    "10111101", -- 1520 - 0x5f0  :  189 - 0xbd -- Sprite 0x5f
    "11111111", -- 1521 - 0x5f1  :  255 - 0xff
    "11111111", -- 1522 - 0x5f2  :  255 - 0xff
    "11111111", -- 1523 - 0x5f3  :  255 - 0xff
    "11111111", -- 1524 - 0x5f4  :  255 - 0xff
    "11111111", -- 1525 - 0x5f5  :  255 - 0xff
    "11111111", -- 1526 - 0x5f6  :  255 - 0xff
    "11111111", -- 1527 - 0x5f7  :  255 - 0xff
    "01111110", -- 1528 - 0x5f8  :  126 - 0x7e
    "01111110", -- 1529 - 0x5f9  :  126 - 0x7e
    "01111110", -- 1530 - 0x5fa  :  126 - 0x7e
    "01111110", -- 1531 - 0x5fb  :  126 - 0x7e
    "01111110", -- 1532 - 0x5fc  :  126 - 0x7e
    "01111110", -- 1533 - 0x5fd  :  126 - 0x7e
    "01111110", -- 1534 - 0x5fe  :  126 - 0x7e
    "01111110", -- 1535 - 0x5ff  :  126 - 0x7e
    "11101110", -- 1536 - 0x600  :  238 - 0xee -- Sprite 0x60
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "11111110", -- 1538 - 0x602  :  254 - 0xfe
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000001", -- 1540 - 0x604  :    1 - 0x1
    "00001111", -- 1541 - 0x605  :   15 - 0xf
    "10001111", -- 1542 - 0x606  :  143 - 0x8f
    "11111111", -- 1543 - 0x607  :  255 - 0xff
    "11101110", -- 1544 - 0x608  :  238 - 0xee
    "11101110", -- 1545 - 0x609  :  238 - 0xee
    "11111110", -- 1546 - 0x60a  :  254 - 0xfe
    "11111100", -- 1547 - 0x60b  :  252 - 0xfc
    "11100000", -- 1548 - 0x60c  :  224 - 0xe0
    "11100000", -- 1549 - 0x60d  :  224 - 0xe0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "11101110", -- 1552 - 0x610  :  238 - 0xee -- Sprite 0x61
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "11111100", -- 1554 - 0x612  :  252 - 0xfc
    "00000001", -- 1555 - 0x613  :    1 - 0x1
    "00000001", -- 1556 - 0x614  :    1 - 0x1
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "10001000", -- 1558 - 0x616  :  136 - 0x88
    "11111111", -- 1559 - 0x617  :  255 - 0xff
    "11101110", -- 1560 - 0x618  :  238 - 0xee
    "11101110", -- 1561 - 0x619  :  238 - 0xee
    "11111100", -- 1562 - 0x61a  :  252 - 0xfc
    "11111100", -- 1563 - 0x61b  :  252 - 0xfc
    "11101110", -- 1564 - 0x61c  :  238 - 0xee
    "11101110", -- 1565 - 0x61d  :  238 - 0xee
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "11100011", -- 1568 - 0x620  :  227 - 0xe3 -- Sprite 0x62
    "00001111", -- 1569 - 0x621  :   15 - 0xf
    "11101111", -- 1570 - 0x622  :  239 - 0xef
    "00001111", -- 1571 - 0x623  :   15 - 0xf
    "00000001", -- 1572 - 0x624  :    1 - 0x1
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "10000000", -- 1574 - 0x626  :  128 - 0x80
    "11111111", -- 1575 - 0x627  :  255 - 0xff
    "11100000", -- 1576 - 0x628  :  224 - 0xe0
    "11100000", -- 1577 - 0x629  :  224 - 0xe0
    "11100000", -- 1578 - 0x62a  :  224 - 0xe0
    "11100000", -- 1579 - 0x62b  :  224 - 0xe0
    "11111110", -- 1580 - 0x62c  :  254 - 0xfe
    "11111110", -- 1581 - 0x62d  :  254 - 0xfe
    "00000000", -- 1582 - 0x62e  :    0 - 0x0
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "11001110", -- 1584 - 0x630  :  206 - 0xce -- Sprite 0x63
    "11110000", -- 1585 - 0x631  :  240 - 0xf0
    "11111110", -- 1586 - 0x632  :  254 - 0xfe
    "00010000", -- 1587 - 0x633  :   16 - 0x10
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "10000000", -- 1589 - 0x635  :  128 - 0x80
    "11000001", -- 1590 - 0x636  :  193 - 0xc1
    "11111111", -- 1591 - 0x637  :  255 - 0xff
    "00001110", -- 1592 - 0x638  :   14 - 0xe
    "00001110", -- 1593 - 0x639  :   14 - 0xe
    "00001110", -- 1594 - 0x63a  :   14 - 0xe
    "11101110", -- 1595 - 0x63b  :  238 - 0xee
    "11111110", -- 1596 - 0x63c  :  254 - 0xfe
    "01111100", -- 1597 - 0x63d  :  124 - 0x7c
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "11111011", -- 1600 - 0x640  :  251 - 0xfb -- Sprite 0x64
    "11000011", -- 1601 - 0x641  :  195 - 0xc3
    "11111011", -- 1602 - 0x642  :  251 - 0xfb
    "11000011", -- 1603 - 0x643  :  195 - 0xc3
    "11000011", -- 1604 - 0x644  :  195 - 0xc3
    "11000011", -- 1605 - 0x645  :  195 - 0xc3
    "11100011", -- 1606 - 0x646  :  227 - 0xe3
    "11111111", -- 1607 - 0x647  :  255 - 0xff
    "00111000", -- 1608 - 0x648  :   56 - 0x38
    "00111000", -- 1609 - 0x649  :   56 - 0x38
    "00111000", -- 1610 - 0x64a  :   56 - 0x38
    "00111000", -- 1611 - 0x64b  :   56 - 0x38
    "00111000", -- 1612 - 0x64c  :   56 - 0x38
    "00111000", -- 1613 - 0x64d  :   56 - 0x38
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "11101110", -- 1616 - 0x650  :  238 - 0xee -- Sprite 0x65
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "11111110", -- 1618 - 0x652  :  254 - 0xfe
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "10001000", -- 1622 - 0x656  :  136 - 0x88
    "11111111", -- 1623 - 0x657  :  255 - 0xff
    "11101110", -- 1624 - 0x658  :  238 - 0xee
    "11101110", -- 1625 - 0x659  :  238 - 0xee
    "11111110", -- 1626 - 0x65a  :  254 - 0xfe
    "11111110", -- 1627 - 0x65b  :  254 - 0xfe
    "11101110", -- 1628 - 0x65c  :  238 - 0xee
    "11101110", -- 1629 - 0x65d  :  238 - 0xee
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "11101111", -- 1632 - 0x660  :  239 - 0xef -- Sprite 0x66
    "00001111", -- 1633 - 0x661  :   15 - 0xf
    "11101111", -- 1634 - 0x662  :  239 - 0xef
    "00000001", -- 1635 - 0x663  :    1 - 0x1
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "10000000", -- 1638 - 0x666  :  128 - 0x80
    "11111111", -- 1639 - 0x667  :  255 - 0xff
    "11100000", -- 1640 - 0x668  :  224 - 0xe0
    "11100000", -- 1641 - 0x669  :  224 - 0xe0
    "11100000", -- 1642 - 0x66a  :  224 - 0xe0
    "11101110", -- 1643 - 0x66b  :  238 - 0xee
    "11111110", -- 1644 - 0x66c  :  254 - 0xfe
    "11111110", -- 1645 - 0x66d  :  254 - 0xfe
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "11101110", -- 1648 - 0x670  :  238 - 0xee -- Sprite 0x67
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "11111110", -- 1650 - 0x672  :  254 - 0xfe
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00001000", -- 1653 - 0x675  :    8 - 0x8
    "10011100", -- 1654 - 0x676  :  156 - 0x9c
    "11111111", -- 1655 - 0x677  :  255 - 0xff
    "11101110", -- 1656 - 0x678  :  238 - 0xee
    "11101110", -- 1657 - 0x679  :  238 - 0xee
    "11111110", -- 1658 - 0x67a  :  254 - 0xfe
    "11111110", -- 1659 - 0x67b  :  254 - 0xfe
    "11101110", -- 1660 - 0x67c  :  238 - 0xee
    "11000110", -- 1661 - 0x67d  :  198 - 0xc6
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "11101110", -- 1664 - 0x680  :  238 - 0xee -- Sprite 0x68
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "11101110", -- 1666 - 0x682  :  238 - 0xee
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "10001000", -- 1670 - 0x686  :  136 - 0x88
    "11111111", -- 1671 - 0x687  :  255 - 0xff
    "11101110", -- 1672 - 0x688  :  238 - 0xee
    "11101110", -- 1673 - 0x689  :  238 - 0xee
    "11101110", -- 1674 - 0x68a  :  238 - 0xee
    "11101110", -- 1675 - 0x68b  :  238 - 0xee
    "11101110", -- 1676 - 0x68c  :  238 - 0xee
    "11101110", -- 1677 - 0x68d  :  238 - 0xee
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "11101110", -- 1680 - 0x690  :  238 - 0xee -- Sprite 0x69
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "11101110", -- 1682 - 0x692  :  238 - 0xee
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00000000", -- 1685 - 0x695  :    0 - 0x0
    "10000001", -- 1686 - 0x696  :  129 - 0x81
    "11111111", -- 1687 - 0x697  :  255 - 0xff
    "11101110", -- 1688 - 0x698  :  238 - 0xee
    "11101110", -- 1689 - 0x699  :  238 - 0xee
    "11101110", -- 1690 - 0x69a  :  238 - 0xee
    "11101110", -- 1691 - 0x69b  :  238 - 0xee
    "11111110", -- 1692 - 0x69c  :  254 - 0xfe
    "11111100", -- 1693 - 0x69d  :  252 - 0xfc
    "00000000", -- 1694 - 0x69e  :    0 - 0x0
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "11101110", -- 1696 - 0x6a0  :  238 - 0xee -- Sprite 0x6a
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "11101110", -- 1698 - 0x6a2  :  238 - 0xee
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "10000000", -- 1701 - 0x6a5  :  128 - 0x80
    "11000001", -- 1702 - 0x6a6  :  193 - 0xc1
    "11111111", -- 1703 - 0x6a7  :  255 - 0xff
    "11101110", -- 1704 - 0x6a8  :  238 - 0xee
    "11101110", -- 1705 - 0x6a9  :  238 - 0xee
    "11101110", -- 1706 - 0x6aa  :  238 - 0xee
    "11101110", -- 1707 - 0x6ab  :  238 - 0xee
    "11111110", -- 1708 - 0x6ac  :  254 - 0xfe
    "01111100", -- 1709 - 0x6ad  :  124 - 0x7c
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "11100011", -- 1712 - 0x6b0  :  227 - 0xe3 -- Sprite 0x6b
    "00001111", -- 1713 - 0x6b1  :   15 - 0xf
    "11101111", -- 1714 - 0x6b2  :  239 - 0xef
    "00001111", -- 1715 - 0x6b3  :   15 - 0xf
    "00000001", -- 1716 - 0x6b4  :    1 - 0x1
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "10000000", -- 1718 - 0x6b6  :  128 - 0x80
    "11111111", -- 1719 - 0x6b7  :  255 - 0xff
    "11100000", -- 1720 - 0x6b8  :  224 - 0xe0
    "11100000", -- 1721 - 0x6b9  :  224 - 0xe0
    "11100000", -- 1722 - 0x6ba  :  224 - 0xe0
    "11100000", -- 1723 - 0x6bb  :  224 - 0xe0
    "11111110", -- 1724 - 0x6bc  :  254 - 0xfe
    "11111110", -- 1725 - 0x6bd  :  254 - 0xfe
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "10011001", -- 1728 - 0x6c0  :  153 - 0x99 -- Sprite 0x6c
    "11100011", -- 1729 - 0x6c1  :  227 - 0xe3
    "11110011", -- 1730 - 0x6c2  :  243 - 0xf3
    "11000111", -- 1731 - 0x6c3  :  199 - 0xc7
    "10000001", -- 1732 - 0x6c4  :  129 - 0x81
    "10001000", -- 1733 - 0x6c5  :  136 - 0x88
    "11001100", -- 1734 - 0x6c6  :  204 - 0xcc
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "00011000", -- 1736 - 0x6c8  :   24 - 0x18
    "00011000", -- 1737 - 0x6c9  :   24 - 0x18
    "00110000", -- 1738 - 0x6ca  :   48 - 0x30
    "00110000", -- 1739 - 0x6cb  :   48 - 0x30
    "01100110", -- 1740 - 0x6cc  :  102 - 0x66
    "01100110", -- 1741 - 0x6cd  :  102 - 0x66
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "11100011", -- 1744 - 0x6d0  :  227 - 0xe3 -- Sprite 0x6d
    "00001111", -- 1745 - 0x6d1  :   15 - 0xf
    "11101111", -- 1746 - 0x6d2  :  239 - 0xef
    "00001111", -- 1747 - 0x6d3  :   15 - 0xf
    "00001111", -- 1748 - 0x6d4  :   15 - 0xf
    "00001111", -- 1749 - 0x6d5  :   15 - 0xf
    "10001111", -- 1750 - 0x6d6  :  143 - 0x8f
    "11111111", -- 1751 - 0x6d7  :  255 - 0xff
    "11100000", -- 1752 - 0x6d8  :  224 - 0xe0
    "11100000", -- 1753 - 0x6d9  :  224 - 0xe0
    "11100000", -- 1754 - 0x6da  :  224 - 0xe0
    "11100000", -- 1755 - 0x6db  :  224 - 0xe0
    "11100000", -- 1756 - 0x6dc  :  224 - 0xe0
    "11100000", -- 1757 - 0x6dd  :  224 - 0xe0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "11101110", -- 1760 - 0x6e0  :  238 - 0xee -- Sprite 0x6e
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "11101110", -- 1762 - 0x6e2  :  238 - 0xee
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "10000000", -- 1765 - 0x6e5  :  128 - 0x80
    "11000001", -- 1766 - 0x6e6  :  193 - 0xc1
    "11111111", -- 1767 - 0x6e7  :  255 - 0xff
    "11101110", -- 1768 - 0x6e8  :  238 - 0xee
    "11101110", -- 1769 - 0x6e9  :  238 - 0xee
    "11101110", -- 1770 - 0x6ea  :  238 - 0xee
    "11101110", -- 1771 - 0x6eb  :  238 - 0xee
    "11111110", -- 1772 - 0x6ec  :  254 - 0xfe
    "01111100", -- 1773 - 0x6ed  :  124 - 0x7c
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "11111111", -- 1776 - 0x6f0  :  255 - 0xff -- Sprite 0x6f
    "11111111", -- 1777 - 0x6f1  :  255 - 0xff
    "11111111", -- 1778 - 0x6f2  :  255 - 0xff
    "10111101", -- 1779 - 0x6f3  :  189 - 0xbd
    "11111111", -- 1780 - 0x6f4  :  255 - 0xff
    "11011011", -- 1781 - 0x6f5  :  219 - 0xdb
    "11111111", -- 1782 - 0x6f6  :  255 - 0xff
    "11111111", -- 1783 - 0x6f7  :  255 - 0xff
    "01111110", -- 1784 - 0x6f8  :  126 - 0x7e
    "01111110", -- 1785 - 0x6f9  :  126 - 0x7e
    "01111110", -- 1786 - 0x6fa  :  126 - 0x7e
    "01111110", -- 1787 - 0x6fb  :  126 - 0x7e
    "00111100", -- 1788 - 0x6fc  :   60 - 0x3c
    "00111100", -- 1789 - 0x6fd  :   60 - 0x3c
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "11111011", -- 1792 - 0x700  :  251 - 0xfb -- Sprite 0x70
    "11101111", -- 1793 - 0x701  :  239 - 0xef
    "11011111", -- 1794 - 0x702  :  223 - 0xdf
    "11111111", -- 1795 - 0x703  :  255 - 0xff
    "10111111", -- 1796 - 0x704  :  191 - 0xbf
    "10111111", -- 1797 - 0x705  :  191 - 0xbf
    "11111110", -- 1798 - 0x706  :  254 - 0xfe
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "00000111", -- 1800 - 0x708  :    7 - 0x7
    "00011111", -- 1801 - 0x709  :   31 - 0x1f
    "00111111", -- 1802 - 0x70a  :   63 - 0x3f
    "00111111", -- 1803 - 0x70b  :   63 - 0x3f
    "01111111", -- 1804 - 0x70c  :  127 - 0x7f
    "01111111", -- 1805 - 0x70d  :  127 - 0x7f
    "01111111", -- 1806 - 0x70e  :  127 - 0x7f
    "01111110", -- 1807 - 0x70f  :  126 - 0x7e
    "11011111", -- 1808 - 0x710  :  223 - 0xdf -- Sprite 0x71
    "11110111", -- 1809 - 0x711  :  247 - 0xf7
    "11111011", -- 1810 - 0x712  :  251 - 0xfb
    "11111111", -- 1811 - 0x713  :  255 - 0xff
    "11111101", -- 1812 - 0x714  :  253 - 0xfd
    "11111101", -- 1813 - 0x715  :  253 - 0xfd
    "01111111", -- 1814 - 0x716  :  127 - 0x7f
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "11100000", -- 1816 - 0x718  :  224 - 0xe0
    "11111000", -- 1817 - 0x719  :  248 - 0xf8
    "11111100", -- 1818 - 0x71a  :  252 - 0xfc
    "11111100", -- 1819 - 0x71b  :  252 - 0xfc
    "11111110", -- 1820 - 0x71c  :  254 - 0xfe
    "11111110", -- 1821 - 0x71d  :  254 - 0xfe
    "11111110", -- 1822 - 0x71e  :  254 - 0xfe
    "01111110", -- 1823 - 0x71f  :  126 - 0x7e
    "11111111", -- 1824 - 0x720  :  255 - 0xff -- Sprite 0x72
    "11111111", -- 1825 - 0x721  :  255 - 0xff
    "11111111", -- 1826 - 0x722  :  255 - 0xff
    "11111111", -- 1827 - 0x723  :  255 - 0xff
    "11111111", -- 1828 - 0x724  :  255 - 0xff
    "11111111", -- 1829 - 0x725  :  255 - 0xff
    "11111111", -- 1830 - 0x726  :  255 - 0xff
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "01111110", -- 1832 - 0x728  :  126 - 0x7e
    "01111110", -- 1833 - 0x729  :  126 - 0x7e
    "01111110", -- 1834 - 0x72a  :  126 - 0x7e
    "01111110", -- 1835 - 0x72b  :  126 - 0x7e
    "01111110", -- 1836 - 0x72c  :  126 - 0x7e
    "01111110", -- 1837 - 0x72d  :  126 - 0x7e
    "01111110", -- 1838 - 0x72e  :  126 - 0x7e
    "01111110", -- 1839 - 0x72f  :  126 - 0x7e
    "11111111", -- 1840 - 0x730  :  255 - 0xff -- Sprite 0x73
    "11111110", -- 1841 - 0x731  :  254 - 0xfe
    "10111111", -- 1842 - 0x732  :  191 - 0xbf
    "10111111", -- 1843 - 0x733  :  191 - 0xbf
    "11111111", -- 1844 - 0x734  :  255 - 0xff
    "11011111", -- 1845 - 0x735  :  223 - 0xdf
    "11101111", -- 1846 - 0x736  :  239 - 0xef
    "11111011", -- 1847 - 0x737  :  251 - 0xfb
    "01111110", -- 1848 - 0x738  :  126 - 0x7e
    "01111111", -- 1849 - 0x739  :  127 - 0x7f
    "01111111", -- 1850 - 0x73a  :  127 - 0x7f
    "01111111", -- 1851 - 0x73b  :  127 - 0x7f
    "00111111", -- 1852 - 0x73c  :   63 - 0x3f
    "00111111", -- 1853 - 0x73d  :   63 - 0x3f
    "00011111", -- 1854 - 0x73e  :   31 - 0x1f
    "00000111", -- 1855 - 0x73f  :    7 - 0x7
    "11111111", -- 1856 - 0x740  :  255 - 0xff -- Sprite 0x74
    "01111111", -- 1857 - 0x741  :  127 - 0x7f
    "11111101", -- 1858 - 0x742  :  253 - 0xfd
    "11111101", -- 1859 - 0x743  :  253 - 0xfd
    "11111111", -- 1860 - 0x744  :  255 - 0xff
    "11111011", -- 1861 - 0x745  :  251 - 0xfb
    "11110111", -- 1862 - 0x746  :  247 - 0xf7
    "11011111", -- 1863 - 0x747  :  223 - 0xdf
    "01111110", -- 1864 - 0x748  :  126 - 0x7e
    "11111110", -- 1865 - 0x749  :  254 - 0xfe
    "11111110", -- 1866 - 0x74a  :  254 - 0xfe
    "11111110", -- 1867 - 0x74b  :  254 - 0xfe
    "11111100", -- 1868 - 0x74c  :  252 - 0xfc
    "11111100", -- 1869 - 0x74d  :  252 - 0xfc
    "11111000", -- 1870 - 0x74e  :  248 - 0xf8
    "11100000", -- 1871 - 0x74f  :  224 - 0xe0
    "11111111", -- 1872 - 0x750  :  255 - 0xff -- Sprite 0x75
    "11111111", -- 1873 - 0x751  :  255 - 0xff
    "11111111", -- 1874 - 0x752  :  255 - 0xff
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "11111111", -- 1876 - 0x754  :  255 - 0xff
    "11111111", -- 1877 - 0x755  :  255 - 0xff
    "11111111", -- 1878 - 0x756  :  255 - 0xff
    "11111111", -- 1879 - 0x757  :  255 - 0xff
    "01111111", -- 1880 - 0x758  :  127 - 0x7f
    "01111111", -- 1881 - 0x759  :  127 - 0x7f
    "01111111", -- 1882 - 0x75a  :  127 - 0x7f
    "01111111", -- 1883 - 0x75b  :  127 - 0x7f
    "01111111", -- 1884 - 0x75c  :  127 - 0x7f
    "01111111", -- 1885 - 0x75d  :  127 - 0x7f
    "00000111", -- 1886 - 0x75e  :    7 - 0x7
    "00000111", -- 1887 - 0x75f  :    7 - 0x7
    "11111111", -- 1888 - 0x760  :  255 - 0xff -- Sprite 0x76
    "11111111", -- 1889 - 0x761  :  255 - 0xff
    "11111111", -- 1890 - 0x762  :  255 - 0xff
    "11111111", -- 1891 - 0x763  :  255 - 0xff
    "11111111", -- 1892 - 0x764  :  255 - 0xff
    "11111111", -- 1893 - 0x765  :  255 - 0xff
    "11111111", -- 1894 - 0x766  :  255 - 0xff
    "11111111", -- 1895 - 0x767  :  255 - 0xff
    "11111110", -- 1896 - 0x768  :  254 - 0xfe
    "11111110", -- 1897 - 0x769  :  254 - 0xfe
    "11111110", -- 1898 - 0x76a  :  254 - 0xfe
    "11111110", -- 1899 - 0x76b  :  254 - 0xfe
    "11111110", -- 1900 - 0x76c  :  254 - 0xfe
    "11111110", -- 1901 - 0x76d  :  254 - 0xfe
    "11100000", -- 1902 - 0x76e  :  224 - 0xe0
    "11100000", -- 1903 - 0x76f  :  224 - 0xe0
    "11111111", -- 1904 - 0x770  :  255 - 0xff -- Sprite 0x77
    "11111111", -- 1905 - 0x771  :  255 - 0xff
    "11111111", -- 1906 - 0x772  :  255 - 0xff
    "11111111", -- 1907 - 0x773  :  255 - 0xff
    "11111111", -- 1908 - 0x774  :  255 - 0xff
    "11111111", -- 1909 - 0x775  :  255 - 0xff
    "11111111", -- 1910 - 0x776  :  255 - 0xff
    "11111111", -- 1911 - 0x777  :  255 - 0xff
    "00000111", -- 1912 - 0x778  :    7 - 0x7
    "00000111", -- 1913 - 0x779  :    7 - 0x7
    "00000111", -- 1914 - 0x77a  :    7 - 0x7
    "00000111", -- 1915 - 0x77b  :    7 - 0x7
    "00000111", -- 1916 - 0x77c  :    7 - 0x7
    "00000111", -- 1917 - 0x77d  :    7 - 0x7
    "00000111", -- 1918 - 0x77e  :    7 - 0x7
    "00000111", -- 1919 - 0x77f  :    7 - 0x7
    "11111111", -- 1920 - 0x780  :  255 - 0xff -- Sprite 0x78
    "11111111", -- 1921 - 0x781  :  255 - 0xff
    "11111111", -- 1922 - 0x782  :  255 - 0xff
    "11111111", -- 1923 - 0x783  :  255 - 0xff
    "11111111", -- 1924 - 0x784  :  255 - 0xff
    "11111111", -- 1925 - 0x785  :  255 - 0xff
    "11111111", -- 1926 - 0x786  :  255 - 0xff
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11100000", -- 1928 - 0x788  :  224 - 0xe0
    "11100000", -- 1929 - 0x789  :  224 - 0xe0
    "11100000", -- 1930 - 0x78a  :  224 - 0xe0
    "11100000", -- 1931 - 0x78b  :  224 - 0xe0
    "11100000", -- 1932 - 0x78c  :  224 - 0xe0
    "11100000", -- 1933 - 0x78d  :  224 - 0xe0
    "11100000", -- 1934 - 0x78e  :  224 - 0xe0
    "11100000", -- 1935 - 0x78f  :  224 - 0xe0
    "11111111", -- 1936 - 0x790  :  255 - 0xff -- Sprite 0x79
    "11111111", -- 1937 - 0x791  :  255 - 0xff
    "11111111", -- 1938 - 0x792  :  255 - 0xff
    "11111111", -- 1939 - 0x793  :  255 - 0xff
    "11111111", -- 1940 - 0x794  :  255 - 0xff
    "11111111", -- 1941 - 0x795  :  255 - 0xff
    "11111111", -- 1942 - 0x796  :  255 - 0xff
    "11111111", -- 1943 - 0x797  :  255 - 0xff
    "01111111", -- 1944 - 0x798  :  127 - 0x7f
    "01111111", -- 1945 - 0x799  :  127 - 0x7f
    "01111111", -- 1946 - 0x79a  :  127 - 0x7f
    "01111111", -- 1947 - 0x79b  :  127 - 0x7f
    "01111111", -- 1948 - 0x79c  :  127 - 0x7f
    "01111111", -- 1949 - 0x79d  :  127 - 0x7f
    "01111110", -- 1950 - 0x79e  :  126 - 0x7e
    "01111110", -- 1951 - 0x79f  :  126 - 0x7e
    "11111111", -- 1952 - 0x7a0  :  255 - 0xff -- Sprite 0x7a
    "11111111", -- 1953 - 0x7a1  :  255 - 0xff
    "11111111", -- 1954 - 0x7a2  :  255 - 0xff
    "11111111", -- 1955 - 0x7a3  :  255 - 0xff
    "11111111", -- 1956 - 0x7a4  :  255 - 0xff
    "11111111", -- 1957 - 0x7a5  :  255 - 0xff
    "11111111", -- 1958 - 0x7a6  :  255 - 0xff
    "11111111", -- 1959 - 0x7a7  :  255 - 0xff
    "11111110", -- 1960 - 0x7a8  :  254 - 0xfe
    "11111110", -- 1961 - 0x7a9  :  254 - 0xfe
    "11111110", -- 1962 - 0x7aa  :  254 - 0xfe
    "11111110", -- 1963 - 0x7ab  :  254 - 0xfe
    "11111110", -- 1964 - 0x7ac  :  254 - 0xfe
    "11111110", -- 1965 - 0x7ad  :  254 - 0xfe
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "11111111", -- 1968 - 0x7b0  :  255 - 0xff -- Sprite 0x7b
    "11111111", -- 1969 - 0x7b1  :  255 - 0xff
    "11111111", -- 1970 - 0x7b2  :  255 - 0xff
    "11111111", -- 1971 - 0x7b3  :  255 - 0xff
    "11111111", -- 1972 - 0x7b4  :  255 - 0xff
    "11111111", -- 1973 - 0x7b5  :  255 - 0xff
    "11111111", -- 1974 - 0x7b6  :  255 - 0xff
    "11111111", -- 1975 - 0x7b7  :  255 - 0xff
    "01111110", -- 1976 - 0x7b8  :  126 - 0x7e
    "01111111", -- 1977 - 0x7b9  :  127 - 0x7f
    "01111111", -- 1978 - 0x7ba  :  127 - 0x7f
    "01111111", -- 1979 - 0x7bb  :  127 - 0x7f
    "01111111", -- 1980 - 0x7bc  :  127 - 0x7f
    "01111111", -- 1981 - 0x7bd  :  127 - 0x7f
    "01111111", -- 1982 - 0x7be  :  127 - 0x7f
    "01111110", -- 1983 - 0x7bf  :  126 - 0x7e
    "11111111", -- 1984 - 0x7c0  :  255 - 0xff -- Sprite 0x7c
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "11111111", -- 1986 - 0x7c2  :  255 - 0xff
    "11111111", -- 1987 - 0x7c3  :  255 - 0xff
    "11111111", -- 1988 - 0x7c4  :  255 - 0xff
    "11111111", -- 1989 - 0x7c5  :  255 - 0xff
    "11111111", -- 1990 - 0x7c6  :  255 - 0xff
    "11111111", -- 1991 - 0x7c7  :  255 - 0xff
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0
    "11110000", -- 1993 - 0x7c9  :  240 - 0xf0
    "11110000", -- 1994 - 0x7ca  :  240 - 0xf0
    "11110000", -- 1995 - 0x7cb  :  240 - 0xf0
    "11110000", -- 1996 - 0x7cc  :  240 - 0xf0
    "11110000", -- 1997 - 0x7cd  :  240 - 0xf0
    "11110000", -- 1998 - 0x7ce  :  240 - 0xf0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "11111111", -- 2000 - 0x7d0  :  255 - 0xff -- Sprite 0x7d
    "11111111", -- 2001 - 0x7d1  :  255 - 0xff
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "11111111", -- 2004 - 0x7d4  :  255 - 0xff
    "11111111", -- 2005 - 0x7d5  :  255 - 0xff
    "11111111", -- 2006 - 0x7d6  :  255 - 0xff
    "11111111", -- 2007 - 0x7d7  :  255 - 0xff
    "01111110", -- 2008 - 0x7d8  :  126 - 0x7e
    "01111110", -- 2009 - 0x7d9  :  126 - 0x7e
    "01111111", -- 2010 - 0x7da  :  127 - 0x7f
    "01111111", -- 2011 - 0x7db  :  127 - 0x7f
    "01111111", -- 2012 - 0x7dc  :  127 - 0x7f
    "01111111", -- 2013 - 0x7dd  :  127 - 0x7f
    "01111111", -- 2014 - 0x7de  :  127 - 0x7f
    "01111111", -- 2015 - 0x7df  :  127 - 0x7f
    "11111111", -- 2016 - 0x7e0  :  255 - 0xff -- Sprite 0x7e
    "11111111", -- 2017 - 0x7e1  :  255 - 0xff
    "11111111", -- 2018 - 0x7e2  :  255 - 0xff
    "11111111", -- 2019 - 0x7e3  :  255 - 0xff
    "11111111", -- 2020 - 0x7e4  :  255 - 0xff
    "11111111", -- 2021 - 0x7e5  :  255 - 0xff
    "11111111", -- 2022 - 0x7e6  :  255 - 0xff
    "11111111", -- 2023 - 0x7e7  :  255 - 0xff
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "11111110", -- 2026 - 0x7ea  :  254 - 0xfe
    "11111110", -- 2027 - 0x7eb  :  254 - 0xfe
    "11111110", -- 2028 - 0x7ec  :  254 - 0xfe
    "11111110", -- 2029 - 0x7ed  :  254 - 0xfe
    "11111110", -- 2030 - 0x7ee  :  254 - 0xfe
    "11111110", -- 2031 - 0x7ef  :  254 - 0xfe
    "11111111", -- 2032 - 0x7f0  :  255 - 0xff -- Sprite 0x7f
    "11111111", -- 2033 - 0x7f1  :  255 - 0xff
    "11111111", -- 2034 - 0x7f2  :  255 - 0xff
    "11111111", -- 2035 - 0x7f3  :  255 - 0xff
    "11111111", -- 2036 - 0x7f4  :  255 - 0xff
    "11111111", -- 2037 - 0x7f5  :  255 - 0xff
    "11111111", -- 2038 - 0x7f6  :  255 - 0xff
    "11111111", -- 2039 - 0x7f7  :  255 - 0xff
    "01111110", -- 2040 - 0x7f8  :  126 - 0x7e
    "11111110", -- 2041 - 0x7f9  :  254 - 0xfe
    "11111110", -- 2042 - 0x7fa  :  254 - 0xfe
    "11111110", -- 2043 - 0x7fb  :  254 - 0xfe
    "11111110", -- 2044 - 0x7fc  :  254 - 0xfe
    "11111110", -- 2045 - 0x7fd  :  254 - 0xfe
    "11111110", -- 2046 - 0x7fe  :  254 - 0xfe
    "01111110", -- 2047 - 0x7ff  :  126 - 0x7e
    "10111111", -- 2048 - 0x800  :  191 - 0xbf -- Sprite 0x80
    "11110111", -- 2049 - 0x801  :  247 - 0xf7
    "11111101", -- 2050 - 0x802  :  253 - 0xfd
    "11011111", -- 2051 - 0x803  :  223 - 0xdf
    "11111011", -- 2052 - 0x804  :  251 - 0xfb
    "10111111", -- 2053 - 0x805  :  191 - 0xbf
    "11111110", -- 2054 - 0x806  :  254 - 0xfe
    "11101111", -- 2055 - 0x807  :  239 - 0xef
    "01000000", -- 2056 - 0x808  :   64 - 0x40
    "00001000", -- 2057 - 0x809  :    8 - 0x8
    "00000010", -- 2058 - 0x80a  :    2 - 0x2
    "00100000", -- 2059 - 0x80b  :   32 - 0x20
    "00000100", -- 2060 - 0x80c  :    4 - 0x4
    "01000000", -- 2061 - 0x80d  :   64 - 0x40
    "00000001", -- 2062 - 0x80e  :    1 - 0x1
    "00010000", -- 2063 - 0x80f  :   16 - 0x10
    "11111111", -- 2064 - 0x810  :  255 - 0xff -- Sprite 0x81
    "11101110", -- 2065 - 0x811  :  238 - 0xee
    "11111111", -- 2066 - 0x812  :  255 - 0xff
    "11011111", -- 2067 - 0x813  :  223 - 0xdf
    "01110111", -- 2068 - 0x814  :  119 - 0x77
    "11111101", -- 2069 - 0x815  :  253 - 0xfd
    "11011111", -- 2070 - 0x816  :  223 - 0xdf
    "10111111", -- 2071 - 0x817  :  191 - 0xbf
    "00000000", -- 2072 - 0x818  :    0 - 0x0
    "00010001", -- 2073 - 0x819  :   17 - 0x11
    "00000000", -- 2074 - 0x81a  :    0 - 0x0
    "00100000", -- 2075 - 0x81b  :   32 - 0x20
    "10001000", -- 2076 - 0x81c  :  136 - 0x88
    "00000010", -- 2077 - 0x81d  :    2 - 0x2
    "00100000", -- 2078 - 0x81e  :   32 - 0x20
    "01000000", -- 2079 - 0x81f  :   64 - 0x40
    "11111110", -- 2080 - 0x820  :  254 - 0xfe -- Sprite 0x82
    "11101111", -- 2081 - 0x821  :  239 - 0xef
    "10111111", -- 2082 - 0x822  :  191 - 0xbf
    "11110111", -- 2083 - 0x823  :  247 - 0xf7
    "11111101", -- 2084 - 0x824  :  253 - 0xfd
    "11011111", -- 2085 - 0x825  :  223 - 0xdf
    "11111011", -- 2086 - 0x826  :  251 - 0xfb
    "10111111", -- 2087 - 0x827  :  191 - 0xbf
    "00000001", -- 2088 - 0x828  :    1 - 0x1
    "00010000", -- 2089 - 0x829  :   16 - 0x10
    "01000000", -- 2090 - 0x82a  :   64 - 0x40
    "00001000", -- 2091 - 0x82b  :    8 - 0x8
    "00000010", -- 2092 - 0x82c  :    2 - 0x2
    "00100000", -- 2093 - 0x82d  :   32 - 0x20
    "00000100", -- 2094 - 0x82e  :    4 - 0x4
    "01000000", -- 2095 - 0x82f  :   64 - 0x40
    "11101111", -- 2096 - 0x830  :  239 - 0xef -- Sprite 0x83
    "11111111", -- 2097 - 0x831  :  255 - 0xff
    "10111011", -- 2098 - 0x832  :  187 - 0xbb
    "11111111", -- 2099 - 0x833  :  255 - 0xff
    "11110111", -- 2100 - 0x834  :  247 - 0xf7
    "11011101", -- 2101 - 0x835  :  221 - 0xdd
    "01111111", -- 2102 - 0x836  :  127 - 0x7f
    "11110111", -- 2103 - 0x837  :  247 - 0xf7
    "00010000", -- 2104 - 0x838  :   16 - 0x10
    "00000000", -- 2105 - 0x839  :    0 - 0x0
    "01000100", -- 2106 - 0x83a  :   68 - 0x44
    "00000000", -- 2107 - 0x83b  :    0 - 0x0
    "00001000", -- 2108 - 0x83c  :    8 - 0x8
    "00100010", -- 2109 - 0x83d  :   34 - 0x22
    "10000000", -- 2110 - 0x83e  :  128 - 0x80
    "00001000", -- 2111 - 0x83f  :    8 - 0x8
    "11111111", -- 2112 - 0x840  :  255 - 0xff -- Sprite 0x84
    "11101110", -- 2113 - 0x841  :  238 - 0xee
    "11111011", -- 2114 - 0x842  :  251 - 0xfb
    "10111111", -- 2115 - 0x843  :  191 - 0xbf
    "01111111", -- 2116 - 0x844  :  127 - 0x7f
    "11101101", -- 2117 - 0x845  :  237 - 0xed
    "11111111", -- 2118 - 0x846  :  255 - 0xff
    "10111111", -- 2119 - 0x847  :  191 - 0xbf
    "00010100", -- 2120 - 0x848  :   20 - 0x14
    "10110101", -- 2121 - 0x849  :  181 - 0xb5
    "01000100", -- 2122 - 0x84a  :   68 - 0x44
    "01001010", -- 2123 - 0x84b  :   74 - 0x4a
    "10010010", -- 2124 - 0x84c  :  146 - 0x92
    "10010010", -- 2125 - 0x84d  :  146 - 0x92
    "01000100", -- 2126 - 0x84e  :   68 - 0x44
    "01001001", -- 2127 - 0x84f  :   73 - 0x49
    "11111111", -- 2128 - 0x850  :  255 - 0xff -- Sprite 0x85
    "10111111", -- 2129 - 0x851  :  191 - 0xbf
    "01111101", -- 2130 - 0x852  :  125 - 0x7d
    "11110111", -- 2131 - 0x853  :  247 - 0xf7
    "11011011", -- 2132 - 0x854  :  219 - 0xdb
    "11111101", -- 2133 - 0x855  :  253 - 0xfd
    "01111110", -- 2134 - 0x856  :  126 - 0x7e
    "11111011", -- 2135 - 0x857  :  251 - 0xfb
    "01000010", -- 2136 - 0x858  :   66 - 0x42
    "01001010", -- 2137 - 0x859  :   74 - 0x4a
    "11001010", -- 2138 - 0x85a  :  202 - 0xca
    "00101001", -- 2139 - 0x85b  :   41 - 0x29
    "10100110", -- 2140 - 0x85c  :  166 - 0xa6
    "10010010", -- 2141 - 0x85d  :  146 - 0x92
    "10001001", -- 2142 - 0x85e  :  137 - 0x89
    "00101101", -- 2143 - 0x85f  :   45 - 0x2d
    "11111111", -- 2144 - 0x860  :  255 - 0xff -- Sprite 0x86
    "11110111", -- 2145 - 0x861  :  247 - 0xf7
    "11111111", -- 2146 - 0x862  :  255 - 0xff
    "11011101", -- 2147 - 0x863  :  221 - 0xdd
    "01111111", -- 2148 - 0x864  :  127 - 0x7f
    "11110111", -- 2149 - 0x865  :  247 - 0xf7
    "11101111", -- 2150 - 0x866  :  239 - 0xef
    "10111101", -- 2151 - 0x867  :  189 - 0xbd
    "10001000", -- 2152 - 0x868  :  136 - 0x88
    "00101001", -- 2153 - 0x869  :   41 - 0x29
    "10000010", -- 2154 - 0x86a  :  130 - 0x82
    "10110110", -- 2155 - 0x86b  :  182 - 0xb6
    "10001000", -- 2156 - 0x86c  :  136 - 0x88
    "01001001", -- 2157 - 0x86d  :   73 - 0x49
    "01010010", -- 2158 - 0x86e  :   82 - 0x52
    "01010010", -- 2159 - 0x86f  :   82 - 0x52
    "01011111", -- 2160 - 0x870  :   95 - 0x5f -- Sprite 0x87
    "11111101", -- 2161 - 0x871  :  253 - 0xfd
    "11110110", -- 2162 - 0x872  :  246 - 0xf6
    "01111111", -- 2163 - 0x873  :  127 - 0x7f
    "10011111", -- 2164 - 0x874  :  159 - 0x9f
    "11111110", -- 2165 - 0x875  :  254 - 0xfe
    "11111111", -- 2166 - 0x876  :  255 - 0xff
    "11101111", -- 2167 - 0x877  :  239 - 0xef
    "10110010", -- 2168 - 0x878  :  178 - 0xb2
    "01001010", -- 2169 - 0x879  :   74 - 0x4a
    "10101001", -- 2170 - 0x87a  :  169 - 0xa9
    "10100100", -- 2171 - 0x87b  :  164 - 0xa4
    "01100010", -- 2172 - 0x87c  :   98 - 0x62
    "01001011", -- 2173 - 0x87d  :   75 - 0x4b
    "10010000", -- 2174 - 0x87e  :  144 - 0x90
    "10010010", -- 2175 - 0x87f  :  146 - 0x92
    "11111111", -- 2176 - 0x880  :  255 - 0xff -- Sprite 0x88
    "11111111", -- 2177 - 0x881  :  255 - 0xff
    "10011111", -- 2178 - 0x882  :  159 - 0x9f
    "10110011", -- 2179 - 0x883  :  179 - 0xb3
    "11110011", -- 2180 - 0x884  :  243 - 0xf3
    "11111111", -- 2181 - 0x885  :  255 - 0xff
    "11111111", -- 2182 - 0x886  :  255 - 0xff
    "11111111", -- 2183 - 0x887  :  255 - 0xff
    "00000000", -- 2184 - 0x888  :    0 - 0x0
    "01100000", -- 2185 - 0x889  :   96 - 0x60
    "11111110", -- 2186 - 0x88a  :  254 - 0xfe
    "11111111", -- 2187 - 0x88b  :  255 - 0xff
    "01111111", -- 2188 - 0x88c  :  127 - 0x7f
    "00011111", -- 2189 - 0x88d  :   31 - 0x1f
    "00001110", -- 2190 - 0x88e  :   14 - 0xe
    "00000000", -- 2191 - 0x88f  :    0 - 0x0
    "11111111", -- 2192 - 0x890  :  255 - 0xff -- Sprite 0x89
    "11001111", -- 2193 - 0x891  :  207 - 0xcf
    "11011111", -- 2194 - 0x892  :  223 - 0xdf
    "11111111", -- 2195 - 0x893  :  255 - 0xff
    "11110011", -- 2196 - 0x894  :  243 - 0xf3
    "11110011", -- 2197 - 0x895  :  243 - 0xf3
    "11111111", -- 2198 - 0x896  :  255 - 0xff
    "11111111", -- 2199 - 0x897  :  255 - 0xff
    "00110000", -- 2200 - 0x898  :   48 - 0x30
    "01111000", -- 2201 - 0x899  :  120 - 0x78
    "01111000", -- 2202 - 0x89a  :  120 - 0x78
    "00111110", -- 2203 - 0x89b  :   62 - 0x3e
    "00011111", -- 2204 - 0x89c  :   31 - 0x1f
    "00011111", -- 2205 - 0x89d  :   31 - 0x1f
    "00011111", -- 2206 - 0x89e  :   31 - 0x1f
    "00001110", -- 2207 - 0x89f  :   14 - 0xe
    "10111111", -- 2208 - 0x8a0  :  191 - 0xbf -- Sprite 0x8a
    "11110111", -- 2209 - 0x8a1  :  247 - 0xf7
    "11111101", -- 2210 - 0x8a2  :  253 - 0xfd
    "11111111", -- 2211 - 0x8a3  :  255 - 0xff
    "11111011", -- 2212 - 0x8a4  :  251 - 0xfb
    "10111111", -- 2213 - 0x8a5  :  191 - 0xbf
    "11111110", -- 2214 - 0x8a6  :  254 - 0xfe
    "11101111", -- 2215 - 0x8a7  :  239 - 0xef
    "01000000", -- 2216 - 0x8a8  :   64 - 0x40
    "00001000", -- 2217 - 0x8a9  :    8 - 0x8
    "00000010", -- 2218 - 0x8aa  :    2 - 0x2
    "00101000", -- 2219 - 0x8ab  :   40 - 0x28
    "00010100", -- 2220 - 0x8ac  :   20 - 0x14
    "01010100", -- 2221 - 0x8ad  :   84 - 0x54
    "00000001", -- 2222 - 0x8ae  :    1 - 0x1
    "00010000", -- 2223 - 0x8af  :   16 - 0x10
    "10111111", -- 2224 - 0x8b0  :  191 - 0xbf -- Sprite 0x8b
    "11111111", -- 2225 - 0x8b1  :  255 - 0xff
    "11101110", -- 2226 - 0x8b2  :  238 - 0xee
    "11111111", -- 2227 - 0x8b3  :  255 - 0xff
    "11011111", -- 2228 - 0x8b4  :  223 - 0xdf
    "01111101", -- 2229 - 0x8b5  :  125 - 0x7d
    "11111111", -- 2230 - 0x8b6  :  255 - 0xff
    "11011111", -- 2231 - 0x8b7  :  223 - 0xdf
    "01000000", -- 2232 - 0x8b8  :   64 - 0x40
    "00000000", -- 2233 - 0x8b9  :    0 - 0x0
    "10010001", -- 2234 - 0x8ba  :  145 - 0x91
    "00010100", -- 2235 - 0x8bb  :   20 - 0x14
    "00101000", -- 2236 - 0x8bc  :   40 - 0x28
    "10001010", -- 2237 - 0x8bd  :  138 - 0x8a
    "01000000", -- 2238 - 0x8be  :   64 - 0x40
    "00100000", -- 2239 - 0x8bf  :   32 - 0x20
    "11111111", -- 2240 - 0x8c0  :  255 - 0xff -- Sprite 0x8c
    "11111000", -- 2241 - 0x8c1  :  248 - 0xf8
    "11100010", -- 2242 - 0x8c2  :  226 - 0xe2
    "11010111", -- 2243 - 0x8c3  :  215 - 0xd7
    "11001111", -- 2244 - 0x8c4  :  207 - 0xcf
    "10011111", -- 2245 - 0x8c5  :  159 - 0x9f
    "10111110", -- 2246 - 0x8c6  :  190 - 0xbe
    "10011101", -- 2247 - 0x8c7  :  157 - 0x9d
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0
    "00000111", -- 2249 - 0x8c9  :    7 - 0x7
    "00011111", -- 2250 - 0x8ca  :   31 - 0x1f
    "00111111", -- 2251 - 0x8cb  :   63 - 0x3f
    "00111111", -- 2252 - 0x8cc  :   63 - 0x3f
    "01111111", -- 2253 - 0x8cd  :  127 - 0x7f
    "01111111", -- 2254 - 0x8ce  :  127 - 0x7f
    "01111111", -- 2255 - 0x8cf  :  127 - 0x7f
    "11111111", -- 2256 - 0x8d0  :  255 - 0xff -- Sprite 0x8d
    "00011111", -- 2257 - 0x8d1  :   31 - 0x1f
    "10100111", -- 2258 - 0x8d2  :  167 - 0xa7
    "11000011", -- 2259 - 0x8d3  :  195 - 0xc3
    "11100011", -- 2260 - 0x8d4  :  227 - 0xe3
    "01000001", -- 2261 - 0x8d5  :   65 - 0x41
    "10100001", -- 2262 - 0x8d6  :  161 - 0xa1
    "00000001", -- 2263 - 0x8d7  :    1 - 0x1
    "00000000", -- 2264 - 0x8d8  :    0 - 0x0
    "11100000", -- 2265 - 0x8d9  :  224 - 0xe0
    "11111000", -- 2266 - 0x8da  :  248 - 0xf8
    "11111000", -- 2267 - 0x8db  :  248 - 0xf8
    "11110000", -- 2268 - 0x8dc  :  240 - 0xf0
    "11111000", -- 2269 - 0x8dd  :  248 - 0xf8
    "11110100", -- 2270 - 0x8de  :  244 - 0xf4
    "11111000", -- 2271 - 0x8df  :  248 - 0xf8
    "10111110", -- 2272 - 0x8e0  :  190 - 0xbe -- Sprite 0x8e
    "11111111", -- 2273 - 0x8e1  :  255 - 0xff
    "11011111", -- 2274 - 0x8e2  :  223 - 0xdf
    "11111111", -- 2275 - 0x8e3  :  255 - 0xff
    "11101111", -- 2276 - 0x8e4  :  239 - 0xef
    "11111111", -- 2277 - 0x8e5  :  255 - 0xff
    "11110111", -- 2278 - 0x8e6  :  247 - 0xf7
    "11111111", -- 2279 - 0x8e7  :  255 - 0xff
    "01111111", -- 2280 - 0x8e8  :  127 - 0x7f
    "00111111", -- 2281 - 0x8e9  :   63 - 0x3f
    "00111111", -- 2282 - 0x8ea  :   63 - 0x3f
    "00011111", -- 2283 - 0x8eb  :   31 - 0x1f
    "00011111", -- 2284 - 0x8ec  :   31 - 0x1f
    "00001111", -- 2285 - 0x8ed  :   15 - 0xf
    "00001111", -- 2286 - 0x8ee  :   15 - 0xf
    "00000111", -- 2287 - 0x8ef  :    7 - 0x7
    "01111101", -- 2288 - 0x8f0  :  125 - 0x7d -- Sprite 0x8f
    "11111111", -- 2289 - 0x8f1  :  255 - 0xff
    "11111011", -- 2290 - 0x8f2  :  251 - 0xfb
    "11111111", -- 2291 - 0x8f3  :  255 - 0xff
    "11110111", -- 2292 - 0x8f4  :  247 - 0xf7
    "11111111", -- 2293 - 0x8f5  :  255 - 0xff
    "11101111", -- 2294 - 0x8f6  :  239 - 0xef
    "11111111", -- 2295 - 0x8f7  :  255 - 0xff
    "11111110", -- 2296 - 0x8f8  :  254 - 0xfe
    "11111100", -- 2297 - 0x8f9  :  252 - 0xfc
    "11111100", -- 2298 - 0x8fa  :  252 - 0xfc
    "11111000", -- 2299 - 0x8fb  :  248 - 0xf8
    "11111000", -- 2300 - 0x8fc  :  248 - 0xf8
    "11110000", -- 2301 - 0x8fd  :  240 - 0xf0
    "11110000", -- 2302 - 0x8fe  :  240 - 0xf0
    "11100000", -- 2303 - 0x8ff  :  224 - 0xe0
    "10111110", -- 2304 - 0x900  :  190 - 0xbe -- Sprite 0x90
    "11110111", -- 2305 - 0x901  :  247 - 0xf7
    "11111111", -- 2306 - 0x902  :  255 - 0xff
    "11011111", -- 2307 - 0x903  :  223 - 0xdf
    "11111011", -- 2308 - 0x904  :  251 - 0xfb
    "11111110", -- 2309 - 0x905  :  254 - 0xfe
    "10111111", -- 2310 - 0x906  :  191 - 0xbf
    "11110111", -- 2311 - 0x907  :  247 - 0xf7
    "01000001", -- 2312 - 0x908  :   65 - 0x41
    "00001000", -- 2313 - 0x909  :    8 - 0x8
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "00100000", -- 2315 - 0x90b  :   32 - 0x20
    "00000100", -- 2316 - 0x90c  :    4 - 0x4
    "00000001", -- 2317 - 0x90d  :    1 - 0x1
    "01000000", -- 2318 - 0x90e  :   64 - 0x40
    "00001000", -- 2319 - 0x90f  :    8 - 0x8
    "11101110", -- 2320 - 0x910  :  238 - 0xee -- Sprite 0x91
    "11111111", -- 2321 - 0x911  :  255 - 0xff
    "01111011", -- 2322 - 0x912  :  123 - 0x7b
    "11111101", -- 2323 - 0x913  :  253 - 0xfd
    "11101111", -- 2324 - 0x914  :  239 - 0xef
    "11111111", -- 2325 - 0x915  :  255 - 0xff
    "10111101", -- 2326 - 0x916  :  189 - 0xbd
    "11111111", -- 2327 - 0x917  :  255 - 0xff
    "00010001", -- 2328 - 0x918  :   17 - 0x11
    "00000000", -- 2329 - 0x919  :    0 - 0x0
    "10000100", -- 2330 - 0x91a  :  132 - 0x84
    "00000010", -- 2331 - 0x91b  :    2 - 0x2
    "00010000", -- 2332 - 0x91c  :   16 - 0x10
    "00000000", -- 2333 - 0x91d  :    0 - 0x0
    "01000010", -- 2334 - 0x91e  :   66 - 0x42
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "11111011", -- 2336 - 0x920  :  251 - 0xfb -- Sprite 0x92
    "10111111", -- 2337 - 0x921  :  191 - 0xbf
    "11101111", -- 2338 - 0x922  :  239 - 0xef
    "11111101", -- 2339 - 0x923  :  253 - 0xfd
    "11111111", -- 2340 - 0x924  :  255 - 0xff
    "10111111", -- 2341 - 0x925  :  191 - 0xbf
    "11111011", -- 2342 - 0x926  :  251 - 0xfb
    "11011111", -- 2343 - 0x927  :  223 - 0xdf
    "00000100", -- 2344 - 0x928  :    4 - 0x4
    "01000000", -- 2345 - 0x929  :   64 - 0x40
    "00010000", -- 2346 - 0x92a  :   16 - 0x10
    "00000010", -- 2347 - 0x92b  :    2 - 0x2
    "00000000", -- 2348 - 0x92c  :    0 - 0x0
    "01000000", -- 2349 - 0x92d  :   64 - 0x40
    "00000100", -- 2350 - 0x92e  :    4 - 0x4
    "00100000", -- 2351 - 0x92f  :   32 - 0x20
    "10111101", -- 2352 - 0x930  :  189 - 0xbd -- Sprite 0x93
    "11111111", -- 2353 - 0x931  :  255 - 0xff
    "01110111", -- 2354 - 0x932  :  119 - 0x77
    "11111110", -- 2355 - 0x933  :  254 - 0xfe
    "11011111", -- 2356 - 0x934  :  223 - 0xdf
    "11111011", -- 2357 - 0x935  :  251 - 0xfb
    "11101111", -- 2358 - 0x936  :  239 - 0xef
    "01111111", -- 2359 - 0x937  :  127 - 0x7f
    "01000010", -- 2360 - 0x938  :   66 - 0x42
    "00000000", -- 2361 - 0x939  :    0 - 0x0
    "10001000", -- 2362 - 0x93a  :  136 - 0x88
    "00000001", -- 2363 - 0x93b  :    1 - 0x1
    "00100000", -- 2364 - 0x93c  :   32 - 0x20
    "00000100", -- 2365 - 0x93d  :    4 - 0x4
    "00010000", -- 2366 - 0x93e  :   16 - 0x10
    "10000000", -- 2367 - 0x93f  :  128 - 0x80
    "01111111", -- 2368 - 0x940  :  127 - 0x7f -- Sprite 0x94
    "11110111", -- 2369 - 0x941  :  247 - 0xf7
    "11011101", -- 2370 - 0x942  :  221 - 0xdd
    "01111011", -- 2371 - 0x943  :  123 - 0x7b
    "11111111", -- 2372 - 0x944  :  255 - 0xff
    "11101110", -- 2373 - 0x945  :  238 - 0xee
    "10111011", -- 2374 - 0x946  :  187 - 0xbb
    "11111101", -- 2375 - 0x947  :  253 - 0xfd
    "11001000", -- 2376 - 0x948  :  200 - 0xc8
    "00101010", -- 2377 - 0x949  :   42 - 0x2a
    "10100010", -- 2378 - 0x94a  :  162 - 0xa2
    "10010100", -- 2379 - 0x94b  :  148 - 0x94
    "10010001", -- 2380 - 0x94c  :  145 - 0x91
    "01010101", -- 2381 - 0x94d  :   85 - 0x55
    "01000100", -- 2382 - 0x94e  :   68 - 0x44
    "00010010", -- 2383 - 0x94f  :   18 - 0x12
    "11010111", -- 2384 - 0x950  :  215 - 0xd7 -- Sprite 0x95
    "01111111", -- 2385 - 0x951  :  127 - 0x7f
    "11111101", -- 2386 - 0x952  :  253 - 0xfd
    "11101110", -- 2387 - 0x953  :  238 - 0xee
    "11110111", -- 2388 - 0x954  :  247 - 0xf7
    "10111011", -- 2389 - 0x955  :  187 - 0xbb
    "11101111", -- 2390 - 0x956  :  239 - 0xef
    "11110111", -- 2391 - 0x957  :  247 - 0xf7
    "10101010", -- 2392 - 0x958  :  170 - 0xaa
    "10100010", -- 2393 - 0x959  :  162 - 0xa2
    "00010010", -- 2394 - 0x95a  :   18 - 0x12
    "01010011", -- 2395 - 0x95b  :   83 - 0x53
    "01001100", -- 2396 - 0x95c  :   76 - 0x4c
    "01010101", -- 2397 - 0x95d  :   85 - 0x55
    "10010001", -- 2398 - 0x95e  :  145 - 0x91
    "01001000", -- 2399 - 0x95f  :   72 - 0x48
    "10111111", -- 2400 - 0x960  :  191 - 0xbf -- Sprite 0x96
    "11101110", -- 2401 - 0x961  :  238 - 0xee
    "11011011", -- 2402 - 0x962  :  219 - 0xdb
    "11111111", -- 2403 - 0x963  :  255 - 0xff
    "01110111", -- 2404 - 0x964  :  119 - 0x77
    "11011101", -- 2405 - 0x965  :  221 - 0xdd
    "11101111", -- 2406 - 0x966  :  239 - 0xef
    "11111011", -- 2407 - 0x967  :  251 - 0xfb
    "01010001", -- 2408 - 0x968  :   81 - 0x51
    "00010101", -- 2409 - 0x969  :   21 - 0x15
    "10100100", -- 2410 - 0x96a  :  164 - 0xa4
    "10001100", -- 2411 - 0x96b  :  140 - 0x8c
    "10101010", -- 2412 - 0x96c  :  170 - 0xaa
    "00100010", -- 2413 - 0x96d  :   34 - 0x22
    "10010000", -- 2414 - 0x96e  :  144 - 0x90
    "01000110", -- 2415 - 0x96f  :   70 - 0x46
    "11111101", -- 2416 - 0x970  :  253 - 0xfd -- Sprite 0x97
    "11101110", -- 2417 - 0x971  :  238 - 0xee
    "11111011", -- 2418 - 0x972  :  251 - 0xfb
    "11111101", -- 2419 - 0x973  :  253 - 0xfd
    "11110101", -- 2420 - 0x974  :  245 - 0xf5
    "11011111", -- 2421 - 0x975  :  223 - 0xdf
    "01111111", -- 2422 - 0x976  :  127 - 0x7f
    "10111011", -- 2423 - 0x977  :  187 - 0xbb
    "00010011", -- 2424 - 0x978  :   19 - 0x13
    "01010101", -- 2425 - 0x979  :   85 - 0x55
    "01100100", -- 2426 - 0x97a  :  100 - 0x64
    "00010010", -- 2427 - 0x97b  :   18 - 0x12
    "10101010", -- 2428 - 0x97c  :  170 - 0xaa
    "10101000", -- 2429 - 0x97d  :  168 - 0xa8
    "10000100", -- 2430 - 0x97e  :  132 - 0x84
    "11010100", -- 2431 - 0x97f  :  212 - 0xd4
    "11111111", -- 2432 - 0x980  :  255 - 0xff -- Sprite 0x98
    "11001111", -- 2433 - 0x981  :  207 - 0xcf
    "11011111", -- 2434 - 0x982  :  223 - 0xdf
    "11111111", -- 2435 - 0x983  :  255 - 0xff
    "11110011", -- 2436 - 0x984  :  243 - 0xf3
    "11110011", -- 2437 - 0x985  :  243 - 0xf3
    "11111111", -- 2438 - 0x986  :  255 - 0xff
    "11111111", -- 2439 - 0x987  :  255 - 0xff
    "00110000", -- 2440 - 0x988  :   48 - 0x30
    "01111000", -- 2441 - 0x989  :  120 - 0x78
    "01111000", -- 2442 - 0x98a  :  120 - 0x78
    "00111110", -- 2443 - 0x98b  :   62 - 0x3e
    "00011111", -- 2444 - 0x98c  :   31 - 0x1f
    "00011111", -- 2445 - 0x98d  :   31 - 0x1f
    "00011111", -- 2446 - 0x98e  :   31 - 0x1f
    "00001110", -- 2447 - 0x98f  :   14 - 0xe
    "11111111", -- 2448 - 0x990  :  255 - 0xff -- Sprite 0x99
    "11111111", -- 2449 - 0x991  :  255 - 0xff
    "10011111", -- 2450 - 0x992  :  159 - 0x9f
    "10110011", -- 2451 - 0x993  :  179 - 0xb3
    "11110011", -- 2452 - 0x994  :  243 - 0xf3
    "11111111", -- 2453 - 0x995  :  255 - 0xff
    "11111111", -- 2454 - 0x996  :  255 - 0xff
    "11111111", -- 2455 - 0x997  :  255 - 0xff
    "00000000", -- 2456 - 0x998  :    0 - 0x0
    "01100000", -- 2457 - 0x999  :   96 - 0x60
    "11111110", -- 2458 - 0x99a  :  254 - 0xfe
    "11111111", -- 2459 - 0x99b  :  255 - 0xff
    "01111111", -- 2460 - 0x99c  :  127 - 0x7f
    "00011111", -- 2461 - 0x99d  :   31 - 0x1f
    "00001110", -- 2462 - 0x99e  :   14 - 0xe
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "10111111", -- 2464 - 0x9a0  :  191 - 0xbf -- Sprite 0x9a
    "11110111", -- 2465 - 0x9a1  :  247 - 0xf7
    "11111111", -- 2466 - 0x9a2  :  255 - 0xff
    "11011111", -- 2467 - 0x9a3  :  223 - 0xdf
    "11111011", -- 2468 - 0x9a4  :  251 - 0xfb
    "11111111", -- 2469 - 0x9a5  :  255 - 0xff
    "10111111", -- 2470 - 0x9a6  :  191 - 0xbf
    "11110111", -- 2471 - 0x9a7  :  247 - 0xf7
    "01000000", -- 2472 - 0x9a8  :   64 - 0x40
    "00001100", -- 2473 - 0x9a9  :   12 - 0xc
    "00000000", -- 2474 - 0x9aa  :    0 - 0x0
    "00101000", -- 2475 - 0x9ab  :   40 - 0x28
    "00101100", -- 2476 - 0x9ac  :   44 - 0x2c
    "00010001", -- 2477 - 0x9ad  :   17 - 0x11
    "01000000", -- 2478 - 0x9ae  :   64 - 0x40
    "00001000", -- 2479 - 0x9af  :    8 - 0x8
    "11011111", -- 2480 - 0x9b0  :  223 - 0xdf -- Sprite 0x9b
    "11111111", -- 2481 - 0x9b1  :  255 - 0xff
    "01111011", -- 2482 - 0x9b2  :  123 - 0x7b
    "11111111", -- 2483 - 0x9b3  :  255 - 0xff
    "11101111", -- 2484 - 0x9b4  :  239 - 0xef
    "11111101", -- 2485 - 0x9b5  :  253 - 0xfd
    "10111111", -- 2486 - 0x9b6  :  191 - 0xbf
    "11111111", -- 2487 - 0x9b7  :  255 - 0xff
    "00100000", -- 2488 - 0x9b8  :   32 - 0x20
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "10010100", -- 2490 - 0x9ba  :  148 - 0x94
    "01001000", -- 2491 - 0x9bb  :   72 - 0x48
    "00011000", -- 2492 - 0x9bc  :   24 - 0x18
    "00000110", -- 2493 - 0x9bd  :    6 - 0x6
    "01000000", -- 2494 - 0x9be  :   64 - 0x40
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "10111010", -- 2496 - 0x9c0  :  186 - 0xba -- Sprite 0x9c
    "10011100", -- 2497 - 0x9c1  :  156 - 0x9c
    "10101010", -- 2498 - 0x9c2  :  170 - 0xaa
    "11000000", -- 2499 - 0x9c3  :  192 - 0xc0
    "11000000", -- 2500 - 0x9c4  :  192 - 0xc0
    "11100000", -- 2501 - 0x9c5  :  224 - 0xe0
    "11111000", -- 2502 - 0x9c6  :  248 - 0xf8
    "11111111", -- 2503 - 0x9c7  :  255 - 0xff
    "01111111", -- 2504 - 0x9c8  :  127 - 0x7f
    "01111111", -- 2505 - 0x9c9  :  127 - 0x7f
    "01111111", -- 2506 - 0x9ca  :  127 - 0x7f
    "00111111", -- 2507 - 0x9cb  :   63 - 0x3f
    "00110101", -- 2508 - 0x9cc  :   53 - 0x35
    "00000010", -- 2509 - 0x9cd  :    2 - 0x2
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000001", -- 2512 - 0x9d0  :    1 - 0x1 -- Sprite 0x9d
    "00000001", -- 2513 - 0x9d1  :    1 - 0x1
    "00000001", -- 2514 - 0x9d2  :    1 - 0x1
    "00000011", -- 2515 - 0x9d3  :    3 - 0x3
    "00000011", -- 2516 - 0x9d4  :    3 - 0x3
    "00000111", -- 2517 - 0x9d5  :    7 - 0x7
    "00011111", -- 2518 - 0x9d6  :   31 - 0x1f
    "11111111", -- 2519 - 0x9d7  :  255 - 0xff
    "11110100", -- 2520 - 0x9d8  :  244 - 0xf4
    "11111000", -- 2521 - 0x9d9  :  248 - 0xf8
    "11110000", -- 2522 - 0x9da  :  240 - 0xf0
    "11101000", -- 2523 - 0x9db  :  232 - 0xe8
    "01010000", -- 2524 - 0x9dc  :   80 - 0x50
    "10000000", -- 2525 - 0x9dd  :  128 - 0x80
    "00000000", -- 2526 - 0x9de  :    0 - 0x0
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "01111101", -- 2528 - 0x9e0  :  125 - 0x7d -- Sprite 0x9e
    "11111111", -- 2529 - 0x9e1  :  255 - 0xff
    "11111011", -- 2530 - 0x9e2  :  251 - 0xfb
    "11111111", -- 2531 - 0x9e3  :  255 - 0xff
    "11111111", -- 2532 - 0x9e4  :  255 - 0xff
    "11111011", -- 2533 - 0x9e5  :  251 - 0xfb
    "11111111", -- 2534 - 0x9e6  :  255 - 0xff
    "01111101", -- 2535 - 0x9e7  :  125 - 0x7d
    "11111110", -- 2536 - 0x9e8  :  254 - 0xfe
    "11111100", -- 2537 - 0x9e9  :  252 - 0xfc
    "11111100", -- 2538 - 0x9ea  :  252 - 0xfc
    "11111000", -- 2539 - 0x9eb  :  248 - 0xf8
    "11111000", -- 2540 - 0x9ec  :  248 - 0xf8
    "11111100", -- 2541 - 0x9ed  :  252 - 0xfc
    "11111100", -- 2542 - 0x9ee  :  252 - 0xfc
    "11111110", -- 2543 - 0x9ef  :  254 - 0xfe
    "11111111", -- 2544 - 0x9f0  :  255 - 0xff -- Sprite 0x9f
    "11111111", -- 2545 - 0x9f1  :  255 - 0xff
    "10111101", -- 2546 - 0x9f2  :  189 - 0xbd
    "11111111", -- 2547 - 0x9f3  :  255 - 0xff
    "11111111", -- 2548 - 0x9f4  :  255 - 0xff
    "11111111", -- 2549 - 0x9f5  :  255 - 0xff
    "11111111", -- 2550 - 0x9f6  :  255 - 0xff
    "10111101", -- 2551 - 0x9f7  :  189 - 0xbd
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "01111110", -- 2554 - 0x9fa  :  126 - 0x7e
    "01111110", -- 2555 - 0x9fb  :  126 - 0x7e
    "01111110", -- 2556 - 0x9fc  :  126 - 0x7e
    "01111110", -- 2557 - 0x9fd  :  126 - 0x7e
    "01111110", -- 2558 - 0x9fe  :  126 - 0x7e
    "01111110", -- 2559 - 0x9ff  :  126 - 0x7e
    "11101111", -- 2560 - 0xa00  :  239 - 0xef -- Sprite 0xa0
    "11000111", -- 2561 - 0xa01  :  199 - 0xc7
    "10000011", -- 2562 - 0xa02  :  131 - 0x83
    "00000111", -- 2563 - 0xa03  :    7 - 0x7
    "10001111", -- 2564 - 0xa04  :  143 - 0x8f
    "11011101", -- 2565 - 0xa05  :  221 - 0xdd
    "11111010", -- 2566 - 0xa06  :  250 - 0xfa
    "11111101", -- 2567 - 0xa07  :  253 - 0xfd
    "00010000", -- 2568 - 0xa08  :   16 - 0x10
    "00111000", -- 2569 - 0xa09  :   56 - 0x38
    "01111100", -- 2570 - 0xa0a  :  124 - 0x7c
    "11111000", -- 2571 - 0xa0b  :  248 - 0xf8
    "01110000", -- 2572 - 0xa0c  :  112 - 0x70
    "00100010", -- 2573 - 0xa0d  :   34 - 0x22
    "00000101", -- 2574 - 0xa0e  :    5 - 0x5
    "00000010", -- 2575 - 0xa0f  :    2 - 0x2
    "11101111", -- 2576 - 0xa10  :  239 - 0xef -- Sprite 0xa1
    "11000111", -- 2577 - 0xa11  :  199 - 0xc7
    "10000011", -- 2578 - 0xa12  :  131 - 0x83
    "00011111", -- 2579 - 0xa13  :   31 - 0x1f
    "10010000", -- 2580 - 0xa14  :  144 - 0x90
    "11010100", -- 2581 - 0xa15  :  212 - 0xd4
    "11110011", -- 2582 - 0xa16  :  243 - 0xf3
    "11110010", -- 2583 - 0xa17  :  242 - 0xf2
    "00010000", -- 2584 - 0xa18  :   16 - 0x10
    "00111000", -- 2585 - 0xa19  :   56 - 0x38
    "01111100", -- 2586 - 0xa1a  :  124 - 0x7c
    "11100000", -- 2587 - 0xa1b  :  224 - 0xe0
    "01100000", -- 2588 - 0xa1c  :   96 - 0x60
    "00100000", -- 2589 - 0xa1d  :   32 - 0x20
    "00000000", -- 2590 - 0xa1e  :    0 - 0x0
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "11101111", -- 2592 - 0xa20  :  239 - 0xef -- Sprite 0xa2
    "11000111", -- 2593 - 0xa21  :  199 - 0xc7
    "10000011", -- 2594 - 0xa22  :  131 - 0x83
    "11111111", -- 2595 - 0xa23  :  255 - 0xff
    "00000000", -- 2596 - 0xa24  :    0 - 0x0
    "00000000", -- 2597 - 0xa25  :    0 - 0x0
    "01010101", -- 2598 - 0xa26  :   85 - 0x55
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00010000", -- 2600 - 0xa28  :   16 - 0x10
    "00111000", -- 2601 - 0xa29  :   56 - 0x38
    "01111100", -- 2602 - 0xa2a  :  124 - 0x7c
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "11110000", -- 2608 - 0xa30  :  240 - 0xf0 -- Sprite 0xa3
    "11010010", -- 2609 - 0xa31  :  210 - 0xd2
    "10010000", -- 2610 - 0xa32  :  144 - 0x90
    "00010010", -- 2611 - 0xa33  :   18 - 0x12
    "10010000", -- 2612 - 0xa34  :  144 - 0x90
    "11010010", -- 2613 - 0xa35  :  210 - 0xd2
    "11110000", -- 2614 - 0xa36  :  240 - 0xf0
    "11110010", -- 2615 - 0xa37  :  242 - 0xf2
    "00000000", -- 2616 - 0xa38  :    0 - 0x0
    "00100000", -- 2617 - 0xa39  :   32 - 0x20
    "01100000", -- 2618 - 0xa3a  :   96 - 0x60
    "11100000", -- 2619 - 0xa3b  :  224 - 0xe0
    "01100000", -- 2620 - 0xa3c  :   96 - 0x60
    "00100000", -- 2621 - 0xa3d  :   32 - 0x20
    "00000000", -- 2622 - 0xa3e  :    0 - 0x0
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "11110000", -- 2624 - 0xa40  :  240 - 0xf0 -- Sprite 0xa4
    "11010011", -- 2625 - 0xa41  :  211 - 0xd3
    "10010100", -- 2626 - 0xa42  :  148 - 0x94
    "00011000", -- 2627 - 0xa43  :   24 - 0x18
    "10011111", -- 2628 - 0xa44  :  159 - 0x9f
    "11011101", -- 2629 - 0xa45  :  221 - 0xdd
    "11111010", -- 2630 - 0xa46  :  250 - 0xfa
    "11111101", -- 2631 - 0xa47  :  253 - 0xfd
    "00000000", -- 2632 - 0xa48  :    0 - 0x0
    "00100000", -- 2633 - 0xa49  :   32 - 0x20
    "01100011", -- 2634 - 0xa4a  :   99 - 0x63
    "11100111", -- 2635 - 0xa4b  :  231 - 0xe7
    "01100000", -- 2636 - 0xa4c  :   96 - 0x60
    "00100010", -- 2637 - 0xa4d  :   34 - 0x22
    "00000101", -- 2638 - 0xa4e  :    5 - 0x5
    "00000010", -- 2639 - 0xa4f  :    2 - 0x2
    "00000000", -- 2640 - 0xa50  :    0 - 0x0 -- Sprite 0xa5
    "11111111", -- 2641 - 0xa51  :  255 - 0xff
    "00000000", -- 2642 - 0xa52  :    0 - 0x0
    "00000000", -- 2643 - 0xa53  :    0 - 0x0
    "11111111", -- 2644 - 0xa54  :  255 - 0xff
    "11011101", -- 2645 - 0xa55  :  221 - 0xdd
    "11111010", -- 2646 - 0xa56  :  250 - 0xfa
    "11111101", -- 2647 - 0xa57  :  253 - 0xfd
    "00000000", -- 2648 - 0xa58  :    0 - 0x0
    "00000000", -- 2649 - 0xa59  :    0 - 0x0
    "11111111", -- 2650 - 0xa5a  :  255 - 0xff
    "11111111", -- 2651 - 0xa5b  :  255 - 0xff
    "00000000", -- 2652 - 0xa5c  :    0 - 0x0
    "00100010", -- 2653 - 0xa5d  :   34 - 0x22
    "00000101", -- 2654 - 0xa5e  :    5 - 0x5
    "00000010", -- 2655 - 0xa5f  :    2 - 0x2
    "11101111", -- 2656 - 0xa60  :  239 - 0xef -- Sprite 0xa6
    "11000111", -- 2657 - 0xa61  :  199 - 0xc7
    "10000011", -- 2658 - 0xa62  :  131 - 0x83
    "11111111", -- 2659 - 0xa63  :  255 - 0xff
    "00011111", -- 2660 - 0xa64  :   31 - 0x1f
    "00101101", -- 2661 - 0xa65  :   45 - 0x2d
    "01001010", -- 2662 - 0xa66  :   74 - 0x4a
    "01001101", -- 2663 - 0xa67  :   77 - 0x4d
    "00010000", -- 2664 - 0xa68  :   16 - 0x10
    "00111000", -- 2665 - 0xa69  :   56 - 0x38
    "01111100", -- 2666 - 0xa6a  :  124 - 0x7c
    "00000000", -- 2667 - 0xa6b  :    0 - 0x0
    "00000000", -- 2668 - 0xa6c  :    0 - 0x0
    "00010010", -- 2669 - 0xa6d  :   18 - 0x12
    "00110101", -- 2670 - 0xa6e  :   53 - 0x35
    "00110010", -- 2671 - 0xa6f  :   50 - 0x32
    "01001111", -- 2672 - 0xa70  :   79 - 0x4f -- Sprite 0xa7
    "01001111", -- 2673 - 0xa71  :   79 - 0x4f
    "01001011", -- 2674 - 0xa72  :   75 - 0x4b
    "01001111", -- 2675 - 0xa73  :   79 - 0x4f
    "01001111", -- 2676 - 0xa74  :   79 - 0x4f
    "01001101", -- 2677 - 0xa75  :   77 - 0x4d
    "01001010", -- 2678 - 0xa76  :   74 - 0x4a
    "01001101", -- 2679 - 0xa77  :   77 - 0x4d
    "00110000", -- 2680 - 0xa78  :   48 - 0x30
    "00110000", -- 2681 - 0xa79  :   48 - 0x30
    "00110100", -- 2682 - 0xa7a  :   52 - 0x34
    "00110000", -- 2683 - 0xa7b  :   48 - 0x30
    "00110000", -- 2684 - 0xa7c  :   48 - 0x30
    "00110010", -- 2685 - 0xa7d  :   50 - 0x32
    "00110101", -- 2686 - 0xa7e  :   53 - 0x35
    "00110010", -- 2687 - 0xa7f  :   50 - 0x32
    "01001111", -- 2688 - 0xa80  :   79 - 0x4f -- Sprite 0xa8
    "11001111", -- 2689 - 0xa81  :  207 - 0xcf
    "00001011", -- 2690 - 0xa82  :   11 - 0xb
    "00001111", -- 2691 - 0xa83  :   15 - 0xf
    "11111111", -- 2692 - 0xa84  :  255 - 0xff
    "11011101", -- 2693 - 0xa85  :  221 - 0xdd
    "11111010", -- 2694 - 0xa86  :  250 - 0xfa
    "11111101", -- 2695 - 0xa87  :  253 - 0xfd
    "00110000", -- 2696 - 0xa88  :   48 - 0x30
    "00110000", -- 2697 - 0xa89  :   48 - 0x30
    "11110100", -- 2698 - 0xa8a  :  244 - 0xf4
    "11110000", -- 2699 - 0xa8b  :  240 - 0xf0
    "00000000", -- 2700 - 0xa8c  :    0 - 0x0
    "00100010", -- 2701 - 0xa8d  :   34 - 0x22
    "00000101", -- 2702 - 0xa8e  :    5 - 0x5
    "00000010", -- 2703 - 0xa8f  :    2 - 0x2
    "11111111", -- 2704 - 0xa90  :  255 - 0xff -- Sprite 0xa9
    "11111111", -- 2705 - 0xa91  :  255 - 0xff
    "11111111", -- 2706 - 0xa92  :  255 - 0xff
    "11111111", -- 2707 - 0xa93  :  255 - 0xff
    "11111111", -- 2708 - 0xa94  :  255 - 0xff
    "11111111", -- 2709 - 0xa95  :  255 - 0xff
    "11111111", -- 2710 - 0xa96  :  255 - 0xff
    "11111111", -- 2711 - 0xa97  :  255 - 0xff
    "00000000", -- 2712 - 0xa98  :    0 - 0x0
    "00000000", -- 2713 - 0xa99  :    0 - 0x0
    "00000000", -- 2714 - 0xa9a  :    0 - 0x0
    "00000000", -- 2715 - 0xa9b  :    0 - 0x0
    "00000000", -- 2716 - 0xa9c  :    0 - 0x0
    "00000000", -- 2717 - 0xa9d  :    0 - 0x0
    "00000000", -- 2718 - 0xa9e  :    0 - 0x0
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "11111111", -- 2720 - 0xaa0  :  255 - 0xff -- Sprite 0xaa
    "11111111", -- 2721 - 0xaa1  :  255 - 0xff
    "10101111", -- 2722 - 0xaa2  :  175 - 0xaf
    "01010111", -- 2723 - 0xaa3  :   87 - 0x57
    "10001111", -- 2724 - 0xaa4  :  143 - 0x8f
    "11011101", -- 2725 - 0xaa5  :  221 - 0xdd
    "11111010", -- 2726 - 0xaa6  :  250 - 0xfa
    "11111101", -- 2727 - 0xaa7  :  253 - 0xfd
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "01010000", -- 2730 - 0xaaa  :   80 - 0x50
    "10101000", -- 2731 - 0xaab  :  168 - 0xa8
    "01110000", -- 2732 - 0xaac  :  112 - 0x70
    "00100010", -- 2733 - 0xaad  :   34 - 0x22
    "00000101", -- 2734 - 0xaae  :    5 - 0x5
    "00000010", -- 2735 - 0xaaf  :    2 - 0x2
    "11111111", -- 2736 - 0xab0  :  255 - 0xff -- Sprite 0xab
    "00000000", -- 2737 - 0xab1  :    0 - 0x0
    "00000000", -- 2738 - 0xab2  :    0 - 0x0
    "00000000", -- 2739 - 0xab3  :    0 - 0x0
    "00000000", -- 2740 - 0xab4  :    0 - 0x0
    "00000000", -- 2741 - 0xab5  :    0 - 0x0
    "00000000", -- 2742 - 0xab6  :    0 - 0x0
    "00000000", -- 2743 - 0xab7  :    0 - 0x0
    "00000000", -- 2744 - 0xab8  :    0 - 0x0
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "00000000", -- 2747 - 0xabb  :    0 - 0x0
    "00000000", -- 2748 - 0xabc  :    0 - 0x0
    "00000000", -- 2749 - 0xabd  :    0 - 0x0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "00000000", -- 2752 - 0xac0  :    0 - 0x0 -- Sprite 0xac
    "00000000", -- 2753 - 0xac1  :    0 - 0x0
    "00000000", -- 2754 - 0xac2  :    0 - 0x0
    "00000000", -- 2755 - 0xac3  :    0 - 0x0
    "00000000", -- 2756 - 0xac4  :    0 - 0x0
    "00000000", -- 2757 - 0xac5  :    0 - 0x0
    "00000000", -- 2758 - 0xac6  :    0 - 0x0
    "00000000", -- 2759 - 0xac7  :    0 - 0x0
    "00000000", -- 2760 - 0xac8  :    0 - 0x0
    "00000000", -- 2761 - 0xac9  :    0 - 0x0
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000000", -- 2763 - 0xacb  :    0 - 0x0
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "00000000", -- 2768 - 0xad0  :    0 - 0x0 -- Sprite 0xad
    "11111111", -- 2769 - 0xad1  :  255 - 0xff
    "00000000", -- 2770 - 0xad2  :    0 - 0x0
    "11111111", -- 2771 - 0xad3  :  255 - 0xff
    "11111111", -- 2772 - 0xad4  :  255 - 0xff
    "11111111", -- 2773 - 0xad5  :  255 - 0xff
    "11111111", -- 2774 - 0xad6  :  255 - 0xff
    "11111111", -- 2775 - 0xad7  :  255 - 0xff
    "00000000", -- 2776 - 0xad8  :    0 - 0x0
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "11111111", -- 2778 - 0xada  :  255 - 0xff
    "00000000", -- 2779 - 0xadb  :    0 - 0x0
    "00000000", -- 2780 - 0xadc  :    0 - 0x0
    "00000000", -- 2781 - 0xadd  :    0 - 0x0
    "00000000", -- 2782 - 0xade  :    0 - 0x0
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "11111111", -- 2784 - 0xae0  :  255 - 0xff -- Sprite 0xae
    "11111111", -- 2785 - 0xae1  :  255 - 0xff
    "11111111", -- 2786 - 0xae2  :  255 - 0xff
    "11111111", -- 2787 - 0xae3  :  255 - 0xff
    "11111111", -- 2788 - 0xae4  :  255 - 0xff
    "00000000", -- 2789 - 0xae5  :    0 - 0x0
    "11111111", -- 2790 - 0xae6  :  255 - 0xff
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "00000000", -- 2792 - 0xae8  :    0 - 0x0
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000000", -- 2794 - 0xaea  :    0 - 0x0
    "00000000", -- 2795 - 0xaeb  :    0 - 0x0
    "00000000", -- 2796 - 0xaec  :    0 - 0x0
    "11111111", -- 2797 - 0xaed  :  255 - 0xff
    "00000000", -- 2798 - 0xaee  :    0 - 0x0
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "11111111", -- 2800 - 0xaf0  :  255 - 0xff -- Sprite 0xaf
    "11111111", -- 2801 - 0xaf1  :  255 - 0xff
    "11111111", -- 2802 - 0xaf2  :  255 - 0xff
    "11111111", -- 2803 - 0xaf3  :  255 - 0xff
    "11111111", -- 2804 - 0xaf4  :  255 - 0xff
    "11111111", -- 2805 - 0xaf5  :  255 - 0xff
    "11111111", -- 2806 - 0xaf6  :  255 - 0xff
    "11111111", -- 2807 - 0xaf7  :  255 - 0xff
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0
    "00000000", -- 2809 - 0xaf9  :    0 - 0x0
    "00000000", -- 2810 - 0xafa  :    0 - 0x0
    "00000000", -- 2811 - 0xafb  :    0 - 0x0
    "00000000", -- 2812 - 0xafc  :    0 - 0x0
    "00000000", -- 2813 - 0xafd  :    0 - 0x0
    "00000000", -- 2814 - 0xafe  :    0 - 0x0
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "00000000", -- 2816 - 0xb00  :    0 - 0x0 -- Sprite 0xb0
    "00011111", -- 2817 - 0xb01  :   31 - 0x1f
    "00010000", -- 2818 - 0xb02  :   16 - 0x10
    "00010000", -- 2819 - 0xb03  :   16 - 0x10
    "00010000", -- 2820 - 0xb04  :   16 - 0x10
    "00010000", -- 2821 - 0xb05  :   16 - 0x10
    "00010000", -- 2822 - 0xb06  :   16 - 0x10
    "00010000", -- 2823 - 0xb07  :   16 - 0x10
    "00000000", -- 2824 - 0xb08  :    0 - 0x0
    "00011111", -- 2825 - 0xb09  :   31 - 0x1f
    "00011111", -- 2826 - 0xb0a  :   31 - 0x1f
    "00011111", -- 2827 - 0xb0b  :   31 - 0x1f
    "00011111", -- 2828 - 0xb0c  :   31 - 0x1f
    "00011111", -- 2829 - 0xb0d  :   31 - 0x1f
    "00011111", -- 2830 - 0xb0e  :   31 - 0x1f
    "00011111", -- 2831 - 0xb0f  :   31 - 0x1f
    "00000000", -- 2832 - 0xb10  :    0 - 0x0 -- Sprite 0xb1
    "11111000", -- 2833 - 0xb11  :  248 - 0xf8
    "00001000", -- 2834 - 0xb12  :    8 - 0x8
    "00001000", -- 2835 - 0xb13  :    8 - 0x8
    "00001000", -- 2836 - 0xb14  :    8 - 0x8
    "00001000", -- 2837 - 0xb15  :    8 - 0x8
    "00001000", -- 2838 - 0xb16  :    8 - 0x8
    "00001000", -- 2839 - 0xb17  :    8 - 0x8
    "00000000", -- 2840 - 0xb18  :    0 - 0x0
    "11110000", -- 2841 - 0xb19  :  240 - 0xf0
    "11110000", -- 2842 - 0xb1a  :  240 - 0xf0
    "11110000", -- 2843 - 0xb1b  :  240 - 0xf0
    "11110000", -- 2844 - 0xb1c  :  240 - 0xf0
    "11110000", -- 2845 - 0xb1d  :  240 - 0xf0
    "11110000", -- 2846 - 0xb1e  :  240 - 0xf0
    "11110000", -- 2847 - 0xb1f  :  240 - 0xf0
    "00010000", -- 2848 - 0xb20  :   16 - 0x10 -- Sprite 0xb2
    "00010000", -- 2849 - 0xb21  :   16 - 0x10
    "00010000", -- 2850 - 0xb22  :   16 - 0x10
    "00010000", -- 2851 - 0xb23  :   16 - 0x10
    "00011111", -- 2852 - 0xb24  :   31 - 0x1f
    "00011111", -- 2853 - 0xb25  :   31 - 0x1f
    "00001111", -- 2854 - 0xb26  :   15 - 0xf
    "00000000", -- 2855 - 0xb27  :    0 - 0x0
    "00011111", -- 2856 - 0xb28  :   31 - 0x1f
    "00011111", -- 2857 - 0xb29  :   31 - 0x1f
    "00011111", -- 2858 - 0xb2a  :   31 - 0x1f
    "00011111", -- 2859 - 0xb2b  :   31 - 0x1f
    "00000000", -- 2860 - 0xb2c  :    0 - 0x0
    "00000000", -- 2861 - 0xb2d  :    0 - 0x0
    "00000000", -- 2862 - 0xb2e  :    0 - 0x0
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "00001000", -- 2864 - 0xb30  :    8 - 0x8 -- Sprite 0xb3
    "00001000", -- 2865 - 0xb31  :    8 - 0x8
    "00001000", -- 2866 - 0xb32  :    8 - 0x8
    "00001000", -- 2867 - 0xb33  :    8 - 0x8
    "11111000", -- 2868 - 0xb34  :  248 - 0xf8
    "11111000", -- 2869 - 0xb35  :  248 - 0xf8
    "11110000", -- 2870 - 0xb36  :  240 - 0xf0
    "00000000", -- 2871 - 0xb37  :    0 - 0x0
    "11110000", -- 2872 - 0xb38  :  240 - 0xf0
    "11110000", -- 2873 - 0xb39  :  240 - 0xf0
    "11110000", -- 2874 - 0xb3a  :  240 - 0xf0
    "11110000", -- 2875 - 0xb3b  :  240 - 0xf0
    "00000000", -- 2876 - 0xb3c  :    0 - 0x0
    "00000000", -- 2877 - 0xb3d  :    0 - 0x0
    "00000000", -- 2878 - 0xb3e  :    0 - 0x0
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "00000000", -- 2880 - 0xb40  :    0 - 0x0 -- Sprite 0xb4
    "00000000", -- 2881 - 0xb41  :    0 - 0x0
    "00111111", -- 2882 - 0xb42  :   63 - 0x3f
    "01100000", -- 2883 - 0xb43  :   96 - 0x60
    "01100000", -- 2884 - 0xb44  :   96 - 0x60
    "01100000", -- 2885 - 0xb45  :   96 - 0x60
    "01100000", -- 2886 - 0xb46  :   96 - 0x60
    "01100000", -- 2887 - 0xb47  :   96 - 0x60
    "00000000", -- 2888 - 0xb48  :    0 - 0x0
    "00000000", -- 2889 - 0xb49  :    0 - 0x0
    "00111111", -- 2890 - 0xb4a  :   63 - 0x3f
    "01111111", -- 2891 - 0xb4b  :  127 - 0x7f
    "01111111", -- 2892 - 0xb4c  :  127 - 0x7f
    "01111111", -- 2893 - 0xb4d  :  127 - 0x7f
    "01111111", -- 2894 - 0xb4e  :  127 - 0x7f
    "01111111", -- 2895 - 0xb4f  :  127 - 0x7f
    "00000000", -- 2896 - 0xb50  :    0 - 0x0 -- Sprite 0xb5
    "00000000", -- 2897 - 0xb51  :    0 - 0x0
    "11111100", -- 2898 - 0xb52  :  252 - 0xfc
    "00000110", -- 2899 - 0xb53  :    6 - 0x6
    "00000110", -- 2900 - 0xb54  :    6 - 0x6
    "00000110", -- 2901 - 0xb55  :    6 - 0x6
    "00000110", -- 2902 - 0xb56  :    6 - 0x6
    "00000110", -- 2903 - 0xb57  :    6 - 0x6
    "00000000", -- 2904 - 0xb58  :    0 - 0x0
    "00000000", -- 2905 - 0xb59  :    0 - 0x0
    "11111000", -- 2906 - 0xb5a  :  248 - 0xf8
    "11111000", -- 2907 - 0xb5b  :  248 - 0xf8
    "11111000", -- 2908 - 0xb5c  :  248 - 0xf8
    "11111000", -- 2909 - 0xb5d  :  248 - 0xf8
    "11111000", -- 2910 - 0xb5e  :  248 - 0xf8
    "11111000", -- 2911 - 0xb5f  :  248 - 0xf8
    "01100000", -- 2912 - 0xb60  :   96 - 0x60 -- Sprite 0xb6
    "01100000", -- 2913 - 0xb61  :   96 - 0x60
    "01100000", -- 2914 - 0xb62  :   96 - 0x60
    "01111111", -- 2915 - 0xb63  :  127 - 0x7f
    "01111111", -- 2916 - 0xb64  :  127 - 0x7f
    "00111111", -- 2917 - 0xb65  :   63 - 0x3f
    "00000000", -- 2918 - 0xb66  :    0 - 0x0
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "01111111", -- 2920 - 0xb68  :  127 - 0x7f
    "01111111", -- 2921 - 0xb69  :  127 - 0x7f
    "01111111", -- 2922 - 0xb6a  :  127 - 0x7f
    "01000000", -- 2923 - 0xb6b  :   64 - 0x40
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00000110", -- 2928 - 0xb70  :    6 - 0x6 -- Sprite 0xb7
    "00000110", -- 2929 - 0xb71  :    6 - 0x6
    "00000110", -- 2930 - 0xb72  :    6 - 0x6
    "11111110", -- 2931 - 0xb73  :  254 - 0xfe
    "11111110", -- 2932 - 0xb74  :  254 - 0xfe
    "11111100", -- 2933 - 0xb75  :  252 - 0xfc
    "00000000", -- 2934 - 0xb76  :    0 - 0x0
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "11111000", -- 2936 - 0xb78  :  248 - 0xf8
    "11111000", -- 2937 - 0xb79  :  248 - 0xf8
    "11111000", -- 2938 - 0xb7a  :  248 - 0xf8
    "00000000", -- 2939 - 0xb7b  :    0 - 0x0
    "00000000", -- 2940 - 0xb7c  :    0 - 0x0
    "00000000", -- 2941 - 0xb7d  :    0 - 0x0
    "00000000", -- 2942 - 0xb7e  :    0 - 0x0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "01100000", -- 2944 - 0xb80  :   96 - 0x60 -- Sprite 0xb8
    "11110011", -- 2945 - 0xb81  :  243 - 0xf3
    "11000111", -- 2946 - 0xb82  :  199 - 0xc7
    "10000110", -- 2947 - 0xb83  :  134 - 0x86
    "00000100", -- 2948 - 0xb84  :    4 - 0x4
    "00000100", -- 2949 - 0xb85  :    4 - 0x4
    "00000111", -- 2950 - 0xb86  :    7 - 0x7
    "00000111", -- 2951 - 0xb87  :    7 - 0x7
    "00000000", -- 2952 - 0xb88  :    0 - 0x0
    "00000011", -- 2953 - 0xb89  :    3 - 0x3
    "00000111", -- 2954 - 0xb8a  :    7 - 0x7
    "00000111", -- 2955 - 0xb8b  :    7 - 0x7
    "00000111", -- 2956 - 0xb8c  :    7 - 0x7
    "00000011", -- 2957 - 0xb8d  :    3 - 0x3
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00000110", -- 2960 - 0xb90  :    6 - 0x6 -- Sprite 0xb9
    "10001111", -- 2961 - 0xb91  :  143 - 0x8f
    "11000101", -- 2962 - 0xb92  :  197 - 0xc5
    "00100011", -- 2963 - 0xb93  :   35 - 0x23
    "00101110", -- 2964 - 0xb94  :   46 - 0x2e
    "01100000", -- 2965 - 0xb95  :   96 - 0x60
    "11100001", -- 2966 - 0xb96  :  225 - 0xe1
    "11100001", -- 2967 - 0xb97  :  225 - 0xe1
    "00000000", -- 2968 - 0xb98  :    0 - 0x0
    "11000001", -- 2969 - 0xb99  :  193 - 0xc1
    "11100010", -- 2970 - 0xb9a  :  226 - 0xe2
    "11001100", -- 2971 - 0xb9b  :  204 - 0xcc
    "11000000", -- 2972 - 0xb9c  :  192 - 0xc0
    "10000000", -- 2973 - 0xb9d  :  128 - 0x80
    "00000001", -- 2974 - 0xb9e  :    1 - 0x1
    "00000010", -- 2975 - 0xb9f  :    2 - 0x2
    "11001000", -- 2976 - 0xba0  :  200 - 0xc8 -- Sprite 0xba
    "11111000", -- 2977 - 0xba1  :  248 - 0xf8
    "10110000", -- 2978 - 0xba2  :  176 - 0xb0
    "00010000", -- 2979 - 0xba3  :   16 - 0x10
    "00110000", -- 2980 - 0xba4  :   48 - 0x30
    "11001000", -- 2981 - 0xba5  :  200 - 0xc8
    "11111000", -- 2982 - 0xba6  :  248 - 0xf8
    "10000000", -- 2983 - 0xba7  :  128 - 0x80
    "11110000", -- 2984 - 0xba8  :  240 - 0xf0
    "00000000", -- 2985 - 0xba9  :    0 - 0x0
    "00100000", -- 2986 - 0xbaa  :   32 - 0x20
    "00100000", -- 2987 - 0xbab  :   32 - 0x20
    "00000000", -- 2988 - 0xbac  :    0 - 0x0
    "11110000", -- 2989 - 0xbad  :  240 - 0xf0
    "00000000", -- 2990 - 0xbae  :    0 - 0x0
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "00000011", -- 2992 - 0xbb0  :    3 - 0x3 -- Sprite 0xbb
    "00000000", -- 2993 - 0xbb1  :    0 - 0x0
    "00000000", -- 2994 - 0xbb2  :    0 - 0x0
    "01100000", -- 2995 - 0xbb3  :   96 - 0x60
    "11110000", -- 2996 - 0xbb4  :  240 - 0xf0
    "11010000", -- 2997 - 0xbb5  :  208 - 0xd0
    "10010000", -- 2998 - 0xbb6  :  144 - 0x90
    "01100000", -- 2999 - 0xbb7  :   96 - 0x60
    "00000000", -- 3000 - 0xbb8  :    0 - 0x0
    "00000000", -- 3001 - 0xbb9  :    0 - 0x0
    "00000000", -- 3002 - 0xbba  :    0 - 0x0
    "00000000", -- 3003 - 0xbbb  :    0 - 0x0
    "00000000", -- 3004 - 0xbbc  :    0 - 0x0
    "01100000", -- 3005 - 0xbbd  :   96 - 0x60
    "01100000", -- 3006 - 0xbbe  :   96 - 0x60
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "11000011", -- 3008 - 0xbc0  :  195 - 0xc3 -- Sprite 0xbc
    "00001110", -- 3009 - 0xbc1  :   14 - 0xe
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000110", -- 3011 - 0xbc3  :    6 - 0x6
    "00001111", -- 3012 - 0xbc4  :   15 - 0xf
    "00001101", -- 3013 - 0xbc5  :   13 - 0xd
    "00001001", -- 3014 - 0xbc6  :    9 - 0x9
    "00000110", -- 3015 - 0xbc7  :    6 - 0x6
    "00001100", -- 3016 - 0xbc8  :   12 - 0xc
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000110", -- 3021 - 0xbcd  :    6 - 0x6
    "00000110", -- 3022 - 0xbce  :    6 - 0x6
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "11100000", -- 3024 - 0xbd0  :  224 - 0xe0 -- Sprite 0xbd
    "01100011", -- 3025 - 0xbd1  :   99 - 0x63
    "11100111", -- 3026 - 0xbd2  :  231 - 0xe7
    "11100110", -- 3027 - 0xbd3  :  230 - 0xe6
    "00000100", -- 3028 - 0xbd4  :    4 - 0x4
    "00000100", -- 3029 - 0xbd5  :    4 - 0x4
    "00000111", -- 3030 - 0xbd6  :    7 - 0x7
    "00000111", -- 3031 - 0xbd7  :    7 - 0x7
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0
    "10000011", -- 3033 - 0xbd9  :  131 - 0x83
    "00000111", -- 3034 - 0xbda  :    7 - 0x7
    "00000111", -- 3035 - 0xbdb  :    7 - 0x7
    "00000111", -- 3036 - 0xbdc  :    7 - 0x7
    "00000011", -- 3037 - 0xbdd  :    3 - 0x3
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000111", -- 3040 - 0xbe0  :    7 - 0x7 -- Sprite 0xbe
    "10000011", -- 3041 - 0xbe1  :  131 - 0x83
    "11000111", -- 3042 - 0xbe2  :  199 - 0xc7
    "00100111", -- 3043 - 0xbe3  :   39 - 0x27
    "00100000", -- 3044 - 0xbe4  :   32 - 0x20
    "01100000", -- 3045 - 0xbe5  :   96 - 0x60
    "11100000", -- 3046 - 0xbe6  :  224 - 0xe0
    "11100000", -- 3047 - 0xbe7  :  224 - 0xe0
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0
    "11000100", -- 3049 - 0xbe9  :  196 - 0xc4
    "11100000", -- 3050 - 0xbea  :  224 - 0xe0
    "11000000", -- 3051 - 0xbeb  :  192 - 0xc0
    "11000000", -- 3052 - 0xbec  :  192 - 0xc0
    "10000000", -- 3053 - 0xbed  :  128 - 0x80
    "00000000", -- 3054 - 0xbee  :    0 - 0x0
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "00000011", -- 3056 - 0xbf0  :    3 - 0x3 -- Sprite 0xbf
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00001100", -- 3058 - 0xbf2  :   12 - 0xc
    "00001100", -- 3059 - 0xbf3  :   12 - 0xc
    "11100100", -- 3060 - 0xbf4  :  228 - 0xe4
    "01101100", -- 3061 - 0xbf5  :  108 - 0x6c
    "11101101", -- 3062 - 0xbf6  :  237 - 0xed
    "11100111", -- 3063 - 0xbf7  :  231 - 0xe7
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0
    "00000000", -- 3065 - 0xbf9  :    0 - 0x0
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00001000", -- 3068 - 0xbfc  :    8 - 0x8
    "10001000", -- 3069 - 0xbfd  :  136 - 0x88
    "00001011", -- 3070 - 0xbfe  :   11 - 0xb
    "00001000", -- 3071 - 0xbff  :    8 - 0x8
    "11000000", -- 3072 - 0xc00  :  192 - 0xc0 -- Sprite 0xc0
    "00000000", -- 3073 - 0xc01  :    0 - 0x0
    "00110000", -- 3074 - 0xc02  :   48 - 0x30
    "00110000", -- 3075 - 0xc03  :   48 - 0x30
    "00010111", -- 3076 - 0xc04  :   23 - 0x17
    "00110011", -- 3077 - 0xc05  :   51 - 0x33
    "01110111", -- 3078 - 0xc06  :  119 - 0x77
    "11010111", -- 3079 - 0xc07  :  215 - 0xd7
    "00000000", -- 3080 - 0xc08  :    0 - 0x0
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "00000000", -- 3083 - 0xc0b  :    0 - 0x0
    "00100000", -- 3084 - 0xc0c  :   32 - 0x20
    "00100100", -- 3085 - 0xc0d  :   36 - 0x24
    "10100000", -- 3086 - 0xc0e  :  160 - 0xa0
    "00100000", -- 3087 - 0xc0f  :   32 - 0x20
    "00001100", -- 3088 - 0xc10  :   12 - 0xc -- Sprite 0xc1
    "00000000", -- 3089 - 0xc11  :    0 - 0x0
    "00000000", -- 3090 - 0xc12  :    0 - 0x0
    "00000000", -- 3091 - 0xc13  :    0 - 0x0
    "00000000", -- 3092 - 0xc14  :    0 - 0x0
    "00000000", -- 3093 - 0xc15  :    0 - 0x0
    "00000000", -- 3094 - 0xc16  :    0 - 0x0
    "00000000", -- 3095 - 0xc17  :    0 - 0x0
    "00000000", -- 3096 - 0xc18  :    0 - 0x0
    "00000000", -- 3097 - 0xc19  :    0 - 0x0
    "00000000", -- 3098 - 0xc1a  :    0 - 0x0
    "00000000", -- 3099 - 0xc1b  :    0 - 0x0
    "00000000", -- 3100 - 0xc1c  :    0 - 0x0
    "00000000", -- 3101 - 0xc1d  :    0 - 0x0
    "00000000", -- 3102 - 0xc1e  :    0 - 0x0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00110000", -- 3104 - 0xc20  :   48 - 0x30 -- Sprite 0xc2
    "00000000", -- 3105 - 0xc21  :    0 - 0x0
    "00000000", -- 3106 - 0xc22  :    0 - 0x0
    "00000000", -- 3107 - 0xc23  :    0 - 0x0
    "00000000", -- 3108 - 0xc24  :    0 - 0x0
    "00000000", -- 3109 - 0xc25  :    0 - 0x0
    "00000000", -- 3110 - 0xc26  :    0 - 0x0
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "00000000", -- 3115 - 0xc2b  :    0 - 0x0
    "00000000", -- 3116 - 0xc2c  :    0 - 0x0
    "00000000", -- 3117 - 0xc2d  :    0 - 0x0
    "00000000", -- 3118 - 0xc2e  :    0 - 0x0
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "00000000", -- 3120 - 0xc30  :    0 - 0x0 -- Sprite 0xc3
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "00000100", -- 3122 - 0xc32  :    4 - 0x4
    "00001101", -- 3123 - 0xc33  :   13 - 0xd
    "00001111", -- 3124 - 0xc34  :   15 - 0xf
    "00001100", -- 3125 - 0xc35  :   12 - 0xc
    "00001100", -- 3126 - 0xc36  :   12 - 0xc
    "00000100", -- 3127 - 0xc37  :    4 - 0x4
    "00000000", -- 3128 - 0xc38  :    0 - 0x0
    "00000000", -- 3129 - 0xc39  :    0 - 0x0
    "00001000", -- 3130 - 0xc3a  :    8 - 0x8
    "00001011", -- 3131 - 0xc3b  :   11 - 0xb
    "00001000", -- 3132 - 0xc3c  :    8 - 0x8
    "00001000", -- 3133 - 0xc3d  :    8 - 0x8
    "00001000", -- 3134 - 0xc3e  :    8 - 0x8
    "00001000", -- 3135 - 0xc3f  :    8 - 0x8
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 3137 - 0xc41  :    0 - 0x0
    "00010000", -- 3138 - 0xc42  :   16 - 0x10
    "01110000", -- 3139 - 0xc43  :  112 - 0x70
    "11110000", -- 3140 - 0xc44  :  240 - 0xf0
    "00110000", -- 3141 - 0xc45  :   48 - 0x30
    "00110000", -- 3142 - 0xc46  :   48 - 0x30
    "00010000", -- 3143 - 0xc47  :   16 - 0x10
    "00000000", -- 3144 - 0xc48  :    0 - 0x0
    "00000000", -- 3145 - 0xc49  :    0 - 0x0
    "00100000", -- 3146 - 0xc4a  :   32 - 0x20
    "10100000", -- 3147 - 0xc4b  :  160 - 0xa0
    "00100000", -- 3148 - 0xc4c  :   32 - 0x20
    "00100000", -- 3149 - 0xc4d  :   32 - 0x20
    "00100000", -- 3150 - 0xc4e  :   32 - 0x20
    "00100000", -- 3151 - 0xc4f  :   32 - 0x20
    "11100100", -- 3152 - 0xc50  :  228 - 0xe4 -- Sprite 0xc5
    "00100100", -- 3153 - 0xc51  :   36 - 0x24
    "11101111", -- 3154 - 0xc52  :  239 - 0xef
    "11100111", -- 3155 - 0xc53  :  231 - 0xe7
    "00000110", -- 3156 - 0xc54  :    6 - 0x6
    "00000100", -- 3157 - 0xc55  :    4 - 0x4
    "00000100", -- 3158 - 0xc56  :    4 - 0x4
    "00000111", -- 3159 - 0xc57  :    7 - 0x7
    "00001000", -- 3160 - 0xc58  :    8 - 0x8
    "11001000", -- 3161 - 0xc59  :  200 - 0xc8
    "00000011", -- 3162 - 0xc5a  :    3 - 0x3
    "00000111", -- 3163 - 0xc5b  :    7 - 0x7
    "00000111", -- 3164 - 0xc5c  :    7 - 0x7
    "00000111", -- 3165 - 0xc5d  :    7 - 0x7
    "00000011", -- 3166 - 0xc5e  :    3 - 0x3
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "00010111", -- 3168 - 0xc60  :   23 - 0x17 -- Sprite 0xc6
    "00010001", -- 3169 - 0xc61  :   17 - 0x11
    "10110111", -- 3170 - 0xc62  :  183 - 0xb7
    "11000111", -- 3171 - 0xc63  :  199 - 0xc7
    "00100000", -- 3172 - 0xc64  :   32 - 0x20
    "00100000", -- 3173 - 0xc65  :   32 - 0x20
    "01100000", -- 3174 - 0xc66  :   96 - 0x60
    "11100000", -- 3175 - 0xc67  :  224 - 0xe0
    "00100000", -- 3176 - 0xc68  :   32 - 0x20
    "00100110", -- 3177 - 0xc69  :   38 - 0x26
    "11000000", -- 3178 - 0xc6a  :  192 - 0xc0
    "11100000", -- 3179 - 0xc6b  :  224 - 0xe0
    "11000000", -- 3180 - 0xc6c  :  192 - 0xc0
    "11000000", -- 3181 - 0xc6d  :  192 - 0xc0
    "10000000", -- 3182 - 0xc6e  :  128 - 0x80
    "00000000", -- 3183 - 0xc6f  :    0 - 0x0
    "00000111", -- 3184 - 0xc70  :    7 - 0x7 -- Sprite 0xc7
    "00000011", -- 3185 - 0xc71  :    3 - 0x3
    "00000000", -- 3186 - 0xc72  :    0 - 0x0
    "00000000", -- 3187 - 0xc73  :    0 - 0x0
    "11100000", -- 3188 - 0xc74  :  224 - 0xe0
    "00100000", -- 3189 - 0xc75  :   32 - 0x20
    "11100000", -- 3190 - 0xc76  :  224 - 0xe0
    "11100000", -- 3191 - 0xc77  :  224 - 0xe0
    "00000000", -- 3192 - 0xc78  :    0 - 0x0
    "00000000", -- 3193 - 0xc79  :    0 - 0x0
    "00000000", -- 3194 - 0xc7a  :    0 - 0x0
    "00000000", -- 3195 - 0xc7b  :    0 - 0x0
    "00000000", -- 3196 - 0xc7c  :    0 - 0x0
    "11000000", -- 3197 - 0xc7d  :  192 - 0xc0
    "00000000", -- 3198 - 0xc7e  :    0 - 0x0
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "11100000", -- 3200 - 0xc80  :  224 - 0xe0 -- Sprite 0xc8
    "11000000", -- 3201 - 0xc81  :  192 - 0xc0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000111", -- 3204 - 0xc84  :    7 - 0x7
    "00000001", -- 3205 - 0xc85  :    1 - 0x1
    "00000111", -- 3206 - 0xc86  :    7 - 0x7
    "00000111", -- 3207 - 0xc87  :    7 - 0x7
    "00000000", -- 3208 - 0xc88  :    0 - 0x0
    "00000000", -- 3209 - 0xc89  :    0 - 0x0
    "00000000", -- 3210 - 0xc8a  :    0 - 0x0
    "00000000", -- 3211 - 0xc8b  :    0 - 0x0
    "00000000", -- 3212 - 0xc8c  :    0 - 0x0
    "00000110", -- 3213 - 0xc8d  :    6 - 0x6
    "00000000", -- 3214 - 0xc8e  :    0 - 0x0
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00010011", -- 3216 - 0xc90  :   19 - 0x13 -- Sprite 0xc9
    "00011111", -- 3217 - 0xc91  :   31 - 0x1f
    "00001101", -- 3218 - 0xc92  :   13 - 0xd
    "00000100", -- 3219 - 0xc93  :    4 - 0x4
    "00001100", -- 3220 - 0xc94  :   12 - 0xc
    "00010011", -- 3221 - 0xc95  :   19 - 0x13
    "00011111", -- 3222 - 0xc96  :   31 - 0x1f
    "00000001", -- 3223 - 0xc97  :    1 - 0x1
    "00001111", -- 3224 - 0xc98  :   15 - 0xf
    "00000000", -- 3225 - 0xc99  :    0 - 0x0
    "00001000", -- 3226 - 0xc9a  :    8 - 0x8
    "00001000", -- 3227 - 0xc9b  :    8 - 0x8
    "00000000", -- 3228 - 0xc9c  :    0 - 0x0
    "00001111", -- 3229 - 0xc9d  :   15 - 0xf
    "00000000", -- 3230 - 0xc9e  :    0 - 0x0
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "01100000", -- 3232 - 0xca0  :   96 - 0x60 -- Sprite 0xca
    "11110011", -- 3233 - 0xca1  :  243 - 0xf3
    "10100111", -- 3234 - 0xca2  :  167 - 0xa7
    "11000110", -- 3235 - 0xca3  :  198 - 0xc6
    "01110100", -- 3236 - 0xca4  :  116 - 0x74
    "00000100", -- 3237 - 0xca5  :    4 - 0x4
    "10000111", -- 3238 - 0xca6  :  135 - 0x87
    "10000111", -- 3239 - 0xca7  :  135 - 0x87
    "00000000", -- 3240 - 0xca8  :    0 - 0x0
    "10000011", -- 3241 - 0xca9  :  131 - 0x83
    "01000111", -- 3242 - 0xcaa  :   71 - 0x47
    "00110111", -- 3243 - 0xcab  :   55 - 0x37
    "00000111", -- 3244 - 0xcac  :    7 - 0x7
    "00000011", -- 3245 - 0xcad  :    3 - 0x3
    "10000000", -- 3246 - 0xcae  :  128 - 0x80
    "01000000", -- 3247 - 0xcaf  :   64 - 0x40
    "00000110", -- 3248 - 0xcb0  :    6 - 0x6 -- Sprite 0xcb
    "10001111", -- 3249 - 0xcb1  :  143 - 0x8f
    "11000011", -- 3250 - 0xcb2  :  195 - 0xc3
    "00100001", -- 3251 - 0xcb3  :   33 - 0x21
    "00100000", -- 3252 - 0xcb4  :   32 - 0x20
    "01100000", -- 3253 - 0xcb5  :   96 - 0x60
    "11100000", -- 3254 - 0xcb6  :  224 - 0xe0
    "11100000", -- 3255 - 0xcb7  :  224 - 0xe0
    "00000000", -- 3256 - 0xcb8  :    0 - 0x0
    "11000000", -- 3257 - 0xcb9  :  192 - 0xc0
    "11100000", -- 3258 - 0xcba  :  224 - 0xe0
    "11000000", -- 3259 - 0xcbb  :  192 - 0xc0
    "11000000", -- 3260 - 0xcbc  :  192 - 0xc0
    "10000000", -- 3261 - 0xcbd  :  128 - 0x80
    "00000000", -- 3262 - 0xcbe  :    0 - 0x0
    "00000000", -- 3263 - 0xcbf  :    0 - 0x0
    "11000011", -- 3264 - 0xcc0  :  195 - 0xc3 -- Sprite 0xcc
    "01110000", -- 3265 - 0xcc1  :  112 - 0x70
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "01100000", -- 3267 - 0xcc3  :   96 - 0x60
    "11110000", -- 3268 - 0xcc4  :  240 - 0xf0
    "11010000", -- 3269 - 0xcc5  :  208 - 0xd0
    "10010000", -- 3270 - 0xcc6  :  144 - 0x90
    "01100000", -- 3271 - 0xcc7  :   96 - 0x60
    "00110000", -- 3272 - 0xcc8  :   48 - 0x30
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000000", -- 3274 - 0xcca  :    0 - 0x0
    "00000000", -- 3275 - 0xccb  :    0 - 0x0
    "00000000", -- 3276 - 0xccc  :    0 - 0x0
    "01100000", -- 3277 - 0xccd  :   96 - 0x60
    "01100000", -- 3278 - 0xcce  :   96 - 0x60
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "11000000", -- 3280 - 0xcd0  :  192 - 0xc0 -- Sprite 0xcd
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00000000", -- 3282 - 0xcd2  :    0 - 0x0
    "00000110", -- 3283 - 0xcd3  :    6 - 0x6
    "00001111", -- 3284 - 0xcd4  :   15 - 0xf
    "00001101", -- 3285 - 0xcd5  :   13 - 0xd
    "00001001", -- 3286 - 0xcd6  :    9 - 0x9
    "00000110", -- 3287 - 0xcd7  :    6 - 0x6
    "00000000", -- 3288 - 0xcd8  :    0 - 0x0
    "00000000", -- 3289 - 0xcd9  :    0 - 0x0
    "00000000", -- 3290 - 0xcda  :    0 - 0x0
    "00000000", -- 3291 - 0xcdb  :    0 - 0x0
    "00000000", -- 3292 - 0xcdc  :    0 - 0x0
    "00000110", -- 3293 - 0xcdd  :    6 - 0x6
    "00000110", -- 3294 - 0xcde  :    6 - 0x6
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "11111100", -- 3296 - 0xce0  :  252 - 0xfc -- Sprite 0xce
    "11000000", -- 3297 - 0xce1  :  192 - 0xc0
    "11010001", -- 3298 - 0xce2  :  209 - 0xd1
    "11000010", -- 3299 - 0xce3  :  194 - 0xc2
    "10011110", -- 3300 - 0xce4  :  158 - 0x9e
    "10111111", -- 3301 - 0xce5  :  191 - 0xbf
    "10110000", -- 3302 - 0xce6  :  176 - 0xb0
    "10110011", -- 3303 - 0xce7  :  179 - 0xb3
    "00000000", -- 3304 - 0xce8  :    0 - 0x0
    "00000001", -- 3305 - 0xce9  :    1 - 0x1
    "00011011", -- 3306 - 0xcea  :   27 - 0x1b
    "00010011", -- 3307 - 0xceb  :   19 - 0x13
    "00011111", -- 3308 - 0xcec  :   31 - 0x1f
    "00111111", -- 3309 - 0xced  :   63 - 0x3f
    "00111111", -- 3310 - 0xcee  :   63 - 0x3f
    "00111111", -- 3311 - 0xcef  :   63 - 0x3f
    "00000111", -- 3312 - 0xcf0  :    7 - 0x7 -- Sprite 0xcf
    "11110011", -- 3313 - 0xcf1  :  243 - 0xf3
    "00001011", -- 3314 - 0xcf2  :   11 - 0xb
    "01111011", -- 3315 - 0xcf3  :  123 - 0x7b
    "01111011", -- 3316 - 0xcf4  :  123 - 0x7b
    "11111001", -- 3317 - 0xcf5  :  249 - 0xf9
    "00001101", -- 3318 - 0xcf6  :   13 - 0xd
    "11101101", -- 3319 - 0xcf7  :  237 - 0xed
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0
    "11111000", -- 3321 - 0xcf9  :  248 - 0xf8
    "00001000", -- 3322 - 0xcfa  :    8 - 0x8
    "00001000", -- 3323 - 0xcfb  :    8 - 0x8
    "00001000", -- 3324 - 0xcfc  :    8 - 0x8
    "11111000", -- 3325 - 0xcfd  :  248 - 0xf8
    "11110000", -- 3326 - 0xcfe  :  240 - 0xf0
    "11010000", -- 3327 - 0xcff  :  208 - 0xd0
    "11111111", -- 3328 - 0xd00  :  255 - 0xff -- Sprite 0xd0
    "11111111", -- 3329 - 0xd01  :  255 - 0xff
    "11111111", -- 3330 - 0xd02  :  255 - 0xff
    "11111111", -- 3331 - 0xd03  :  255 - 0xff
    "11101110", -- 3332 - 0xd04  :  238 - 0xee
    "11101110", -- 3333 - 0xd05  :  238 - 0xee
    "11101110", -- 3334 - 0xd06  :  238 - 0xee
    "11101110", -- 3335 - 0xd07  :  238 - 0xee
    "00000000", -- 3336 - 0xd08  :    0 - 0x0
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "01111100", -- 3338 - 0xd0a  :  124 - 0x7c
    "11111110", -- 3339 - 0xd0b  :  254 - 0xfe
    "11101110", -- 3340 - 0xd0c  :  238 - 0xee
    "11101110", -- 3341 - 0xd0d  :  238 - 0xee
    "11101110", -- 3342 - 0xd0e  :  238 - 0xee
    "11101110", -- 3343 - 0xd0f  :  238 - 0xee
    "11111111", -- 3344 - 0xd10  :  255 - 0xff -- Sprite 0xd1
    "11111111", -- 3345 - 0xd11  :  255 - 0xff
    "11111111", -- 3346 - 0xd12  :  255 - 0xff
    "11111011", -- 3347 - 0xd13  :  251 - 0xfb
    "11111011", -- 3348 - 0xd14  :  251 - 0xfb
    "11111011", -- 3349 - 0xd15  :  251 - 0xfb
    "11111011", -- 3350 - 0xd16  :  251 - 0xfb
    "11111011", -- 3351 - 0xd17  :  251 - 0xfb
    "00000000", -- 3352 - 0xd18  :    0 - 0x0
    "00000000", -- 3353 - 0xd19  :    0 - 0x0
    "00111000", -- 3354 - 0xd1a  :   56 - 0x38
    "01111000", -- 3355 - 0xd1b  :  120 - 0x78
    "01111000", -- 3356 - 0xd1c  :  120 - 0x78
    "00111000", -- 3357 - 0xd1d  :   56 - 0x38
    "00111000", -- 3358 - 0xd1e  :   56 - 0x38
    "00111000", -- 3359 - 0xd1f  :   56 - 0x38
    "11111111", -- 3360 - 0xd20  :  255 - 0xff -- Sprite 0xd2
    "11111111", -- 3361 - 0xd21  :  255 - 0xff
    "11111111", -- 3362 - 0xd22  :  255 - 0xff
    "11111111", -- 3363 - 0xd23  :  255 - 0xff
    "11101110", -- 3364 - 0xd24  :  238 - 0xee
    "10001110", -- 3365 - 0xd25  :  142 - 0x8e
    "11111110", -- 3366 - 0xd26  :  254 - 0xfe
    "11111110", -- 3367 - 0xd27  :  254 - 0xfe
    "00000000", -- 3368 - 0xd28  :    0 - 0x0
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "01111100", -- 3370 - 0xd2a  :  124 - 0x7c
    "11111110", -- 3371 - 0xd2b  :  254 - 0xfe
    "11101110", -- 3372 - 0xd2c  :  238 - 0xee
    "00001110", -- 3373 - 0xd2d  :   14 - 0xe
    "00001110", -- 3374 - 0xd2e  :   14 - 0xe
    "01111110", -- 3375 - 0xd2f  :  126 - 0x7e
    "11111111", -- 3376 - 0xd30  :  255 - 0xff -- Sprite 0xd3
    "11111111", -- 3377 - 0xd31  :  255 - 0xff
    "11111111", -- 3378 - 0xd32  :  255 - 0xff
    "11111111", -- 3379 - 0xd33  :  255 - 0xff
    "11101110", -- 3380 - 0xd34  :  238 - 0xee
    "10001110", -- 3381 - 0xd35  :  142 - 0x8e
    "11111100", -- 3382 - 0xd36  :  252 - 0xfc
    "11111101", -- 3383 - 0xd37  :  253 - 0xfd
    "00000000", -- 3384 - 0xd38  :    0 - 0x0
    "00000000", -- 3385 - 0xd39  :    0 - 0x0
    "01111100", -- 3386 - 0xd3a  :  124 - 0x7c
    "11111110", -- 3387 - 0xd3b  :  254 - 0xfe
    "11101110", -- 3388 - 0xd3c  :  238 - 0xee
    "00001110", -- 3389 - 0xd3d  :   14 - 0xe
    "00111100", -- 3390 - 0xd3e  :   60 - 0x3c
    "00111100", -- 3391 - 0xd3f  :   60 - 0x3c
    "11111111", -- 3392 - 0xd40  :  255 - 0xff -- Sprite 0xd4
    "11111111", -- 3393 - 0xd41  :  255 - 0xff
    "11111111", -- 3394 - 0xd42  :  255 - 0xff
    "11111110", -- 3395 - 0xd43  :  254 - 0xfe
    "11101110", -- 3396 - 0xd44  :  238 - 0xee
    "11101110", -- 3397 - 0xd45  :  238 - 0xee
    "11101110", -- 3398 - 0xd46  :  238 - 0xee
    "11101110", -- 3399 - 0xd47  :  238 - 0xee
    "00000000", -- 3400 - 0xd48  :    0 - 0x0
    "00000000", -- 3401 - 0xd49  :    0 - 0x0
    "00111110", -- 3402 - 0xd4a  :   62 - 0x3e
    "01111110", -- 3403 - 0xd4b  :  126 - 0x7e
    "11101110", -- 3404 - 0xd4c  :  238 - 0xee
    "11101110", -- 3405 - 0xd4d  :  238 - 0xee
    "11101110", -- 3406 - 0xd4e  :  238 - 0xee
    "11101110", -- 3407 - 0xd4f  :  238 - 0xee
    "11111111", -- 3408 - 0xd50  :  255 - 0xff -- Sprite 0xd5
    "11111111", -- 3409 - 0xd51  :  255 - 0xff
    "11111111", -- 3410 - 0xd52  :  255 - 0xff
    "11111101", -- 3411 - 0xd53  :  253 - 0xfd
    "11100001", -- 3412 - 0xd54  :  225 - 0xe1
    "11101111", -- 3413 - 0xd55  :  239 - 0xef
    "11111111", -- 3414 - 0xd56  :  255 - 0xff
    "11111111", -- 3415 - 0xd57  :  255 - 0xff
    "00000000", -- 3416 - 0xd58  :    0 - 0x0
    "00000000", -- 3417 - 0xd59  :    0 - 0x0
    "11111100", -- 3418 - 0xd5a  :  252 - 0xfc
    "11111100", -- 3419 - 0xd5b  :  252 - 0xfc
    "11100000", -- 3420 - 0xd5c  :  224 - 0xe0
    "11100000", -- 3421 - 0xd5d  :  224 - 0xe0
    "11111100", -- 3422 - 0xd5e  :  252 - 0xfc
    "11111110", -- 3423 - 0xd5f  :  254 - 0xfe
    "11111111", -- 3424 - 0xd60  :  255 - 0xff -- Sprite 0xd6
    "11111111", -- 3425 - 0xd61  :  255 - 0xff
    "11111111", -- 3426 - 0xd62  :  255 - 0xff
    "11111101", -- 3427 - 0xd63  :  253 - 0xfd
    "11100001", -- 3428 - 0xd64  :  225 - 0xe1
    "11101111", -- 3429 - 0xd65  :  239 - 0xef
    "11111111", -- 3430 - 0xd66  :  255 - 0xff
    "11111111", -- 3431 - 0xd67  :  255 - 0xff
    "00000000", -- 3432 - 0xd68  :    0 - 0x0
    "00000000", -- 3433 - 0xd69  :    0 - 0x0
    "01111100", -- 3434 - 0xd6a  :  124 - 0x7c
    "11111100", -- 3435 - 0xd6b  :  252 - 0xfc
    "11100000", -- 3436 - 0xd6c  :  224 - 0xe0
    "11100000", -- 3437 - 0xd6d  :  224 - 0xe0
    "11111100", -- 3438 - 0xd6e  :  252 - 0xfc
    "11111110", -- 3439 - 0xd6f  :  254 - 0xfe
    "11111111", -- 3440 - 0xd70  :  255 - 0xff -- Sprite 0xd7
    "11111111", -- 3441 - 0xd71  :  255 - 0xff
    "11111111", -- 3442 - 0xd72  :  255 - 0xff
    "11111110", -- 3443 - 0xd73  :  254 - 0xfe
    "11101110", -- 3444 - 0xd74  :  238 - 0xee
    "10001110", -- 3445 - 0xd75  :  142 - 0x8e
    "11111110", -- 3446 - 0xd76  :  254 - 0xfe
    "11111100", -- 3447 - 0xd77  :  252 - 0xfc
    "00000000", -- 3448 - 0xd78  :    0 - 0x0
    "00000000", -- 3449 - 0xd79  :    0 - 0x0
    "11111110", -- 3450 - 0xd7a  :  254 - 0xfe
    "11111110", -- 3451 - 0xd7b  :  254 - 0xfe
    "11101110", -- 3452 - 0xd7c  :  238 - 0xee
    "00001110", -- 3453 - 0xd7d  :   14 - 0xe
    "00001110", -- 3454 - 0xd7e  :   14 - 0xe
    "00011100", -- 3455 - 0xd7f  :   28 - 0x1c
    "11111111", -- 3456 - 0xd80  :  255 - 0xff -- Sprite 0xd8
    "11111111", -- 3457 - 0xd81  :  255 - 0xff
    "11111111", -- 3458 - 0xd82  :  255 - 0xff
    "11111111", -- 3459 - 0xd83  :  255 - 0xff
    "11101110", -- 3460 - 0xd84  :  238 - 0xee
    "11101110", -- 3461 - 0xd85  :  238 - 0xee
    "11111100", -- 3462 - 0xd86  :  252 - 0xfc
    "11111111", -- 3463 - 0xd87  :  255 - 0xff
    "00000000", -- 3464 - 0xd88  :    0 - 0x0
    "00000000", -- 3465 - 0xd89  :    0 - 0x0
    "01111100", -- 3466 - 0xd8a  :  124 - 0x7c
    "11111110", -- 3467 - 0xd8b  :  254 - 0xfe
    "11101110", -- 3468 - 0xd8c  :  238 - 0xee
    "11101110", -- 3469 - 0xd8d  :  238 - 0xee
    "01111100", -- 3470 - 0xd8e  :  124 - 0x7c
    "11111110", -- 3471 - 0xd8f  :  254 - 0xfe
    "11111111", -- 3472 - 0xd90  :  255 - 0xff -- Sprite 0xd9
    "11111111", -- 3473 - 0xd91  :  255 - 0xff
    "11111111", -- 3474 - 0xd92  :  255 - 0xff
    "11111111", -- 3475 - 0xd93  :  255 - 0xff
    "11101110", -- 3476 - 0xd94  :  238 - 0xee
    "11101110", -- 3477 - 0xd95  :  238 - 0xee
    "11101110", -- 3478 - 0xd96  :  238 - 0xee
    "11101110", -- 3479 - 0xd97  :  238 - 0xee
    "00000000", -- 3480 - 0xd98  :    0 - 0x0
    "00000000", -- 3481 - 0xd99  :    0 - 0x0
    "01111100", -- 3482 - 0xd9a  :  124 - 0x7c
    "11111110", -- 3483 - 0xd9b  :  254 - 0xfe
    "11101110", -- 3484 - 0xd9c  :  238 - 0xee
    "11101110", -- 3485 - 0xd9d  :  238 - 0xee
    "11101110", -- 3486 - 0xd9e  :  238 - 0xee
    "11101110", -- 3487 - 0xd9f  :  238 - 0xee
    "00000000", -- 3488 - 0xda0  :    0 - 0x0 -- Sprite 0xda
    "00000000", -- 3489 - 0xda1  :    0 - 0x0
    "00000000", -- 3490 - 0xda2  :    0 - 0x0
    "10000000", -- 3491 - 0xda3  :  128 - 0x80
    "00000000", -- 3492 - 0xda4  :    0 - 0x0
    "00000000", -- 3493 - 0xda5  :    0 - 0x0
    "00000100", -- 3494 - 0xda6  :    4 - 0x4
    "00000000", -- 3495 - 0xda7  :    0 - 0x0
    "00000000", -- 3496 - 0xda8  :    0 - 0x0
    "00100000", -- 3497 - 0xda9  :   32 - 0x20
    "00000000", -- 3498 - 0xdaa  :    0 - 0x0
    "00000010", -- 3499 - 0xdab  :    2 - 0x2
    "00000000", -- 3500 - 0xdac  :    0 - 0x0
    "00100000", -- 3501 - 0xdad  :   32 - 0x20
    "00000000", -- 3502 - 0xdae  :    0 - 0x0
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00000000", -- 3504 - 0xdb0  :    0 - 0x0 -- Sprite 0xdb
    "00000100", -- 3505 - 0xdb1  :    4 - 0x4
    "00000000", -- 3506 - 0xdb2  :    0 - 0x0
    "00010001", -- 3507 - 0xdb3  :   17 - 0x11
    "00000000", -- 3508 - 0xdb4  :    0 - 0x0
    "00000000", -- 3509 - 0xdb5  :    0 - 0x0
    "00000000", -- 3510 - 0xdb6  :    0 - 0x0
    "00100000", -- 3511 - 0xdb7  :   32 - 0x20
    "00100000", -- 3512 - 0xdb8  :   32 - 0x20
    "00000000", -- 3513 - 0xdb9  :    0 - 0x0
    "00000000", -- 3514 - 0xdba  :    0 - 0x0
    "00000000", -- 3515 - 0xdbb  :    0 - 0x0
    "10000000", -- 3516 - 0xdbc  :  128 - 0x80
    "00000000", -- 3517 - 0xdbd  :    0 - 0x0
    "00000100", -- 3518 - 0xdbe  :    4 - 0x4
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0 -- Sprite 0xdc
    "00000000", -- 3521 - 0xdc1  :    0 - 0x0
    "00000000", -- 3522 - 0xdc2  :    0 - 0x0
    "00100000", -- 3523 - 0xdc3  :   32 - 0x20
    "00000000", -- 3524 - 0xdc4  :    0 - 0x0
    "00000000", -- 3525 - 0xdc5  :    0 - 0x0
    "00000000", -- 3526 - 0xdc6  :    0 - 0x0
    "00000100", -- 3527 - 0xdc7  :    4 - 0x4
    "00000000", -- 3528 - 0xdc8  :    0 - 0x0
    "00001000", -- 3529 - 0xdc9  :    8 - 0x8
    "00000000", -- 3530 - 0xdca  :    0 - 0x0
    "00000000", -- 3531 - 0xdcb  :    0 - 0x0
    "00000010", -- 3532 - 0xdcc  :    2 - 0x2
    "00000000", -- 3533 - 0xdcd  :    0 - 0x0
    "01000000", -- 3534 - 0xdce  :   64 - 0x40
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "00000000", -- 3536 - 0xdd0  :    0 - 0x0 -- Sprite 0xdd
    "00000000", -- 3537 - 0xdd1  :    0 - 0x0
    "00010001", -- 3538 - 0xdd2  :   17 - 0x11
    "00000000", -- 3539 - 0xdd3  :    0 - 0x0
    "00000000", -- 3540 - 0xdd4  :    0 - 0x0
    "10000000", -- 3541 - 0xdd5  :  128 - 0x80
    "00000000", -- 3542 - 0xdd6  :    0 - 0x0
    "00000000", -- 3543 - 0xdd7  :    0 - 0x0
    "00000000", -- 3544 - 0xdd8  :    0 - 0x0
    "01000000", -- 3545 - 0xdd9  :   64 - 0x40
    "00000000", -- 3546 - 0xdda  :    0 - 0x0
    "00000000", -- 3547 - 0xddb  :    0 - 0x0
    "00000000", -- 3548 - 0xddc  :    0 - 0x0
    "00000000", -- 3549 - 0xddd  :    0 - 0x0
    "00000010", -- 3550 - 0xdde  :    2 - 0x2
    "00100000", -- 3551 - 0xddf  :   32 - 0x20
    "10110011", -- 3552 - 0xde0  :  179 - 0xb3 -- Sprite 0xde
    "10110011", -- 3553 - 0xde1  :  179 - 0xb3
    "10110011", -- 3554 - 0xde2  :  179 - 0xb3
    "10110011", -- 3555 - 0xde3  :  179 - 0xb3
    "10110000", -- 3556 - 0xde4  :  176 - 0xb0
    "10101111", -- 3557 - 0xde5  :  175 - 0xaf
    "10011111", -- 3558 - 0xde6  :  159 - 0x9f
    "11000000", -- 3559 - 0xde7  :  192 - 0xc0
    "00111110", -- 3560 - 0xde8  :   62 - 0x3e
    "00111111", -- 3561 - 0xde9  :   63 - 0x3f
    "00111110", -- 3562 - 0xdea  :   62 - 0x3e
    "00111100", -- 3563 - 0xdeb  :   60 - 0x3c
    "00111111", -- 3564 - 0xdec  :   63 - 0x3f
    "00110000", -- 3565 - 0xded  :   48 - 0x30
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "11101101", -- 3568 - 0xdf0  :  237 - 0xed -- Sprite 0xdf
    "11001101", -- 3569 - 0xdf1  :  205 - 0xcd
    "11001101", -- 3570 - 0xdf2  :  205 - 0xcd
    "00001101", -- 3571 - 0xdf3  :   13 - 0xd
    "00001101", -- 3572 - 0xdf4  :   13 - 0xd
    "11111101", -- 3573 - 0xdf5  :  253 - 0xfd
    "11111101", -- 3574 - 0xdf6  :  253 - 0xfd
    "00000011", -- 3575 - 0xdf7  :    3 - 0x3
    "00010000", -- 3576 - 0xdf8  :   16 - 0x10
    "10110000", -- 3577 - 0xdf9  :  176 - 0xb0
    "00110000", -- 3578 - 0xdfa  :   48 - 0x30
    "11110000", -- 3579 - 0xdfb  :  240 - 0xf0
    "11110000", -- 3580 - 0xdfc  :  240 - 0xf0
    "00000000", -- 3581 - 0xdfd  :    0 - 0x0
    "00000000", -- 3582 - 0xdfe  :    0 - 0x0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "11101110", -- 3584 - 0xe00  :  238 - 0xee -- Sprite 0xe0
    "11101110", -- 3585 - 0xe01  :  238 - 0xee
    "11101110", -- 3586 - 0xe02  :  238 - 0xee
    "11101110", -- 3587 - 0xe03  :  238 - 0xee
    "11111110", -- 3588 - 0xe04  :  254 - 0xfe
    "11111100", -- 3589 - 0xe05  :  252 - 0xfc
    "11000001", -- 3590 - 0xe06  :  193 - 0xc1
    "11111111", -- 3591 - 0xe07  :  255 - 0xff
    "11101110", -- 3592 - 0xe08  :  238 - 0xee
    "11101110", -- 3593 - 0xe09  :  238 - 0xee
    "11101110", -- 3594 - 0xe0a  :  238 - 0xee
    "11101110", -- 3595 - 0xe0b  :  238 - 0xee
    "11111110", -- 3596 - 0xe0c  :  254 - 0xfe
    "01111100", -- 3597 - 0xe0d  :  124 - 0x7c
    "00000000", -- 3598 - 0xe0e  :    0 - 0x0
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "11111011", -- 3600 - 0xe10  :  251 - 0xfb -- Sprite 0xe1
    "11111011", -- 3601 - 0xe11  :  251 - 0xfb
    "11111011", -- 3602 - 0xe12  :  251 - 0xfb
    "11111011", -- 3603 - 0xe13  :  251 - 0xfb
    "11111111", -- 3604 - 0xe14  :  255 - 0xff
    "11111101", -- 3605 - 0xe15  :  253 - 0xfd
    "11000001", -- 3606 - 0xe16  :  193 - 0xc1
    "11111111", -- 3607 - 0xe17  :  255 - 0xff
    "00111000", -- 3608 - 0xe18  :   56 - 0x38
    "00111000", -- 3609 - 0xe19  :   56 - 0x38
    "00111000", -- 3610 - 0xe1a  :   56 - 0x38
    "00111000", -- 3611 - 0xe1b  :   56 - 0x38
    "01111100", -- 3612 - 0xe1c  :  124 - 0x7c
    "01111100", -- 3613 - 0xe1d  :  124 - 0x7c
    "00000000", -- 3614 - 0xe1e  :    0 - 0x0
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "11111100", -- 3616 - 0xe20  :  252 - 0xfc -- Sprite 0xe2
    "11100001", -- 3617 - 0xe21  :  225 - 0xe1
    "11101111", -- 3618 - 0xe22  :  239 - 0xef
    "11101111", -- 3619 - 0xe23  :  239 - 0xef
    "11111111", -- 3620 - 0xe24  :  255 - 0xff
    "11111110", -- 3621 - 0xe25  :  254 - 0xfe
    "10000000", -- 3622 - 0xe26  :  128 - 0x80
    "11111111", -- 3623 - 0xe27  :  255 - 0xff
    "11111100", -- 3624 - 0xe28  :  252 - 0xfc
    "11100000", -- 3625 - 0xe29  :  224 - 0xe0
    "11100000", -- 3626 - 0xe2a  :  224 - 0xe0
    "11100000", -- 3627 - 0xe2b  :  224 - 0xe0
    "11111110", -- 3628 - 0xe2c  :  254 - 0xfe
    "11111110", -- 3629 - 0xe2d  :  254 - 0xfe
    "00000000", -- 3630 - 0xe2e  :    0 - 0x0
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "11101110", -- 3632 - 0xe30  :  238 - 0xee -- Sprite 0xe3
    "11111110", -- 3633 - 0xe31  :  254 - 0xfe
    "11111110", -- 3634 - 0xe32  :  254 - 0xfe
    "11111110", -- 3635 - 0xe33  :  254 - 0xfe
    "11111110", -- 3636 - 0xe34  :  254 - 0xfe
    "11111100", -- 3637 - 0xe35  :  252 - 0xfc
    "11000001", -- 3638 - 0xe36  :  193 - 0xc1
    "11111111", -- 3639 - 0xe37  :  255 - 0xff
    "00001110", -- 3640 - 0xe38  :   14 - 0xe
    "00001110", -- 3641 - 0xe39  :   14 - 0xe
    "00001110", -- 3642 - 0xe3a  :   14 - 0xe
    "11101110", -- 3643 - 0xe3b  :  238 - 0xee
    "11111110", -- 3644 - 0xe3c  :  254 - 0xfe
    "01111100", -- 3645 - 0xe3d  :  124 - 0x7c
    "00000000", -- 3646 - 0xe3e  :    0 - 0x0
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "11101110", -- 3648 - 0xe40  :  238 - 0xee -- Sprite 0xe4
    "11101110", -- 3649 - 0xe41  :  238 - 0xee
    "11111110", -- 3650 - 0xe42  :  254 - 0xfe
    "11111110", -- 3651 - 0xe43  :  254 - 0xfe
    "10001110", -- 3652 - 0xe44  :  142 - 0x8e
    "11111110", -- 3653 - 0xe45  :  254 - 0xfe
    "11111000", -- 3654 - 0xe46  :  248 - 0xf8
    "11111111", -- 3655 - 0xe47  :  255 - 0xff
    "11101110", -- 3656 - 0xe48  :  238 - 0xee
    "11101110", -- 3657 - 0xe49  :  238 - 0xee
    "11111110", -- 3658 - 0xe4a  :  254 - 0xfe
    "11111110", -- 3659 - 0xe4b  :  254 - 0xfe
    "00001110", -- 3660 - 0xe4c  :   14 - 0xe
    "00001110", -- 3661 - 0xe4d  :   14 - 0xe
    "00000000", -- 3662 - 0xe4e  :    0 - 0x0
    "00000000", -- 3663 - 0xe4f  :    0 - 0x0
    "10001110", -- 3664 - 0xe50  :  142 - 0x8e -- Sprite 0xe5
    "11111110", -- 3665 - 0xe51  :  254 - 0xfe
    "11111110", -- 3666 - 0xe52  :  254 - 0xfe
    "11111110", -- 3667 - 0xe53  :  254 - 0xfe
    "11111110", -- 3668 - 0xe54  :  254 - 0xfe
    "11111100", -- 3669 - 0xe55  :  252 - 0xfc
    "11000001", -- 3670 - 0xe56  :  193 - 0xc1
    "11111111", -- 3671 - 0xe57  :  255 - 0xff
    "00001110", -- 3672 - 0xe58  :   14 - 0xe
    "00001110", -- 3673 - 0xe59  :   14 - 0xe
    "00001110", -- 3674 - 0xe5a  :   14 - 0xe
    "11101110", -- 3675 - 0xe5b  :  238 - 0xee
    "11111110", -- 3676 - 0xe5c  :  254 - 0xfe
    "01111100", -- 3677 - 0xe5d  :  124 - 0x7c
    "00000000", -- 3678 - 0xe5e  :    0 - 0x0
    "00000000", -- 3679 - 0xe5f  :    0 - 0x0
    "11101110", -- 3680 - 0xe60  :  238 - 0xee -- Sprite 0xe6
    "11101110", -- 3681 - 0xe61  :  238 - 0xee
    "11101110", -- 3682 - 0xe62  :  238 - 0xee
    "11101110", -- 3683 - 0xe63  :  238 - 0xee
    "11111110", -- 3684 - 0xe64  :  254 - 0xfe
    "11111100", -- 3685 - 0xe65  :  252 - 0xfc
    "11000001", -- 3686 - 0xe66  :  193 - 0xc1
    "11111111", -- 3687 - 0xe67  :  255 - 0xff
    "11101110", -- 3688 - 0xe68  :  238 - 0xee
    "11101110", -- 3689 - 0xe69  :  238 - 0xee
    "11101110", -- 3690 - 0xe6a  :  238 - 0xee
    "11101110", -- 3691 - 0xe6b  :  238 - 0xee
    "11111110", -- 3692 - 0xe6c  :  254 - 0xfe
    "01111100", -- 3693 - 0xe6d  :  124 - 0x7c
    "00000000", -- 3694 - 0xe6e  :    0 - 0x0
    "00000000", -- 3695 - 0xe6f  :    0 - 0x0
    "11111101", -- 3696 - 0xe70  :  253 - 0xfd -- Sprite 0xe7
    "11111101", -- 3697 - 0xe71  :  253 - 0xfd
    "11111001", -- 3698 - 0xe72  :  249 - 0xf9
    "11111011", -- 3699 - 0xe73  :  251 - 0xfb
    "11111011", -- 3700 - 0xe74  :  251 - 0xfb
    "11111011", -- 3701 - 0xe75  :  251 - 0xfb
    "11100011", -- 3702 - 0xe76  :  227 - 0xe3
    "11111111", -- 3703 - 0xe77  :  255 - 0xff
    "00011100", -- 3704 - 0xe78  :   28 - 0x1c
    "00011100", -- 3705 - 0xe79  :   28 - 0x1c
    "00111000", -- 3706 - 0xe7a  :   56 - 0x38
    "00111000", -- 3707 - 0xe7b  :   56 - 0x38
    "00111000", -- 3708 - 0xe7c  :   56 - 0x38
    "00111000", -- 3709 - 0xe7d  :   56 - 0x38
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "11101110", -- 3712 - 0xe80  :  238 - 0xee -- Sprite 0xe8
    "11101110", -- 3713 - 0xe81  :  238 - 0xee
    "11101110", -- 3714 - 0xe82  :  238 - 0xee
    "11101110", -- 3715 - 0xe83  :  238 - 0xee
    "11111110", -- 3716 - 0xe84  :  254 - 0xfe
    "11111100", -- 3717 - 0xe85  :  252 - 0xfc
    "11000001", -- 3718 - 0xe86  :  193 - 0xc1
    "11111111", -- 3719 - 0xe87  :  255 - 0xff
    "11101110", -- 3720 - 0xe88  :  238 - 0xee
    "11101110", -- 3721 - 0xe89  :  238 - 0xee
    "11101110", -- 3722 - 0xe8a  :  238 - 0xee
    "11101110", -- 3723 - 0xe8b  :  238 - 0xee
    "11111110", -- 3724 - 0xe8c  :  254 - 0xfe
    "01111100", -- 3725 - 0xe8d  :  124 - 0x7c
    "00000000", -- 3726 - 0xe8e  :    0 - 0x0
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "11111110", -- 3728 - 0xe90  :  254 - 0xfe -- Sprite 0xe9
    "11111110", -- 3729 - 0xe91  :  254 - 0xfe
    "11001110", -- 3730 - 0xe92  :  206 - 0xce
    "11111110", -- 3731 - 0xe93  :  254 - 0xfe
    "11111110", -- 3732 - 0xe94  :  254 - 0xfe
    "11111100", -- 3733 - 0xe95  :  252 - 0xfc
    "11000001", -- 3734 - 0xe96  :  193 - 0xc1
    "11111111", -- 3735 - 0xe97  :  255 - 0xff
    "11111110", -- 3736 - 0xe98  :  254 - 0xfe
    "01111110", -- 3737 - 0xe99  :  126 - 0x7e
    "00001110", -- 3738 - 0xe9a  :   14 - 0xe
    "00001110", -- 3739 - 0xe9b  :   14 - 0xe
    "01111110", -- 3740 - 0xe9c  :  126 - 0x7e
    "01111100", -- 3741 - 0xe9d  :  124 - 0x7c
    "00000000", -- 3742 - 0xe9e  :    0 - 0x0
    "00000000", -- 3743 - 0xe9f  :    0 - 0x0
    "00000000", -- 3744 - 0xea0  :    0 - 0x0 -- Sprite 0xea
    "01110000", -- 3745 - 0xea1  :  112 - 0x70
    "00111000", -- 3746 - 0xea2  :   56 - 0x38
    "00000000", -- 3747 - 0xea3  :    0 - 0x0
    "00000010", -- 3748 - 0xea4  :    2 - 0x2
    "00000111", -- 3749 - 0xea5  :    7 - 0x7
    "00000011", -- 3750 - 0xea6  :    3 - 0x3
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "00000000", -- 3752 - 0xea8  :    0 - 0x0
    "01110000", -- 3753 - 0xea9  :  112 - 0x70
    "00111000", -- 3754 - 0xeaa  :   56 - 0x38
    "00000000", -- 3755 - 0xeab  :    0 - 0x0
    "00000010", -- 3756 - 0xeac  :    2 - 0x2
    "00000111", -- 3757 - 0xead  :    7 - 0x7
    "00000011", -- 3758 - 0xeae  :    3 - 0x3
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0 -- Sprite 0xeb
    "00001100", -- 3761 - 0xeb1  :   12 - 0xc
    "00000110", -- 3762 - 0xeb2  :    6 - 0x6
    "00000110", -- 3763 - 0xeb3  :    6 - 0x6
    "01100000", -- 3764 - 0xeb4  :   96 - 0x60
    "01110000", -- 3765 - 0xeb5  :  112 - 0x70
    "00110000", -- 3766 - 0xeb6  :   48 - 0x30
    "00000000", -- 3767 - 0xeb7  :    0 - 0x0
    "00000000", -- 3768 - 0xeb8  :    0 - 0x0
    "00001100", -- 3769 - 0xeb9  :   12 - 0xc
    "00000110", -- 3770 - 0xeba  :    6 - 0x6
    "00000110", -- 3771 - 0xebb  :    6 - 0x6
    "01100000", -- 3772 - 0xebc  :   96 - 0x60
    "01110000", -- 3773 - 0xebd  :  112 - 0x70
    "00110000", -- 3774 - 0xebe  :   48 - 0x30
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Sprite 0xec
    "11000000", -- 3777 - 0xec1  :  192 - 0xc0
    "11100000", -- 3778 - 0xec2  :  224 - 0xe0
    "01100000", -- 3779 - 0xec3  :   96 - 0x60
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00001100", -- 3781 - 0xec5  :   12 - 0xc
    "00001110", -- 3782 - 0xec6  :   14 - 0xe
    "00000110", -- 3783 - 0xec7  :    6 - 0x6
    "00000000", -- 3784 - 0xec8  :    0 - 0x0
    "11000000", -- 3785 - 0xec9  :  192 - 0xc0
    "11100000", -- 3786 - 0xeca  :  224 - 0xe0
    "01100000", -- 3787 - 0xecb  :   96 - 0x60
    "00000000", -- 3788 - 0xecc  :    0 - 0x0
    "00001100", -- 3789 - 0xecd  :   12 - 0xc
    "00001110", -- 3790 - 0xece  :   14 - 0xe
    "00000110", -- 3791 - 0xecf  :    6 - 0x6
    "01100000", -- 3792 - 0xed0  :   96 - 0x60 -- Sprite 0xed
    "01110000", -- 3793 - 0xed1  :  112 - 0x70
    "00110000", -- 3794 - 0xed2  :   48 - 0x30
    "00000000", -- 3795 - 0xed3  :    0 - 0x0
    "00000000", -- 3796 - 0xed4  :    0 - 0x0
    "00001100", -- 3797 - 0xed5  :   12 - 0xc
    "00001110", -- 3798 - 0xed6  :   14 - 0xe
    "00000110", -- 3799 - 0xed7  :    6 - 0x6
    "01100000", -- 3800 - 0xed8  :   96 - 0x60
    "01110000", -- 3801 - 0xed9  :  112 - 0x70
    "00110000", -- 3802 - 0xeda  :   48 - 0x30
    "00000000", -- 3803 - 0xedb  :    0 - 0x0
    "00000000", -- 3804 - 0xedc  :    0 - 0x0
    "00001100", -- 3805 - 0xedd  :   12 - 0xc
    "00001110", -- 3806 - 0xede  :   14 - 0xe
    "00000110", -- 3807 - 0xedf  :    6 - 0x6
    "11111111", -- 3808 - 0xee0  :  255 - 0xff -- Sprite 0xee
    "11111111", -- 3809 - 0xee1  :  255 - 0xff
    "10111101", -- 3810 - 0xee2  :  189 - 0xbd
    "11111111", -- 3811 - 0xee3  :  255 - 0xff
    "11111111", -- 3812 - 0xee4  :  255 - 0xff
    "11111011", -- 3813 - 0xee5  :  251 - 0xfb
    "11111111", -- 3814 - 0xee6  :  255 - 0xff
    "11111111", -- 3815 - 0xee7  :  255 - 0xff
    "00000000", -- 3816 - 0xee8  :    0 - 0x0
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "01000010", -- 3818 - 0xeea  :   66 - 0x42
    "00000000", -- 3819 - 0xeeb  :    0 - 0x0
    "00000000", -- 3820 - 0xeec  :    0 - 0x0
    "00000100", -- 3821 - 0xeed  :    4 - 0x4
    "00000000", -- 3822 - 0xeee  :    0 - 0x0
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "11111111", -- 3824 - 0xef0  :  255 - 0xff -- Sprite 0xef
    "11111111", -- 3825 - 0xef1  :  255 - 0xff
    "11111011", -- 3826 - 0xef2  :  251 - 0xfb
    "11111111", -- 3827 - 0xef3  :  255 - 0xff
    "11011111", -- 3828 - 0xef4  :  223 - 0xdf
    "11111111", -- 3829 - 0xef5  :  255 - 0xff
    "11111111", -- 3830 - 0xef6  :  255 - 0xff
    "11111111", -- 3831 - 0xef7  :  255 - 0xff
    "00000000", -- 3832 - 0xef8  :    0 - 0x0
    "00000000", -- 3833 - 0xef9  :    0 - 0x0
    "00000100", -- 3834 - 0xefa  :    4 - 0x4
    "00000000", -- 3835 - 0xefb  :    0 - 0x0
    "00100000", -- 3836 - 0xefc  :   32 - 0x20
    "00000000", -- 3837 - 0xefd  :    0 - 0x0
    "00000000", -- 3838 - 0xefe  :    0 - 0x0
    "00000000", -- 3839 - 0xeff  :    0 - 0x0
    "00000000", -- 3840 - 0xf00  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 3841 - 0xf01  :    0 - 0x0
    "00000000", -- 3842 - 0xf02  :    0 - 0x0
    "00000000", -- 3843 - 0xf03  :    0 - 0x0
    "00000000", -- 3844 - 0xf04  :    0 - 0x0
    "00000000", -- 3845 - 0xf05  :    0 - 0x0
    "00000000", -- 3846 - 0xf06  :    0 - 0x0
    "00000000", -- 3847 - 0xf07  :    0 - 0x0
    "00000000", -- 3848 - 0xf08  :    0 - 0x0
    "00000000", -- 3849 - 0xf09  :    0 - 0x0
    "00000000", -- 3850 - 0xf0a  :    0 - 0x0
    "00000000", -- 3851 - 0xf0b  :    0 - 0x0
    "00000000", -- 3852 - 0xf0c  :    0 - 0x0
    "00000000", -- 3853 - 0xf0d  :    0 - 0x0
    "00000000", -- 3854 - 0xf0e  :    0 - 0x0
    "00000000", -- 3855 - 0xf0f  :    0 - 0x0
    "00000000", -- 3856 - 0xf10  :    0 - 0x0 -- Sprite 0xf1
    "10000000", -- 3857 - 0xf11  :  128 - 0x80
    "00000000", -- 3858 - 0xf12  :    0 - 0x0
    "00000000", -- 3859 - 0xf13  :    0 - 0x0
    "00000000", -- 3860 - 0xf14  :    0 - 0x0
    "00000000", -- 3861 - 0xf15  :    0 - 0x0
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "10000000", -- 3864 - 0xf18  :  128 - 0x80
    "10000000", -- 3865 - 0xf19  :  128 - 0x80
    "10000000", -- 3866 - 0xf1a  :  128 - 0x80
    "10000000", -- 3867 - 0xf1b  :  128 - 0x80
    "00000000", -- 3868 - 0xf1c  :    0 - 0x0
    "00000000", -- 3869 - 0xf1d  :    0 - 0x0
    "00000000", -- 3870 - 0xf1e  :    0 - 0x0
    "00000000", -- 3871 - 0xf1f  :    0 - 0x0
    "00000000", -- 3872 - 0xf20  :    0 - 0x0 -- Sprite 0xf2
    "11000000", -- 3873 - 0xf21  :  192 - 0xc0
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000000", -- 3876 - 0xf24  :    0 - 0x0
    "00000000", -- 3877 - 0xf25  :    0 - 0x0
    "00000000", -- 3878 - 0xf26  :    0 - 0x0
    "00000000", -- 3879 - 0xf27  :    0 - 0x0
    "11000000", -- 3880 - 0xf28  :  192 - 0xc0
    "11000000", -- 3881 - 0xf29  :  192 - 0xc0
    "11000000", -- 3882 - 0xf2a  :  192 - 0xc0
    "11000000", -- 3883 - 0xf2b  :  192 - 0xc0
    "00000000", -- 3884 - 0xf2c  :    0 - 0x0
    "00000000", -- 3885 - 0xf2d  :    0 - 0x0
    "00000000", -- 3886 - 0xf2e  :    0 - 0x0
    "00000000", -- 3887 - 0xf2f  :    0 - 0x0
    "00000000", -- 3888 - 0xf30  :    0 - 0x0 -- Sprite 0xf3
    "11100000", -- 3889 - 0xf31  :  224 - 0xe0
    "00000000", -- 3890 - 0xf32  :    0 - 0x0
    "00000000", -- 3891 - 0xf33  :    0 - 0x0
    "00000000", -- 3892 - 0xf34  :    0 - 0x0
    "00000000", -- 3893 - 0xf35  :    0 - 0x0
    "00000000", -- 3894 - 0xf36  :    0 - 0x0
    "00000000", -- 3895 - 0xf37  :    0 - 0x0
    "11100000", -- 3896 - 0xf38  :  224 - 0xe0
    "11100000", -- 3897 - 0xf39  :  224 - 0xe0
    "11100000", -- 3898 - 0xf3a  :  224 - 0xe0
    "11100000", -- 3899 - 0xf3b  :  224 - 0xe0
    "00000000", -- 3900 - 0xf3c  :    0 - 0x0
    "00000000", -- 3901 - 0xf3d  :    0 - 0x0
    "00000000", -- 3902 - 0xf3e  :    0 - 0x0
    "00000000", -- 3903 - 0xf3f  :    0 - 0x0
    "00000000", -- 3904 - 0xf40  :    0 - 0x0 -- Sprite 0xf4
    "11110000", -- 3905 - 0xf41  :  240 - 0xf0
    "00000000", -- 3906 - 0xf42  :    0 - 0x0
    "00000000", -- 3907 - 0xf43  :    0 - 0x0
    "00000000", -- 3908 - 0xf44  :    0 - 0x0
    "00000000", -- 3909 - 0xf45  :    0 - 0x0
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "00000000", -- 3911 - 0xf47  :    0 - 0x0
    "11110000", -- 3912 - 0xf48  :  240 - 0xf0
    "11110000", -- 3913 - 0xf49  :  240 - 0xf0
    "11110000", -- 3914 - 0xf4a  :  240 - 0xf0
    "11110000", -- 3915 - 0xf4b  :  240 - 0xf0
    "00000000", -- 3916 - 0xf4c  :    0 - 0x0
    "00000000", -- 3917 - 0xf4d  :    0 - 0x0
    "00000000", -- 3918 - 0xf4e  :    0 - 0x0
    "00000000", -- 3919 - 0xf4f  :    0 - 0x0
    "00000000", -- 3920 - 0xf50  :    0 - 0x0 -- Sprite 0xf5
    "11111000", -- 3921 - 0xf51  :  248 - 0xf8
    "00000000", -- 3922 - 0xf52  :    0 - 0x0
    "00000000", -- 3923 - 0xf53  :    0 - 0x0
    "00000000", -- 3924 - 0xf54  :    0 - 0x0
    "00000000", -- 3925 - 0xf55  :    0 - 0x0
    "00000000", -- 3926 - 0xf56  :    0 - 0x0
    "00000000", -- 3927 - 0xf57  :    0 - 0x0
    "11111000", -- 3928 - 0xf58  :  248 - 0xf8
    "11111000", -- 3929 - 0xf59  :  248 - 0xf8
    "11111000", -- 3930 - 0xf5a  :  248 - 0xf8
    "11111000", -- 3931 - 0xf5b  :  248 - 0xf8
    "00000000", -- 3932 - 0xf5c  :    0 - 0x0
    "00000000", -- 3933 - 0xf5d  :    0 - 0x0
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Sprite 0xf6
    "11111100", -- 3937 - 0xf61  :  252 - 0xfc
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00000000", -- 3941 - 0xf65  :    0 - 0x0
    "00000000", -- 3942 - 0xf66  :    0 - 0x0
    "00000000", -- 3943 - 0xf67  :    0 - 0x0
    "11111100", -- 3944 - 0xf68  :  252 - 0xfc
    "11111100", -- 3945 - 0xf69  :  252 - 0xfc
    "11111100", -- 3946 - 0xf6a  :  252 - 0xfc
    "11111100", -- 3947 - 0xf6b  :  252 - 0xfc
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "00000000", -- 3949 - 0xf6d  :    0 - 0x0
    "00000000", -- 3950 - 0xf6e  :    0 - 0x0
    "00000000", -- 3951 - 0xf6f  :    0 - 0x0
    "00000000", -- 3952 - 0xf70  :    0 - 0x0 -- Sprite 0xf7
    "11111110", -- 3953 - 0xf71  :  254 - 0xfe
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00000000", -- 3958 - 0xf76  :    0 - 0x0
    "00000000", -- 3959 - 0xf77  :    0 - 0x0
    "11111110", -- 3960 - 0xf78  :  254 - 0xfe
    "11111110", -- 3961 - 0xf79  :  254 - 0xfe
    "11111110", -- 3962 - 0xf7a  :  254 - 0xfe
    "11111110", -- 3963 - 0xf7b  :  254 - 0xfe
    "00000000", -- 3964 - 0xf7c  :    0 - 0x0
    "00000000", -- 3965 - 0xf7d  :    0 - 0x0
    "00000000", -- 3966 - 0xf7e  :    0 - 0x0
    "00000000", -- 3967 - 0xf7f  :    0 - 0x0
    "00000000", -- 3968 - 0xf80  :    0 - 0x0 -- Sprite 0xf8
    "11111111", -- 3969 - 0xf81  :  255 - 0xff
    "00000000", -- 3970 - 0xf82  :    0 - 0x0
    "00000000", -- 3971 - 0xf83  :    0 - 0x0
    "00000000", -- 3972 - 0xf84  :    0 - 0x0
    "00000000", -- 3973 - 0xf85  :    0 - 0x0
    "00000000", -- 3974 - 0xf86  :    0 - 0x0
    "00000000", -- 3975 - 0xf87  :    0 - 0x0
    "11111111", -- 3976 - 0xf88  :  255 - 0xff
    "11111111", -- 3977 - 0xf89  :  255 - 0xff
    "11111111", -- 3978 - 0xf8a  :  255 - 0xff
    "11111111", -- 3979 - 0xf8b  :  255 - 0xff
    "00000000", -- 3980 - 0xf8c  :    0 - 0x0
    "00000000", -- 3981 - 0xf8d  :    0 - 0x0
    "00000000", -- 3982 - 0xf8e  :    0 - 0x0
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "11111111", -- 3984 - 0xf90  :  255 - 0xff -- Sprite 0xf9
    "11111111", -- 3985 - 0xf91  :  255 - 0xff
    "11111111", -- 3986 - 0xf92  :  255 - 0xff
    "11111111", -- 3987 - 0xf93  :  255 - 0xff
    "10000000", -- 3988 - 0xf94  :  128 - 0x80
    "10000000", -- 3989 - 0xf95  :  128 - 0x80
    "11000000", -- 3990 - 0xf96  :  192 - 0xc0
    "11000000", -- 3991 - 0xf97  :  192 - 0xc0
    "00000000", -- 3992 - 0xf98  :    0 - 0x0
    "00000000", -- 3993 - 0xf99  :    0 - 0x0
    "00000000", -- 3994 - 0xf9a  :    0 - 0x0
    "00000000", -- 3995 - 0xf9b  :    0 - 0x0
    "01111111", -- 3996 - 0xf9c  :  127 - 0x7f
    "01000000", -- 3997 - 0xf9d  :   64 - 0x40
    "01000000", -- 3998 - 0xf9e  :   64 - 0x40
    "01000000", -- 3999 - 0xf9f  :   64 - 0x40
    "11111111", -- 4000 - 0xfa0  :  255 - 0xff -- Sprite 0xfa
    "11111111", -- 4001 - 0xfa1  :  255 - 0xff
    "11111111", -- 4002 - 0xfa2  :  255 - 0xff
    "11111111", -- 4003 - 0xfa3  :  255 - 0xff
    "00000000", -- 4004 - 0xfa4  :    0 - 0x0
    "00000000", -- 4005 - 0xfa5  :    0 - 0x0
    "00000000", -- 4006 - 0xfa6  :    0 - 0x0
    "00000000", -- 4007 - 0xfa7  :    0 - 0x0
    "00000000", -- 4008 - 0xfa8  :    0 - 0x0
    "00000000", -- 4009 - 0xfa9  :    0 - 0x0
    "00000000", -- 4010 - 0xfaa  :    0 - 0x0
    "00000000", -- 4011 - 0xfab  :    0 - 0x0
    "11111111", -- 4012 - 0xfac  :  255 - 0xff
    "00000000", -- 4013 - 0xfad  :    0 - 0x0
    "00000000", -- 4014 - 0xfae  :    0 - 0x0
    "00000000", -- 4015 - 0xfaf  :    0 - 0x0
    "11111111", -- 4016 - 0xfb0  :  255 - 0xff -- Sprite 0xfb
    "11111111", -- 4017 - 0xfb1  :  255 - 0xff
    "11111111", -- 4018 - 0xfb2  :  255 - 0xff
    "11111111", -- 4019 - 0xfb3  :  255 - 0xff
    "00000001", -- 4020 - 0xfb4  :    1 - 0x1
    "00000000", -- 4021 - 0xfb5  :    0 - 0x0
    "00000010", -- 4022 - 0xfb6  :    2 - 0x2
    "00000010", -- 4023 - 0xfb7  :    2 - 0x2
    "00000000", -- 4024 - 0xfb8  :    0 - 0x0
    "00000000", -- 4025 - 0xfb9  :    0 - 0x0
    "00000000", -- 4026 - 0xfba  :    0 - 0x0
    "00000000", -- 4027 - 0xfbb  :    0 - 0x0
    "11111110", -- 4028 - 0xfbc  :  254 - 0xfe
    "00000010", -- 4029 - 0xfbd  :    2 - 0x2
    "00000010", -- 4030 - 0xfbe  :    2 - 0x2
    "00000010", -- 4031 - 0xfbf  :    2 - 0x2
    "11000000", -- 4032 - 0xfc0  :  192 - 0xc0 -- Sprite 0xfc
    "11000000", -- 4033 - 0xfc1  :  192 - 0xc0
    "10000000", -- 4034 - 0xfc2  :  128 - 0x80
    "10000000", -- 4035 - 0xfc3  :  128 - 0x80
    "11000000", -- 4036 - 0xfc4  :  192 - 0xc0
    "11111111", -- 4037 - 0xfc5  :  255 - 0xff
    "11111111", -- 4038 - 0xfc6  :  255 - 0xff
    "11111111", -- 4039 - 0xfc7  :  255 - 0xff
    "01000000", -- 4040 - 0xfc8  :   64 - 0x40
    "01000000", -- 4041 - 0xfc9  :   64 - 0x40
    "01000000", -- 4042 - 0xfca  :   64 - 0x40
    "01111111", -- 4043 - 0xfcb  :  127 - 0x7f
    "00000000", -- 4044 - 0xfcc  :    0 - 0x0
    "00000000", -- 4045 - 0xfcd  :    0 - 0x0
    "00000000", -- 4046 - 0xfce  :    0 - 0x0
    "00000000", -- 4047 - 0xfcf  :    0 - 0x0
    "00000000", -- 4048 - 0xfd0  :    0 - 0x0 -- Sprite 0xfd
    "00000000", -- 4049 - 0xfd1  :    0 - 0x0
    "00000000", -- 4050 - 0xfd2  :    0 - 0x0
    "00000000", -- 4051 - 0xfd3  :    0 - 0x0
    "00000000", -- 4052 - 0xfd4  :    0 - 0x0
    "11111111", -- 4053 - 0xfd5  :  255 - 0xff
    "11111111", -- 4054 - 0xfd6  :  255 - 0xff
    "11111111", -- 4055 - 0xfd7  :  255 - 0xff
    "00000000", -- 4056 - 0xfd8  :    0 - 0x0
    "00000000", -- 4057 - 0xfd9  :    0 - 0x0
    "00000000", -- 4058 - 0xfda  :    0 - 0x0
    "11111111", -- 4059 - 0xfdb  :  255 - 0xff
    "00000000", -- 4060 - 0xfdc  :    0 - 0x0
    "00000000", -- 4061 - 0xfdd  :    0 - 0x0
    "00000000", -- 4062 - 0xfde  :    0 - 0x0
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00000010", -- 4064 - 0xfe0  :    2 - 0x2 -- Sprite 0xfe
    "00000010", -- 4065 - 0xfe1  :    2 - 0x2
    "00000000", -- 4066 - 0xfe2  :    0 - 0x0
    "00000000", -- 4067 - 0xfe3  :    0 - 0x0
    "00000000", -- 4068 - 0xfe4  :    0 - 0x0
    "11111111", -- 4069 - 0xfe5  :  255 - 0xff
    "11111111", -- 4070 - 0xfe6  :  255 - 0xff
    "11111111", -- 4071 - 0xfe7  :  255 - 0xff
    "00000010", -- 4072 - 0xfe8  :    2 - 0x2
    "00000010", -- 4073 - 0xfe9  :    2 - 0x2
    "00000010", -- 4074 - 0xfea  :    2 - 0x2
    "11111110", -- 4075 - 0xfeb  :  254 - 0xfe
    "00000000", -- 4076 - 0xfec  :    0 - 0x0
    "00000000", -- 4077 - 0xfed  :    0 - 0x0
    "00000000", -- 4078 - 0xfee  :    0 - 0x0
    "00000000", -- 4079 - 0xfef  :    0 - 0x0
    "11111111", -- 4080 - 0xff0  :  255 - 0xff -- Sprite 0xff
    "11111111", -- 4081 - 0xff1  :  255 - 0xff
    "11111111", -- 4082 - 0xff2  :  255 - 0xff
    "11111111", -- 4083 - 0xff3  :  255 - 0xff
    "11111111", -- 4084 - 0xff4  :  255 - 0xff
    "11111111", -- 4085 - 0xff5  :  255 - 0xff
    "11111111", -- 4086 - 0xff6  :  255 - 0xff
    "11111111", -- 4087 - 0xff7  :  255 - 0xff
    "00000000", -- 4088 - 0xff8  :    0 - 0x0
    "00000000", -- 4089 - 0xff9  :    0 - 0x0
    "00000000", -- 4090 - 0xffa  :    0 - 0x0
    "00000000", -- 4091 - 0xffb  :    0 - 0x0
    "00000000", -- 4092 - 0xffc  :    0 - 0x0
    "00000000", -- 4093 - 0xffd  :    0 - 0x0
    "00000000", -- 4094 - 0xffe  :    0 - 0x0
    "00000000", -- 4095 - 0xfff  :    0 - 0x0
          -- Pattern Table 1---------
    "00000000", -- 4096 - 0x1000  :    0 - 0x0 -- Background 0x0
    "00000000", -- 4097 - 0x1001  :    0 - 0x0
    "00000000", -- 4098 - 0x1002  :    0 - 0x0
    "00000000", -- 4099 - 0x1003  :    0 - 0x0
    "00000000", -- 4100 - 0x1004  :    0 - 0x0
    "00000000", -- 4101 - 0x1005  :    0 - 0x0
    "00000000", -- 4102 - 0x1006  :    0 - 0x0
    "00000000", -- 4103 - 0x1007  :    0 - 0x0
    "00000101", -- 4104 - 0x1008  :    5 - 0x5
    "01010101", -- 4105 - 0x1009  :   85 - 0x55
    "01010101", -- 4106 - 0x100a  :   85 - 0x55
    "01010000", -- 4107 - 0x100b  :   80 - 0x50
    "00000000", -- 4108 - 0x100c  :    0 - 0x0
    "00000000", -- 4109 - 0x100d  :    0 - 0x0
    "00000000", -- 4110 - 0x100e  :    0 - 0x0
    "00000000", -- 4111 - 0x100f  :    0 - 0x0
    "00000101", -- 4112 - 0x1010  :    5 - 0x5 -- Background 0x1
    "01010101", -- 4113 - 0x1011  :   85 - 0x55
    "01010101", -- 4114 - 0x1012  :   85 - 0x55
    "01010000", -- 4115 - 0x1013  :   80 - 0x50
    "00000000", -- 4116 - 0x1014  :    0 - 0x0
    "00000000", -- 4117 - 0x1015  :    0 - 0x0
    "00000000", -- 4118 - 0x1016  :    0 - 0x0
    "00000000", -- 4119 - 0x1017  :    0 - 0x0
    "00000101", -- 4120 - 0x1018  :    5 - 0x5
    "01010101", -- 4121 - 0x1019  :   85 - 0x55
    "01010101", -- 4122 - 0x101a  :   85 - 0x55
    "01010000", -- 4123 - 0x101b  :   80 - 0x50
    "00000000", -- 4124 - 0x101c  :    0 - 0x0
    "00000000", -- 4125 - 0x101d  :    0 - 0x0
    "00000000", -- 4126 - 0x101e  :    0 - 0x0
    "00000000", -- 4127 - 0x101f  :    0 - 0x0
    "00000101", -- 4128 - 0x1020  :    5 - 0x5 -- Background 0x2
    "01010000", -- 4129 - 0x1021  :   80 - 0x50
    "00000101", -- 4130 - 0x1022  :    5 - 0x5
    "01010000", -- 4131 - 0x1023  :   80 - 0x50
    "00000000", -- 4132 - 0x1024  :    0 - 0x0
    "00000000", -- 4133 - 0x1025  :    0 - 0x0
    "00000000", -- 4134 - 0x1026  :    0 - 0x0
    "00000000", -- 4135 - 0x1027  :    0 - 0x0
    "00000101", -- 4136 - 0x1028  :    5 - 0x5
    "01010000", -- 4137 - 0x1029  :   80 - 0x50
    "00000101", -- 4138 - 0x102a  :    5 - 0x5
    "01010000", -- 4139 - 0x102b  :   80 - 0x50
    "00000000", -- 4140 - 0x102c  :    0 - 0x0
    "00000000", -- 4141 - 0x102d  :    0 - 0x0
    "00000000", -- 4142 - 0x102e  :    0 - 0x0
    "00000000", -- 4143 - 0x102f  :    0 - 0x0
    "00000101", -- 4144 - 0x1030  :    5 - 0x5 -- Background 0x3
    "01010000", -- 4145 - 0x1031  :   80 - 0x50
    "00000101", -- 4146 - 0x1032  :    5 - 0x5
    "01010000", -- 4147 - 0x1033  :   80 - 0x50
    "00000000", -- 4148 - 0x1034  :    0 - 0x0
    "00000000", -- 4149 - 0x1035  :    0 - 0x0
    "00000000", -- 4150 - 0x1036  :    0 - 0x0
    "00000000", -- 4151 - 0x1037  :    0 - 0x0
    "00000101", -- 4152 - 0x1038  :    5 - 0x5
    "01010101", -- 4153 - 0x1039  :   85 - 0x55
    "01010101", -- 4154 - 0x103a  :   85 - 0x55
    "01010000", -- 4155 - 0x103b  :   80 - 0x50
    "00000000", -- 4156 - 0x103c  :    0 - 0x0
    "00000000", -- 4157 - 0x103d  :    0 - 0x0
    "00000000", -- 4158 - 0x103e  :    0 - 0x0
    "00000000", -- 4159 - 0x103f  :    0 - 0x0
    "00000101", -- 4160 - 0x1040  :    5 - 0x5 -- Background 0x4
    "01010101", -- 4161 - 0x1041  :   85 - 0x55
    "01010101", -- 4162 - 0x1042  :   85 - 0x55
    "01010000", -- 4163 - 0x1043  :   80 - 0x50
    "00000000", -- 4164 - 0x1044  :    0 - 0x0
    "00000000", -- 4165 - 0x1045  :    0 - 0x0
    "00000000", -- 4166 - 0x1046  :    0 - 0x0
    "00000000", -- 4167 - 0x1047  :    0 - 0x0
    "00000101", -- 4168 - 0x1048  :    5 - 0x5
    "01010101", -- 4169 - 0x1049  :   85 - 0x55
    "01010101", -- 4170 - 0x104a  :   85 - 0x55
    "01010000", -- 4171 - 0x104b  :   80 - 0x50
    "00000000", -- 4172 - 0x104c  :    0 - 0x0
    "00000000", -- 4173 - 0x104d  :    0 - 0x0
    "00000000", -- 4174 - 0x104e  :    0 - 0x0
    "00000000", -- 4175 - 0x104f  :    0 - 0x0
    "00000000", -- 4176 - 0x1050  :    0 - 0x0 -- Background 0x5
    "00000000", -- 4177 - 0x1051  :    0 - 0x0
    "00000000", -- 4178 - 0x1052  :    0 - 0x0
    "00000000", -- 4179 - 0x1053  :    0 - 0x0
    "00000000", -- 4180 - 0x1054  :    0 - 0x0
    "00000000", -- 4181 - 0x1055  :    0 - 0x0
    "00000000", -- 4182 - 0x1056  :    0 - 0x0
    "00000000", -- 4183 - 0x1057  :    0 - 0x0
    "00001110", -- 4184 - 0x1058  :   14 - 0xe
    "00000111", -- 4185 - 0x1059  :    7 - 0x7
    "00001000", -- 4186 - 0x105a  :    8 - 0x8
    "01100000", -- 4187 - 0x105b  :   96 - 0x60
    "00000000", -- 4188 - 0x105c  :    0 - 0x0
    "00001010", -- 4189 - 0x105d  :   10 - 0xa
    "00000001", -- 4190 - 0x105e  :    1 - 0x1
    "00010101", -- 4191 - 0x105f  :   21 - 0x15
    "01010101", -- 4192 - 0x1060  :   85 - 0x55 -- Background 0x6
    "01010101", -- 4193 - 0x1061  :   85 - 0x55
    "01010100", -- 4194 - 0x1062  :   84 - 0x54
    "00000000", -- 4195 - 0x1063  :    0 - 0x0
    "00000000", -- 4196 - 0x1064  :    0 - 0x0
    "00000000", -- 4197 - 0x1065  :    0 - 0x0
    "00000000", -- 4198 - 0x1066  :    0 - 0x0
    "00010101", -- 4199 - 0x1067  :   21 - 0x15
    "01010101", -- 4200 - 0x1068  :   85 - 0x55
    "01010101", -- 4201 - 0x1069  :   85 - 0x55
    "01010100", -- 4202 - 0x106a  :   84 - 0x54
    "00000000", -- 4203 - 0x106b  :    0 - 0x0
    "00000000", -- 4204 - 0x106c  :    0 - 0x0
    "00000000", -- 4205 - 0x106d  :    0 - 0x0
    "00000000", -- 4206 - 0x106e  :    0 - 0x0
    "00010110", -- 4207 - 0x106f  :   22 - 0x16
    "10101010", -- 4208 - 0x1070  :  170 - 0xaa -- Background 0x7
    "10011010", -- 4209 - 0x1071  :  154 - 0x9a
    "10010100", -- 4210 - 0x1072  :  148 - 0x94
    "00000000", -- 4211 - 0x1073  :    0 - 0x0
    "00000000", -- 4212 - 0x1074  :    0 - 0x0
    "00000000", -- 4213 - 0x1075  :    0 - 0x0
    "00000000", -- 4214 - 0x1076  :    0 - 0x0
    "00010110", -- 4215 - 0x1077  :   22 - 0x16
    "01010101", -- 4216 - 0x1078  :   85 - 0x55
    "01010101", -- 4217 - 0x1079  :   85 - 0x55
    "10010100", -- 4218 - 0x107a  :  148 - 0x94
    "00000000", -- 4219 - 0x107b  :    0 - 0x0
    "00000000", -- 4220 - 0x107c  :    0 - 0x0
    "00000000", -- 4221 - 0x107d  :    0 - 0x0
    "00000000", -- 4222 - 0x107e  :    0 - 0x0
    "00010110", -- 4223 - 0x107f  :   22 - 0x16
    "01010000", -- 4224 - 0x1080  :   80 - 0x50 -- Background 0x8
    "00000101", -- 4225 - 0x1081  :    5 - 0x5
    "10010100", -- 4226 - 0x1082  :  148 - 0x94
    "00000000", -- 4227 - 0x1083  :    0 - 0x0
    "00000000", -- 4228 - 0x1084  :    0 - 0x0
    "00000000", -- 4229 - 0x1085  :    0 - 0x0
    "00000000", -- 4230 - 0x1086  :    0 - 0x0
    "00010101", -- 4231 - 0x1087  :   21 - 0x15
    "01010000", -- 4232 - 0x1088  :   80 - 0x50
    "00000101", -- 4233 - 0x1089  :    5 - 0x5
    "01010100", -- 4234 - 0x108a  :   84 - 0x54
    "00000000", -- 4235 - 0x108b  :    0 - 0x0
    "00000000", -- 4236 - 0x108c  :    0 - 0x0
    "00000000", -- 4237 - 0x108d  :    0 - 0x0
    "00000000", -- 4238 - 0x108e  :    0 - 0x0
    "00010110", -- 4239 - 0x108f  :   22 - 0x16
    "01010000", -- 4240 - 0x1090  :   80 - 0x50 -- Background 0x9
    "00000101", -- 4241 - 0x1091  :    5 - 0x5
    "10010100", -- 4242 - 0x1092  :  148 - 0x94
    "00000000", -- 4243 - 0x1093  :    0 - 0x0
    "00000000", -- 4244 - 0x1094  :    0 - 0x0
    "00000000", -- 4245 - 0x1095  :    0 - 0x0
    "00000000", -- 4246 - 0x1096  :    0 - 0x0
    "00010110", -- 4247 - 0x1097  :   22 - 0x16
    "01010101", -- 4248 - 0x1098  :   85 - 0x55
    "01010101", -- 4249 - 0x1099  :   85 - 0x55
    "10010100", -- 4250 - 0x109a  :  148 - 0x94
    "00000000", -- 4251 - 0x109b  :    0 - 0x0
    "00000000", -- 4252 - 0x109c  :    0 - 0x0
    "00000000", -- 4253 - 0x109d  :    0 - 0x0
    "00000000", -- 4254 - 0x109e  :    0 - 0x0
    "00010110", -- 4255 - 0x109f  :   22 - 0x16
    "10100110", -- 4256 - 0x10a0  :  166 - 0xa6 -- Background 0xa
    "10101010", -- 4257 - 0x10a1  :  170 - 0xaa
    "10010100", -- 4258 - 0x10a2  :  148 - 0x94
    "00000000", -- 4259 - 0x10a3  :    0 - 0x0
    "00000000", -- 4260 - 0x10a4  :    0 - 0x0
    "00000000", -- 4261 - 0x10a5  :    0 - 0x0
    "00000000", -- 4262 - 0x10a6  :    0 - 0x0
    "00010101", -- 4263 - 0x10a7  :   21 - 0x15
    "01010101", -- 4264 - 0x10a8  :   85 - 0x55
    "01010101", -- 4265 - 0x10a9  :   85 - 0x55
    "01010100", -- 4266 - 0x10aa  :   84 - 0x54
    "00000000", -- 4267 - 0x10ab  :    0 - 0x0
    "00000000", -- 4268 - 0x10ac  :    0 - 0x0
    "00000000", -- 4269 - 0x10ad  :    0 - 0x0
    "00000000", -- 4270 - 0x10ae  :    0 - 0x0
    "00010101", -- 4271 - 0x10af  :   21 - 0x15
    "01010101", -- 4272 - 0x10b0  :   85 - 0x55 -- Background 0xb
    "01010101", -- 4273 - 0x10b1  :   85 - 0x55
    "01010100", -- 4274 - 0x10b2  :   84 - 0x54
    "00000000", -- 4275 - 0x10b3  :    0 - 0x0
    "00000000", -- 4276 - 0x10b4  :    0 - 0x0
    "00000000", -- 4277 - 0x10b5  :    0 - 0x0
    "00000000", -- 4278 - 0x10b6  :    0 - 0x0
    "00001110", -- 4279 - 0x10b7  :   14 - 0xe
    "00000111", -- 4280 - 0x10b8  :    7 - 0x7
    "00001000", -- 4281 - 0x10b9  :    8 - 0x8
    "01110100", -- 4282 - 0x10ba  :  116 - 0x74
    "00000000", -- 4283 - 0x10bb  :    0 - 0x0
    "11011100", -- 4284 - 0x10bc  :  220 - 0xdc
    "00000000", -- 4285 - 0x10bd  :    0 - 0x0
    "00010101", -- 4286 - 0x10be  :   21 - 0x15
    "01010101", -- 4287 - 0x10bf  :   85 - 0x55
    "01010101", -- 4288 - 0x10c0  :   85 - 0x55 -- Background 0xc
    "01010100", -- 4289 - 0x10c1  :   84 - 0x54
    "00000000", -- 4290 - 0x10c2  :    0 - 0x0
    "00000000", -- 4291 - 0x10c3  :    0 - 0x0
    "00000000", -- 4292 - 0x10c4  :    0 - 0x0
    "00000000", -- 4293 - 0x10c5  :    0 - 0x0
    "00011010", -- 4294 - 0x10c6  :   26 - 0x1a
    "10011101", -- 4295 - 0x10c7  :  157 - 0x9d
    "01110110", -- 4296 - 0x10c8  :  118 - 0x76
    "10100100", -- 4297 - 0x10c9  :  164 - 0xa4
    "00000000", -- 4298 - 0x10ca  :    0 - 0x0
    "00000000", -- 4299 - 0x10cb  :    0 - 0x0
    "00000000", -- 4300 - 0x10cc  :    0 - 0x0
    "00000000", -- 4301 - 0x10cd  :    0 - 0x0
    "00010101", -- 4302 - 0x10ce  :   21 - 0x15
    "01010101", -- 4303 - 0x10cf  :   85 - 0x55
    "01010101", -- 4304 - 0x10d0  :   85 - 0x55 -- Background 0xd
    "01010100", -- 4305 - 0x10d1  :   84 - 0x54
    "00000000", -- 4306 - 0x10d2  :    0 - 0x0
    "00000000", -- 4307 - 0x10d3  :    0 - 0x0
    "00000000", -- 4308 - 0x10d4  :    0 - 0x0
    "00000000", -- 4309 - 0x10d5  :    0 - 0x0
    "00010111", -- 4310 - 0x10d6  :   23 - 0x17
    "01010101", -- 4311 - 0x10d7  :   85 - 0x55
    "01010101", -- 4312 - 0x10d8  :   85 - 0x55
    "11010100", -- 4313 - 0x10d9  :  212 - 0xd4
    "00000000", -- 4314 - 0x10da  :    0 - 0x0
    "00000000", -- 4315 - 0x10db  :    0 - 0x0
    "00000000", -- 4316 - 0x10dc  :    0 - 0x0
    "00000000", -- 4317 - 0x10dd  :    0 - 0x0
    "00010101", -- 4318 - 0x10de  :   21 - 0x15
    "01010000", -- 4319 - 0x10df  :   80 - 0x50
    "00000101", -- 4320 - 0x10e0  :    5 - 0x5 -- Background 0xe
    "01010100", -- 4321 - 0x10e1  :   84 - 0x54
    "00000000", -- 4322 - 0x10e2  :    0 - 0x0
    "00000000", -- 4323 - 0x10e3  :    0 - 0x0
    "00000000", -- 4324 - 0x10e4  :    0 - 0x0
    "00000000", -- 4325 - 0x10e5  :    0 - 0x0
    "00010101", -- 4326 - 0x10e6  :   21 - 0x15
    "01010000", -- 4327 - 0x10e7  :   80 - 0x50
    "00000101", -- 4328 - 0x10e8  :    5 - 0x5
    "01010100", -- 4329 - 0x10e9  :   84 - 0x54
    "00000000", -- 4330 - 0x10ea  :    0 - 0x0
    "00000000", -- 4331 - 0x10eb  :    0 - 0x0
    "00000000", -- 4332 - 0x10ec  :    0 - 0x0
    "00000000", -- 4333 - 0x10ed  :    0 - 0x0
    "00010101", -- 4334 - 0x10ee  :   21 - 0x15
    "01010000", -- 4335 - 0x10ef  :   80 - 0x50
    "00000101", -- 4336 - 0x10f0  :    5 - 0x5 -- Background 0xf
    "01010100", -- 4337 - 0x10f1  :   84 - 0x54
    "00000000", -- 4338 - 0x10f2  :    0 - 0x0
    "00000000", -- 4339 - 0x10f3  :    0 - 0x0
    "00000000", -- 4340 - 0x10f4  :    0 - 0x0
    "00000000", -- 4341 - 0x10f5  :    0 - 0x0
    "00010111", -- 4342 - 0x10f6  :   23 - 0x17
    "01010101", -- 4343 - 0x10f7  :   85 - 0x55
    "01010101", -- 4344 - 0x10f8  :   85 - 0x55
    "11010100", -- 4345 - 0x10f9  :  212 - 0xd4
    "00000000", -- 4346 - 0x10fa  :    0 - 0x0
    "00000000", -- 4347 - 0x10fb  :    0 - 0x0
    "00000000", -- 4348 - 0x10fc  :    0 - 0x0
    "00000000", -- 4349 - 0x10fd  :    0 - 0x0
    "00010101", -- 4350 - 0x10fe  :   21 - 0x15
    "01010101", -- 4351 - 0x10ff  :   85 - 0x55
    "01010101", -- 4352 - 0x1100  :   85 - 0x55 -- Background 0x10
    "01010100", -- 4353 - 0x1101  :   84 - 0x54
    "00000000", -- 4354 - 0x1102  :    0 - 0x0
    "00000000", -- 4355 - 0x1103  :    0 - 0x0
    "00000000", -- 4356 - 0x1104  :    0 - 0x0
    "00000000", -- 4357 - 0x1105  :    0 - 0x0
    "00011010", -- 4358 - 0x1106  :   26 - 0x1a
    "10011101", -- 4359 - 0x1107  :  157 - 0x9d
    "01110110", -- 4360 - 0x1108  :  118 - 0x76
    "10100100", -- 4361 - 0x1109  :  164 - 0xa4
    "00000000", -- 4362 - 0x110a  :    0 - 0x0
    "00000000", -- 4363 - 0x110b  :    0 - 0x0
    "00000000", -- 4364 - 0x110c  :    0 - 0x0
    "00000000", -- 4365 - 0x110d  :    0 - 0x0
    "00010101", -- 4366 - 0x110e  :   21 - 0x15
    "01010101", -- 4367 - 0x110f  :   85 - 0x55
    "01010101", -- 4368 - 0x1110  :   85 - 0x55 -- Background 0x11
    "01010100", -- 4369 - 0x1111  :   84 - 0x54
    "00000000", -- 4370 - 0x1112  :    0 - 0x0
    "00000000", -- 4371 - 0x1113  :    0 - 0x0
    "00000000", -- 4372 - 0x1114  :    0 - 0x0
    "00000000", -- 4373 - 0x1115  :    0 - 0x0
    "00001110", -- 4374 - 0x1116  :   14 - 0xe
    "00000111", -- 4375 - 0x1117  :    7 - 0x7
    "00001000", -- 4376 - 0x1118  :    8 - 0x8
    "01111010", -- 4377 - 0x1119  :  122 - 0x7a
    "00000000", -- 4378 - 0x111a  :    0 - 0x0
    "11010001", -- 4379 - 0x111b  :  209 - 0xd1
    "00000000", -- 4380 - 0x111c  :    0 - 0x0
    "00010101", -- 4381 - 0x111d  :   21 - 0x15
    "01010101", -- 4382 - 0x111e  :   85 - 0x55
    "01010101", -- 4383 - 0x111f  :   85 - 0x55
    "01010101", -- 4384 - 0x1120  :   85 - 0x55 -- Background 0x12
    "01010101", -- 4385 - 0x1121  :   85 - 0x55
    "01000000", -- 4386 - 0x1122  :   64 - 0x40
    "00000000", -- 4387 - 0x1123  :    0 - 0x0
    "00000000", -- 4388 - 0x1124  :    0 - 0x0
    "00010101", -- 4389 - 0x1125  :   21 - 0x15
    "01010101", -- 4390 - 0x1126  :   85 - 0x55
    "01010101", -- 4391 - 0x1127  :   85 - 0x55
    "01010101", -- 4392 - 0x1128  :   85 - 0x55
    "01010101", -- 4393 - 0x1129  :   85 - 0x55
    "01000000", -- 4394 - 0x112a  :   64 - 0x40
    "00000000", -- 4395 - 0x112b  :    0 - 0x0
    "00000000", -- 4396 - 0x112c  :    0 - 0x0
    "00010110", -- 4397 - 0x112d  :   22 - 0x16
    "10100101", -- 4398 - 0x112e  :  165 - 0xa5
    "01010101", -- 4399 - 0x112f  :   85 - 0x55
    "01010101", -- 4400 - 0x1130  :   85 - 0x55 -- Background 0x13
    "10101001", -- 4401 - 0x1131  :  169 - 0xa9
    "01000000", -- 4402 - 0x1132  :   64 - 0x40
    "00000000", -- 4403 - 0x1133  :    0 - 0x0
    "00000000", -- 4404 - 0x1134  :    0 - 0x0
    "00010110", -- 4405 - 0x1135  :   22 - 0x16
    "01010101", -- 4406 - 0x1136  :   85 - 0x55
    "01101010", -- 4407 - 0x1137  :  106 - 0x6a
    "10010101", -- 4408 - 0x1138  :  149 - 0x95
    "01011001", -- 4409 - 0x1139  :   89 - 0x59
    "01000000", -- 4410 - 0x113a  :   64 - 0x40
    "00000000", -- 4411 - 0x113b  :    0 - 0x0
    "00000000", -- 4412 - 0x113c  :    0 - 0x0
    "00010110", -- 4413 - 0x113d  :   22 - 0x16
    "01000000", -- 4414 - 0x113e  :   64 - 0x40
    "01010101", -- 4415 - 0x113f  :   85 - 0x55
    "01010101", -- 4416 - 0x1140  :   85 - 0x55 -- Background 0x14
    "01011001", -- 4417 - 0x1141  :   89 - 0x59
    "01000000", -- 4418 - 0x1142  :   64 - 0x40
    "00000000", -- 4419 - 0x1143  :    0 - 0x0
    "00000000", -- 4420 - 0x1144  :    0 - 0x0
    "00010101", -- 4421 - 0x1145  :   21 - 0x15
    "01000000", -- 4422 - 0x1146  :   64 - 0x40
    "01010101", -- 4423 - 0x1147  :   85 - 0x55
    "01010101", -- 4424 - 0x1148  :   85 - 0x55
    "01010101", -- 4425 - 0x1149  :   85 - 0x55
    "01000000", -- 4426 - 0x114a  :   64 - 0x40
    "00000000", -- 4427 - 0x114b  :    0 - 0x0
    "00000000", -- 4428 - 0x114c  :    0 - 0x0
    "00010110", -- 4429 - 0x114d  :   22 - 0x16
    "01000000", -- 4430 - 0x114e  :   64 - 0x40
    "01010101", -- 4431 - 0x114f  :   85 - 0x55
    "01010101", -- 4432 - 0x1150  :   85 - 0x55 -- Background 0x15
    "01011001", -- 4433 - 0x1151  :   89 - 0x59
    "01000000", -- 4434 - 0x1152  :   64 - 0x40
    "00000000", -- 4435 - 0x1153  :    0 - 0x0
    "00000000", -- 4436 - 0x1154  :    0 - 0x0
    "00010110", -- 4437 - 0x1155  :   22 - 0x16
    "01010101", -- 4438 - 0x1156  :   85 - 0x55
    "01101010", -- 4439 - 0x1157  :  106 - 0x6a
    "10010101", -- 4440 - 0x1158  :  149 - 0x95
    "01011001", -- 4441 - 0x1159  :   89 - 0x59
    "01000000", -- 4442 - 0x115a  :   64 - 0x40
    "00000000", -- 4443 - 0x115b  :    0 - 0x0
    "00000000", -- 4444 - 0x115c  :    0 - 0x0
    "00010110", -- 4445 - 0x115d  :   22 - 0x16
    "10100101", -- 4446 - 0x115e  :  165 - 0xa5
    "01010101", -- 4447 - 0x115f  :   85 - 0x55
    "01010101", -- 4448 - 0x1160  :   85 - 0x55 -- Background 0x16
    "10101001", -- 4449 - 0x1161  :  169 - 0xa9
    "01000000", -- 4450 - 0x1162  :   64 - 0x40
    "00000000", -- 4451 - 0x1163  :    0 - 0x0
    "00000000", -- 4452 - 0x1164  :    0 - 0x0
    "00010101", -- 4453 - 0x1165  :   21 - 0x15
    "01010101", -- 4454 - 0x1166  :   85 - 0x55
    "01010101", -- 4455 - 0x1167  :   85 - 0x55
    "01010101", -- 4456 - 0x1168  :   85 - 0x55
    "01010101", -- 4457 - 0x1169  :   85 - 0x55
    "01000000", -- 4458 - 0x116a  :   64 - 0x40
    "00000000", -- 4459 - 0x116b  :    0 - 0x0
    "00000000", -- 4460 - 0x116c  :    0 - 0x0
    "00010101", -- 4461 - 0x116d  :   21 - 0x15
    "01010101", -- 4462 - 0x116e  :   85 - 0x55
    "01010101", -- 4463 - 0x116f  :   85 - 0x55
    "01010101", -- 4464 - 0x1170  :   85 - 0x55 -- Background 0x17
    "01010101", -- 4465 - 0x1171  :   85 - 0x55
    "01000000", -- 4466 - 0x1172  :   64 - 0x40
    "00000000", -- 4467 - 0x1173  :    0 - 0x0
    "00000000", -- 4468 - 0x1174  :    0 - 0x0
    "00010100", -- 4469 - 0x1175  :   20 - 0x14
    "00000110", -- 4470 - 0x1176  :    6 - 0x6
    "00001000", -- 4471 - 0x1177  :    8 - 0x8
    "10110111", -- 4472 - 0x1178  :  183 - 0xb7
    "00000000", -- 4473 - 0x1179  :    0 - 0x0
    "10001011", -- 4474 - 0x117a  :  139 - 0x8b
    "00000000", -- 4475 - 0x117b  :    0 - 0x0
    "00010101", -- 4476 - 0x117c  :   21 - 0x15
    "01010101", -- 4477 - 0x117d  :   85 - 0x55
    "01010101", -- 4478 - 0x117e  :   85 - 0x55
    "01010101", -- 4479 - 0x117f  :   85 - 0x55
    "01010101", -- 4480 - 0x1180  :   85 - 0x55 -- Background 0x18
    "01000000", -- 4481 - 0x1181  :   64 - 0x40
    "00000000", -- 4482 - 0x1182  :    0 - 0x0
    "00000000", -- 4483 - 0x1183  :    0 - 0x0
    "00011010", -- 4484 - 0x1184  :   26 - 0x1a
    "01010111", -- 4485 - 0x1185  :   87 - 0x57
    "01010101", -- 4486 - 0x1186  :   85 - 0x55
    "01011101", -- 4487 - 0x1187  :   93 - 0x5d
    "01011010", -- 4488 - 0x1188  :   90 - 0x5a
    "01000000", -- 4489 - 0x1189  :   64 - 0x40
    "00000000", -- 4490 - 0x118a  :    0 - 0x0
    "00000000", -- 4491 - 0x118b  :    0 - 0x0
    "00011010", -- 4492 - 0x118c  :   26 - 0x1a
    "01010111", -- 4493 - 0x118d  :   87 - 0x57
    "01010101", -- 4494 - 0x118e  :   85 - 0x55
    "01011101", -- 4495 - 0x118f  :   93 - 0x5d
    "01011010", -- 4496 - 0x1190  :   90 - 0x5a -- Background 0x19
    "01000000", -- 4497 - 0x1191  :   64 - 0x40
    "00000000", -- 4498 - 0x1192  :    0 - 0x0
    "00000000", -- 4499 - 0x1193  :    0 - 0x0
    "00010101", -- 4500 - 0x1194  :   21 - 0x15
    "01010111", -- 4501 - 0x1195  :   87 - 0x57
    "01011010", -- 4502 - 0x1196  :   90 - 0x5a
    "01011101", -- 4503 - 0x1197  :   93 - 0x5d
    "01010101", -- 4504 - 0x1198  :   85 - 0x55
    "01000000", -- 4505 - 0x1199  :   64 - 0x40
    "00000000", -- 4506 - 0x119a  :    0 - 0x0
    "00000000", -- 4507 - 0x119b  :    0 - 0x0
    "00010000", -- 4508 - 0x119c  :   16 - 0x10
    "00010101", -- 4509 - 0x119d  :   21 - 0x15
    "01011010", -- 4510 - 0x119e  :   90 - 0x5a
    "01010101", -- 4511 - 0x119f  :   85 - 0x55
    "01010101", -- 4512 - 0x11a0  :   85 - 0x55 -- Background 0x1a
    "01000000", -- 4513 - 0x11a1  :   64 - 0x40
    "00000000", -- 4514 - 0x11a2  :    0 - 0x0
    "00000000", -- 4515 - 0x11a3  :    0 - 0x0
    "00010000", -- 4516 - 0x11a4  :   16 - 0x10
    "00010101", -- 4517 - 0x11a5  :   21 - 0x15
    "01011010", -- 4518 - 0x11a6  :   90 - 0x5a
    "01010101", -- 4519 - 0x11a7  :   85 - 0x55
    "01010101", -- 4520 - 0x11a8  :   85 - 0x55
    "01000000", -- 4521 - 0x11a9  :   64 - 0x40
    "00000000", -- 4522 - 0x11aa  :    0 - 0x0
    "00000000", -- 4523 - 0x11ab  :    0 - 0x0
    "00010000", -- 4524 - 0x11ac  :   16 - 0x10
    "00010101", -- 4525 - 0x11ad  :   21 - 0x15
    "01011010", -- 4526 - 0x11ae  :   90 - 0x5a
    "01010101", -- 4527 - 0x11af  :   85 - 0x55
    "01010101", -- 4528 - 0x11b0  :   85 - 0x55 -- Background 0x1b
    "01000000", -- 4529 - 0x11b1  :   64 - 0x40
    "00000000", -- 4530 - 0x11b2  :    0 - 0x0
    "00000000", -- 4531 - 0x11b3  :    0 - 0x0
    "00010101", -- 4532 - 0x11b4  :   21 - 0x15
    "01010111", -- 4533 - 0x11b5  :   87 - 0x57
    "01011010", -- 4534 - 0x11b6  :   90 - 0x5a
    "01011101", -- 4535 - 0x11b7  :   93 - 0x5d
    "01010101", -- 4536 - 0x11b8  :   85 - 0x55
    "01000000", -- 4537 - 0x11b9  :   64 - 0x40
    "00000000", -- 4538 - 0x11ba  :    0 - 0x0
    "00000000", -- 4539 - 0x11bb  :    0 - 0x0
    "00011010", -- 4540 - 0x11bc  :   26 - 0x1a
    "01010111", -- 4541 - 0x11bd  :   87 - 0x57
    "01010101", -- 4542 - 0x11be  :   85 - 0x55
    "01011101", -- 4543 - 0x11bf  :   93 - 0x5d
    "01011010", -- 4544 - 0x11c0  :   90 - 0x5a -- Background 0x1c
    "01000000", -- 4545 - 0x11c1  :   64 - 0x40
    "00000000", -- 4546 - 0x11c2  :    0 - 0x0
    "00000000", -- 4547 - 0x11c3  :    0 - 0x0
    "00011010", -- 4548 - 0x11c4  :   26 - 0x1a
    "01010111", -- 4549 - 0x11c5  :   87 - 0x57
    "01010101", -- 4550 - 0x11c6  :   85 - 0x55
    "01011101", -- 4551 - 0x11c7  :   93 - 0x5d
    "01011010", -- 4552 - 0x11c8  :   90 - 0x5a
    "01000000", -- 4553 - 0x11c9  :   64 - 0x40
    "00000000", -- 4554 - 0x11ca  :    0 - 0x0
    "00000000", -- 4555 - 0x11cb  :    0 - 0x0
    "00010101", -- 4556 - 0x11cc  :   21 - 0x15
    "01010101", -- 4557 - 0x11cd  :   85 - 0x55
    "01010101", -- 4558 - 0x11ce  :   85 - 0x55
    "01010101", -- 4559 - 0x11cf  :   85 - 0x55
    "01010101", -- 4560 - 0x11d0  :   85 - 0x55 -- Background 0x1d
    "01000000", -- 4561 - 0x11d1  :   64 - 0x40
    "00000000", -- 4562 - 0x11d2  :    0 - 0x0
    "00000000", -- 4563 - 0x11d3  :    0 - 0x0
    "00010100", -- 4564 - 0x11d4  :   20 - 0x14
    "00000011", -- 4565 - 0x11d5  :    3 - 0x3
    "00001000", -- 4566 - 0x11d6  :    8 - 0x8
    "10101101", -- 4567 - 0x11d7  :  173 - 0xad
    "00000000", -- 4568 - 0x11d8  :    0 - 0x0
    "10010011", -- 4569 - 0x11d9  :  147 - 0x93
    "00000000", -- 4570 - 0x11da  :    0 - 0x0
    "00010101", -- 4571 - 0x11db  :   21 - 0x15
    "01010101", -- 4572 - 0x11dc  :   85 - 0x55
    "01010101", -- 4573 - 0x11dd  :   85 - 0x55
    "01010101", -- 4574 - 0x11de  :   85 - 0x55
    "01010101", -- 4575 - 0x11df  :   85 - 0x55
    "01010101", -- 4576 - 0x11e0  :   85 - 0x55 -- Background 0x1e
    "01010000", -- 4577 - 0x11e1  :   80 - 0x50
    "00000000", -- 4578 - 0x11e2  :    0 - 0x0
    "00010101", -- 4579 - 0x11e3  :   21 - 0x15
    "01110101", -- 4580 - 0x11e4  :  117 - 0x75
    "01010101", -- 4581 - 0x11e5  :   85 - 0x55
    "01010111", -- 4582 - 0x11e6  :   87 - 0x57
    "01010101", -- 4583 - 0x11e7  :   85 - 0x55
    "01010111", -- 4584 - 0x11e8  :   87 - 0x57
    "01010000", -- 4585 - 0x11e9  :   80 - 0x50
    "00000000", -- 4586 - 0x11ea  :    0 - 0x0
    "00011101", -- 4587 - 0x11eb  :   29 - 0x1d
    "01010101", -- 4588 - 0x11ec  :   85 - 0x55
    "01110101", -- 4589 - 0x11ed  :  117 - 0x75
    "01010101", -- 4590 - 0x11ee  :   85 - 0x55
    "01011101", -- 4591 - 0x11ef  :   93 - 0x5d
    "01010101", -- 4592 - 0x11f0  :   85 - 0x55 -- Background 0x1f
    "01010000", -- 4593 - 0x11f1  :   80 - 0x50
    "00000000", -- 4594 - 0x11f2  :    0 - 0x0
    "00010101", -- 4595 - 0x11f3  :   21 - 0x15
    "01010111", -- 4596 - 0x11f4  :   87 - 0x57
    "01010101", -- 4597 - 0x11f5  :   85 - 0x55
    "01010101", -- 4598 - 0x11f6  :   85 - 0x55
    "01010101", -- 4599 - 0x11f7  :   85 - 0x55
    "01110101", -- 4600 - 0x11f8  :  117 - 0x75
    "01010000", -- 4601 - 0x11f9  :   80 - 0x50
    "00000000", -- 4602 - 0x11fa  :    0 - 0x0
    "00010101", -- 4603 - 0x11fb  :   21 - 0x15
    "01010101", -- 4604 - 0x11fc  :   85 - 0x55
    "01010101", -- 4605 - 0x11fd  :   85 - 0x55
    "00000001", -- 4606 - 0x11fe  :    1 - 0x1
    "01010101", -- 4607 - 0x11ff  :   85 - 0x55
    "01010101", -- 4608 - 0x1200  :   85 - 0x55 -- Background 0x20
    "11010000", -- 4609 - 0x1201  :  208 - 0xd0
    "00000000", -- 4610 - 0x1202  :    0 - 0x0
    "00010111", -- 4611 - 0x1203  :   23 - 0x17
    "01010101", -- 4612 - 0x1204  :   85 - 0x55
    "01010101", -- 4613 - 0x1205  :   85 - 0x55
    "00000001", -- 4614 - 0x1206  :    1 - 0x1
    "01010111", -- 4615 - 0x1207  :   87 - 0x57
    "01010101", -- 4616 - 0x1208  :   85 - 0x55
    "01010000", -- 4617 - 0x1209  :   80 - 0x50
    "00000000", -- 4618 - 0x120a  :    0 - 0x0
    "00010101", -- 4619 - 0x120b  :   21 - 0x15
    "01011101", -- 4620 - 0x120c  :   93 - 0x5d
    "01010101", -- 4621 - 0x120d  :   85 - 0x55
    "00000001", -- 4622 - 0x120e  :    1 - 0x1
    "01010101", -- 4623 - 0x120f  :   85 - 0x55
    "01010101", -- 4624 - 0x1210  :   85 - 0x55 -- Background 0x21
    "01010000", -- 4625 - 0x1211  :   80 - 0x50
    "00000000", -- 4626 - 0x1212  :    0 - 0x0
    "00010101", -- 4627 - 0x1213  :   21 - 0x15
    "01010101", -- 4628 - 0x1214  :   85 - 0x55
    "01110101", -- 4629 - 0x1215  :  117 - 0x75
    "01010101", -- 4630 - 0x1216  :   85 - 0x55
    "01010101", -- 4631 - 0x1217  :   85 - 0x55
    "01110101", -- 4632 - 0x1218  :  117 - 0x75
    "01010000", -- 4633 - 0x1219  :   80 - 0x50
    "00000000", -- 4634 - 0x121a  :    0 - 0x0
    "00011101", -- 4635 - 0x121b  :   29 - 0x1d
    "01010101", -- 4636 - 0x121c  :   85 - 0x55
    "01010101", -- 4637 - 0x121d  :   85 - 0x55
    "01010101", -- 4638 - 0x121e  :   85 - 0x55
    "01110101", -- 4639 - 0x121f  :  117 - 0x75
    "01010101", -- 4640 - 0x1220  :   85 - 0x55 -- Background 0x22
    "01010000", -- 4641 - 0x1221  :   80 - 0x50
    "00000000", -- 4642 - 0x1222  :    0 - 0x0
    "00010101", -- 4643 - 0x1223  :   21 - 0x15
    "01110101", -- 4644 - 0x1224  :  117 - 0x75
    "01010101", -- 4645 - 0x1225  :   85 - 0x55
    "11010101", -- 4646 - 0x1226  :  213 - 0xd5
    "01010101", -- 4647 - 0x1227  :   85 - 0x55
    "01010111", -- 4648 - 0x1228  :   87 - 0x57
    "01010000", -- 4649 - 0x1229  :   80 - 0x50
    "00000000", -- 4650 - 0x122a  :    0 - 0x0
    "00010101", -- 4651 - 0x122b  :   21 - 0x15
    "01010101", -- 4652 - 0x122c  :   85 - 0x55
    "01010101", -- 4653 - 0x122d  :   85 - 0x55
    "01010101", -- 4654 - 0x122e  :   85 - 0x55
    "01010101", -- 4655 - 0x122f  :   85 - 0x55
    "01010101", -- 4656 - 0x1230  :   85 - 0x55 -- Background 0x23
    "01010000", -- 4657 - 0x1231  :   80 - 0x50
    "00000000", -- 4658 - 0x1232  :    0 - 0x0
    "00011001", -- 4659 - 0x1233  :   25 - 0x19
    "00001101", -- 4660 - 0x1234  :   13 - 0xd
    "00001000", -- 4661 - 0x1235  :    8 - 0x8
    "11110111", -- 4662 - 0x1236  :  247 - 0xf7
    "00000000", -- 4663 - 0x1237  :    0 - 0x0
    "01100111", -- 4664 - 0x1238  :  103 - 0x67
    "00000000", -- 4665 - 0x1239  :    0 - 0x0
    "00010101", -- 4666 - 0x123a  :   21 - 0x15
    "01010101", -- 4667 - 0x123b  :   85 - 0x55
    "01010101", -- 4668 - 0x123c  :   85 - 0x55
    "01010101", -- 4669 - 0x123d  :   85 - 0x55
    "01010101", -- 4670 - 0x123e  :   85 - 0x55
    "01010101", -- 4671 - 0x123f  :   85 - 0x55
    "01010000", -- 4672 - 0x1240  :   80 - 0x50 -- Background 0x24
    "00000000", -- 4673 - 0x1241  :    0 - 0x0
    "00011010", -- 4674 - 0x1242  :   26 - 0x1a
    "10101001", -- 4675 - 0x1243  :  169 - 0xa9
    "10101010", -- 4676 - 0x1244  :  170 - 0xaa
    "10011001", -- 4677 - 0x1245  :  153 - 0x99
    "01011001", -- 4678 - 0x1246  :   89 - 0x59
    "10101010", -- 4679 - 0x1247  :  170 - 0xaa
    "10010000", -- 4680 - 0x1248  :  144 - 0x90
    "00000000", -- 4681 - 0x1249  :    0 - 0x0
    "00011001", -- 4682 - 0x124a  :   25 - 0x19
    "01011001", -- 4683 - 0x124b  :   89 - 0x59
    "10010101", -- 4684 - 0x124c  :  149 - 0x95
    "10011001", -- 4685 - 0x124d  :  153 - 0x99
    "01011001", -- 4686 - 0x124e  :   89 - 0x59
    "10010101", -- 4687 - 0x124f  :  149 - 0x95
    "10010000", -- 4688 - 0x1250  :  144 - 0x90 -- Background 0x25
    "00000000", -- 4689 - 0x1251  :    0 - 0x0
    "00010101", -- 4690 - 0x1252  :   21 - 0x15
    "01011001", -- 4691 - 0x1253  :   89 - 0x59
    "10010101", -- 4692 - 0x1254  :  149 - 0x95
    "10011001", -- 4693 - 0x1255  :  153 - 0x99
    "01011001", -- 4694 - 0x1256  :   89 - 0x59
    "10010101", -- 4695 - 0x1257  :  149 - 0x95
    "01010000", -- 4696 - 0x1258  :   80 - 0x50
    "00000000", -- 4697 - 0x1259  :    0 - 0x0
    "00010000", -- 4698 - 0x125a  :   16 - 0x10
    "00010101", -- 4699 - 0x125b  :   21 - 0x15
    "10010101", -- 4700 - 0x125c  :  149 - 0x95
    "10011010", -- 4701 - 0x125d  :  154 - 0x9a
    "10101001", -- 4702 - 0x125e  :  169 - 0xa9
    "01010101", -- 4703 - 0x125f  :   85 - 0x55
    "01010000", -- 4704 - 0x1260  :   80 - 0x50 -- Background 0x26
    "00000000", -- 4705 - 0x1261  :    0 - 0x0
    "00010000", -- 4706 - 0x1262  :   16 - 0x10
    "00010101", -- 4707 - 0x1263  :   21 - 0x15
    "01010101", -- 4708 - 0x1264  :   85 - 0x55
    "01010101", -- 4709 - 0x1265  :   85 - 0x55
    "01010101", -- 4710 - 0x1266  :   85 - 0x55
    "01010101", -- 4711 - 0x1267  :   85 - 0x55
    "01010000", -- 4712 - 0x1268  :   80 - 0x50
    "00000000", -- 4713 - 0x1269  :    0 - 0x0
    "00010000", -- 4714 - 0x126a  :   16 - 0x10
    "00010101", -- 4715 - 0x126b  :   21 - 0x15
    "10101010", -- 4716 - 0x126c  :  170 - 0xaa
    "10011001", -- 4717 - 0x126d  :  153 - 0x99
    "01011001", -- 4718 - 0x126e  :   89 - 0x59
    "01010101", -- 4719 - 0x126f  :   85 - 0x55
    "01010000", -- 4720 - 0x1270  :   80 - 0x50 -- Background 0x27
    "00000000", -- 4721 - 0x1271  :    0 - 0x0
    "00010101", -- 4722 - 0x1272  :   21 - 0x15
    "01011001", -- 4723 - 0x1273  :   89 - 0x59
    "10010101", -- 4724 - 0x1274  :  149 - 0x95
    "10011001", -- 4725 - 0x1275  :  153 - 0x99
    "01011001", -- 4726 - 0x1276  :   89 - 0x59
    "10010101", -- 4727 - 0x1277  :  149 - 0x95
    "01010000", -- 4728 - 0x1278  :   80 - 0x50
    "00000000", -- 4729 - 0x1279  :    0 - 0x0
    "00011001", -- 4730 - 0x127a  :   25 - 0x19
    "01011001", -- 4731 - 0x127b  :   89 - 0x59
    "10010101", -- 4732 - 0x127c  :  149 - 0x95
    "10011001", -- 4733 - 0x127d  :  153 - 0x99
    "01011001", -- 4734 - 0x127e  :   89 - 0x59
    "10010101", -- 4735 - 0x127f  :  149 - 0x95
    "10010000", -- 4736 - 0x1280  :  144 - 0x90 -- Background 0x28
    "00000000", -- 4737 - 0x1281  :    0 - 0x0
    "00011010", -- 4738 - 0x1282  :   26 - 0x1a
    "10101001", -- 4739 - 0x1283  :  169 - 0xa9
    "10010101", -- 4740 - 0x1284  :  149 - 0x95
    "10011010", -- 4741 - 0x1285  :  154 - 0x9a
    "10101001", -- 4742 - 0x1286  :  169 - 0xa9
    "10101010", -- 4743 - 0x1287  :  170 - 0xaa
    "10010000", -- 4744 - 0x1288  :  144 - 0x90
    "00000000", -- 4745 - 0x1289  :    0 - 0x0
    "00010101", -- 4746 - 0x128a  :   21 - 0x15
    "01010101", -- 4747 - 0x128b  :   85 - 0x55
    "01010101", -- 4748 - 0x128c  :   85 - 0x55
    "01010101", -- 4749 - 0x128d  :   85 - 0x55
    "01010101", -- 4750 - 0x128e  :   85 - 0x55
    "01010101", -- 4751 - 0x128f  :   85 - 0x55
    "01010000", -- 4752 - 0x1290  :   80 - 0x50 -- Background 0x29
    "00000000", -- 4753 - 0x1291  :    0 - 0x0
    "00011001", -- 4754 - 0x1292  :   25 - 0x19
    "00000011", -- 4755 - 0x1293  :    3 - 0x3
    "00001000", -- 4756 - 0x1294  :    8 - 0x8
    "10111110", -- 4757 - 0x1295  :  190 - 0xbe
    "00000000", -- 4758 - 0x1296  :    0 - 0x0
    "10000110", -- 4759 - 0x1297  :  134 - 0x86
    "00000000", -- 4760 - 0x1298  :    0 - 0x0
    "00010101", -- 4761 - 0x1299  :   21 - 0x15
    "01010111", -- 4762 - 0x129a  :   87 - 0x57
    "01010101", -- 4763 - 0x129b  :   85 - 0x55
    "01010101", -- 4764 - 0x129c  :   85 - 0x55
    "01010111", -- 4765 - 0x129d  :   87 - 0x57
    "01010101", -- 4766 - 0x129e  :   85 - 0x55
    "01010000", -- 4767 - 0x129f  :   80 - 0x50
    "00000000", -- 4768 - 0x12a0  :    0 - 0x0 -- Background 0x2a
    "00010101", -- 4769 - 0x12a1  :   21 - 0x15
    "01010111", -- 4770 - 0x12a2  :   87 - 0x57
    "01101010", -- 4771 - 0x12a3  :  106 - 0x6a
    "01010110", -- 4772 - 0x12a4  :   86 - 0x56
    "10100111", -- 4773 - 0x12a5  :  167 - 0xa7
    "01010101", -- 4774 - 0x12a6  :   85 - 0x55
    "01010000", -- 4775 - 0x12a7  :   80 - 0x50
    "00000000", -- 4776 - 0x12a8  :    0 - 0x0
    "00010101", -- 4777 - 0x12a9  :   21 - 0x15
    "01010111", -- 4778 - 0x12aa  :   87 - 0x57
    "01101010", -- 4779 - 0x12ab  :  106 - 0x6a
    "01010110", -- 4780 - 0x12ac  :   86 - 0x56
    "10100111", -- 4781 - 0x12ad  :  167 - 0xa7
    "01010101", -- 4782 - 0x12ae  :   85 - 0x55
    "01010000", -- 4783 - 0x12af  :   80 - 0x50
    "00000000", -- 4784 - 0x12b0  :    0 - 0x0 -- Background 0x2b
    "00010101", -- 4785 - 0x12b1  :   21 - 0x15
    "01010111", -- 4786 - 0x12b2  :   87 - 0x57
    "01010101", -- 4787 - 0x12b3  :   85 - 0x55
    "01110101", -- 4788 - 0x12b4  :  117 - 0x75
    "01010111", -- 4789 - 0x12b5  :   87 - 0x57
    "01010101", -- 4790 - 0x12b6  :   85 - 0x55
    "01010000", -- 4791 - 0x12b7  :   80 - 0x50
    "00000000", -- 4792 - 0x12b8  :    0 - 0x0
    "00010000", -- 4793 - 0x12b9  :   16 - 0x10
    "00010101", -- 4794 - 0x12ba  :   21 - 0x15
    "01010101", -- 4795 - 0x12bb  :   85 - 0x55
    "01110101", -- 4796 - 0x12bc  :  117 - 0x75
    "01010101", -- 4797 - 0x12bd  :   85 - 0x55
    "01010101", -- 4798 - 0x12be  :   85 - 0x55
    "01010000", -- 4799 - 0x12bf  :   80 - 0x50
    "00000000", -- 4800 - 0x12c0  :    0 - 0x0 -- Background 0x2c
    "00010000", -- 4801 - 0x12c1  :   16 - 0x10
    "00010101", -- 4802 - 0x12c2  :   21 - 0x15
    "01010101", -- 4803 - 0x12c3  :   85 - 0x55
    "01110101", -- 4804 - 0x12c4  :  117 - 0x75
    "01010101", -- 4805 - 0x12c5  :   85 - 0x55
    "01010101", -- 4806 - 0x12c6  :   85 - 0x55
    "01010000", -- 4807 - 0x12c7  :   80 - 0x50
    "00000000", -- 4808 - 0x12c8  :    0 - 0x0
    "00010000", -- 4809 - 0x12c9  :   16 - 0x10
    "00010101", -- 4810 - 0x12ca  :   21 - 0x15
    "01010101", -- 4811 - 0x12cb  :   85 - 0x55
    "01110101", -- 4812 - 0x12cc  :  117 - 0x75
    "01010101", -- 4813 - 0x12cd  :   85 - 0x55
    "01010101", -- 4814 - 0x12ce  :   85 - 0x55
    "01010000", -- 4815 - 0x12cf  :   80 - 0x50
    "00000000", -- 4816 - 0x12d0  :    0 - 0x0 -- Background 0x2d
    "00010101", -- 4817 - 0x12d1  :   21 - 0x15
    "01010111", -- 4818 - 0x12d2  :   87 - 0x57
    "01010101", -- 4819 - 0x12d3  :   85 - 0x55
    "01110101", -- 4820 - 0x12d4  :  117 - 0x75
    "01010111", -- 4821 - 0x12d5  :   87 - 0x57
    "01010101", -- 4822 - 0x12d6  :   85 - 0x55
    "01010000", -- 4823 - 0x12d7  :   80 - 0x50
    "00000000", -- 4824 - 0x12d8  :    0 - 0x0
    "00010101", -- 4825 - 0x12d9  :   21 - 0x15
    "01010111", -- 4826 - 0x12da  :   87 - 0x57
    "01101010", -- 4827 - 0x12db  :  106 - 0x6a
    "01010110", -- 4828 - 0x12dc  :   86 - 0x56
    "10100111", -- 4829 - 0x12dd  :  167 - 0xa7
    "01010101", -- 4830 - 0x12de  :   85 - 0x55
    "01010000", -- 4831 - 0x12df  :   80 - 0x50
    "00000000", -- 4832 - 0x12e0  :    0 - 0x0 -- Background 0x2e
    "00010101", -- 4833 - 0x12e1  :   21 - 0x15
    "01010111", -- 4834 - 0x12e2  :   87 - 0x57
    "01101010", -- 4835 - 0x12e3  :  106 - 0x6a
    "01010110", -- 4836 - 0x12e4  :   86 - 0x56
    "10100111", -- 4837 - 0x12e5  :  167 - 0xa7
    "01010101", -- 4838 - 0x12e6  :   85 - 0x55
    "01010000", -- 4839 - 0x12e7  :   80 - 0x50
    "00000000", -- 4840 - 0x12e8  :    0 - 0x0
    "00010101", -- 4841 - 0x12e9  :   21 - 0x15
    "01010111", -- 4842 - 0x12ea  :   87 - 0x57
    "01010101", -- 4843 - 0x12eb  :   85 - 0x55
    "01010101", -- 4844 - 0x12ec  :   85 - 0x55
    "01010111", -- 4845 - 0x12ed  :   87 - 0x57
    "01010101", -- 4846 - 0x12ee  :   85 - 0x55
    "01010000", -- 4847 - 0x12ef  :   80 - 0x50
    "00000000", -- 4848 - 0x12f0  :    0 - 0x0 -- Background 0x2f
    "00011001", -- 4849 - 0x12f1  :   25 - 0x19
    "00000011", -- 4850 - 0x12f2  :    3 - 0x3
    "00001000", -- 4851 - 0x12f3  :    8 - 0x8
    "11011101", -- 4852 - 0x12f4  :  221 - 0xdd
    "00000000", -- 4853 - 0x12f5  :    0 - 0x0
    "01110011", -- 4854 - 0x12f6  :  115 - 0x73
    "00000000", -- 4855 - 0x12f7  :    0 - 0x0
    "00010101", -- 4856 - 0x12f8  :   21 - 0x15
    "01010101", -- 4857 - 0x12f9  :   85 - 0x55
    "01010101", -- 4858 - 0x12fa  :   85 - 0x55
    "01010101", -- 4859 - 0x12fb  :   85 - 0x55
    "01010101", -- 4860 - 0x12fc  :   85 - 0x55
    "01010101", -- 4861 - 0x12fd  :   85 - 0x55
    "01010101", -- 4862 - 0x12fe  :   85 - 0x55
    "01010100", -- 4863 - 0x12ff  :   84 - 0x54
    "00011001", -- 4864 - 0x1300  :   25 - 0x19 -- Background 0x30
    "01100101", -- 4865 - 0x1301  :  101 - 0x65
    "10010110", -- 4866 - 0x1302  :  150 - 0x96
    "10100101", -- 4867 - 0x1303  :  165 - 0xa5
    "01011010", -- 4868 - 0x1304  :   90 - 0x5a
    "10010110", -- 4869 - 0x1305  :  150 - 0x96
    "01011001", -- 4870 - 0x1306  :   89 - 0x59
    "01100100", -- 4871 - 0x1307  :  100 - 0x64
    "00011001", -- 4872 - 0x1308  :   25 - 0x19
    "01100101", -- 4873 - 0x1309  :  101 - 0x65
    "10010101", -- 4874 - 0x130a  :  149 - 0x95
    "01010101", -- 4875 - 0x130b  :   85 - 0x55
    "01010101", -- 4876 - 0x130c  :   85 - 0x55
    "01010110", -- 4877 - 0x130d  :   86 - 0x56
    "01011001", -- 4878 - 0x130e  :   89 - 0x59
    "01100100", -- 4879 - 0x130f  :  100 - 0x64
    "00011001", -- 4880 - 0x1310  :   25 - 0x19 -- Background 0x31
    "01100101", -- 4881 - 0x1311  :  101 - 0x65
    "10010110", -- 4882 - 0x1312  :  150 - 0x96
    "10100101", -- 4883 - 0x1313  :  165 - 0xa5
    "01011010", -- 4884 - 0x1314  :   90 - 0x5a
    "10010110", -- 4885 - 0x1315  :  150 - 0x96
    "01011001", -- 4886 - 0x1316  :   89 - 0x59
    "01100100", -- 4887 - 0x1317  :  100 - 0x64
    "00010101", -- 4888 - 0x1318  :   21 - 0x15
    "01010101", -- 4889 - 0x1319  :   85 - 0x55
    "01010101", -- 4890 - 0x131a  :   85 - 0x55
    "01010000", -- 4891 - 0x131b  :   80 - 0x50
    "00000101", -- 4892 - 0x131c  :    5 - 0x5
    "01010101", -- 4893 - 0x131d  :   85 - 0x55
    "01010101", -- 4894 - 0x131e  :   85 - 0x55
    "01010100", -- 4895 - 0x131f  :   84 - 0x54
    "00011111", -- 4896 - 0x1320  :   31 - 0x1f -- Background 0x32
    "01111101", -- 4897 - 0x1321  :  125 - 0x7d
    "11010101", -- 4898 - 0x1322  :  213 - 0xd5
    "01010000", -- 4899 - 0x1323  :   80 - 0x50
    "00000101", -- 4900 - 0x1324  :    5 - 0x5
    "01010111", -- 4901 - 0x1325  :   87 - 0x57
    "11111111", -- 4902 - 0x1326  :  255 - 0xff
    "01110100", -- 4903 - 0x1327  :  116 - 0x74
    "00010101", -- 4904 - 0x1328  :   21 - 0x15
    "01010101", -- 4905 - 0x1329  :   85 - 0x55
    "01010101", -- 4906 - 0x132a  :   85 - 0x55
    "01010000", -- 4907 - 0x132b  :   80 - 0x50
    "00000101", -- 4908 - 0x132c  :    5 - 0x5
    "01010101", -- 4909 - 0x132d  :   85 - 0x55
    "01010101", -- 4910 - 0x132e  :   85 - 0x55
    "01010100", -- 4911 - 0x132f  :   84 - 0x54
    "00011001", -- 4912 - 0x1330  :   25 - 0x19 -- Background 0x33
    "01100101", -- 4913 - 0x1331  :  101 - 0x65
    "10010110", -- 4914 - 0x1332  :  150 - 0x96
    "10100101", -- 4915 - 0x1333  :  165 - 0xa5
    "01011010", -- 4916 - 0x1334  :   90 - 0x5a
    "10010110", -- 4917 - 0x1335  :  150 - 0x96
    "01011001", -- 4918 - 0x1336  :   89 - 0x59
    "01100100", -- 4919 - 0x1337  :  100 - 0x64
    "00011001", -- 4920 - 0x1338  :   25 - 0x19
    "01100101", -- 4921 - 0x1339  :  101 - 0x65
    "10010101", -- 4922 - 0x133a  :  149 - 0x95
    "01010101", -- 4923 - 0x133b  :   85 - 0x55
    "01010101", -- 4924 - 0x133c  :   85 - 0x55
    "01010110", -- 4925 - 0x133d  :   86 - 0x56
    "01011001", -- 4926 - 0x133e  :   89 - 0x59
    "01100100", -- 4927 - 0x133f  :  100 - 0x64
    "00011001", -- 4928 - 0x1340  :   25 - 0x19 -- Background 0x34
    "01100101", -- 4929 - 0x1341  :  101 - 0x65
    "10010110", -- 4930 - 0x1342  :  150 - 0x96
    "10100101", -- 4931 - 0x1343  :  165 - 0xa5
    "01011010", -- 4932 - 0x1344  :   90 - 0x5a
    "10010110", -- 4933 - 0x1345  :  150 - 0x96
    "01011001", -- 4934 - 0x1346  :   89 - 0x59
    "01100100", -- 4935 - 0x1347  :  100 - 0x64
    "00010101", -- 4936 - 0x1348  :   21 - 0x15
    "01010101", -- 4937 - 0x1349  :   85 - 0x55
    "01010101", -- 4938 - 0x134a  :   85 - 0x55
    "01010101", -- 4939 - 0x134b  :   85 - 0x55
    "01010101", -- 4940 - 0x134c  :   85 - 0x55
    "01010101", -- 4941 - 0x134d  :   85 - 0x55
    "01010101", -- 4942 - 0x134e  :   85 - 0x55
    "01010100", -- 4943 - 0x134f  :   84 - 0x54
    "00011110", -- 4944 - 0x1350  :   30 - 0x1e -- Background 0x35
    "00001111", -- 4945 - 0x1351  :   15 - 0xf
    "00001000", -- 4946 - 0x1352  :    8 - 0x8
    "11110111", -- 4947 - 0x1353  :  247 - 0xf7
    "00000000", -- 4948 - 0x1354  :    0 - 0x0
    "01100111", -- 4949 - 0x1355  :  103 - 0x67
    "00000000", -- 4950 - 0x1356  :    0 - 0x0
    "00010101", -- 4951 - 0x1357  :   21 - 0x15
    "01010101", -- 4952 - 0x1358  :   85 - 0x55
    "01010101", -- 4953 - 0x1359  :   85 - 0x55
    "01010101", -- 4954 - 0x135a  :   85 - 0x55
    "01010101", -- 4955 - 0x135b  :   85 - 0x55
    "01010101", -- 4956 - 0x135c  :   85 - 0x55
    "01010101", -- 4957 - 0x135d  :   85 - 0x55
    "01010100", -- 4958 - 0x135e  :   84 - 0x54
    "00010111", -- 4959 - 0x135f  :   23 - 0x17
    "01110101", -- 4960 - 0x1360  :  117 - 0x75 -- Background 0x36
    "01010110", -- 4961 - 0x1361  :   86 - 0x56
    "10100101", -- 4962 - 0x1362  :  165 - 0xa5
    "01011010", -- 4963 - 0x1363  :   90 - 0x5a
    "10010101", -- 4964 - 0x1364  :  149 - 0x95
    "01011101", -- 4965 - 0x1365  :   93 - 0x5d
    "11010100", -- 4966 - 0x1366  :  212 - 0xd4
    "00010101", -- 4967 - 0x1367  :   21 - 0x15
    "01010101", -- 4968 - 0x1368  :   85 - 0x55
    "01110110", -- 4969 - 0x1369  :  118 - 0x76
    "10100101", -- 4970 - 0x136a  :  165 - 0xa5
    "01011010", -- 4971 - 0x136b  :   90 - 0x5a
    "10011101", -- 4972 - 0x136c  :  157 - 0x9d
    "01010101", -- 4973 - 0x136d  :   85 - 0x55
    "01010100", -- 4974 - 0x136e  :   84 - 0x54
    "00010111", -- 4975 - 0x136f  :   23 - 0x17
    "01010101", -- 4976 - 0x1370  :   85 - 0x55 -- Background 0x37
    "01110101", -- 4977 - 0x1371  :  117 - 0x75
    "01010101", -- 4978 - 0x1372  :   85 - 0x55
    "01010101", -- 4979 - 0x1373  :   85 - 0x55
    "01011101", -- 4980 - 0x1374  :   93 - 0x5d
    "01010101", -- 4981 - 0x1375  :   85 - 0x55
    "11010100", -- 4982 - 0x1376  :  212 - 0xd4
    "00010101", -- 4983 - 0x1377  :   21 - 0x15
    "01101010", -- 4984 - 0x1378  :  106 - 0x6a
    "01110101", -- 4985 - 0x1379  :  117 - 0x75
    "01010000", -- 4986 - 0x137a  :   80 - 0x50
    "00000101", -- 4987 - 0x137b  :    5 - 0x5
    "01011101", -- 4988 - 0x137c  :   93 - 0x5d
    "10101001", -- 4989 - 0x137d  :  169 - 0xa9
    "01010100", -- 4990 - 0x137e  :   84 - 0x54
    "00010101", -- 4991 - 0x137f  :   21 - 0x15
    "01101110", -- 4992 - 0x1380  :  110 - 0x6e -- Background 0x38
    "01110101", -- 4993 - 0x1381  :  117 - 0x75
    "01010000", -- 4994 - 0x1382  :   80 - 0x50
    "00000101", -- 4995 - 0x1383  :    5 - 0x5
    "01011101", -- 4996 - 0x1384  :   93 - 0x5d
    "10111001", -- 4997 - 0x1385  :  185 - 0xb9
    "01010100", -- 4998 - 0x1386  :   84 - 0x54
    "00010101", -- 4999 - 0x1387  :   21 - 0x15
    "01101010", -- 5000 - 0x1388  :  106 - 0x6a
    "01110101", -- 5001 - 0x1389  :  117 - 0x75
    "01010000", -- 5002 - 0x138a  :   80 - 0x50
    "00000101", -- 5003 - 0x138b  :    5 - 0x5
    "01011101", -- 5004 - 0x138c  :   93 - 0x5d
    "10101001", -- 5005 - 0x138d  :  169 - 0xa9
    "01010100", -- 5006 - 0x138e  :   84 - 0x54
    "00010111", -- 5007 - 0x138f  :   23 - 0x17
    "01010101", -- 5008 - 0x1390  :   85 - 0x55 -- Background 0x39
    "01110101", -- 5009 - 0x1391  :  117 - 0x75
    "01010101", -- 5010 - 0x1392  :   85 - 0x55
    "01010101", -- 5011 - 0x1393  :   85 - 0x55
    "01011101", -- 5012 - 0x1394  :   93 - 0x5d
    "01010101", -- 5013 - 0x1395  :   85 - 0x55
    "11010100", -- 5014 - 0x1396  :  212 - 0xd4
    "00010101", -- 5015 - 0x1397  :   21 - 0x15
    "01010101", -- 5016 - 0x1398  :   85 - 0x55
    "01110101", -- 5017 - 0x1399  :  117 - 0x75
    "10101010", -- 5018 - 0x139a  :  170 - 0xaa
    "10101010", -- 5019 - 0x139b  :  170 - 0xaa
    "01011101", -- 5020 - 0x139c  :   93 - 0x5d
    "01010101", -- 5021 - 0x139d  :   85 - 0x55
    "01010100", -- 5022 - 0x139e  :   84 - 0x54
    "00010111", -- 5023 - 0x139f  :   23 - 0x17
    "01110101", -- 5024 - 0x13a0  :  117 - 0x75 -- Background 0x3a
    "01010101", -- 5025 - 0x13a1  :   85 - 0x55
    "01101010", -- 5026 - 0x13a2  :  106 - 0x6a
    "10101001", -- 5027 - 0x13a3  :  169 - 0xa9
    "01010101", -- 5028 - 0x13a4  :   85 - 0x55
    "01011101", -- 5029 - 0x13a5  :   93 - 0x5d
    "11010100", -- 5030 - 0x13a6  :  212 - 0xd4
    "00010101", -- 5031 - 0x13a7  :   21 - 0x15
    "01010101", -- 5032 - 0x13a8  :   85 - 0x55
    "01010101", -- 5033 - 0x13a9  :   85 - 0x55
    "01010101", -- 5034 - 0x13aa  :   85 - 0x55
    "01010101", -- 5035 - 0x13ab  :   85 - 0x55
    "01010101", -- 5036 - 0x13ac  :   85 - 0x55
    "01010101", -- 5037 - 0x13ad  :   85 - 0x55
    "01010100", -- 5038 - 0x13ae  :   84 - 0x54
    "00011110", -- 5039 - 0x13af  :   30 - 0x1e
    "00001111", -- 5040 - 0x13b0  :   15 - 0xf -- Background 0x3b
    "00001000", -- 5041 - 0x13b1  :    8 - 0x8
    "11111000", -- 5042 - 0x13b2  :  248 - 0xf8
    "00000000", -- 5043 - 0x13b3  :    0 - 0x0
    "01100111", -- 5044 - 0x13b4  :  103 - 0x67
    "00000000", -- 5045 - 0x13b5  :    0 - 0x0
    "00000000", -- 5046 - 0x13b6  :    0 - 0x0
    "00000000", -- 5047 - 0x13b7  :    0 - 0x0
    "00000000", -- 5048 - 0x13b8  :    0 - 0x0
    "00000000", -- 5049 - 0x13b9  :    0 - 0x0
    "00000000", -- 5050 - 0x13ba  :    0 - 0x0
    "00000000", -- 5051 - 0x13bb  :    0 - 0x0
    "00000000", -- 5052 - 0x13bc  :    0 - 0x0
    "00000000", -- 5053 - 0x13bd  :    0 - 0x0
    "00000000", -- 5054 - 0x13be  :    0 - 0x0
    "00000000", -- 5055 - 0x13bf  :    0 - 0x0
    "00000000", -- 5056 - 0x13c0  :    0 - 0x0 -- Background 0x3c
    "00000000", -- 5057 - 0x13c1  :    0 - 0x0
    "00000000", -- 5058 - 0x13c2  :    0 - 0x0
    "00000000", -- 5059 - 0x13c3  :    0 - 0x0
    "00000000", -- 5060 - 0x13c4  :    0 - 0x0
    "00000000", -- 5061 - 0x13c5  :    0 - 0x0
    "00000000", -- 5062 - 0x13c6  :    0 - 0x0
    "00000000", -- 5063 - 0x13c7  :    0 - 0x0
    "00000000", -- 5064 - 0x13c8  :    0 - 0x0
    "00000000", -- 5065 - 0x13c9  :    0 - 0x0
    "00000000", -- 5066 - 0x13ca  :    0 - 0x0
    "00000000", -- 5067 - 0x13cb  :    0 - 0x0
    "00000000", -- 5068 - 0x13cc  :    0 - 0x0
    "00000000", -- 5069 - 0x13cd  :    0 - 0x0
    "00000000", -- 5070 - 0x13ce  :    0 - 0x0
    "00000000", -- 5071 - 0x13cf  :    0 - 0x0
    "00000000", -- 5072 - 0x13d0  :    0 - 0x0 -- Background 0x3d
    "00000000", -- 5073 - 0x13d1  :    0 - 0x0
    "00000000", -- 5074 - 0x13d2  :    0 - 0x0
    "00000000", -- 5075 - 0x13d3  :    0 - 0x0
    "00000000", -- 5076 - 0x13d4  :    0 - 0x0
    "00000000", -- 5077 - 0x13d5  :    0 - 0x0
    "00000000", -- 5078 - 0x13d6  :    0 - 0x0
    "00000000", -- 5079 - 0x13d7  :    0 - 0x0
    "00000000", -- 5080 - 0x13d8  :    0 - 0x0
    "00000000", -- 5081 - 0x13d9  :    0 - 0x0
    "00000000", -- 5082 - 0x13da  :    0 - 0x0
    "00000000", -- 5083 - 0x13db  :    0 - 0x0
    "00000000", -- 5084 - 0x13dc  :    0 - 0x0
    "00000000", -- 5085 - 0x13dd  :    0 - 0x0
    "00000000", -- 5086 - 0x13de  :    0 - 0x0
    "00000000", -- 5087 - 0x13df  :    0 - 0x0
    "00000000", -- 5088 - 0x13e0  :    0 - 0x0 -- Background 0x3e
    "00000000", -- 5089 - 0x13e1  :    0 - 0x0
    "00000000", -- 5090 - 0x13e2  :    0 - 0x0
    "00000000", -- 5091 - 0x13e3  :    0 - 0x0
    "00000000", -- 5092 - 0x13e4  :    0 - 0x0
    "00000000", -- 5093 - 0x13e5  :    0 - 0x0
    "00000000", -- 5094 - 0x13e6  :    0 - 0x0
    "00000000", -- 5095 - 0x13e7  :    0 - 0x0
    "00000000", -- 5096 - 0x13e8  :    0 - 0x0
    "00000000", -- 5097 - 0x13e9  :    0 - 0x0
    "00000000", -- 5098 - 0x13ea  :    0 - 0x0
    "00000000", -- 5099 - 0x13eb  :    0 - 0x0
    "00000000", -- 5100 - 0x13ec  :    0 - 0x0
    "00000000", -- 5101 - 0x13ed  :    0 - 0x0
    "00000000", -- 5102 - 0x13ee  :    0 - 0x0
    "00000000", -- 5103 - 0x13ef  :    0 - 0x0
    "00000000", -- 5104 - 0x13f0  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 5105 - 0x13f1  :    0 - 0x0
    "00000000", -- 5106 - 0x13f2  :    0 - 0x0
    "00000000", -- 5107 - 0x13f3  :    0 - 0x0
    "00000000", -- 5108 - 0x13f4  :    0 - 0x0
    "00000000", -- 5109 - 0x13f5  :    0 - 0x0
    "00000000", -- 5110 - 0x13f6  :    0 - 0x0
    "00000000", -- 5111 - 0x13f7  :    0 - 0x0
    "00000000", -- 5112 - 0x13f8  :    0 - 0x0
    "00000000", -- 5113 - 0x13f9  :    0 - 0x0
    "00000000", -- 5114 - 0x13fa  :    0 - 0x0
    "00000000", -- 5115 - 0x13fb  :    0 - 0x0
    "00000000", -- 5116 - 0x13fc  :    0 - 0x0
    "00000000", -- 5117 - 0x13fd  :    0 - 0x0
    "00000000", -- 5118 - 0x13fe  :    0 - 0x0
    "00000000", -- 5119 - 0x13ff  :    0 - 0x0
    "00000000", -- 5120 - 0x1400  :    0 - 0x0 -- Background 0x40
    "00000000", -- 5121 - 0x1401  :    0 - 0x0
    "00000000", -- 5122 - 0x1402  :    0 - 0x0
    "00000000", -- 5123 - 0x1403  :    0 - 0x0
    "00000000", -- 5124 - 0x1404  :    0 - 0x0
    "00000000", -- 5125 - 0x1405  :    0 - 0x0
    "00000000", -- 5126 - 0x1406  :    0 - 0x0
    "00000000", -- 5127 - 0x1407  :    0 - 0x0
    "00000000", -- 5128 - 0x1408  :    0 - 0x0
    "00000000", -- 5129 - 0x1409  :    0 - 0x0
    "00000000", -- 5130 - 0x140a  :    0 - 0x0
    "00000000", -- 5131 - 0x140b  :    0 - 0x0
    "00000000", -- 5132 - 0x140c  :    0 - 0x0
    "00000000", -- 5133 - 0x140d  :    0 - 0x0
    "00000000", -- 5134 - 0x140e  :    0 - 0x0
    "00000000", -- 5135 - 0x140f  :    0 - 0x0
    "00000000", -- 5136 - 0x1410  :    0 - 0x0 -- Background 0x41
    "00000000", -- 5137 - 0x1411  :    0 - 0x0
    "00000000", -- 5138 - 0x1412  :    0 - 0x0
    "00000000", -- 5139 - 0x1413  :    0 - 0x0
    "00000000", -- 5140 - 0x1414  :    0 - 0x0
    "00000000", -- 5141 - 0x1415  :    0 - 0x0
    "00000000", -- 5142 - 0x1416  :    0 - 0x0
    "00000000", -- 5143 - 0x1417  :    0 - 0x0
    "00000000", -- 5144 - 0x1418  :    0 - 0x0
    "00000000", -- 5145 - 0x1419  :    0 - 0x0
    "00000000", -- 5146 - 0x141a  :    0 - 0x0
    "00000000", -- 5147 - 0x141b  :    0 - 0x0
    "00000000", -- 5148 - 0x141c  :    0 - 0x0
    "00000000", -- 5149 - 0x141d  :    0 - 0x0
    "00000000", -- 5150 - 0x141e  :    0 - 0x0
    "00000000", -- 5151 - 0x141f  :    0 - 0x0
    "00000000", -- 5152 - 0x1420  :    0 - 0x0 -- Background 0x42
    "00000000", -- 5153 - 0x1421  :    0 - 0x0
    "00000000", -- 5154 - 0x1422  :    0 - 0x0
    "00000000", -- 5155 - 0x1423  :    0 - 0x0
    "00000000", -- 5156 - 0x1424  :    0 - 0x0
    "00000000", -- 5157 - 0x1425  :    0 - 0x0
    "00000000", -- 5158 - 0x1426  :    0 - 0x0
    "00000000", -- 5159 - 0x1427  :    0 - 0x0
    "00000000", -- 5160 - 0x1428  :    0 - 0x0
    "00000000", -- 5161 - 0x1429  :    0 - 0x0
    "00000000", -- 5162 - 0x142a  :    0 - 0x0
    "00000000", -- 5163 - 0x142b  :    0 - 0x0
    "00000000", -- 5164 - 0x142c  :    0 - 0x0
    "00000000", -- 5165 - 0x142d  :    0 - 0x0
    "00000000", -- 5166 - 0x142e  :    0 - 0x0
    "00000000", -- 5167 - 0x142f  :    0 - 0x0
    "00000000", -- 5168 - 0x1430  :    0 - 0x0 -- Background 0x43
    "00000000", -- 5169 - 0x1431  :    0 - 0x0
    "00000000", -- 5170 - 0x1432  :    0 - 0x0
    "00000000", -- 5171 - 0x1433  :    0 - 0x0
    "00000000", -- 5172 - 0x1434  :    0 - 0x0
    "00000000", -- 5173 - 0x1435  :    0 - 0x0
    "00000000", -- 5174 - 0x1436  :    0 - 0x0
    "00000000", -- 5175 - 0x1437  :    0 - 0x0
    "00000000", -- 5176 - 0x1438  :    0 - 0x0
    "00000000", -- 5177 - 0x1439  :    0 - 0x0
    "00000000", -- 5178 - 0x143a  :    0 - 0x0
    "00000000", -- 5179 - 0x143b  :    0 - 0x0
    "00000000", -- 5180 - 0x143c  :    0 - 0x0
    "00000000", -- 5181 - 0x143d  :    0 - 0x0
    "00000000", -- 5182 - 0x143e  :    0 - 0x0
    "00000000", -- 5183 - 0x143f  :    0 - 0x0
    "00000000", -- 5184 - 0x1440  :    0 - 0x0 -- Background 0x44
    "00000000", -- 5185 - 0x1441  :    0 - 0x0
    "00000000", -- 5186 - 0x1442  :    0 - 0x0
    "00000000", -- 5187 - 0x1443  :    0 - 0x0
    "00000000", -- 5188 - 0x1444  :    0 - 0x0
    "00000000", -- 5189 - 0x1445  :    0 - 0x0
    "00000000", -- 5190 - 0x1446  :    0 - 0x0
    "00000000", -- 5191 - 0x1447  :    0 - 0x0
    "00000000", -- 5192 - 0x1448  :    0 - 0x0
    "00000000", -- 5193 - 0x1449  :    0 - 0x0
    "00000000", -- 5194 - 0x144a  :    0 - 0x0
    "00000000", -- 5195 - 0x144b  :    0 - 0x0
    "00000000", -- 5196 - 0x144c  :    0 - 0x0
    "00000000", -- 5197 - 0x144d  :    0 - 0x0
    "00000000", -- 5198 - 0x144e  :    0 - 0x0
    "00000000", -- 5199 - 0x144f  :    0 - 0x0
    "00000000", -- 5200 - 0x1450  :    0 - 0x0 -- Background 0x45
    "00000000", -- 5201 - 0x1451  :    0 - 0x0
    "00000000", -- 5202 - 0x1452  :    0 - 0x0
    "00000000", -- 5203 - 0x1453  :    0 - 0x0
    "00000000", -- 5204 - 0x1454  :    0 - 0x0
    "00000000", -- 5205 - 0x1455  :    0 - 0x0
    "00000000", -- 5206 - 0x1456  :    0 - 0x0
    "00000000", -- 5207 - 0x1457  :    0 - 0x0
    "00000000", -- 5208 - 0x1458  :    0 - 0x0
    "00000000", -- 5209 - 0x1459  :    0 - 0x0
    "00000000", -- 5210 - 0x145a  :    0 - 0x0
    "00000000", -- 5211 - 0x145b  :    0 - 0x0
    "00000000", -- 5212 - 0x145c  :    0 - 0x0
    "00000000", -- 5213 - 0x145d  :    0 - 0x0
    "00000000", -- 5214 - 0x145e  :    0 - 0x0
    "00000000", -- 5215 - 0x145f  :    0 - 0x0
    "00000000", -- 5216 - 0x1460  :    0 - 0x0 -- Background 0x46
    "00000000", -- 5217 - 0x1461  :    0 - 0x0
    "00000000", -- 5218 - 0x1462  :    0 - 0x0
    "00000000", -- 5219 - 0x1463  :    0 - 0x0
    "00000000", -- 5220 - 0x1464  :    0 - 0x0
    "00000000", -- 5221 - 0x1465  :    0 - 0x0
    "00000000", -- 5222 - 0x1466  :    0 - 0x0
    "00000000", -- 5223 - 0x1467  :    0 - 0x0
    "00000000", -- 5224 - 0x1468  :    0 - 0x0
    "00000000", -- 5225 - 0x1469  :    0 - 0x0
    "00000000", -- 5226 - 0x146a  :    0 - 0x0
    "00000000", -- 5227 - 0x146b  :    0 - 0x0
    "00000000", -- 5228 - 0x146c  :    0 - 0x0
    "00000000", -- 5229 - 0x146d  :    0 - 0x0
    "00000000", -- 5230 - 0x146e  :    0 - 0x0
    "00000000", -- 5231 - 0x146f  :    0 - 0x0
    "00000000", -- 5232 - 0x1470  :    0 - 0x0 -- Background 0x47
    "00000000", -- 5233 - 0x1471  :    0 - 0x0
    "00000000", -- 5234 - 0x1472  :    0 - 0x0
    "00000000", -- 5235 - 0x1473  :    0 - 0x0
    "00000000", -- 5236 - 0x1474  :    0 - 0x0
    "00000000", -- 5237 - 0x1475  :    0 - 0x0
    "00000000", -- 5238 - 0x1476  :    0 - 0x0
    "00000000", -- 5239 - 0x1477  :    0 - 0x0
    "00000000", -- 5240 - 0x1478  :    0 - 0x0
    "00000000", -- 5241 - 0x1479  :    0 - 0x0
    "00000000", -- 5242 - 0x147a  :    0 - 0x0
    "00000000", -- 5243 - 0x147b  :    0 - 0x0
    "00000000", -- 5244 - 0x147c  :    0 - 0x0
    "00000000", -- 5245 - 0x147d  :    0 - 0x0
    "00000000", -- 5246 - 0x147e  :    0 - 0x0
    "00000000", -- 5247 - 0x147f  :    0 - 0x0
    "00000000", -- 5248 - 0x1480  :    0 - 0x0 -- Background 0x48
    "00000000", -- 5249 - 0x1481  :    0 - 0x0
    "00000000", -- 5250 - 0x1482  :    0 - 0x0
    "00000000", -- 5251 - 0x1483  :    0 - 0x0
    "00000000", -- 5252 - 0x1484  :    0 - 0x0
    "00000000", -- 5253 - 0x1485  :    0 - 0x0
    "00000000", -- 5254 - 0x1486  :    0 - 0x0
    "00000000", -- 5255 - 0x1487  :    0 - 0x0
    "00000000", -- 5256 - 0x1488  :    0 - 0x0
    "00000000", -- 5257 - 0x1489  :    0 - 0x0
    "00000000", -- 5258 - 0x148a  :    0 - 0x0
    "00000000", -- 5259 - 0x148b  :    0 - 0x0
    "00000000", -- 5260 - 0x148c  :    0 - 0x0
    "00000000", -- 5261 - 0x148d  :    0 - 0x0
    "00000000", -- 5262 - 0x148e  :    0 - 0x0
    "00000000", -- 5263 - 0x148f  :    0 - 0x0
    "00000000", -- 5264 - 0x1490  :    0 - 0x0 -- Background 0x49
    "00000000", -- 5265 - 0x1491  :    0 - 0x0
    "00000000", -- 5266 - 0x1492  :    0 - 0x0
    "00000000", -- 5267 - 0x1493  :    0 - 0x0
    "00000000", -- 5268 - 0x1494  :    0 - 0x0
    "00000000", -- 5269 - 0x1495  :    0 - 0x0
    "00000000", -- 5270 - 0x1496  :    0 - 0x0
    "00000000", -- 5271 - 0x1497  :    0 - 0x0
    "00000000", -- 5272 - 0x1498  :    0 - 0x0
    "00000000", -- 5273 - 0x1499  :    0 - 0x0
    "00000000", -- 5274 - 0x149a  :    0 - 0x0
    "00000000", -- 5275 - 0x149b  :    0 - 0x0
    "00000000", -- 5276 - 0x149c  :    0 - 0x0
    "00000000", -- 5277 - 0x149d  :    0 - 0x0
    "00000000", -- 5278 - 0x149e  :    0 - 0x0
    "00000000", -- 5279 - 0x149f  :    0 - 0x0
    "00000000", -- 5280 - 0x14a0  :    0 - 0x0 -- Background 0x4a
    "00000000", -- 5281 - 0x14a1  :    0 - 0x0
    "00000000", -- 5282 - 0x14a2  :    0 - 0x0
    "00000000", -- 5283 - 0x14a3  :    0 - 0x0
    "00000000", -- 5284 - 0x14a4  :    0 - 0x0
    "00000000", -- 5285 - 0x14a5  :    0 - 0x0
    "00000000", -- 5286 - 0x14a6  :    0 - 0x0
    "00000000", -- 5287 - 0x14a7  :    0 - 0x0
    "00000000", -- 5288 - 0x14a8  :    0 - 0x0
    "00000000", -- 5289 - 0x14a9  :    0 - 0x0
    "00000000", -- 5290 - 0x14aa  :    0 - 0x0
    "00000000", -- 5291 - 0x14ab  :    0 - 0x0
    "00000000", -- 5292 - 0x14ac  :    0 - 0x0
    "00000000", -- 5293 - 0x14ad  :    0 - 0x0
    "00000000", -- 5294 - 0x14ae  :    0 - 0x0
    "00000000", -- 5295 - 0x14af  :    0 - 0x0
    "00000000", -- 5296 - 0x14b0  :    0 - 0x0 -- Background 0x4b
    "00000000", -- 5297 - 0x14b1  :    0 - 0x0
    "00000000", -- 5298 - 0x14b2  :    0 - 0x0
    "00000000", -- 5299 - 0x14b3  :    0 - 0x0
    "00000000", -- 5300 - 0x14b4  :    0 - 0x0
    "00000000", -- 5301 - 0x14b5  :    0 - 0x0
    "00000000", -- 5302 - 0x14b6  :    0 - 0x0
    "00000000", -- 5303 - 0x14b7  :    0 - 0x0
    "00000000", -- 5304 - 0x14b8  :    0 - 0x0
    "00000000", -- 5305 - 0x14b9  :    0 - 0x0
    "00000000", -- 5306 - 0x14ba  :    0 - 0x0
    "00000000", -- 5307 - 0x14bb  :    0 - 0x0
    "00000000", -- 5308 - 0x14bc  :    0 - 0x0
    "00000000", -- 5309 - 0x14bd  :    0 - 0x0
    "00000000", -- 5310 - 0x14be  :    0 - 0x0
    "00000000", -- 5311 - 0x14bf  :    0 - 0x0
    "00000000", -- 5312 - 0x14c0  :    0 - 0x0 -- Background 0x4c
    "00000000", -- 5313 - 0x14c1  :    0 - 0x0
    "00000000", -- 5314 - 0x14c2  :    0 - 0x0
    "00000000", -- 5315 - 0x14c3  :    0 - 0x0
    "00000000", -- 5316 - 0x14c4  :    0 - 0x0
    "00000000", -- 5317 - 0x14c5  :    0 - 0x0
    "00000000", -- 5318 - 0x14c6  :    0 - 0x0
    "00000000", -- 5319 - 0x14c7  :    0 - 0x0
    "00000000", -- 5320 - 0x14c8  :    0 - 0x0
    "00000000", -- 5321 - 0x14c9  :    0 - 0x0
    "00000000", -- 5322 - 0x14ca  :    0 - 0x0
    "00000000", -- 5323 - 0x14cb  :    0 - 0x0
    "00000000", -- 5324 - 0x14cc  :    0 - 0x0
    "00000000", -- 5325 - 0x14cd  :    0 - 0x0
    "00000000", -- 5326 - 0x14ce  :    0 - 0x0
    "00000000", -- 5327 - 0x14cf  :    0 - 0x0
    "00000000", -- 5328 - 0x14d0  :    0 - 0x0 -- Background 0x4d
    "00000000", -- 5329 - 0x14d1  :    0 - 0x0
    "00000000", -- 5330 - 0x14d2  :    0 - 0x0
    "00000000", -- 5331 - 0x14d3  :    0 - 0x0
    "00000000", -- 5332 - 0x14d4  :    0 - 0x0
    "00000000", -- 5333 - 0x14d5  :    0 - 0x0
    "00000000", -- 5334 - 0x14d6  :    0 - 0x0
    "00000000", -- 5335 - 0x14d7  :    0 - 0x0
    "00000000", -- 5336 - 0x14d8  :    0 - 0x0
    "00000000", -- 5337 - 0x14d9  :    0 - 0x0
    "00000000", -- 5338 - 0x14da  :    0 - 0x0
    "00000000", -- 5339 - 0x14db  :    0 - 0x0
    "00000000", -- 5340 - 0x14dc  :    0 - 0x0
    "00000000", -- 5341 - 0x14dd  :    0 - 0x0
    "00000000", -- 5342 - 0x14de  :    0 - 0x0
    "00000000", -- 5343 - 0x14df  :    0 - 0x0
    "00000000", -- 5344 - 0x14e0  :    0 - 0x0 -- Background 0x4e
    "00000000", -- 5345 - 0x14e1  :    0 - 0x0
    "00000000", -- 5346 - 0x14e2  :    0 - 0x0
    "00000000", -- 5347 - 0x14e3  :    0 - 0x0
    "00000000", -- 5348 - 0x14e4  :    0 - 0x0
    "00000000", -- 5349 - 0x14e5  :    0 - 0x0
    "00000000", -- 5350 - 0x14e6  :    0 - 0x0
    "00000000", -- 5351 - 0x14e7  :    0 - 0x0
    "00000000", -- 5352 - 0x14e8  :    0 - 0x0
    "00000000", -- 5353 - 0x14e9  :    0 - 0x0
    "00000000", -- 5354 - 0x14ea  :    0 - 0x0
    "00000000", -- 5355 - 0x14eb  :    0 - 0x0
    "00000000", -- 5356 - 0x14ec  :    0 - 0x0
    "00000000", -- 5357 - 0x14ed  :    0 - 0x0
    "00000000", -- 5358 - 0x14ee  :    0 - 0x0
    "00000000", -- 5359 - 0x14ef  :    0 - 0x0
    "00000000", -- 5360 - 0x14f0  :    0 - 0x0 -- Background 0x4f
    "00000000", -- 5361 - 0x14f1  :    0 - 0x0
    "00000000", -- 5362 - 0x14f2  :    0 - 0x0
    "00000000", -- 5363 - 0x14f3  :    0 - 0x0
    "00000000", -- 5364 - 0x14f4  :    0 - 0x0
    "00000000", -- 5365 - 0x14f5  :    0 - 0x0
    "00000000", -- 5366 - 0x14f6  :    0 - 0x0
    "00000000", -- 5367 - 0x14f7  :    0 - 0x0
    "00000000", -- 5368 - 0x14f8  :    0 - 0x0
    "00000000", -- 5369 - 0x14f9  :    0 - 0x0
    "00000000", -- 5370 - 0x14fa  :    0 - 0x0
    "00000000", -- 5371 - 0x14fb  :    0 - 0x0
    "00000000", -- 5372 - 0x14fc  :    0 - 0x0
    "00000000", -- 5373 - 0x14fd  :    0 - 0x0
    "00000000", -- 5374 - 0x14fe  :    0 - 0x0
    "00000000", -- 5375 - 0x14ff  :    0 - 0x0
    "00000000", -- 5376 - 0x1500  :    0 - 0x0 -- Background 0x50
    "00000000", -- 5377 - 0x1501  :    0 - 0x0
    "00000000", -- 5378 - 0x1502  :    0 - 0x0
    "00000000", -- 5379 - 0x1503  :    0 - 0x0
    "00000000", -- 5380 - 0x1504  :    0 - 0x0
    "00000000", -- 5381 - 0x1505  :    0 - 0x0
    "00000000", -- 5382 - 0x1506  :    0 - 0x0
    "00000000", -- 5383 - 0x1507  :    0 - 0x0
    "00000000", -- 5384 - 0x1508  :    0 - 0x0
    "00000000", -- 5385 - 0x1509  :    0 - 0x0
    "00000000", -- 5386 - 0x150a  :    0 - 0x0
    "00000000", -- 5387 - 0x150b  :    0 - 0x0
    "00000000", -- 5388 - 0x150c  :    0 - 0x0
    "00000000", -- 5389 - 0x150d  :    0 - 0x0
    "00000000", -- 5390 - 0x150e  :    0 - 0x0
    "00000000", -- 5391 - 0x150f  :    0 - 0x0
    "00000000", -- 5392 - 0x1510  :    0 - 0x0 -- Background 0x51
    "00000000", -- 5393 - 0x1511  :    0 - 0x0
    "00000000", -- 5394 - 0x1512  :    0 - 0x0
    "00000000", -- 5395 - 0x1513  :    0 - 0x0
    "00000000", -- 5396 - 0x1514  :    0 - 0x0
    "00000000", -- 5397 - 0x1515  :    0 - 0x0
    "00000000", -- 5398 - 0x1516  :    0 - 0x0
    "00000000", -- 5399 - 0x1517  :    0 - 0x0
    "00000000", -- 5400 - 0x1518  :    0 - 0x0
    "00000000", -- 5401 - 0x1519  :    0 - 0x0
    "00000000", -- 5402 - 0x151a  :    0 - 0x0
    "00000000", -- 5403 - 0x151b  :    0 - 0x0
    "00000000", -- 5404 - 0x151c  :    0 - 0x0
    "00000000", -- 5405 - 0x151d  :    0 - 0x0
    "00000000", -- 5406 - 0x151e  :    0 - 0x0
    "00000000", -- 5407 - 0x151f  :    0 - 0x0
    "00000000", -- 5408 - 0x1520  :    0 - 0x0 -- Background 0x52
    "00000000", -- 5409 - 0x1521  :    0 - 0x0
    "00000000", -- 5410 - 0x1522  :    0 - 0x0
    "00000000", -- 5411 - 0x1523  :    0 - 0x0
    "00000000", -- 5412 - 0x1524  :    0 - 0x0
    "00000000", -- 5413 - 0x1525  :    0 - 0x0
    "00000000", -- 5414 - 0x1526  :    0 - 0x0
    "00000000", -- 5415 - 0x1527  :    0 - 0x0
    "00000000", -- 5416 - 0x1528  :    0 - 0x0
    "00000000", -- 5417 - 0x1529  :    0 - 0x0
    "00000000", -- 5418 - 0x152a  :    0 - 0x0
    "00000000", -- 5419 - 0x152b  :    0 - 0x0
    "00000000", -- 5420 - 0x152c  :    0 - 0x0
    "00000000", -- 5421 - 0x152d  :    0 - 0x0
    "00000000", -- 5422 - 0x152e  :    0 - 0x0
    "00000000", -- 5423 - 0x152f  :    0 - 0x0
    "00000000", -- 5424 - 0x1530  :    0 - 0x0 -- Background 0x53
    "00000000", -- 5425 - 0x1531  :    0 - 0x0
    "00000000", -- 5426 - 0x1532  :    0 - 0x0
    "00000000", -- 5427 - 0x1533  :    0 - 0x0
    "00000000", -- 5428 - 0x1534  :    0 - 0x0
    "00000000", -- 5429 - 0x1535  :    0 - 0x0
    "00000000", -- 5430 - 0x1536  :    0 - 0x0
    "00000000", -- 5431 - 0x1537  :    0 - 0x0
    "00000000", -- 5432 - 0x1538  :    0 - 0x0
    "00000000", -- 5433 - 0x1539  :    0 - 0x0
    "00000000", -- 5434 - 0x153a  :    0 - 0x0
    "00000000", -- 5435 - 0x153b  :    0 - 0x0
    "00000000", -- 5436 - 0x153c  :    0 - 0x0
    "00000000", -- 5437 - 0x153d  :    0 - 0x0
    "00000000", -- 5438 - 0x153e  :    0 - 0x0
    "00000000", -- 5439 - 0x153f  :    0 - 0x0
    "00000000", -- 5440 - 0x1540  :    0 - 0x0 -- Background 0x54
    "00000000", -- 5441 - 0x1541  :    0 - 0x0
    "00000000", -- 5442 - 0x1542  :    0 - 0x0
    "00000000", -- 5443 - 0x1543  :    0 - 0x0
    "00000000", -- 5444 - 0x1544  :    0 - 0x0
    "00000000", -- 5445 - 0x1545  :    0 - 0x0
    "00000000", -- 5446 - 0x1546  :    0 - 0x0
    "00000000", -- 5447 - 0x1547  :    0 - 0x0
    "00000000", -- 5448 - 0x1548  :    0 - 0x0
    "00000000", -- 5449 - 0x1549  :    0 - 0x0
    "00000000", -- 5450 - 0x154a  :    0 - 0x0
    "00000000", -- 5451 - 0x154b  :    0 - 0x0
    "00000000", -- 5452 - 0x154c  :    0 - 0x0
    "00000000", -- 5453 - 0x154d  :    0 - 0x0
    "00000000", -- 5454 - 0x154e  :    0 - 0x0
    "00000000", -- 5455 - 0x154f  :    0 - 0x0
    "00000000", -- 5456 - 0x1550  :    0 - 0x0 -- Background 0x55
    "00000000", -- 5457 - 0x1551  :    0 - 0x0
    "00000000", -- 5458 - 0x1552  :    0 - 0x0
    "00000000", -- 5459 - 0x1553  :    0 - 0x0
    "00000000", -- 5460 - 0x1554  :    0 - 0x0
    "00000000", -- 5461 - 0x1555  :    0 - 0x0
    "00000000", -- 5462 - 0x1556  :    0 - 0x0
    "00000000", -- 5463 - 0x1557  :    0 - 0x0
    "00000000", -- 5464 - 0x1558  :    0 - 0x0
    "00000000", -- 5465 - 0x1559  :    0 - 0x0
    "00000000", -- 5466 - 0x155a  :    0 - 0x0
    "00000000", -- 5467 - 0x155b  :    0 - 0x0
    "00000000", -- 5468 - 0x155c  :    0 - 0x0
    "00000000", -- 5469 - 0x155d  :    0 - 0x0
    "00000000", -- 5470 - 0x155e  :    0 - 0x0
    "00000000", -- 5471 - 0x155f  :    0 - 0x0
    "00000000", -- 5472 - 0x1560  :    0 - 0x0 -- Background 0x56
    "00000000", -- 5473 - 0x1561  :    0 - 0x0
    "00000000", -- 5474 - 0x1562  :    0 - 0x0
    "00000000", -- 5475 - 0x1563  :    0 - 0x0
    "00000000", -- 5476 - 0x1564  :    0 - 0x0
    "00000000", -- 5477 - 0x1565  :    0 - 0x0
    "00000000", -- 5478 - 0x1566  :    0 - 0x0
    "00000000", -- 5479 - 0x1567  :    0 - 0x0
    "00000000", -- 5480 - 0x1568  :    0 - 0x0
    "00000000", -- 5481 - 0x1569  :    0 - 0x0
    "00000000", -- 5482 - 0x156a  :    0 - 0x0
    "00000000", -- 5483 - 0x156b  :    0 - 0x0
    "00000000", -- 5484 - 0x156c  :    0 - 0x0
    "00000000", -- 5485 - 0x156d  :    0 - 0x0
    "00000000", -- 5486 - 0x156e  :    0 - 0x0
    "00000000", -- 5487 - 0x156f  :    0 - 0x0
    "00000000", -- 5488 - 0x1570  :    0 - 0x0 -- Background 0x57
    "00000000", -- 5489 - 0x1571  :    0 - 0x0
    "00000000", -- 5490 - 0x1572  :    0 - 0x0
    "00000000", -- 5491 - 0x1573  :    0 - 0x0
    "00000000", -- 5492 - 0x1574  :    0 - 0x0
    "00000000", -- 5493 - 0x1575  :    0 - 0x0
    "00000000", -- 5494 - 0x1576  :    0 - 0x0
    "00000000", -- 5495 - 0x1577  :    0 - 0x0
    "00000000", -- 5496 - 0x1578  :    0 - 0x0
    "00000000", -- 5497 - 0x1579  :    0 - 0x0
    "00000000", -- 5498 - 0x157a  :    0 - 0x0
    "00000000", -- 5499 - 0x157b  :    0 - 0x0
    "00000000", -- 5500 - 0x157c  :    0 - 0x0
    "00000000", -- 5501 - 0x157d  :    0 - 0x0
    "00000000", -- 5502 - 0x157e  :    0 - 0x0
    "00000000", -- 5503 - 0x157f  :    0 - 0x0
    "00000000", -- 5504 - 0x1580  :    0 - 0x0 -- Background 0x58
    "00000000", -- 5505 - 0x1581  :    0 - 0x0
    "00000000", -- 5506 - 0x1582  :    0 - 0x0
    "00000000", -- 5507 - 0x1583  :    0 - 0x0
    "00000000", -- 5508 - 0x1584  :    0 - 0x0
    "00000000", -- 5509 - 0x1585  :    0 - 0x0
    "00000000", -- 5510 - 0x1586  :    0 - 0x0
    "00000000", -- 5511 - 0x1587  :    0 - 0x0
    "00000000", -- 5512 - 0x1588  :    0 - 0x0
    "00000000", -- 5513 - 0x1589  :    0 - 0x0
    "00000000", -- 5514 - 0x158a  :    0 - 0x0
    "00000000", -- 5515 - 0x158b  :    0 - 0x0
    "00000000", -- 5516 - 0x158c  :    0 - 0x0
    "00000000", -- 5517 - 0x158d  :    0 - 0x0
    "00000000", -- 5518 - 0x158e  :    0 - 0x0
    "00000000", -- 5519 - 0x158f  :    0 - 0x0
    "00000000", -- 5520 - 0x1590  :    0 - 0x0 -- Background 0x59
    "00000000", -- 5521 - 0x1591  :    0 - 0x0
    "00000000", -- 5522 - 0x1592  :    0 - 0x0
    "00000000", -- 5523 - 0x1593  :    0 - 0x0
    "00000000", -- 5524 - 0x1594  :    0 - 0x0
    "00000000", -- 5525 - 0x1595  :    0 - 0x0
    "00000000", -- 5526 - 0x1596  :    0 - 0x0
    "00000000", -- 5527 - 0x1597  :    0 - 0x0
    "00000000", -- 5528 - 0x1598  :    0 - 0x0
    "00000000", -- 5529 - 0x1599  :    0 - 0x0
    "00000000", -- 5530 - 0x159a  :    0 - 0x0
    "00000000", -- 5531 - 0x159b  :    0 - 0x0
    "00000000", -- 5532 - 0x159c  :    0 - 0x0
    "00000000", -- 5533 - 0x159d  :    0 - 0x0
    "00000000", -- 5534 - 0x159e  :    0 - 0x0
    "00000000", -- 5535 - 0x159f  :    0 - 0x0
    "00000000", -- 5536 - 0x15a0  :    0 - 0x0 -- Background 0x5a
    "00000000", -- 5537 - 0x15a1  :    0 - 0x0
    "00000000", -- 5538 - 0x15a2  :    0 - 0x0
    "00000000", -- 5539 - 0x15a3  :    0 - 0x0
    "00000000", -- 5540 - 0x15a4  :    0 - 0x0
    "00000000", -- 5541 - 0x15a5  :    0 - 0x0
    "00000000", -- 5542 - 0x15a6  :    0 - 0x0
    "00000000", -- 5543 - 0x15a7  :    0 - 0x0
    "00000000", -- 5544 - 0x15a8  :    0 - 0x0
    "00000000", -- 5545 - 0x15a9  :    0 - 0x0
    "00000000", -- 5546 - 0x15aa  :    0 - 0x0
    "00000000", -- 5547 - 0x15ab  :    0 - 0x0
    "00000000", -- 5548 - 0x15ac  :    0 - 0x0
    "00000000", -- 5549 - 0x15ad  :    0 - 0x0
    "00000000", -- 5550 - 0x15ae  :    0 - 0x0
    "00000000", -- 5551 - 0x15af  :    0 - 0x0
    "00000000", -- 5552 - 0x15b0  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 5553 - 0x15b1  :    0 - 0x0
    "00000000", -- 5554 - 0x15b2  :    0 - 0x0
    "00000000", -- 5555 - 0x15b3  :    0 - 0x0
    "00000000", -- 5556 - 0x15b4  :    0 - 0x0
    "00000000", -- 5557 - 0x15b5  :    0 - 0x0
    "00000000", -- 5558 - 0x15b6  :    0 - 0x0
    "00000000", -- 5559 - 0x15b7  :    0 - 0x0
    "00000000", -- 5560 - 0x15b8  :    0 - 0x0
    "00000000", -- 5561 - 0x15b9  :    0 - 0x0
    "00000000", -- 5562 - 0x15ba  :    0 - 0x0
    "00000000", -- 5563 - 0x15bb  :    0 - 0x0
    "00000000", -- 5564 - 0x15bc  :    0 - 0x0
    "00000000", -- 5565 - 0x15bd  :    0 - 0x0
    "00000000", -- 5566 - 0x15be  :    0 - 0x0
    "00000000", -- 5567 - 0x15bf  :    0 - 0x0
    "00000000", -- 5568 - 0x15c0  :    0 - 0x0 -- Background 0x5c
    "00000000", -- 5569 - 0x15c1  :    0 - 0x0
    "00000000", -- 5570 - 0x15c2  :    0 - 0x0
    "00000000", -- 5571 - 0x15c3  :    0 - 0x0
    "00000000", -- 5572 - 0x15c4  :    0 - 0x0
    "00000000", -- 5573 - 0x15c5  :    0 - 0x0
    "00000000", -- 5574 - 0x15c6  :    0 - 0x0
    "00000000", -- 5575 - 0x15c7  :    0 - 0x0
    "00000000", -- 5576 - 0x15c8  :    0 - 0x0
    "00000000", -- 5577 - 0x15c9  :    0 - 0x0
    "00000000", -- 5578 - 0x15ca  :    0 - 0x0
    "00000000", -- 5579 - 0x15cb  :    0 - 0x0
    "00000000", -- 5580 - 0x15cc  :    0 - 0x0
    "00000000", -- 5581 - 0x15cd  :    0 - 0x0
    "00000000", -- 5582 - 0x15ce  :    0 - 0x0
    "00000000", -- 5583 - 0x15cf  :    0 - 0x0
    "00000000", -- 5584 - 0x15d0  :    0 - 0x0 -- Background 0x5d
    "00000000", -- 5585 - 0x15d1  :    0 - 0x0
    "00000000", -- 5586 - 0x15d2  :    0 - 0x0
    "00000000", -- 5587 - 0x15d3  :    0 - 0x0
    "00000000", -- 5588 - 0x15d4  :    0 - 0x0
    "00000000", -- 5589 - 0x15d5  :    0 - 0x0
    "00000000", -- 5590 - 0x15d6  :    0 - 0x0
    "00000000", -- 5591 - 0x15d7  :    0 - 0x0
    "00000000", -- 5592 - 0x15d8  :    0 - 0x0
    "00000000", -- 5593 - 0x15d9  :    0 - 0x0
    "00000000", -- 5594 - 0x15da  :    0 - 0x0
    "00000000", -- 5595 - 0x15db  :    0 - 0x0
    "00000000", -- 5596 - 0x15dc  :    0 - 0x0
    "00000000", -- 5597 - 0x15dd  :    0 - 0x0
    "00000000", -- 5598 - 0x15de  :    0 - 0x0
    "00000000", -- 5599 - 0x15df  :    0 - 0x0
    "00000000", -- 5600 - 0x15e0  :    0 - 0x0 -- Background 0x5e
    "00000000", -- 5601 - 0x15e1  :    0 - 0x0
    "00000000", -- 5602 - 0x15e2  :    0 - 0x0
    "00000000", -- 5603 - 0x15e3  :    0 - 0x0
    "00000000", -- 5604 - 0x15e4  :    0 - 0x0
    "00000000", -- 5605 - 0x15e5  :    0 - 0x0
    "00000000", -- 5606 - 0x15e6  :    0 - 0x0
    "00000000", -- 5607 - 0x15e7  :    0 - 0x0
    "00000000", -- 5608 - 0x15e8  :    0 - 0x0
    "00000000", -- 5609 - 0x15e9  :    0 - 0x0
    "00000000", -- 5610 - 0x15ea  :    0 - 0x0
    "00000000", -- 5611 - 0x15eb  :    0 - 0x0
    "00000000", -- 5612 - 0x15ec  :    0 - 0x0
    "00000000", -- 5613 - 0x15ed  :    0 - 0x0
    "00000000", -- 5614 - 0x15ee  :    0 - 0x0
    "00000000", -- 5615 - 0x15ef  :    0 - 0x0
    "00000000", -- 5616 - 0x15f0  :    0 - 0x0 -- Background 0x5f
    "00000000", -- 5617 - 0x15f1  :    0 - 0x0
    "00000000", -- 5618 - 0x15f2  :    0 - 0x0
    "00000000", -- 5619 - 0x15f3  :    0 - 0x0
    "00000000", -- 5620 - 0x15f4  :    0 - 0x0
    "00000000", -- 5621 - 0x15f5  :    0 - 0x0
    "00000000", -- 5622 - 0x15f6  :    0 - 0x0
    "00000000", -- 5623 - 0x15f7  :    0 - 0x0
    "00000000", -- 5624 - 0x15f8  :    0 - 0x0
    "00000000", -- 5625 - 0x15f9  :    0 - 0x0
    "00000000", -- 5626 - 0x15fa  :    0 - 0x0
    "00000000", -- 5627 - 0x15fb  :    0 - 0x0
    "00000000", -- 5628 - 0x15fc  :    0 - 0x0
    "00000000", -- 5629 - 0x15fd  :    0 - 0x0
    "00000000", -- 5630 - 0x15fe  :    0 - 0x0
    "00000000", -- 5631 - 0x15ff  :    0 - 0x0
    "00000000", -- 5632 - 0x1600  :    0 - 0x0 -- Background 0x60
    "00000000", -- 5633 - 0x1601  :    0 - 0x0
    "00000000", -- 5634 - 0x1602  :    0 - 0x0
    "00000000", -- 5635 - 0x1603  :    0 - 0x0
    "00000000", -- 5636 - 0x1604  :    0 - 0x0
    "00000000", -- 5637 - 0x1605  :    0 - 0x0
    "00000000", -- 5638 - 0x1606  :    0 - 0x0
    "00000000", -- 5639 - 0x1607  :    0 - 0x0
    "00000000", -- 5640 - 0x1608  :    0 - 0x0
    "00000000", -- 5641 - 0x1609  :    0 - 0x0
    "00000000", -- 5642 - 0x160a  :    0 - 0x0
    "00000000", -- 5643 - 0x160b  :    0 - 0x0
    "00000000", -- 5644 - 0x160c  :    0 - 0x0
    "00000000", -- 5645 - 0x160d  :    0 - 0x0
    "00000000", -- 5646 - 0x160e  :    0 - 0x0
    "00000000", -- 5647 - 0x160f  :    0 - 0x0
    "00000000", -- 5648 - 0x1610  :    0 - 0x0 -- Background 0x61
    "00000000", -- 5649 - 0x1611  :    0 - 0x0
    "00000000", -- 5650 - 0x1612  :    0 - 0x0
    "00000000", -- 5651 - 0x1613  :    0 - 0x0
    "00000000", -- 5652 - 0x1614  :    0 - 0x0
    "00000000", -- 5653 - 0x1615  :    0 - 0x0
    "00000000", -- 5654 - 0x1616  :    0 - 0x0
    "00000000", -- 5655 - 0x1617  :    0 - 0x0
    "00000000", -- 5656 - 0x1618  :    0 - 0x0
    "00000000", -- 5657 - 0x1619  :    0 - 0x0
    "00000000", -- 5658 - 0x161a  :    0 - 0x0
    "00000000", -- 5659 - 0x161b  :    0 - 0x0
    "00000000", -- 5660 - 0x161c  :    0 - 0x0
    "00000000", -- 5661 - 0x161d  :    0 - 0x0
    "00000000", -- 5662 - 0x161e  :    0 - 0x0
    "00000000", -- 5663 - 0x161f  :    0 - 0x0
    "00000000", -- 5664 - 0x1620  :    0 - 0x0 -- Background 0x62
    "00000000", -- 5665 - 0x1621  :    0 - 0x0
    "00000000", -- 5666 - 0x1622  :    0 - 0x0
    "00000000", -- 5667 - 0x1623  :    0 - 0x0
    "00000000", -- 5668 - 0x1624  :    0 - 0x0
    "00000000", -- 5669 - 0x1625  :    0 - 0x0
    "00000000", -- 5670 - 0x1626  :    0 - 0x0
    "00000000", -- 5671 - 0x1627  :    0 - 0x0
    "00000000", -- 5672 - 0x1628  :    0 - 0x0
    "00000000", -- 5673 - 0x1629  :    0 - 0x0
    "00000000", -- 5674 - 0x162a  :    0 - 0x0
    "00000000", -- 5675 - 0x162b  :    0 - 0x0
    "00000000", -- 5676 - 0x162c  :    0 - 0x0
    "00000000", -- 5677 - 0x162d  :    0 - 0x0
    "00000000", -- 5678 - 0x162e  :    0 - 0x0
    "00000000", -- 5679 - 0x162f  :    0 - 0x0
    "00000000", -- 5680 - 0x1630  :    0 - 0x0 -- Background 0x63
    "00000000", -- 5681 - 0x1631  :    0 - 0x0
    "00000000", -- 5682 - 0x1632  :    0 - 0x0
    "00000000", -- 5683 - 0x1633  :    0 - 0x0
    "00000000", -- 5684 - 0x1634  :    0 - 0x0
    "00000000", -- 5685 - 0x1635  :    0 - 0x0
    "00000000", -- 5686 - 0x1636  :    0 - 0x0
    "00000000", -- 5687 - 0x1637  :    0 - 0x0
    "00000000", -- 5688 - 0x1638  :    0 - 0x0
    "00000000", -- 5689 - 0x1639  :    0 - 0x0
    "00000000", -- 5690 - 0x163a  :    0 - 0x0
    "00000000", -- 5691 - 0x163b  :    0 - 0x0
    "00000000", -- 5692 - 0x163c  :    0 - 0x0
    "00000000", -- 5693 - 0x163d  :    0 - 0x0
    "00000000", -- 5694 - 0x163e  :    0 - 0x0
    "00000000", -- 5695 - 0x163f  :    0 - 0x0
    "00000000", -- 5696 - 0x1640  :    0 - 0x0 -- Background 0x64
    "00000000", -- 5697 - 0x1641  :    0 - 0x0
    "00000000", -- 5698 - 0x1642  :    0 - 0x0
    "00000000", -- 5699 - 0x1643  :    0 - 0x0
    "00000000", -- 5700 - 0x1644  :    0 - 0x0
    "00000000", -- 5701 - 0x1645  :    0 - 0x0
    "00000000", -- 5702 - 0x1646  :    0 - 0x0
    "00000000", -- 5703 - 0x1647  :    0 - 0x0
    "00000000", -- 5704 - 0x1648  :    0 - 0x0
    "00000000", -- 5705 - 0x1649  :    0 - 0x0
    "00000000", -- 5706 - 0x164a  :    0 - 0x0
    "00000000", -- 5707 - 0x164b  :    0 - 0x0
    "00000000", -- 5708 - 0x164c  :    0 - 0x0
    "00000000", -- 5709 - 0x164d  :    0 - 0x0
    "00000000", -- 5710 - 0x164e  :    0 - 0x0
    "00000000", -- 5711 - 0x164f  :    0 - 0x0
    "00000000", -- 5712 - 0x1650  :    0 - 0x0 -- Background 0x65
    "00000000", -- 5713 - 0x1651  :    0 - 0x0
    "00000000", -- 5714 - 0x1652  :    0 - 0x0
    "00000000", -- 5715 - 0x1653  :    0 - 0x0
    "00000000", -- 5716 - 0x1654  :    0 - 0x0
    "00000000", -- 5717 - 0x1655  :    0 - 0x0
    "00000000", -- 5718 - 0x1656  :    0 - 0x0
    "00000000", -- 5719 - 0x1657  :    0 - 0x0
    "00000000", -- 5720 - 0x1658  :    0 - 0x0
    "00000000", -- 5721 - 0x1659  :    0 - 0x0
    "00000000", -- 5722 - 0x165a  :    0 - 0x0
    "00000000", -- 5723 - 0x165b  :    0 - 0x0
    "00000000", -- 5724 - 0x165c  :    0 - 0x0
    "00000000", -- 5725 - 0x165d  :    0 - 0x0
    "00000000", -- 5726 - 0x165e  :    0 - 0x0
    "00000000", -- 5727 - 0x165f  :    0 - 0x0
    "00000000", -- 5728 - 0x1660  :    0 - 0x0 -- Background 0x66
    "00000000", -- 5729 - 0x1661  :    0 - 0x0
    "00000000", -- 5730 - 0x1662  :    0 - 0x0
    "00000000", -- 5731 - 0x1663  :    0 - 0x0
    "00000000", -- 5732 - 0x1664  :    0 - 0x0
    "00000000", -- 5733 - 0x1665  :    0 - 0x0
    "00000000", -- 5734 - 0x1666  :    0 - 0x0
    "00000000", -- 5735 - 0x1667  :    0 - 0x0
    "00000000", -- 5736 - 0x1668  :    0 - 0x0
    "00000000", -- 5737 - 0x1669  :    0 - 0x0
    "00000000", -- 5738 - 0x166a  :    0 - 0x0
    "00000000", -- 5739 - 0x166b  :    0 - 0x0
    "00000000", -- 5740 - 0x166c  :    0 - 0x0
    "00000000", -- 5741 - 0x166d  :    0 - 0x0
    "00000000", -- 5742 - 0x166e  :    0 - 0x0
    "00000000", -- 5743 - 0x166f  :    0 - 0x0
    "00000000", -- 5744 - 0x1670  :    0 - 0x0 -- Background 0x67
    "00000000", -- 5745 - 0x1671  :    0 - 0x0
    "00000000", -- 5746 - 0x1672  :    0 - 0x0
    "00000000", -- 5747 - 0x1673  :    0 - 0x0
    "00000000", -- 5748 - 0x1674  :    0 - 0x0
    "00000000", -- 5749 - 0x1675  :    0 - 0x0
    "00000000", -- 5750 - 0x1676  :    0 - 0x0
    "00000000", -- 5751 - 0x1677  :    0 - 0x0
    "00000000", -- 5752 - 0x1678  :    0 - 0x0
    "00000000", -- 5753 - 0x1679  :    0 - 0x0
    "00000000", -- 5754 - 0x167a  :    0 - 0x0
    "00000000", -- 5755 - 0x167b  :    0 - 0x0
    "00000000", -- 5756 - 0x167c  :    0 - 0x0
    "00000000", -- 5757 - 0x167d  :    0 - 0x0
    "00000000", -- 5758 - 0x167e  :    0 - 0x0
    "00000000", -- 5759 - 0x167f  :    0 - 0x0
    "00000000", -- 5760 - 0x1680  :    0 - 0x0 -- Background 0x68
    "00000000", -- 5761 - 0x1681  :    0 - 0x0
    "00000000", -- 5762 - 0x1682  :    0 - 0x0
    "00000000", -- 5763 - 0x1683  :    0 - 0x0
    "00000000", -- 5764 - 0x1684  :    0 - 0x0
    "00000000", -- 5765 - 0x1685  :    0 - 0x0
    "00000000", -- 5766 - 0x1686  :    0 - 0x0
    "00000000", -- 5767 - 0x1687  :    0 - 0x0
    "00000000", -- 5768 - 0x1688  :    0 - 0x0
    "00000000", -- 5769 - 0x1689  :    0 - 0x0
    "00000000", -- 5770 - 0x168a  :    0 - 0x0
    "00000000", -- 5771 - 0x168b  :    0 - 0x0
    "00000000", -- 5772 - 0x168c  :    0 - 0x0
    "00000000", -- 5773 - 0x168d  :    0 - 0x0
    "00000000", -- 5774 - 0x168e  :    0 - 0x0
    "00000000", -- 5775 - 0x168f  :    0 - 0x0
    "00000000", -- 5776 - 0x1690  :    0 - 0x0 -- Background 0x69
    "00000000", -- 5777 - 0x1691  :    0 - 0x0
    "00000000", -- 5778 - 0x1692  :    0 - 0x0
    "00000000", -- 5779 - 0x1693  :    0 - 0x0
    "00000000", -- 5780 - 0x1694  :    0 - 0x0
    "00000000", -- 5781 - 0x1695  :    0 - 0x0
    "00000000", -- 5782 - 0x1696  :    0 - 0x0
    "00000000", -- 5783 - 0x1697  :    0 - 0x0
    "00000000", -- 5784 - 0x1698  :    0 - 0x0
    "00000000", -- 5785 - 0x1699  :    0 - 0x0
    "00000000", -- 5786 - 0x169a  :    0 - 0x0
    "00000000", -- 5787 - 0x169b  :    0 - 0x0
    "00000000", -- 5788 - 0x169c  :    0 - 0x0
    "00000000", -- 5789 - 0x169d  :    0 - 0x0
    "00000000", -- 5790 - 0x169e  :    0 - 0x0
    "00000000", -- 5791 - 0x169f  :    0 - 0x0
    "00000000", -- 5792 - 0x16a0  :    0 - 0x0 -- Background 0x6a
    "00000000", -- 5793 - 0x16a1  :    0 - 0x0
    "00000000", -- 5794 - 0x16a2  :    0 - 0x0
    "00000000", -- 5795 - 0x16a3  :    0 - 0x0
    "00000000", -- 5796 - 0x16a4  :    0 - 0x0
    "00000000", -- 5797 - 0x16a5  :    0 - 0x0
    "00000000", -- 5798 - 0x16a6  :    0 - 0x0
    "00000000", -- 5799 - 0x16a7  :    0 - 0x0
    "00000000", -- 5800 - 0x16a8  :    0 - 0x0
    "00000000", -- 5801 - 0x16a9  :    0 - 0x0
    "00000000", -- 5802 - 0x16aa  :    0 - 0x0
    "00000000", -- 5803 - 0x16ab  :    0 - 0x0
    "00000000", -- 5804 - 0x16ac  :    0 - 0x0
    "00000000", -- 5805 - 0x16ad  :    0 - 0x0
    "00000000", -- 5806 - 0x16ae  :    0 - 0x0
    "00000000", -- 5807 - 0x16af  :    0 - 0x0
    "00000000", -- 5808 - 0x16b0  :    0 - 0x0 -- Background 0x6b
    "00000000", -- 5809 - 0x16b1  :    0 - 0x0
    "00000000", -- 5810 - 0x16b2  :    0 - 0x0
    "00000000", -- 5811 - 0x16b3  :    0 - 0x0
    "00000000", -- 5812 - 0x16b4  :    0 - 0x0
    "00000000", -- 5813 - 0x16b5  :    0 - 0x0
    "00000000", -- 5814 - 0x16b6  :    0 - 0x0
    "00000000", -- 5815 - 0x16b7  :    0 - 0x0
    "00000000", -- 5816 - 0x16b8  :    0 - 0x0
    "00000000", -- 5817 - 0x16b9  :    0 - 0x0
    "00000000", -- 5818 - 0x16ba  :    0 - 0x0
    "00000000", -- 5819 - 0x16bb  :    0 - 0x0
    "00000000", -- 5820 - 0x16bc  :    0 - 0x0
    "00000000", -- 5821 - 0x16bd  :    0 - 0x0
    "00000000", -- 5822 - 0x16be  :    0 - 0x0
    "00000000", -- 5823 - 0x16bf  :    0 - 0x0
    "00000000", -- 5824 - 0x16c0  :    0 - 0x0 -- Background 0x6c
    "00000000", -- 5825 - 0x16c1  :    0 - 0x0
    "00000000", -- 5826 - 0x16c2  :    0 - 0x0
    "00000000", -- 5827 - 0x16c3  :    0 - 0x0
    "00000000", -- 5828 - 0x16c4  :    0 - 0x0
    "00000000", -- 5829 - 0x16c5  :    0 - 0x0
    "00000000", -- 5830 - 0x16c6  :    0 - 0x0
    "00000000", -- 5831 - 0x16c7  :    0 - 0x0
    "00000000", -- 5832 - 0x16c8  :    0 - 0x0
    "00000000", -- 5833 - 0x16c9  :    0 - 0x0
    "00000000", -- 5834 - 0x16ca  :    0 - 0x0
    "00000000", -- 5835 - 0x16cb  :    0 - 0x0
    "00000000", -- 5836 - 0x16cc  :    0 - 0x0
    "00000000", -- 5837 - 0x16cd  :    0 - 0x0
    "00000000", -- 5838 - 0x16ce  :    0 - 0x0
    "00000000", -- 5839 - 0x16cf  :    0 - 0x0
    "00000000", -- 5840 - 0x16d0  :    0 - 0x0 -- Background 0x6d
    "00000000", -- 5841 - 0x16d1  :    0 - 0x0
    "00000000", -- 5842 - 0x16d2  :    0 - 0x0
    "00000000", -- 5843 - 0x16d3  :    0 - 0x0
    "00000000", -- 5844 - 0x16d4  :    0 - 0x0
    "00000000", -- 5845 - 0x16d5  :    0 - 0x0
    "00000000", -- 5846 - 0x16d6  :    0 - 0x0
    "00000000", -- 5847 - 0x16d7  :    0 - 0x0
    "00000000", -- 5848 - 0x16d8  :    0 - 0x0
    "00000000", -- 5849 - 0x16d9  :    0 - 0x0
    "00000000", -- 5850 - 0x16da  :    0 - 0x0
    "00000000", -- 5851 - 0x16db  :    0 - 0x0
    "00000000", -- 5852 - 0x16dc  :    0 - 0x0
    "00000000", -- 5853 - 0x16dd  :    0 - 0x0
    "00000000", -- 5854 - 0x16de  :    0 - 0x0
    "00000000", -- 5855 - 0x16df  :    0 - 0x0
    "00000000", -- 5856 - 0x16e0  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 5857 - 0x16e1  :    0 - 0x0
    "00000000", -- 5858 - 0x16e2  :    0 - 0x0
    "00000000", -- 5859 - 0x16e3  :    0 - 0x0
    "00000000", -- 5860 - 0x16e4  :    0 - 0x0
    "00000000", -- 5861 - 0x16e5  :    0 - 0x0
    "00000000", -- 5862 - 0x16e6  :    0 - 0x0
    "00000000", -- 5863 - 0x16e7  :    0 - 0x0
    "00000000", -- 5864 - 0x16e8  :    0 - 0x0
    "00000000", -- 5865 - 0x16e9  :    0 - 0x0
    "00000000", -- 5866 - 0x16ea  :    0 - 0x0
    "00000000", -- 5867 - 0x16eb  :    0 - 0x0
    "00000000", -- 5868 - 0x16ec  :    0 - 0x0
    "00000000", -- 5869 - 0x16ed  :    0 - 0x0
    "00000000", -- 5870 - 0x16ee  :    0 - 0x0
    "00000000", -- 5871 - 0x16ef  :    0 - 0x0
    "00000000", -- 5872 - 0x16f0  :    0 - 0x0 -- Background 0x6f
    "00000000", -- 5873 - 0x16f1  :    0 - 0x0
    "00000000", -- 5874 - 0x16f2  :    0 - 0x0
    "00000000", -- 5875 - 0x16f3  :    0 - 0x0
    "00000000", -- 5876 - 0x16f4  :    0 - 0x0
    "00000000", -- 5877 - 0x16f5  :    0 - 0x0
    "00000000", -- 5878 - 0x16f6  :    0 - 0x0
    "00000000", -- 5879 - 0x16f7  :    0 - 0x0
    "00000000", -- 5880 - 0x16f8  :    0 - 0x0
    "00000000", -- 5881 - 0x16f9  :    0 - 0x0
    "00000000", -- 5882 - 0x16fa  :    0 - 0x0
    "00000000", -- 5883 - 0x16fb  :    0 - 0x0
    "00000000", -- 5884 - 0x16fc  :    0 - 0x0
    "00000000", -- 5885 - 0x16fd  :    0 - 0x0
    "00000000", -- 5886 - 0x16fe  :    0 - 0x0
    "00000000", -- 5887 - 0x16ff  :    0 - 0x0
    "00000000", -- 5888 - 0x1700  :    0 - 0x0 -- Background 0x70
    "00000000", -- 5889 - 0x1701  :    0 - 0x0
    "00000000", -- 5890 - 0x1702  :    0 - 0x0
    "00000000", -- 5891 - 0x1703  :    0 - 0x0
    "00000000", -- 5892 - 0x1704  :    0 - 0x0
    "00000000", -- 5893 - 0x1705  :    0 - 0x0
    "00000000", -- 5894 - 0x1706  :    0 - 0x0
    "00000000", -- 5895 - 0x1707  :    0 - 0x0
    "00000000", -- 5896 - 0x1708  :    0 - 0x0
    "00000000", -- 5897 - 0x1709  :    0 - 0x0
    "00000000", -- 5898 - 0x170a  :    0 - 0x0
    "00000000", -- 5899 - 0x170b  :    0 - 0x0
    "00000000", -- 5900 - 0x170c  :    0 - 0x0
    "00000000", -- 5901 - 0x170d  :    0 - 0x0
    "00000000", -- 5902 - 0x170e  :    0 - 0x0
    "00000000", -- 5903 - 0x170f  :    0 - 0x0
    "00000000", -- 5904 - 0x1710  :    0 - 0x0 -- Background 0x71
    "00000000", -- 5905 - 0x1711  :    0 - 0x0
    "00000000", -- 5906 - 0x1712  :    0 - 0x0
    "00000000", -- 5907 - 0x1713  :    0 - 0x0
    "00000000", -- 5908 - 0x1714  :    0 - 0x0
    "00000000", -- 5909 - 0x1715  :    0 - 0x0
    "00000000", -- 5910 - 0x1716  :    0 - 0x0
    "00000000", -- 5911 - 0x1717  :    0 - 0x0
    "00000000", -- 5912 - 0x1718  :    0 - 0x0
    "00000000", -- 5913 - 0x1719  :    0 - 0x0
    "00000000", -- 5914 - 0x171a  :    0 - 0x0
    "00000000", -- 5915 - 0x171b  :    0 - 0x0
    "00000000", -- 5916 - 0x171c  :    0 - 0x0
    "00000000", -- 5917 - 0x171d  :    0 - 0x0
    "00000000", -- 5918 - 0x171e  :    0 - 0x0
    "00000000", -- 5919 - 0x171f  :    0 - 0x0
    "00000000", -- 5920 - 0x1720  :    0 - 0x0 -- Background 0x72
    "00000000", -- 5921 - 0x1721  :    0 - 0x0
    "00000000", -- 5922 - 0x1722  :    0 - 0x0
    "00000000", -- 5923 - 0x1723  :    0 - 0x0
    "00000000", -- 5924 - 0x1724  :    0 - 0x0
    "00000000", -- 5925 - 0x1725  :    0 - 0x0
    "00000000", -- 5926 - 0x1726  :    0 - 0x0
    "00000000", -- 5927 - 0x1727  :    0 - 0x0
    "00000000", -- 5928 - 0x1728  :    0 - 0x0
    "00000000", -- 5929 - 0x1729  :    0 - 0x0
    "00000000", -- 5930 - 0x172a  :    0 - 0x0
    "00000000", -- 5931 - 0x172b  :    0 - 0x0
    "00000000", -- 5932 - 0x172c  :    0 - 0x0
    "00000000", -- 5933 - 0x172d  :    0 - 0x0
    "00000000", -- 5934 - 0x172e  :    0 - 0x0
    "00000000", -- 5935 - 0x172f  :    0 - 0x0
    "00000000", -- 5936 - 0x1730  :    0 - 0x0 -- Background 0x73
    "00000000", -- 5937 - 0x1731  :    0 - 0x0
    "00000000", -- 5938 - 0x1732  :    0 - 0x0
    "00000000", -- 5939 - 0x1733  :    0 - 0x0
    "00000000", -- 5940 - 0x1734  :    0 - 0x0
    "00000000", -- 5941 - 0x1735  :    0 - 0x0
    "00000000", -- 5942 - 0x1736  :    0 - 0x0
    "00000000", -- 5943 - 0x1737  :    0 - 0x0
    "00000000", -- 5944 - 0x1738  :    0 - 0x0
    "00000000", -- 5945 - 0x1739  :    0 - 0x0
    "00000000", -- 5946 - 0x173a  :    0 - 0x0
    "00000000", -- 5947 - 0x173b  :    0 - 0x0
    "00000000", -- 5948 - 0x173c  :    0 - 0x0
    "00000000", -- 5949 - 0x173d  :    0 - 0x0
    "00000000", -- 5950 - 0x173e  :    0 - 0x0
    "00000000", -- 5951 - 0x173f  :    0 - 0x0
    "00000000", -- 5952 - 0x1740  :    0 - 0x0 -- Background 0x74
    "00000000", -- 5953 - 0x1741  :    0 - 0x0
    "00000000", -- 5954 - 0x1742  :    0 - 0x0
    "00000000", -- 5955 - 0x1743  :    0 - 0x0
    "00000000", -- 5956 - 0x1744  :    0 - 0x0
    "00000000", -- 5957 - 0x1745  :    0 - 0x0
    "00000000", -- 5958 - 0x1746  :    0 - 0x0
    "00000000", -- 5959 - 0x1747  :    0 - 0x0
    "00000000", -- 5960 - 0x1748  :    0 - 0x0
    "00000000", -- 5961 - 0x1749  :    0 - 0x0
    "00000000", -- 5962 - 0x174a  :    0 - 0x0
    "00000000", -- 5963 - 0x174b  :    0 - 0x0
    "00000000", -- 5964 - 0x174c  :    0 - 0x0
    "00000000", -- 5965 - 0x174d  :    0 - 0x0
    "00000000", -- 5966 - 0x174e  :    0 - 0x0
    "00000000", -- 5967 - 0x174f  :    0 - 0x0
    "00000000", -- 5968 - 0x1750  :    0 - 0x0 -- Background 0x75
    "00000000", -- 5969 - 0x1751  :    0 - 0x0
    "00000000", -- 5970 - 0x1752  :    0 - 0x0
    "00000000", -- 5971 - 0x1753  :    0 - 0x0
    "00000000", -- 5972 - 0x1754  :    0 - 0x0
    "00000000", -- 5973 - 0x1755  :    0 - 0x0
    "00000000", -- 5974 - 0x1756  :    0 - 0x0
    "00000000", -- 5975 - 0x1757  :    0 - 0x0
    "00000000", -- 5976 - 0x1758  :    0 - 0x0
    "00000000", -- 5977 - 0x1759  :    0 - 0x0
    "00000000", -- 5978 - 0x175a  :    0 - 0x0
    "00000000", -- 5979 - 0x175b  :    0 - 0x0
    "00000000", -- 5980 - 0x175c  :    0 - 0x0
    "00000000", -- 5981 - 0x175d  :    0 - 0x0
    "00000000", -- 5982 - 0x175e  :    0 - 0x0
    "00000000", -- 5983 - 0x175f  :    0 - 0x0
    "00000000", -- 5984 - 0x1760  :    0 - 0x0 -- Background 0x76
    "00000000", -- 5985 - 0x1761  :    0 - 0x0
    "00000000", -- 5986 - 0x1762  :    0 - 0x0
    "00000000", -- 5987 - 0x1763  :    0 - 0x0
    "00000000", -- 5988 - 0x1764  :    0 - 0x0
    "00000000", -- 5989 - 0x1765  :    0 - 0x0
    "00000000", -- 5990 - 0x1766  :    0 - 0x0
    "00000000", -- 5991 - 0x1767  :    0 - 0x0
    "00000000", -- 5992 - 0x1768  :    0 - 0x0
    "00000000", -- 5993 - 0x1769  :    0 - 0x0
    "00000000", -- 5994 - 0x176a  :    0 - 0x0
    "00000000", -- 5995 - 0x176b  :    0 - 0x0
    "00000000", -- 5996 - 0x176c  :    0 - 0x0
    "00000000", -- 5997 - 0x176d  :    0 - 0x0
    "00000000", -- 5998 - 0x176e  :    0 - 0x0
    "00000000", -- 5999 - 0x176f  :    0 - 0x0
    "00000000", -- 6000 - 0x1770  :    0 - 0x0 -- Background 0x77
    "00000000", -- 6001 - 0x1771  :    0 - 0x0
    "00000000", -- 6002 - 0x1772  :    0 - 0x0
    "00000000", -- 6003 - 0x1773  :    0 - 0x0
    "00000000", -- 6004 - 0x1774  :    0 - 0x0
    "00000000", -- 6005 - 0x1775  :    0 - 0x0
    "00000000", -- 6006 - 0x1776  :    0 - 0x0
    "00000000", -- 6007 - 0x1777  :    0 - 0x0
    "00000000", -- 6008 - 0x1778  :    0 - 0x0
    "00000000", -- 6009 - 0x1779  :    0 - 0x0
    "00000000", -- 6010 - 0x177a  :    0 - 0x0
    "00000000", -- 6011 - 0x177b  :    0 - 0x0
    "00000000", -- 6012 - 0x177c  :    0 - 0x0
    "00000000", -- 6013 - 0x177d  :    0 - 0x0
    "00000000", -- 6014 - 0x177e  :    0 - 0x0
    "00000000", -- 6015 - 0x177f  :    0 - 0x0
    "00000000", -- 6016 - 0x1780  :    0 - 0x0 -- Background 0x78
    "00000000", -- 6017 - 0x1781  :    0 - 0x0
    "00000000", -- 6018 - 0x1782  :    0 - 0x0
    "00000000", -- 6019 - 0x1783  :    0 - 0x0
    "00000000", -- 6020 - 0x1784  :    0 - 0x0
    "00000000", -- 6021 - 0x1785  :    0 - 0x0
    "00000000", -- 6022 - 0x1786  :    0 - 0x0
    "00000000", -- 6023 - 0x1787  :    0 - 0x0
    "00000000", -- 6024 - 0x1788  :    0 - 0x0
    "00000000", -- 6025 - 0x1789  :    0 - 0x0
    "00000000", -- 6026 - 0x178a  :    0 - 0x0
    "00000000", -- 6027 - 0x178b  :    0 - 0x0
    "00000000", -- 6028 - 0x178c  :    0 - 0x0
    "00000000", -- 6029 - 0x178d  :    0 - 0x0
    "00000000", -- 6030 - 0x178e  :    0 - 0x0
    "00000000", -- 6031 - 0x178f  :    0 - 0x0
    "00000000", -- 6032 - 0x1790  :    0 - 0x0 -- Background 0x79
    "00000000", -- 6033 - 0x1791  :    0 - 0x0
    "00000000", -- 6034 - 0x1792  :    0 - 0x0
    "00000000", -- 6035 - 0x1793  :    0 - 0x0
    "00000000", -- 6036 - 0x1794  :    0 - 0x0
    "00000000", -- 6037 - 0x1795  :    0 - 0x0
    "00000000", -- 6038 - 0x1796  :    0 - 0x0
    "00000000", -- 6039 - 0x1797  :    0 - 0x0
    "00000000", -- 6040 - 0x1798  :    0 - 0x0
    "00000000", -- 6041 - 0x1799  :    0 - 0x0
    "00000000", -- 6042 - 0x179a  :    0 - 0x0
    "00000000", -- 6043 - 0x179b  :    0 - 0x0
    "00000000", -- 6044 - 0x179c  :    0 - 0x0
    "00000000", -- 6045 - 0x179d  :    0 - 0x0
    "00000000", -- 6046 - 0x179e  :    0 - 0x0
    "00000000", -- 6047 - 0x179f  :    0 - 0x0
    "00000000", -- 6048 - 0x17a0  :    0 - 0x0 -- Background 0x7a
    "00000000", -- 6049 - 0x17a1  :    0 - 0x0
    "00000000", -- 6050 - 0x17a2  :    0 - 0x0
    "00000000", -- 6051 - 0x17a3  :    0 - 0x0
    "00000000", -- 6052 - 0x17a4  :    0 - 0x0
    "00000000", -- 6053 - 0x17a5  :    0 - 0x0
    "00000000", -- 6054 - 0x17a6  :    0 - 0x0
    "00000000", -- 6055 - 0x17a7  :    0 - 0x0
    "00000000", -- 6056 - 0x17a8  :    0 - 0x0
    "00000000", -- 6057 - 0x17a9  :    0 - 0x0
    "00000000", -- 6058 - 0x17aa  :    0 - 0x0
    "00000000", -- 6059 - 0x17ab  :    0 - 0x0
    "00000000", -- 6060 - 0x17ac  :    0 - 0x0
    "00000000", -- 6061 - 0x17ad  :    0 - 0x0
    "00000000", -- 6062 - 0x17ae  :    0 - 0x0
    "00000000", -- 6063 - 0x17af  :    0 - 0x0
    "00000000", -- 6064 - 0x17b0  :    0 - 0x0 -- Background 0x7b
    "00000000", -- 6065 - 0x17b1  :    0 - 0x0
    "00000000", -- 6066 - 0x17b2  :    0 - 0x0
    "00000000", -- 6067 - 0x17b3  :    0 - 0x0
    "00000000", -- 6068 - 0x17b4  :    0 - 0x0
    "00000000", -- 6069 - 0x17b5  :    0 - 0x0
    "00000000", -- 6070 - 0x17b6  :    0 - 0x0
    "00000000", -- 6071 - 0x17b7  :    0 - 0x0
    "00000000", -- 6072 - 0x17b8  :    0 - 0x0
    "00000000", -- 6073 - 0x17b9  :    0 - 0x0
    "00000000", -- 6074 - 0x17ba  :    0 - 0x0
    "00000000", -- 6075 - 0x17bb  :    0 - 0x0
    "00000000", -- 6076 - 0x17bc  :    0 - 0x0
    "00000000", -- 6077 - 0x17bd  :    0 - 0x0
    "00000000", -- 6078 - 0x17be  :    0 - 0x0
    "00000000", -- 6079 - 0x17bf  :    0 - 0x0
    "00000000", -- 6080 - 0x17c0  :    0 - 0x0 -- Background 0x7c
    "00000000", -- 6081 - 0x17c1  :    0 - 0x0
    "00000000", -- 6082 - 0x17c2  :    0 - 0x0
    "00000000", -- 6083 - 0x17c3  :    0 - 0x0
    "00000000", -- 6084 - 0x17c4  :    0 - 0x0
    "00000000", -- 6085 - 0x17c5  :    0 - 0x0
    "00000000", -- 6086 - 0x17c6  :    0 - 0x0
    "00000000", -- 6087 - 0x17c7  :    0 - 0x0
    "00000000", -- 6088 - 0x17c8  :    0 - 0x0
    "00000000", -- 6089 - 0x17c9  :    0 - 0x0
    "00000000", -- 6090 - 0x17ca  :    0 - 0x0
    "00000000", -- 6091 - 0x17cb  :    0 - 0x0
    "00000000", -- 6092 - 0x17cc  :    0 - 0x0
    "00000000", -- 6093 - 0x17cd  :    0 - 0x0
    "00000000", -- 6094 - 0x17ce  :    0 - 0x0
    "00000000", -- 6095 - 0x17cf  :    0 - 0x0
    "00000000", -- 6096 - 0x17d0  :    0 - 0x0 -- Background 0x7d
    "00000000", -- 6097 - 0x17d1  :    0 - 0x0
    "00000000", -- 6098 - 0x17d2  :    0 - 0x0
    "00000000", -- 6099 - 0x17d3  :    0 - 0x0
    "00000000", -- 6100 - 0x17d4  :    0 - 0x0
    "00000000", -- 6101 - 0x17d5  :    0 - 0x0
    "00000000", -- 6102 - 0x17d6  :    0 - 0x0
    "00000000", -- 6103 - 0x17d7  :    0 - 0x0
    "00000000", -- 6104 - 0x17d8  :    0 - 0x0
    "00000000", -- 6105 - 0x17d9  :    0 - 0x0
    "00000000", -- 6106 - 0x17da  :    0 - 0x0
    "00000000", -- 6107 - 0x17db  :    0 - 0x0
    "00000000", -- 6108 - 0x17dc  :    0 - 0x0
    "00000000", -- 6109 - 0x17dd  :    0 - 0x0
    "00000000", -- 6110 - 0x17de  :    0 - 0x0
    "00000000", -- 6111 - 0x17df  :    0 - 0x0
    "00000000", -- 6112 - 0x17e0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 6113 - 0x17e1  :    0 - 0x0
    "00000000", -- 6114 - 0x17e2  :    0 - 0x0
    "00000000", -- 6115 - 0x17e3  :    0 - 0x0
    "00000000", -- 6116 - 0x17e4  :    0 - 0x0
    "00000000", -- 6117 - 0x17e5  :    0 - 0x0
    "00000000", -- 6118 - 0x17e6  :    0 - 0x0
    "00000000", -- 6119 - 0x17e7  :    0 - 0x0
    "00000000", -- 6120 - 0x17e8  :    0 - 0x0
    "00000000", -- 6121 - 0x17e9  :    0 - 0x0
    "00000000", -- 6122 - 0x17ea  :    0 - 0x0
    "00000000", -- 6123 - 0x17eb  :    0 - 0x0
    "00000000", -- 6124 - 0x17ec  :    0 - 0x0
    "00000000", -- 6125 - 0x17ed  :    0 - 0x0
    "00000000", -- 6126 - 0x17ee  :    0 - 0x0
    "00000000", -- 6127 - 0x17ef  :    0 - 0x0
    "00000000", -- 6128 - 0x17f0  :    0 - 0x0 -- Background 0x7f
    "00000000", -- 6129 - 0x17f1  :    0 - 0x0
    "00000000", -- 6130 - 0x17f2  :    0 - 0x0
    "00000000", -- 6131 - 0x17f3  :    0 - 0x0
    "00000000", -- 6132 - 0x17f4  :    0 - 0x0
    "00000000", -- 6133 - 0x17f5  :    0 - 0x0
    "00000000", -- 6134 - 0x17f6  :    0 - 0x0
    "00000000", -- 6135 - 0x17f7  :    0 - 0x0
    "00000000", -- 6136 - 0x17f8  :    0 - 0x0
    "00000000", -- 6137 - 0x17f9  :    0 - 0x0
    "00000000", -- 6138 - 0x17fa  :    0 - 0x0
    "00000000", -- 6139 - 0x17fb  :    0 - 0x0
    "00000000", -- 6140 - 0x17fc  :    0 - 0x0
    "00000000", -- 6141 - 0x17fd  :    0 - 0x0
    "00000000", -- 6142 - 0x17fe  :    0 - 0x0
    "00000000", -- 6143 - 0x17ff  :    0 - 0x0
    "10111111", -- 6144 - 0x1800  :  191 - 0xbf -- Background 0x80
    "11110111", -- 6145 - 0x1801  :  247 - 0xf7
    "11111101", -- 6146 - 0x1802  :  253 - 0xfd
    "11011111", -- 6147 - 0x1803  :  223 - 0xdf
    "11111011", -- 6148 - 0x1804  :  251 - 0xfb
    "10111111", -- 6149 - 0x1805  :  191 - 0xbf
    "11111110", -- 6150 - 0x1806  :  254 - 0xfe
    "11101111", -- 6151 - 0x1807  :  239 - 0xef
    "01000000", -- 6152 - 0x1808  :   64 - 0x40
    "00001000", -- 6153 - 0x1809  :    8 - 0x8
    "00000010", -- 6154 - 0x180a  :    2 - 0x2
    "00100000", -- 6155 - 0x180b  :   32 - 0x20
    "00000100", -- 6156 - 0x180c  :    4 - 0x4
    "01000000", -- 6157 - 0x180d  :   64 - 0x40
    "00000001", -- 6158 - 0x180e  :    1 - 0x1
    "00010000", -- 6159 - 0x180f  :   16 - 0x10
    "11111111", -- 6160 - 0x1810  :  255 - 0xff -- Background 0x81
    "11101110", -- 6161 - 0x1811  :  238 - 0xee
    "11111111", -- 6162 - 0x1812  :  255 - 0xff
    "11011111", -- 6163 - 0x1813  :  223 - 0xdf
    "01110111", -- 6164 - 0x1814  :  119 - 0x77
    "11111101", -- 6165 - 0x1815  :  253 - 0xfd
    "11011111", -- 6166 - 0x1816  :  223 - 0xdf
    "10111111", -- 6167 - 0x1817  :  191 - 0xbf
    "00000000", -- 6168 - 0x1818  :    0 - 0x0
    "00010001", -- 6169 - 0x1819  :   17 - 0x11
    "00000000", -- 6170 - 0x181a  :    0 - 0x0
    "00100000", -- 6171 - 0x181b  :   32 - 0x20
    "10001000", -- 6172 - 0x181c  :  136 - 0x88
    "00000010", -- 6173 - 0x181d  :    2 - 0x2
    "00100000", -- 6174 - 0x181e  :   32 - 0x20
    "01000000", -- 6175 - 0x181f  :   64 - 0x40
    "11111110", -- 6176 - 0x1820  :  254 - 0xfe -- Background 0x82
    "11101111", -- 6177 - 0x1821  :  239 - 0xef
    "10111111", -- 6178 - 0x1822  :  191 - 0xbf
    "11110111", -- 6179 - 0x1823  :  247 - 0xf7
    "11111101", -- 6180 - 0x1824  :  253 - 0xfd
    "11011111", -- 6181 - 0x1825  :  223 - 0xdf
    "11111011", -- 6182 - 0x1826  :  251 - 0xfb
    "10111111", -- 6183 - 0x1827  :  191 - 0xbf
    "00000001", -- 6184 - 0x1828  :    1 - 0x1
    "00010000", -- 6185 - 0x1829  :   16 - 0x10
    "01000000", -- 6186 - 0x182a  :   64 - 0x40
    "00001000", -- 6187 - 0x182b  :    8 - 0x8
    "00000010", -- 6188 - 0x182c  :    2 - 0x2
    "00100000", -- 6189 - 0x182d  :   32 - 0x20
    "00000100", -- 6190 - 0x182e  :    4 - 0x4
    "01000000", -- 6191 - 0x182f  :   64 - 0x40
    "11101111", -- 6192 - 0x1830  :  239 - 0xef -- Background 0x83
    "11111111", -- 6193 - 0x1831  :  255 - 0xff
    "10111011", -- 6194 - 0x1832  :  187 - 0xbb
    "11111111", -- 6195 - 0x1833  :  255 - 0xff
    "11110111", -- 6196 - 0x1834  :  247 - 0xf7
    "11011101", -- 6197 - 0x1835  :  221 - 0xdd
    "01111111", -- 6198 - 0x1836  :  127 - 0x7f
    "11110111", -- 6199 - 0x1837  :  247 - 0xf7
    "00010000", -- 6200 - 0x1838  :   16 - 0x10
    "00000000", -- 6201 - 0x1839  :    0 - 0x0
    "01000100", -- 6202 - 0x183a  :   68 - 0x44
    "00000000", -- 6203 - 0x183b  :    0 - 0x0
    "00001000", -- 6204 - 0x183c  :    8 - 0x8
    "00100010", -- 6205 - 0x183d  :   34 - 0x22
    "10000000", -- 6206 - 0x183e  :  128 - 0x80
    "00001000", -- 6207 - 0x183f  :    8 - 0x8
    "11111111", -- 6208 - 0x1840  :  255 - 0xff -- Background 0x84
    "11101110", -- 6209 - 0x1841  :  238 - 0xee
    "11111011", -- 6210 - 0x1842  :  251 - 0xfb
    "10111111", -- 6211 - 0x1843  :  191 - 0xbf
    "01111111", -- 6212 - 0x1844  :  127 - 0x7f
    "11101101", -- 6213 - 0x1845  :  237 - 0xed
    "11111111", -- 6214 - 0x1846  :  255 - 0xff
    "10111111", -- 6215 - 0x1847  :  191 - 0xbf
    "00010100", -- 6216 - 0x1848  :   20 - 0x14
    "10110101", -- 6217 - 0x1849  :  181 - 0xb5
    "01000100", -- 6218 - 0x184a  :   68 - 0x44
    "01001010", -- 6219 - 0x184b  :   74 - 0x4a
    "10010010", -- 6220 - 0x184c  :  146 - 0x92
    "10010010", -- 6221 - 0x184d  :  146 - 0x92
    "01000100", -- 6222 - 0x184e  :   68 - 0x44
    "01001001", -- 6223 - 0x184f  :   73 - 0x49
    "11111111", -- 6224 - 0x1850  :  255 - 0xff -- Background 0x85
    "10111111", -- 6225 - 0x1851  :  191 - 0xbf
    "01111101", -- 6226 - 0x1852  :  125 - 0x7d
    "11110111", -- 6227 - 0x1853  :  247 - 0xf7
    "11011011", -- 6228 - 0x1854  :  219 - 0xdb
    "11111101", -- 6229 - 0x1855  :  253 - 0xfd
    "01111110", -- 6230 - 0x1856  :  126 - 0x7e
    "11111011", -- 6231 - 0x1857  :  251 - 0xfb
    "01000010", -- 6232 - 0x1858  :   66 - 0x42
    "01001010", -- 6233 - 0x1859  :   74 - 0x4a
    "11001010", -- 6234 - 0x185a  :  202 - 0xca
    "00101001", -- 6235 - 0x185b  :   41 - 0x29
    "10100110", -- 6236 - 0x185c  :  166 - 0xa6
    "10010010", -- 6237 - 0x185d  :  146 - 0x92
    "10001001", -- 6238 - 0x185e  :  137 - 0x89
    "00101101", -- 6239 - 0x185f  :   45 - 0x2d
    "11111111", -- 6240 - 0x1860  :  255 - 0xff -- Background 0x86
    "11110111", -- 6241 - 0x1861  :  247 - 0xf7
    "11111111", -- 6242 - 0x1862  :  255 - 0xff
    "11011101", -- 6243 - 0x1863  :  221 - 0xdd
    "01111111", -- 6244 - 0x1864  :  127 - 0x7f
    "11110111", -- 6245 - 0x1865  :  247 - 0xf7
    "11101111", -- 6246 - 0x1866  :  239 - 0xef
    "10111101", -- 6247 - 0x1867  :  189 - 0xbd
    "10001000", -- 6248 - 0x1868  :  136 - 0x88
    "00101001", -- 6249 - 0x1869  :   41 - 0x29
    "10000010", -- 6250 - 0x186a  :  130 - 0x82
    "10110110", -- 6251 - 0x186b  :  182 - 0xb6
    "10001000", -- 6252 - 0x186c  :  136 - 0x88
    "01001001", -- 6253 - 0x186d  :   73 - 0x49
    "01010010", -- 6254 - 0x186e  :   82 - 0x52
    "01010010", -- 6255 - 0x186f  :   82 - 0x52
    "01011111", -- 6256 - 0x1870  :   95 - 0x5f -- Background 0x87
    "11111101", -- 6257 - 0x1871  :  253 - 0xfd
    "11110110", -- 6258 - 0x1872  :  246 - 0xf6
    "01111111", -- 6259 - 0x1873  :  127 - 0x7f
    "10011111", -- 6260 - 0x1874  :  159 - 0x9f
    "11111110", -- 6261 - 0x1875  :  254 - 0xfe
    "11111111", -- 6262 - 0x1876  :  255 - 0xff
    "11101111", -- 6263 - 0x1877  :  239 - 0xef
    "10110010", -- 6264 - 0x1878  :  178 - 0xb2
    "01001010", -- 6265 - 0x1879  :   74 - 0x4a
    "10101001", -- 6266 - 0x187a  :  169 - 0xa9
    "10100100", -- 6267 - 0x187b  :  164 - 0xa4
    "01100010", -- 6268 - 0x187c  :   98 - 0x62
    "01001011", -- 6269 - 0x187d  :   75 - 0x4b
    "10010000", -- 6270 - 0x187e  :  144 - 0x90
    "10010010", -- 6271 - 0x187f  :  146 - 0x92
    "11111111", -- 6272 - 0x1880  :  255 - 0xff -- Background 0x88
    "10011111", -- 6273 - 0x1881  :  159 - 0x9f
    "10111111", -- 6274 - 0x1882  :  191 - 0xbf
    "11111111", -- 6275 - 0x1883  :  255 - 0xff
    "11110011", -- 6276 - 0x1884  :  243 - 0xf3
    "11110011", -- 6277 - 0x1885  :  243 - 0xf3
    "11111111", -- 6278 - 0x1886  :  255 - 0xff
    "11111111", -- 6279 - 0x1887  :  255 - 0xff
    "01100000", -- 6280 - 0x1888  :   96 - 0x60
    "11110000", -- 6281 - 0x1889  :  240 - 0xf0
    "11110000", -- 6282 - 0x188a  :  240 - 0xf0
    "01101110", -- 6283 - 0x188b  :  110 - 0x6e
    "00011111", -- 6284 - 0x188c  :   31 - 0x1f
    "00011111", -- 6285 - 0x188d  :   31 - 0x1f
    "00011111", -- 6286 - 0x188e  :   31 - 0x1f
    "00001110", -- 6287 - 0x188f  :   14 - 0xe
    "11111111", -- 6288 - 0x1890  :  255 - 0xff -- Background 0x89
    "10011111", -- 6289 - 0x1891  :  159 - 0x9f
    "10111111", -- 6290 - 0x1892  :  191 - 0xbf
    "11110011", -- 6291 - 0x1893  :  243 - 0xf3
    "11110011", -- 6292 - 0x1894  :  243 - 0xf3
    "11111111", -- 6293 - 0x1895  :  255 - 0xff
    "11111111", -- 6294 - 0x1896  :  255 - 0xff
    "11111111", -- 6295 - 0x1897  :  255 - 0xff
    "01100000", -- 6296 - 0x1898  :   96 - 0x60
    "11110000", -- 6297 - 0x1899  :  240 - 0xf0
    "11111110", -- 6298 - 0x189a  :  254 - 0xfe
    "01111111", -- 6299 - 0x189b  :  127 - 0x7f
    "00011111", -- 6300 - 0x189c  :   31 - 0x1f
    "00011111", -- 6301 - 0x189d  :   31 - 0x1f
    "00001110", -- 6302 - 0x189e  :   14 - 0xe
    "00000000", -- 6303 - 0x189f  :    0 - 0x0
    "10111111", -- 6304 - 0x18a0  :  191 - 0xbf -- Background 0x8a
    "11110111", -- 6305 - 0x18a1  :  247 - 0xf7
    "11111101", -- 6306 - 0x18a2  :  253 - 0xfd
    "11111111", -- 6307 - 0x18a3  :  255 - 0xff
    "11111011", -- 6308 - 0x18a4  :  251 - 0xfb
    "10111111", -- 6309 - 0x18a5  :  191 - 0xbf
    "11111110", -- 6310 - 0x18a6  :  254 - 0xfe
    "11101111", -- 6311 - 0x18a7  :  239 - 0xef
    "01000000", -- 6312 - 0x18a8  :   64 - 0x40
    "00001000", -- 6313 - 0x18a9  :    8 - 0x8
    "00000010", -- 6314 - 0x18aa  :    2 - 0x2
    "00101000", -- 6315 - 0x18ab  :   40 - 0x28
    "00010100", -- 6316 - 0x18ac  :   20 - 0x14
    "01010100", -- 6317 - 0x18ad  :   84 - 0x54
    "00000001", -- 6318 - 0x18ae  :    1 - 0x1
    "00010000", -- 6319 - 0x18af  :   16 - 0x10
    "10111111", -- 6320 - 0x18b0  :  191 - 0xbf -- Background 0x8b
    "11111111", -- 6321 - 0x18b1  :  255 - 0xff
    "11101110", -- 6322 - 0x18b2  :  238 - 0xee
    "11111111", -- 6323 - 0x18b3  :  255 - 0xff
    "11011111", -- 6324 - 0x18b4  :  223 - 0xdf
    "01111101", -- 6325 - 0x18b5  :  125 - 0x7d
    "11111111", -- 6326 - 0x18b6  :  255 - 0xff
    "11011111", -- 6327 - 0x18b7  :  223 - 0xdf
    "01000000", -- 6328 - 0x18b8  :   64 - 0x40
    "00000000", -- 6329 - 0x18b9  :    0 - 0x0
    "10010001", -- 6330 - 0x18ba  :  145 - 0x91
    "00010100", -- 6331 - 0x18bb  :   20 - 0x14
    "00101000", -- 6332 - 0x18bc  :   40 - 0x28
    "10001010", -- 6333 - 0x18bd  :  138 - 0x8a
    "01000000", -- 6334 - 0x18be  :   64 - 0x40
    "00100000", -- 6335 - 0x18bf  :   32 - 0x20
    "11111111", -- 6336 - 0x18c0  :  255 - 0xff -- Background 0x8c
    "11111000", -- 6337 - 0x18c1  :  248 - 0xf8
    "11100010", -- 6338 - 0x18c2  :  226 - 0xe2
    "11010111", -- 6339 - 0x18c3  :  215 - 0xd7
    "11001111", -- 6340 - 0x18c4  :  207 - 0xcf
    "10011111", -- 6341 - 0x18c5  :  159 - 0x9f
    "10111110", -- 6342 - 0x18c6  :  190 - 0xbe
    "10011101", -- 6343 - 0x18c7  :  157 - 0x9d
    "00000000", -- 6344 - 0x18c8  :    0 - 0x0
    "00000111", -- 6345 - 0x18c9  :    7 - 0x7
    "00011111", -- 6346 - 0x18ca  :   31 - 0x1f
    "00111111", -- 6347 - 0x18cb  :   63 - 0x3f
    "00111111", -- 6348 - 0x18cc  :   63 - 0x3f
    "01111111", -- 6349 - 0x18cd  :  127 - 0x7f
    "01111111", -- 6350 - 0x18ce  :  127 - 0x7f
    "01111111", -- 6351 - 0x18cf  :  127 - 0x7f
    "11111111", -- 6352 - 0x18d0  :  255 - 0xff -- Background 0x8d
    "00011111", -- 6353 - 0x18d1  :   31 - 0x1f
    "10100111", -- 6354 - 0x18d2  :  167 - 0xa7
    "11000011", -- 6355 - 0x18d3  :  195 - 0xc3
    "11100011", -- 6356 - 0x18d4  :  227 - 0xe3
    "01000001", -- 6357 - 0x18d5  :   65 - 0x41
    "10100001", -- 6358 - 0x18d6  :  161 - 0xa1
    "00000001", -- 6359 - 0x18d7  :    1 - 0x1
    "00000000", -- 6360 - 0x18d8  :    0 - 0x0
    "11100000", -- 6361 - 0x18d9  :  224 - 0xe0
    "11111000", -- 6362 - 0x18da  :  248 - 0xf8
    "11111000", -- 6363 - 0x18db  :  248 - 0xf8
    "11110000", -- 6364 - 0x18dc  :  240 - 0xf0
    "11111000", -- 6365 - 0x18dd  :  248 - 0xf8
    "11110100", -- 6366 - 0x18de  :  244 - 0xf4
    "11111000", -- 6367 - 0x18df  :  248 - 0xf8
    "10111110", -- 6368 - 0x18e0  :  190 - 0xbe -- Background 0x8e
    "11111111", -- 6369 - 0x18e1  :  255 - 0xff
    "11011111", -- 6370 - 0x18e2  :  223 - 0xdf
    "11111111", -- 6371 - 0x18e3  :  255 - 0xff
    "11101111", -- 6372 - 0x18e4  :  239 - 0xef
    "11111111", -- 6373 - 0x18e5  :  255 - 0xff
    "11110111", -- 6374 - 0x18e6  :  247 - 0xf7
    "11111111", -- 6375 - 0x18e7  :  255 - 0xff
    "01111111", -- 6376 - 0x18e8  :  127 - 0x7f
    "00111111", -- 6377 - 0x18e9  :   63 - 0x3f
    "00111111", -- 6378 - 0x18ea  :   63 - 0x3f
    "00011111", -- 6379 - 0x18eb  :   31 - 0x1f
    "00011111", -- 6380 - 0x18ec  :   31 - 0x1f
    "00001111", -- 6381 - 0x18ed  :   15 - 0xf
    "00001111", -- 6382 - 0x18ee  :   15 - 0xf
    "00000111", -- 6383 - 0x18ef  :    7 - 0x7
    "01111101", -- 6384 - 0x18f0  :  125 - 0x7d -- Background 0x8f
    "11111111", -- 6385 - 0x18f1  :  255 - 0xff
    "11111011", -- 6386 - 0x18f2  :  251 - 0xfb
    "11111111", -- 6387 - 0x18f3  :  255 - 0xff
    "11110111", -- 6388 - 0x18f4  :  247 - 0xf7
    "11111111", -- 6389 - 0x18f5  :  255 - 0xff
    "11101111", -- 6390 - 0x18f6  :  239 - 0xef
    "11111111", -- 6391 - 0x18f7  :  255 - 0xff
    "11111110", -- 6392 - 0x18f8  :  254 - 0xfe
    "11111100", -- 6393 - 0x18f9  :  252 - 0xfc
    "11111100", -- 6394 - 0x18fa  :  252 - 0xfc
    "11111000", -- 6395 - 0x18fb  :  248 - 0xf8
    "11111000", -- 6396 - 0x18fc  :  248 - 0xf8
    "11110000", -- 6397 - 0x18fd  :  240 - 0xf0
    "11110000", -- 6398 - 0x18fe  :  240 - 0xf0
    "11100000", -- 6399 - 0x18ff  :  224 - 0xe0
    "10111110", -- 6400 - 0x1900  :  190 - 0xbe -- Background 0x90
    "11110111", -- 6401 - 0x1901  :  247 - 0xf7
    "11111111", -- 6402 - 0x1902  :  255 - 0xff
    "11011111", -- 6403 - 0x1903  :  223 - 0xdf
    "11111011", -- 6404 - 0x1904  :  251 - 0xfb
    "11111110", -- 6405 - 0x1905  :  254 - 0xfe
    "10111111", -- 6406 - 0x1906  :  191 - 0xbf
    "11110111", -- 6407 - 0x1907  :  247 - 0xf7
    "01000001", -- 6408 - 0x1908  :   65 - 0x41
    "00001000", -- 6409 - 0x1909  :    8 - 0x8
    "00000000", -- 6410 - 0x190a  :    0 - 0x0
    "00100000", -- 6411 - 0x190b  :   32 - 0x20
    "00000100", -- 6412 - 0x190c  :    4 - 0x4
    "00000001", -- 6413 - 0x190d  :    1 - 0x1
    "01000000", -- 6414 - 0x190e  :   64 - 0x40
    "00001000", -- 6415 - 0x190f  :    8 - 0x8
    "11101110", -- 6416 - 0x1910  :  238 - 0xee -- Background 0x91
    "11111111", -- 6417 - 0x1911  :  255 - 0xff
    "01111011", -- 6418 - 0x1912  :  123 - 0x7b
    "11111101", -- 6419 - 0x1913  :  253 - 0xfd
    "11101111", -- 6420 - 0x1914  :  239 - 0xef
    "11111111", -- 6421 - 0x1915  :  255 - 0xff
    "10111101", -- 6422 - 0x1916  :  189 - 0xbd
    "11111111", -- 6423 - 0x1917  :  255 - 0xff
    "00010001", -- 6424 - 0x1918  :   17 - 0x11
    "00000000", -- 6425 - 0x1919  :    0 - 0x0
    "10000100", -- 6426 - 0x191a  :  132 - 0x84
    "00000010", -- 6427 - 0x191b  :    2 - 0x2
    "00010000", -- 6428 - 0x191c  :   16 - 0x10
    "00000000", -- 6429 - 0x191d  :    0 - 0x0
    "01000010", -- 6430 - 0x191e  :   66 - 0x42
    "00000000", -- 6431 - 0x191f  :    0 - 0x0
    "11111011", -- 6432 - 0x1920  :  251 - 0xfb -- Background 0x92
    "10111111", -- 6433 - 0x1921  :  191 - 0xbf
    "11101111", -- 6434 - 0x1922  :  239 - 0xef
    "11111101", -- 6435 - 0x1923  :  253 - 0xfd
    "11111111", -- 6436 - 0x1924  :  255 - 0xff
    "10111111", -- 6437 - 0x1925  :  191 - 0xbf
    "11111011", -- 6438 - 0x1926  :  251 - 0xfb
    "11011111", -- 6439 - 0x1927  :  223 - 0xdf
    "00000100", -- 6440 - 0x1928  :    4 - 0x4
    "01000000", -- 6441 - 0x1929  :   64 - 0x40
    "00010000", -- 6442 - 0x192a  :   16 - 0x10
    "00000010", -- 6443 - 0x192b  :    2 - 0x2
    "00000000", -- 6444 - 0x192c  :    0 - 0x0
    "01000000", -- 6445 - 0x192d  :   64 - 0x40
    "00000100", -- 6446 - 0x192e  :    4 - 0x4
    "00100000", -- 6447 - 0x192f  :   32 - 0x20
    "10111101", -- 6448 - 0x1930  :  189 - 0xbd -- Background 0x93
    "11111111", -- 6449 - 0x1931  :  255 - 0xff
    "01110111", -- 6450 - 0x1932  :  119 - 0x77
    "11111110", -- 6451 - 0x1933  :  254 - 0xfe
    "11011111", -- 6452 - 0x1934  :  223 - 0xdf
    "11111011", -- 6453 - 0x1935  :  251 - 0xfb
    "11101111", -- 6454 - 0x1936  :  239 - 0xef
    "01111111", -- 6455 - 0x1937  :  127 - 0x7f
    "01000010", -- 6456 - 0x1938  :   66 - 0x42
    "00000000", -- 6457 - 0x1939  :    0 - 0x0
    "10001000", -- 6458 - 0x193a  :  136 - 0x88
    "00000001", -- 6459 - 0x193b  :    1 - 0x1
    "00100000", -- 6460 - 0x193c  :   32 - 0x20
    "00000100", -- 6461 - 0x193d  :    4 - 0x4
    "00010000", -- 6462 - 0x193e  :   16 - 0x10
    "10000000", -- 6463 - 0x193f  :  128 - 0x80
    "01111111", -- 6464 - 0x1940  :  127 - 0x7f -- Background 0x94
    "11110111", -- 6465 - 0x1941  :  247 - 0xf7
    "11011101", -- 6466 - 0x1942  :  221 - 0xdd
    "01111011", -- 6467 - 0x1943  :  123 - 0x7b
    "11111111", -- 6468 - 0x1944  :  255 - 0xff
    "11101110", -- 6469 - 0x1945  :  238 - 0xee
    "10111011", -- 6470 - 0x1946  :  187 - 0xbb
    "11111101", -- 6471 - 0x1947  :  253 - 0xfd
    "11001000", -- 6472 - 0x1948  :  200 - 0xc8
    "00101010", -- 6473 - 0x1949  :   42 - 0x2a
    "10100010", -- 6474 - 0x194a  :  162 - 0xa2
    "10010100", -- 6475 - 0x194b  :  148 - 0x94
    "10010001", -- 6476 - 0x194c  :  145 - 0x91
    "01010101", -- 6477 - 0x194d  :   85 - 0x55
    "01000100", -- 6478 - 0x194e  :   68 - 0x44
    "00010010", -- 6479 - 0x194f  :   18 - 0x12
    "11010111", -- 6480 - 0x1950  :  215 - 0xd7 -- Background 0x95
    "01111111", -- 6481 - 0x1951  :  127 - 0x7f
    "11111101", -- 6482 - 0x1952  :  253 - 0xfd
    "11101110", -- 6483 - 0x1953  :  238 - 0xee
    "11110111", -- 6484 - 0x1954  :  247 - 0xf7
    "10111011", -- 6485 - 0x1955  :  187 - 0xbb
    "11101111", -- 6486 - 0x1956  :  239 - 0xef
    "11110111", -- 6487 - 0x1957  :  247 - 0xf7
    "10101010", -- 6488 - 0x1958  :  170 - 0xaa
    "10100010", -- 6489 - 0x1959  :  162 - 0xa2
    "00010010", -- 6490 - 0x195a  :   18 - 0x12
    "01010011", -- 6491 - 0x195b  :   83 - 0x53
    "01001100", -- 6492 - 0x195c  :   76 - 0x4c
    "01010101", -- 6493 - 0x195d  :   85 - 0x55
    "10010001", -- 6494 - 0x195e  :  145 - 0x91
    "01001000", -- 6495 - 0x195f  :   72 - 0x48
    "10111111", -- 6496 - 0x1960  :  191 - 0xbf -- Background 0x96
    "11101110", -- 6497 - 0x1961  :  238 - 0xee
    "11011011", -- 6498 - 0x1962  :  219 - 0xdb
    "11111111", -- 6499 - 0x1963  :  255 - 0xff
    "01110111", -- 6500 - 0x1964  :  119 - 0x77
    "11011101", -- 6501 - 0x1965  :  221 - 0xdd
    "11101111", -- 6502 - 0x1966  :  239 - 0xef
    "11111011", -- 6503 - 0x1967  :  251 - 0xfb
    "01010001", -- 6504 - 0x1968  :   81 - 0x51
    "00010101", -- 6505 - 0x1969  :   21 - 0x15
    "10100100", -- 6506 - 0x196a  :  164 - 0xa4
    "10001100", -- 6507 - 0x196b  :  140 - 0x8c
    "10101010", -- 6508 - 0x196c  :  170 - 0xaa
    "00100010", -- 6509 - 0x196d  :   34 - 0x22
    "10010000", -- 6510 - 0x196e  :  144 - 0x90
    "01000110", -- 6511 - 0x196f  :   70 - 0x46
    "11111101", -- 6512 - 0x1970  :  253 - 0xfd -- Background 0x97
    "11101110", -- 6513 - 0x1971  :  238 - 0xee
    "11111011", -- 6514 - 0x1972  :  251 - 0xfb
    "11111101", -- 6515 - 0x1973  :  253 - 0xfd
    "11110101", -- 6516 - 0x1974  :  245 - 0xf5
    "11011111", -- 6517 - 0x1975  :  223 - 0xdf
    "01111111", -- 6518 - 0x1976  :  127 - 0x7f
    "10111011", -- 6519 - 0x1977  :  187 - 0xbb
    "00010011", -- 6520 - 0x1978  :   19 - 0x13
    "01010101", -- 6521 - 0x1979  :   85 - 0x55
    "01100100", -- 6522 - 0x197a  :  100 - 0x64
    "00010010", -- 6523 - 0x197b  :   18 - 0x12
    "10101010", -- 6524 - 0x197c  :  170 - 0xaa
    "10101000", -- 6525 - 0x197d  :  168 - 0xa8
    "10000100", -- 6526 - 0x197e  :  132 - 0x84
    "11010100", -- 6527 - 0x197f  :  212 - 0xd4
    "11111111", -- 6528 - 0x1980  :  255 - 0xff -- Background 0x98
    "10011111", -- 6529 - 0x1981  :  159 - 0x9f
    "10111111", -- 6530 - 0x1982  :  191 - 0xbf
    "11110011", -- 6531 - 0x1983  :  243 - 0xf3
    "11110011", -- 6532 - 0x1984  :  243 - 0xf3
    "11111111", -- 6533 - 0x1985  :  255 - 0xff
    "11111111", -- 6534 - 0x1986  :  255 - 0xff
    "11111111", -- 6535 - 0x1987  :  255 - 0xff
    "01100000", -- 6536 - 0x1988  :   96 - 0x60
    "11110000", -- 6537 - 0x1989  :  240 - 0xf0
    "11111110", -- 6538 - 0x198a  :  254 - 0xfe
    "01111111", -- 6539 - 0x198b  :  127 - 0x7f
    "00011111", -- 6540 - 0x198c  :   31 - 0x1f
    "00011111", -- 6541 - 0x198d  :   31 - 0x1f
    "00001110", -- 6542 - 0x198e  :   14 - 0xe
    "00000000", -- 6543 - 0x198f  :    0 - 0x0
    "11111111", -- 6544 - 0x1990  :  255 - 0xff -- Background 0x99
    "10011111", -- 6545 - 0x1991  :  159 - 0x9f
    "10111111", -- 6546 - 0x1992  :  191 - 0xbf
    "11111111", -- 6547 - 0x1993  :  255 - 0xff
    "11110011", -- 6548 - 0x1994  :  243 - 0xf3
    "11110011", -- 6549 - 0x1995  :  243 - 0xf3
    "11111111", -- 6550 - 0x1996  :  255 - 0xff
    "11111111", -- 6551 - 0x1997  :  255 - 0xff
    "01100000", -- 6552 - 0x1998  :   96 - 0x60
    "11110000", -- 6553 - 0x1999  :  240 - 0xf0
    "11110000", -- 6554 - 0x199a  :  240 - 0xf0
    "01101110", -- 6555 - 0x199b  :  110 - 0x6e
    "00011111", -- 6556 - 0x199c  :   31 - 0x1f
    "00011111", -- 6557 - 0x199d  :   31 - 0x1f
    "00011111", -- 6558 - 0x199e  :   31 - 0x1f
    "00001110", -- 6559 - 0x199f  :   14 - 0xe
    "10111111", -- 6560 - 0x19a0  :  191 - 0xbf -- Background 0x9a
    "11110111", -- 6561 - 0x19a1  :  247 - 0xf7
    "11111111", -- 6562 - 0x19a2  :  255 - 0xff
    "11011111", -- 6563 - 0x19a3  :  223 - 0xdf
    "11111011", -- 6564 - 0x19a4  :  251 - 0xfb
    "11111111", -- 6565 - 0x19a5  :  255 - 0xff
    "10111111", -- 6566 - 0x19a6  :  191 - 0xbf
    "11110111", -- 6567 - 0x19a7  :  247 - 0xf7
    "01000000", -- 6568 - 0x19a8  :   64 - 0x40
    "00001100", -- 6569 - 0x19a9  :   12 - 0xc
    "00000000", -- 6570 - 0x19aa  :    0 - 0x0
    "00101000", -- 6571 - 0x19ab  :   40 - 0x28
    "00101100", -- 6572 - 0x19ac  :   44 - 0x2c
    "00010001", -- 6573 - 0x19ad  :   17 - 0x11
    "01000000", -- 6574 - 0x19ae  :   64 - 0x40
    "00001000", -- 6575 - 0x19af  :    8 - 0x8
    "11011111", -- 6576 - 0x19b0  :  223 - 0xdf -- Background 0x9b
    "11111111", -- 6577 - 0x19b1  :  255 - 0xff
    "01111011", -- 6578 - 0x19b2  :  123 - 0x7b
    "11111111", -- 6579 - 0x19b3  :  255 - 0xff
    "11101111", -- 6580 - 0x19b4  :  239 - 0xef
    "11111101", -- 6581 - 0x19b5  :  253 - 0xfd
    "10111111", -- 6582 - 0x19b6  :  191 - 0xbf
    "11111111", -- 6583 - 0x19b7  :  255 - 0xff
    "00100000", -- 6584 - 0x19b8  :   32 - 0x20
    "00000000", -- 6585 - 0x19b9  :    0 - 0x0
    "10010100", -- 6586 - 0x19ba  :  148 - 0x94
    "01001000", -- 6587 - 0x19bb  :   72 - 0x48
    "00011000", -- 6588 - 0x19bc  :   24 - 0x18
    "00000110", -- 6589 - 0x19bd  :    6 - 0x6
    "01000000", -- 6590 - 0x19be  :   64 - 0x40
    "00000000", -- 6591 - 0x19bf  :    0 - 0x0
    "10111010", -- 6592 - 0x19c0  :  186 - 0xba -- Background 0x9c
    "10011100", -- 6593 - 0x19c1  :  156 - 0x9c
    "10101010", -- 6594 - 0x19c2  :  170 - 0xaa
    "11000000", -- 6595 - 0x19c3  :  192 - 0xc0
    "11000000", -- 6596 - 0x19c4  :  192 - 0xc0
    "11100000", -- 6597 - 0x19c5  :  224 - 0xe0
    "11111000", -- 6598 - 0x19c6  :  248 - 0xf8
    "11111111", -- 6599 - 0x19c7  :  255 - 0xff
    "01111111", -- 6600 - 0x19c8  :  127 - 0x7f
    "01111111", -- 6601 - 0x19c9  :  127 - 0x7f
    "01111111", -- 6602 - 0x19ca  :  127 - 0x7f
    "00111111", -- 6603 - 0x19cb  :   63 - 0x3f
    "00110101", -- 6604 - 0x19cc  :   53 - 0x35
    "00000010", -- 6605 - 0x19cd  :    2 - 0x2
    "00000000", -- 6606 - 0x19ce  :    0 - 0x0
    "00000000", -- 6607 - 0x19cf  :    0 - 0x0
    "00000001", -- 6608 - 0x19d0  :    1 - 0x1 -- Background 0x9d
    "00000001", -- 6609 - 0x19d1  :    1 - 0x1
    "00000001", -- 6610 - 0x19d2  :    1 - 0x1
    "00000011", -- 6611 - 0x19d3  :    3 - 0x3
    "00000011", -- 6612 - 0x19d4  :    3 - 0x3
    "00000111", -- 6613 - 0x19d5  :    7 - 0x7
    "00011111", -- 6614 - 0x19d6  :   31 - 0x1f
    "11111111", -- 6615 - 0x19d7  :  255 - 0xff
    "11110100", -- 6616 - 0x19d8  :  244 - 0xf4
    "11111000", -- 6617 - 0x19d9  :  248 - 0xf8
    "11110000", -- 6618 - 0x19da  :  240 - 0xf0
    "11101000", -- 6619 - 0x19db  :  232 - 0xe8
    "01010000", -- 6620 - 0x19dc  :   80 - 0x50
    "10000000", -- 6621 - 0x19dd  :  128 - 0x80
    "00000000", -- 6622 - 0x19de  :    0 - 0x0
    "00000000", -- 6623 - 0x19df  :    0 - 0x0
    "01111101", -- 6624 - 0x19e0  :  125 - 0x7d -- Background 0x9e
    "11111111", -- 6625 - 0x19e1  :  255 - 0xff
    "11111011", -- 6626 - 0x19e2  :  251 - 0xfb
    "11111111", -- 6627 - 0x19e3  :  255 - 0xff
    "11111111", -- 6628 - 0x19e4  :  255 - 0xff
    "11111011", -- 6629 - 0x19e5  :  251 - 0xfb
    "11111111", -- 6630 - 0x19e6  :  255 - 0xff
    "01111101", -- 6631 - 0x19e7  :  125 - 0x7d
    "11111110", -- 6632 - 0x19e8  :  254 - 0xfe
    "11111100", -- 6633 - 0x19e9  :  252 - 0xfc
    "11111100", -- 6634 - 0x19ea  :  252 - 0xfc
    "11111000", -- 6635 - 0x19eb  :  248 - 0xf8
    "11111000", -- 6636 - 0x19ec  :  248 - 0xf8
    "11111100", -- 6637 - 0x19ed  :  252 - 0xfc
    "11111100", -- 6638 - 0x19ee  :  252 - 0xfc
    "11111110", -- 6639 - 0x19ef  :  254 - 0xfe
    "11111111", -- 6640 - 0x19f0  :  255 - 0xff -- Background 0x9f
    "11111111", -- 6641 - 0x19f1  :  255 - 0xff
    "10111101", -- 6642 - 0x19f2  :  189 - 0xbd
    "11111111", -- 6643 - 0x19f3  :  255 - 0xff
    "11111111", -- 6644 - 0x19f4  :  255 - 0xff
    "11111111", -- 6645 - 0x19f5  :  255 - 0xff
    "11111111", -- 6646 - 0x19f6  :  255 - 0xff
    "10111101", -- 6647 - 0x19f7  :  189 - 0xbd
    "00000000", -- 6648 - 0x19f8  :    0 - 0x0
    "00000000", -- 6649 - 0x19f9  :    0 - 0x0
    "01111110", -- 6650 - 0x19fa  :  126 - 0x7e
    "01111110", -- 6651 - 0x19fb  :  126 - 0x7e
    "01111110", -- 6652 - 0x19fc  :  126 - 0x7e
    "01111110", -- 6653 - 0x19fd  :  126 - 0x7e
    "01111110", -- 6654 - 0x19fe  :  126 - 0x7e
    "01111110", -- 6655 - 0x19ff  :  126 - 0x7e
    "11101111", -- 6656 - 0x1a00  :  239 - 0xef -- Background 0xa0
    "11000111", -- 6657 - 0x1a01  :  199 - 0xc7
    "10000011", -- 6658 - 0x1a02  :  131 - 0x83
    "00000111", -- 6659 - 0x1a03  :    7 - 0x7
    "10001111", -- 6660 - 0x1a04  :  143 - 0x8f
    "11011101", -- 6661 - 0x1a05  :  221 - 0xdd
    "11111010", -- 6662 - 0x1a06  :  250 - 0xfa
    "11111101", -- 6663 - 0x1a07  :  253 - 0xfd
    "00010000", -- 6664 - 0x1a08  :   16 - 0x10
    "00111000", -- 6665 - 0x1a09  :   56 - 0x38
    "01111100", -- 6666 - 0x1a0a  :  124 - 0x7c
    "11111000", -- 6667 - 0x1a0b  :  248 - 0xf8
    "01110000", -- 6668 - 0x1a0c  :  112 - 0x70
    "00100010", -- 6669 - 0x1a0d  :   34 - 0x22
    "00000101", -- 6670 - 0x1a0e  :    5 - 0x5
    "00000010", -- 6671 - 0x1a0f  :    2 - 0x2
    "11101111", -- 6672 - 0x1a10  :  239 - 0xef -- Background 0xa1
    "11000111", -- 6673 - 0x1a11  :  199 - 0xc7
    "10000011", -- 6674 - 0x1a12  :  131 - 0x83
    "00011111", -- 6675 - 0x1a13  :   31 - 0x1f
    "10010000", -- 6676 - 0x1a14  :  144 - 0x90
    "11010100", -- 6677 - 0x1a15  :  212 - 0xd4
    "11110011", -- 6678 - 0x1a16  :  243 - 0xf3
    "11110010", -- 6679 - 0x1a17  :  242 - 0xf2
    "00010000", -- 6680 - 0x1a18  :   16 - 0x10
    "00111000", -- 6681 - 0x1a19  :   56 - 0x38
    "01111100", -- 6682 - 0x1a1a  :  124 - 0x7c
    "11100000", -- 6683 - 0x1a1b  :  224 - 0xe0
    "01100000", -- 6684 - 0x1a1c  :   96 - 0x60
    "00100000", -- 6685 - 0x1a1d  :   32 - 0x20
    "00000000", -- 6686 - 0x1a1e  :    0 - 0x0
    "00000000", -- 6687 - 0x1a1f  :    0 - 0x0
    "11101111", -- 6688 - 0x1a20  :  239 - 0xef -- Background 0xa2
    "11000111", -- 6689 - 0x1a21  :  199 - 0xc7
    "10000011", -- 6690 - 0x1a22  :  131 - 0x83
    "11111111", -- 6691 - 0x1a23  :  255 - 0xff
    "00000000", -- 6692 - 0x1a24  :    0 - 0x0
    "00000000", -- 6693 - 0x1a25  :    0 - 0x0
    "01010101", -- 6694 - 0x1a26  :   85 - 0x55
    "00000000", -- 6695 - 0x1a27  :    0 - 0x0
    "00010000", -- 6696 - 0x1a28  :   16 - 0x10
    "00111000", -- 6697 - 0x1a29  :   56 - 0x38
    "01111100", -- 6698 - 0x1a2a  :  124 - 0x7c
    "00000000", -- 6699 - 0x1a2b  :    0 - 0x0
    "00000000", -- 6700 - 0x1a2c  :    0 - 0x0
    "00000000", -- 6701 - 0x1a2d  :    0 - 0x0
    "00000000", -- 6702 - 0x1a2e  :    0 - 0x0
    "00000000", -- 6703 - 0x1a2f  :    0 - 0x0
    "11110000", -- 6704 - 0x1a30  :  240 - 0xf0 -- Background 0xa3
    "11010010", -- 6705 - 0x1a31  :  210 - 0xd2
    "10010000", -- 6706 - 0x1a32  :  144 - 0x90
    "00010010", -- 6707 - 0x1a33  :   18 - 0x12
    "10010000", -- 6708 - 0x1a34  :  144 - 0x90
    "11010010", -- 6709 - 0x1a35  :  210 - 0xd2
    "11110000", -- 6710 - 0x1a36  :  240 - 0xf0
    "11110010", -- 6711 - 0x1a37  :  242 - 0xf2
    "00000000", -- 6712 - 0x1a38  :    0 - 0x0
    "00100000", -- 6713 - 0x1a39  :   32 - 0x20
    "01100000", -- 6714 - 0x1a3a  :   96 - 0x60
    "11100000", -- 6715 - 0x1a3b  :  224 - 0xe0
    "01100000", -- 6716 - 0x1a3c  :   96 - 0x60
    "00100000", -- 6717 - 0x1a3d  :   32 - 0x20
    "00000000", -- 6718 - 0x1a3e  :    0 - 0x0
    "00000000", -- 6719 - 0x1a3f  :    0 - 0x0
    "11110000", -- 6720 - 0x1a40  :  240 - 0xf0 -- Background 0xa4
    "11010011", -- 6721 - 0x1a41  :  211 - 0xd3
    "10010100", -- 6722 - 0x1a42  :  148 - 0x94
    "00011000", -- 6723 - 0x1a43  :   24 - 0x18
    "10011111", -- 6724 - 0x1a44  :  159 - 0x9f
    "11011101", -- 6725 - 0x1a45  :  221 - 0xdd
    "11111010", -- 6726 - 0x1a46  :  250 - 0xfa
    "11111101", -- 6727 - 0x1a47  :  253 - 0xfd
    "00000000", -- 6728 - 0x1a48  :    0 - 0x0
    "00100000", -- 6729 - 0x1a49  :   32 - 0x20
    "01100011", -- 6730 - 0x1a4a  :   99 - 0x63
    "11100111", -- 6731 - 0x1a4b  :  231 - 0xe7
    "01100000", -- 6732 - 0x1a4c  :   96 - 0x60
    "00100010", -- 6733 - 0x1a4d  :   34 - 0x22
    "00000101", -- 6734 - 0x1a4e  :    5 - 0x5
    "00000010", -- 6735 - 0x1a4f  :    2 - 0x2
    "00000000", -- 6736 - 0x1a50  :    0 - 0x0 -- Background 0xa5
    "11111111", -- 6737 - 0x1a51  :  255 - 0xff
    "00000000", -- 6738 - 0x1a52  :    0 - 0x0
    "00000000", -- 6739 - 0x1a53  :    0 - 0x0
    "11111111", -- 6740 - 0x1a54  :  255 - 0xff
    "11011101", -- 6741 - 0x1a55  :  221 - 0xdd
    "11111010", -- 6742 - 0x1a56  :  250 - 0xfa
    "11111101", -- 6743 - 0x1a57  :  253 - 0xfd
    "00000000", -- 6744 - 0x1a58  :    0 - 0x0
    "00000000", -- 6745 - 0x1a59  :    0 - 0x0
    "11111111", -- 6746 - 0x1a5a  :  255 - 0xff
    "11111111", -- 6747 - 0x1a5b  :  255 - 0xff
    "00000000", -- 6748 - 0x1a5c  :    0 - 0x0
    "00100010", -- 6749 - 0x1a5d  :   34 - 0x22
    "00000101", -- 6750 - 0x1a5e  :    5 - 0x5
    "00000010", -- 6751 - 0x1a5f  :    2 - 0x2
    "11101111", -- 6752 - 0x1a60  :  239 - 0xef -- Background 0xa6
    "11000111", -- 6753 - 0x1a61  :  199 - 0xc7
    "10000011", -- 6754 - 0x1a62  :  131 - 0x83
    "11111111", -- 6755 - 0x1a63  :  255 - 0xff
    "00011111", -- 6756 - 0x1a64  :   31 - 0x1f
    "00101101", -- 6757 - 0x1a65  :   45 - 0x2d
    "01001010", -- 6758 - 0x1a66  :   74 - 0x4a
    "01001101", -- 6759 - 0x1a67  :   77 - 0x4d
    "00010000", -- 6760 - 0x1a68  :   16 - 0x10
    "00111000", -- 6761 - 0x1a69  :   56 - 0x38
    "01111100", -- 6762 - 0x1a6a  :  124 - 0x7c
    "00000000", -- 6763 - 0x1a6b  :    0 - 0x0
    "00000000", -- 6764 - 0x1a6c  :    0 - 0x0
    "00010010", -- 6765 - 0x1a6d  :   18 - 0x12
    "00110101", -- 6766 - 0x1a6e  :   53 - 0x35
    "00110010", -- 6767 - 0x1a6f  :   50 - 0x32
    "01001111", -- 6768 - 0x1a70  :   79 - 0x4f -- Background 0xa7
    "01001111", -- 6769 - 0x1a71  :   79 - 0x4f
    "01001011", -- 6770 - 0x1a72  :   75 - 0x4b
    "01001111", -- 6771 - 0x1a73  :   79 - 0x4f
    "01001111", -- 6772 - 0x1a74  :   79 - 0x4f
    "01001101", -- 6773 - 0x1a75  :   77 - 0x4d
    "01001010", -- 6774 - 0x1a76  :   74 - 0x4a
    "01001101", -- 6775 - 0x1a77  :   77 - 0x4d
    "00110000", -- 6776 - 0x1a78  :   48 - 0x30
    "00110000", -- 6777 - 0x1a79  :   48 - 0x30
    "00110100", -- 6778 - 0x1a7a  :   52 - 0x34
    "00110000", -- 6779 - 0x1a7b  :   48 - 0x30
    "00110000", -- 6780 - 0x1a7c  :   48 - 0x30
    "00110010", -- 6781 - 0x1a7d  :   50 - 0x32
    "00110101", -- 6782 - 0x1a7e  :   53 - 0x35
    "00110010", -- 6783 - 0x1a7f  :   50 - 0x32
    "01001111", -- 6784 - 0x1a80  :   79 - 0x4f -- Background 0xa8
    "11001111", -- 6785 - 0x1a81  :  207 - 0xcf
    "00001011", -- 6786 - 0x1a82  :   11 - 0xb
    "00001111", -- 6787 - 0x1a83  :   15 - 0xf
    "11111111", -- 6788 - 0x1a84  :  255 - 0xff
    "11011101", -- 6789 - 0x1a85  :  221 - 0xdd
    "11111010", -- 6790 - 0x1a86  :  250 - 0xfa
    "11111101", -- 6791 - 0x1a87  :  253 - 0xfd
    "00110000", -- 6792 - 0x1a88  :   48 - 0x30
    "00110000", -- 6793 - 0x1a89  :   48 - 0x30
    "11110100", -- 6794 - 0x1a8a  :  244 - 0xf4
    "11110000", -- 6795 - 0x1a8b  :  240 - 0xf0
    "00000000", -- 6796 - 0x1a8c  :    0 - 0x0
    "00100010", -- 6797 - 0x1a8d  :   34 - 0x22
    "00000101", -- 6798 - 0x1a8e  :    5 - 0x5
    "00000010", -- 6799 - 0x1a8f  :    2 - 0x2
    "11111111", -- 6800 - 0x1a90  :  255 - 0xff -- Background 0xa9
    "11111111", -- 6801 - 0x1a91  :  255 - 0xff
    "11111111", -- 6802 - 0x1a92  :  255 - 0xff
    "11111111", -- 6803 - 0x1a93  :  255 - 0xff
    "11111111", -- 6804 - 0x1a94  :  255 - 0xff
    "11111111", -- 6805 - 0x1a95  :  255 - 0xff
    "11111111", -- 6806 - 0x1a96  :  255 - 0xff
    "11111111", -- 6807 - 0x1a97  :  255 - 0xff
    "00000000", -- 6808 - 0x1a98  :    0 - 0x0
    "00000000", -- 6809 - 0x1a99  :    0 - 0x0
    "00000000", -- 6810 - 0x1a9a  :    0 - 0x0
    "00000000", -- 6811 - 0x1a9b  :    0 - 0x0
    "00000000", -- 6812 - 0x1a9c  :    0 - 0x0
    "00000000", -- 6813 - 0x1a9d  :    0 - 0x0
    "00000000", -- 6814 - 0x1a9e  :    0 - 0x0
    "00000000", -- 6815 - 0x1a9f  :    0 - 0x0
    "11111111", -- 6816 - 0x1aa0  :  255 - 0xff -- Background 0xaa
    "11111111", -- 6817 - 0x1aa1  :  255 - 0xff
    "10101111", -- 6818 - 0x1aa2  :  175 - 0xaf
    "01010111", -- 6819 - 0x1aa3  :   87 - 0x57
    "10001111", -- 6820 - 0x1aa4  :  143 - 0x8f
    "11011101", -- 6821 - 0x1aa5  :  221 - 0xdd
    "11111010", -- 6822 - 0x1aa6  :  250 - 0xfa
    "11111101", -- 6823 - 0x1aa7  :  253 - 0xfd
    "00000000", -- 6824 - 0x1aa8  :    0 - 0x0
    "00000000", -- 6825 - 0x1aa9  :    0 - 0x0
    "01010000", -- 6826 - 0x1aaa  :   80 - 0x50
    "10101000", -- 6827 - 0x1aab  :  168 - 0xa8
    "01110000", -- 6828 - 0x1aac  :  112 - 0x70
    "00100010", -- 6829 - 0x1aad  :   34 - 0x22
    "00000101", -- 6830 - 0x1aae  :    5 - 0x5
    "00000010", -- 6831 - 0x1aaf  :    2 - 0x2
    "11111111", -- 6832 - 0x1ab0  :  255 - 0xff -- Background 0xab
    "00000000", -- 6833 - 0x1ab1  :    0 - 0x0
    "00000000", -- 6834 - 0x1ab2  :    0 - 0x0
    "00000000", -- 6835 - 0x1ab3  :    0 - 0x0
    "00000000", -- 6836 - 0x1ab4  :    0 - 0x0
    "00000000", -- 6837 - 0x1ab5  :    0 - 0x0
    "00000000", -- 6838 - 0x1ab6  :    0 - 0x0
    "00000000", -- 6839 - 0x1ab7  :    0 - 0x0
    "00000000", -- 6840 - 0x1ab8  :    0 - 0x0
    "00000000", -- 6841 - 0x1ab9  :    0 - 0x0
    "00000000", -- 6842 - 0x1aba  :    0 - 0x0
    "00000000", -- 6843 - 0x1abb  :    0 - 0x0
    "00000000", -- 6844 - 0x1abc  :    0 - 0x0
    "00000000", -- 6845 - 0x1abd  :    0 - 0x0
    "00000000", -- 6846 - 0x1abe  :    0 - 0x0
    "00000000", -- 6847 - 0x1abf  :    0 - 0x0
    "00000000", -- 6848 - 0x1ac0  :    0 - 0x0 -- Background 0xac
    "00000000", -- 6849 - 0x1ac1  :    0 - 0x0
    "00000000", -- 6850 - 0x1ac2  :    0 - 0x0
    "00000000", -- 6851 - 0x1ac3  :    0 - 0x0
    "00000000", -- 6852 - 0x1ac4  :    0 - 0x0
    "00000000", -- 6853 - 0x1ac5  :    0 - 0x0
    "00000000", -- 6854 - 0x1ac6  :    0 - 0x0
    "00000000", -- 6855 - 0x1ac7  :    0 - 0x0
    "00000000", -- 6856 - 0x1ac8  :    0 - 0x0
    "00000000", -- 6857 - 0x1ac9  :    0 - 0x0
    "00000000", -- 6858 - 0x1aca  :    0 - 0x0
    "00000000", -- 6859 - 0x1acb  :    0 - 0x0
    "00000000", -- 6860 - 0x1acc  :    0 - 0x0
    "00000000", -- 6861 - 0x1acd  :    0 - 0x0
    "00000000", -- 6862 - 0x1ace  :    0 - 0x0
    "00000000", -- 6863 - 0x1acf  :    0 - 0x0
    "00000000", -- 6864 - 0x1ad0  :    0 - 0x0 -- Background 0xad
    "11111111", -- 6865 - 0x1ad1  :  255 - 0xff
    "00000000", -- 6866 - 0x1ad2  :    0 - 0x0
    "11111111", -- 6867 - 0x1ad3  :  255 - 0xff
    "11111111", -- 6868 - 0x1ad4  :  255 - 0xff
    "11111111", -- 6869 - 0x1ad5  :  255 - 0xff
    "11111111", -- 6870 - 0x1ad6  :  255 - 0xff
    "11111111", -- 6871 - 0x1ad7  :  255 - 0xff
    "00000000", -- 6872 - 0x1ad8  :    0 - 0x0
    "00000000", -- 6873 - 0x1ad9  :    0 - 0x0
    "11111111", -- 6874 - 0x1ada  :  255 - 0xff
    "00000000", -- 6875 - 0x1adb  :    0 - 0x0
    "00000000", -- 6876 - 0x1adc  :    0 - 0x0
    "00000000", -- 6877 - 0x1add  :    0 - 0x0
    "00000000", -- 6878 - 0x1ade  :    0 - 0x0
    "00000000", -- 6879 - 0x1adf  :    0 - 0x0
    "11111111", -- 6880 - 0x1ae0  :  255 - 0xff -- Background 0xae
    "11111111", -- 6881 - 0x1ae1  :  255 - 0xff
    "11111111", -- 6882 - 0x1ae2  :  255 - 0xff
    "11111111", -- 6883 - 0x1ae3  :  255 - 0xff
    "11111111", -- 6884 - 0x1ae4  :  255 - 0xff
    "00000000", -- 6885 - 0x1ae5  :    0 - 0x0
    "11111111", -- 6886 - 0x1ae6  :  255 - 0xff
    "00000000", -- 6887 - 0x1ae7  :    0 - 0x0
    "00000000", -- 6888 - 0x1ae8  :    0 - 0x0
    "00000000", -- 6889 - 0x1ae9  :    0 - 0x0
    "00000000", -- 6890 - 0x1aea  :    0 - 0x0
    "00000000", -- 6891 - 0x1aeb  :    0 - 0x0
    "00000000", -- 6892 - 0x1aec  :    0 - 0x0
    "11111111", -- 6893 - 0x1aed  :  255 - 0xff
    "00000000", -- 6894 - 0x1aee  :    0 - 0x0
    "00000000", -- 6895 - 0x1aef  :    0 - 0x0
    "11111111", -- 6896 - 0x1af0  :  255 - 0xff -- Background 0xaf
    "11111111", -- 6897 - 0x1af1  :  255 - 0xff
    "11111111", -- 6898 - 0x1af2  :  255 - 0xff
    "11111111", -- 6899 - 0x1af3  :  255 - 0xff
    "11111111", -- 6900 - 0x1af4  :  255 - 0xff
    "11111111", -- 6901 - 0x1af5  :  255 - 0xff
    "11111111", -- 6902 - 0x1af6  :  255 - 0xff
    "11111111", -- 6903 - 0x1af7  :  255 - 0xff
    "00000000", -- 6904 - 0x1af8  :    0 - 0x0
    "00000000", -- 6905 - 0x1af9  :    0 - 0x0
    "00000000", -- 6906 - 0x1afa  :    0 - 0x0
    "00000000", -- 6907 - 0x1afb  :    0 - 0x0
    "00000000", -- 6908 - 0x1afc  :    0 - 0x0
    "00000000", -- 6909 - 0x1afd  :    0 - 0x0
    "00000000", -- 6910 - 0x1afe  :    0 - 0x0
    "00000000", -- 6911 - 0x1aff  :    0 - 0x0
    "00000000", -- 6912 - 0x1b00  :    0 - 0x0 -- Background 0xb0
    "00000000", -- 6913 - 0x1b01  :    0 - 0x0
    "00011111", -- 6914 - 0x1b02  :   31 - 0x1f
    "00010000", -- 6915 - 0x1b03  :   16 - 0x10
    "00010000", -- 6916 - 0x1b04  :   16 - 0x10
    "00010000", -- 6917 - 0x1b05  :   16 - 0x10
    "00010000", -- 6918 - 0x1b06  :   16 - 0x10
    "00010000", -- 6919 - 0x1b07  :   16 - 0x10
    "00000000", -- 6920 - 0x1b08  :    0 - 0x0
    "00000000", -- 6921 - 0x1b09  :    0 - 0x0
    "00011111", -- 6922 - 0x1b0a  :   31 - 0x1f
    "00011111", -- 6923 - 0x1b0b  :   31 - 0x1f
    "00011111", -- 6924 - 0x1b0c  :   31 - 0x1f
    "00011111", -- 6925 - 0x1b0d  :   31 - 0x1f
    "00011111", -- 6926 - 0x1b0e  :   31 - 0x1f
    "00011111", -- 6927 - 0x1b0f  :   31 - 0x1f
    "00000000", -- 6928 - 0x1b10  :    0 - 0x0 -- Background 0xb1
    "00000000", -- 6929 - 0x1b11  :    0 - 0x0
    "11111000", -- 6930 - 0x1b12  :  248 - 0xf8
    "00001000", -- 6931 - 0x1b13  :    8 - 0x8
    "00001000", -- 6932 - 0x1b14  :    8 - 0x8
    "00001000", -- 6933 - 0x1b15  :    8 - 0x8
    "00001000", -- 6934 - 0x1b16  :    8 - 0x8
    "00001000", -- 6935 - 0x1b17  :    8 - 0x8
    "00000000", -- 6936 - 0x1b18  :    0 - 0x0
    "00000000", -- 6937 - 0x1b19  :    0 - 0x0
    "11110000", -- 6938 - 0x1b1a  :  240 - 0xf0
    "11110000", -- 6939 - 0x1b1b  :  240 - 0xf0
    "11110000", -- 6940 - 0x1b1c  :  240 - 0xf0
    "11110000", -- 6941 - 0x1b1d  :  240 - 0xf0
    "11110000", -- 6942 - 0x1b1e  :  240 - 0xf0
    "11110000", -- 6943 - 0x1b1f  :  240 - 0xf0
    "00010000", -- 6944 - 0x1b20  :   16 - 0x10 -- Background 0xb2
    "00010000", -- 6945 - 0x1b21  :   16 - 0x10
    "00010000", -- 6946 - 0x1b22  :   16 - 0x10
    "00010000", -- 6947 - 0x1b23  :   16 - 0x10
    "00010000", -- 6948 - 0x1b24  :   16 - 0x10
    "00011111", -- 6949 - 0x1b25  :   31 - 0x1f
    "00011111", -- 6950 - 0x1b26  :   31 - 0x1f
    "00001111", -- 6951 - 0x1b27  :   15 - 0xf
    "00011111", -- 6952 - 0x1b28  :   31 - 0x1f
    "00011111", -- 6953 - 0x1b29  :   31 - 0x1f
    "00011111", -- 6954 - 0x1b2a  :   31 - 0x1f
    "00011111", -- 6955 - 0x1b2b  :   31 - 0x1f
    "00011111", -- 6956 - 0x1b2c  :   31 - 0x1f
    "00000000", -- 6957 - 0x1b2d  :    0 - 0x0
    "00000000", -- 6958 - 0x1b2e  :    0 - 0x0
    "00000000", -- 6959 - 0x1b2f  :    0 - 0x0
    "00001000", -- 6960 - 0x1b30  :    8 - 0x8 -- Background 0xb3
    "00001000", -- 6961 - 0x1b31  :    8 - 0x8
    "00001000", -- 6962 - 0x1b32  :    8 - 0x8
    "00001000", -- 6963 - 0x1b33  :    8 - 0x8
    "00001000", -- 6964 - 0x1b34  :    8 - 0x8
    "11111000", -- 6965 - 0x1b35  :  248 - 0xf8
    "11111000", -- 6966 - 0x1b36  :  248 - 0xf8
    "11110000", -- 6967 - 0x1b37  :  240 - 0xf0
    "11110000", -- 6968 - 0x1b38  :  240 - 0xf0
    "11110000", -- 6969 - 0x1b39  :  240 - 0xf0
    "11110000", -- 6970 - 0x1b3a  :  240 - 0xf0
    "11110000", -- 6971 - 0x1b3b  :  240 - 0xf0
    "11110000", -- 6972 - 0x1b3c  :  240 - 0xf0
    "00000000", -- 6973 - 0x1b3d  :    0 - 0x0
    "00000000", -- 6974 - 0x1b3e  :    0 - 0x0
    "00000000", -- 6975 - 0x1b3f  :    0 - 0x0
    "00000000", -- 6976 - 0x1b40  :    0 - 0x0 -- Background 0xb4
    "00000000", -- 6977 - 0x1b41  :    0 - 0x0
    "00000000", -- 6978 - 0x1b42  :    0 - 0x0
    "00111111", -- 6979 - 0x1b43  :   63 - 0x3f
    "01100000", -- 6980 - 0x1b44  :   96 - 0x60
    "01100000", -- 6981 - 0x1b45  :   96 - 0x60
    "01100000", -- 6982 - 0x1b46  :   96 - 0x60
    "01100000", -- 6983 - 0x1b47  :   96 - 0x60
    "00000000", -- 6984 - 0x1b48  :    0 - 0x0
    "00000000", -- 6985 - 0x1b49  :    0 - 0x0
    "00000000", -- 6986 - 0x1b4a  :    0 - 0x0
    "00111111", -- 6987 - 0x1b4b  :   63 - 0x3f
    "01111111", -- 6988 - 0x1b4c  :  127 - 0x7f
    "01111111", -- 6989 - 0x1b4d  :  127 - 0x7f
    "01111111", -- 6990 - 0x1b4e  :  127 - 0x7f
    "01111111", -- 6991 - 0x1b4f  :  127 - 0x7f
    "00000000", -- 6992 - 0x1b50  :    0 - 0x0 -- Background 0xb5
    "00000000", -- 6993 - 0x1b51  :    0 - 0x0
    "00000000", -- 6994 - 0x1b52  :    0 - 0x0
    "11111100", -- 6995 - 0x1b53  :  252 - 0xfc
    "00000110", -- 6996 - 0x1b54  :    6 - 0x6
    "00000110", -- 6997 - 0x1b55  :    6 - 0x6
    "00000110", -- 6998 - 0x1b56  :    6 - 0x6
    "00000110", -- 6999 - 0x1b57  :    6 - 0x6
    "00000000", -- 7000 - 0x1b58  :    0 - 0x0
    "00000000", -- 7001 - 0x1b59  :    0 - 0x0
    "00000000", -- 7002 - 0x1b5a  :    0 - 0x0
    "11111000", -- 7003 - 0x1b5b  :  248 - 0xf8
    "11111000", -- 7004 - 0x1b5c  :  248 - 0xf8
    "11111000", -- 7005 - 0x1b5d  :  248 - 0xf8
    "11111000", -- 7006 - 0x1b5e  :  248 - 0xf8
    "11111000", -- 7007 - 0x1b5f  :  248 - 0xf8
    "01100000", -- 7008 - 0x1b60  :   96 - 0x60 -- Background 0xb6
    "01100000", -- 7009 - 0x1b61  :   96 - 0x60
    "01100000", -- 7010 - 0x1b62  :   96 - 0x60
    "01100000", -- 7011 - 0x1b63  :   96 - 0x60
    "01111111", -- 7012 - 0x1b64  :  127 - 0x7f
    "01111111", -- 7013 - 0x1b65  :  127 - 0x7f
    "00111111", -- 7014 - 0x1b66  :   63 - 0x3f
    "00000000", -- 7015 - 0x1b67  :    0 - 0x0
    "01111111", -- 7016 - 0x1b68  :  127 - 0x7f
    "01111111", -- 7017 - 0x1b69  :  127 - 0x7f
    "01111111", -- 7018 - 0x1b6a  :  127 - 0x7f
    "01111111", -- 7019 - 0x1b6b  :  127 - 0x7f
    "01000000", -- 7020 - 0x1b6c  :   64 - 0x40
    "00000000", -- 7021 - 0x1b6d  :    0 - 0x0
    "00000000", -- 7022 - 0x1b6e  :    0 - 0x0
    "00000000", -- 7023 - 0x1b6f  :    0 - 0x0
    "00000110", -- 7024 - 0x1b70  :    6 - 0x6 -- Background 0xb7
    "00000110", -- 7025 - 0x1b71  :    6 - 0x6
    "00000110", -- 7026 - 0x1b72  :    6 - 0x6
    "00000110", -- 7027 - 0x1b73  :    6 - 0x6
    "11111110", -- 7028 - 0x1b74  :  254 - 0xfe
    "11111110", -- 7029 - 0x1b75  :  254 - 0xfe
    "11111100", -- 7030 - 0x1b76  :  252 - 0xfc
    "00000000", -- 7031 - 0x1b77  :    0 - 0x0
    "11111000", -- 7032 - 0x1b78  :  248 - 0xf8
    "11111000", -- 7033 - 0x1b79  :  248 - 0xf8
    "11111000", -- 7034 - 0x1b7a  :  248 - 0xf8
    "11111000", -- 7035 - 0x1b7b  :  248 - 0xf8
    "00000000", -- 7036 - 0x1b7c  :    0 - 0x0
    "00000000", -- 7037 - 0x1b7d  :    0 - 0x0
    "00000000", -- 7038 - 0x1b7e  :    0 - 0x0
    "00000000", -- 7039 - 0x1b7f  :    0 - 0x0
    "01100000", -- 7040 - 0x1b80  :   96 - 0x60 -- Background 0xb8
    "11110000", -- 7041 - 0x1b81  :  240 - 0xf0
    "11000011", -- 7042 - 0x1b82  :  195 - 0xc3
    "10000111", -- 7043 - 0x1b83  :  135 - 0x87
    "00000110", -- 7044 - 0x1b84  :    6 - 0x6
    "00000100", -- 7045 - 0x1b85  :    4 - 0x4
    "00000100", -- 7046 - 0x1b86  :    4 - 0x4
    "00000111", -- 7047 - 0x1b87  :    7 - 0x7
    "00000000", -- 7048 - 0x1b88  :    0 - 0x0
    "00000000", -- 7049 - 0x1b89  :    0 - 0x0
    "00000011", -- 7050 - 0x1b8a  :    3 - 0x3
    "00000111", -- 7051 - 0x1b8b  :    7 - 0x7
    "00000111", -- 7052 - 0x1b8c  :    7 - 0x7
    "00000111", -- 7053 - 0x1b8d  :    7 - 0x7
    "00000011", -- 7054 - 0x1b8e  :    3 - 0x3
    "00000000", -- 7055 - 0x1b8f  :    0 - 0x0
    "00000110", -- 7056 - 0x1b90  :    6 - 0x6 -- Background 0xb9
    "00001111", -- 7057 - 0x1b91  :   15 - 0xf
    "10000111", -- 7058 - 0x1b92  :  135 - 0x87
    "11000001", -- 7059 - 0x1b93  :  193 - 0xc1
    "00100011", -- 7060 - 0x1b94  :   35 - 0x23
    "00101110", -- 7061 - 0x1b95  :   46 - 0x2e
    "01100000", -- 7062 - 0x1b96  :   96 - 0x60
    "11100001", -- 7063 - 0x1b97  :  225 - 0xe1
    "00000000", -- 7064 - 0x1b98  :    0 - 0x0
    "00000000", -- 7065 - 0x1b99  :    0 - 0x0
    "11000001", -- 7066 - 0x1b9a  :  193 - 0xc1
    "11100010", -- 7067 - 0x1b9b  :  226 - 0xe2
    "11001100", -- 7068 - 0x1b9c  :  204 - 0xcc
    "11000000", -- 7069 - 0x1b9d  :  192 - 0xc0
    "10000000", -- 7070 - 0x1b9e  :  128 - 0x80
    "00000001", -- 7071 - 0x1b9f  :    1 - 0x1
    "00000000", -- 7072 - 0x1ba0  :    0 - 0x0 -- Background 0xba
    "11001000", -- 7073 - 0x1ba1  :  200 - 0xc8
    "11111000", -- 7074 - 0x1ba2  :  248 - 0xf8
    "10110000", -- 7075 - 0x1ba3  :  176 - 0xb0
    "00010000", -- 7076 - 0x1ba4  :   16 - 0x10
    "00110000", -- 7077 - 0x1ba5  :   48 - 0x30
    "11001000", -- 7078 - 0x1ba6  :  200 - 0xc8
    "11111000", -- 7079 - 0x1ba7  :  248 - 0xf8
    "00000000", -- 7080 - 0x1ba8  :    0 - 0x0
    "11110000", -- 7081 - 0x1ba9  :  240 - 0xf0
    "00000000", -- 7082 - 0x1baa  :    0 - 0x0
    "00100000", -- 7083 - 0x1bab  :   32 - 0x20
    "00100000", -- 7084 - 0x1bac  :   32 - 0x20
    "00000000", -- 7085 - 0x1bad  :    0 - 0x0
    "11110000", -- 7086 - 0x1bae  :  240 - 0xf0
    "00000000", -- 7087 - 0x1baf  :    0 - 0x0
    "00000111", -- 7088 - 0x1bb0  :    7 - 0x7 -- Background 0xbb
    "00000011", -- 7089 - 0x1bb1  :    3 - 0x3
    "00000000", -- 7090 - 0x1bb2  :    0 - 0x0
    "01100000", -- 7091 - 0x1bb3  :   96 - 0x60
    "11110000", -- 7092 - 0x1bb4  :  240 - 0xf0
    "11010000", -- 7093 - 0x1bb5  :  208 - 0xd0
    "10010000", -- 7094 - 0x1bb6  :  144 - 0x90
    "01100000", -- 7095 - 0x1bb7  :   96 - 0x60
    "00000000", -- 7096 - 0x1bb8  :    0 - 0x0
    "00000000", -- 7097 - 0x1bb9  :    0 - 0x0
    "00000000", -- 7098 - 0x1bba  :    0 - 0x0
    "00000000", -- 7099 - 0x1bbb  :    0 - 0x0
    "00000000", -- 7100 - 0x1bbc  :    0 - 0x0
    "01100000", -- 7101 - 0x1bbd  :   96 - 0x60
    "01100000", -- 7102 - 0x1bbe  :   96 - 0x60
    "00000000", -- 7103 - 0x1bbf  :    0 - 0x0
    "11100001", -- 7104 - 0x1bc0  :  225 - 0xe1 -- Background 0xbc
    "11000011", -- 7105 - 0x1bc1  :  195 - 0xc3
    "00001110", -- 7106 - 0x1bc2  :   14 - 0xe
    "00000110", -- 7107 - 0x1bc3  :    6 - 0x6
    "00001111", -- 7108 - 0x1bc4  :   15 - 0xf
    "00001101", -- 7109 - 0x1bc5  :   13 - 0xd
    "00001001", -- 7110 - 0x1bc6  :    9 - 0x9
    "00000110", -- 7111 - 0x1bc7  :    6 - 0x6
    "00000010", -- 7112 - 0x1bc8  :    2 - 0x2
    "00001100", -- 7113 - 0x1bc9  :   12 - 0xc
    "00000000", -- 7114 - 0x1bca  :    0 - 0x0
    "00000000", -- 7115 - 0x1bcb  :    0 - 0x0
    "00000000", -- 7116 - 0x1bcc  :    0 - 0x0
    "00000110", -- 7117 - 0x1bcd  :    6 - 0x6
    "00000110", -- 7118 - 0x1bce  :    6 - 0x6
    "00000000", -- 7119 - 0x1bcf  :    0 - 0x0
    "11100000", -- 7120 - 0x1bd0  :  224 - 0xe0 -- Background 0xbd
    "01100000", -- 7121 - 0x1bd1  :   96 - 0x60
    "11100011", -- 7122 - 0x1bd2  :  227 - 0xe3
    "11100111", -- 7123 - 0x1bd3  :  231 - 0xe7
    "00000110", -- 7124 - 0x1bd4  :    6 - 0x6
    "00000100", -- 7125 - 0x1bd5  :    4 - 0x4
    "00000100", -- 7126 - 0x1bd6  :    4 - 0x4
    "00000111", -- 7127 - 0x1bd7  :    7 - 0x7
    "00000000", -- 7128 - 0x1bd8  :    0 - 0x0
    "10000000", -- 7129 - 0x1bd9  :  128 - 0x80
    "00000011", -- 7130 - 0x1bda  :    3 - 0x3
    "00000111", -- 7131 - 0x1bdb  :    7 - 0x7
    "00000111", -- 7132 - 0x1bdc  :    7 - 0x7
    "00000111", -- 7133 - 0x1bdd  :    7 - 0x7
    "00000011", -- 7134 - 0x1bde  :    3 - 0x3
    "00000000", -- 7135 - 0x1bdf  :    0 - 0x0
    "00000111", -- 7136 - 0x1be0  :    7 - 0x7 -- Background 0xbe
    "00000011", -- 7137 - 0x1be1  :    3 - 0x3
    "10000111", -- 7138 - 0x1be2  :  135 - 0x87
    "11000111", -- 7139 - 0x1be3  :  199 - 0xc7
    "00100000", -- 7140 - 0x1be4  :   32 - 0x20
    "00100000", -- 7141 - 0x1be5  :   32 - 0x20
    "01100000", -- 7142 - 0x1be6  :   96 - 0x60
    "11100000", -- 7143 - 0x1be7  :  224 - 0xe0
    "00000000", -- 7144 - 0x1be8  :    0 - 0x0
    "00000100", -- 7145 - 0x1be9  :    4 - 0x4
    "11000000", -- 7146 - 0x1bea  :  192 - 0xc0
    "11100000", -- 7147 - 0x1beb  :  224 - 0xe0
    "11000000", -- 7148 - 0x1bec  :  192 - 0xc0
    "11000000", -- 7149 - 0x1bed  :  192 - 0xc0
    "10000000", -- 7150 - 0x1bee  :  128 - 0x80
    "00000000", -- 7151 - 0x1bef  :    0 - 0x0
    "00000111", -- 7152 - 0x1bf0  :    7 - 0x7 -- Background 0xbf
    "00000011", -- 7153 - 0x1bf1  :    3 - 0x3
    "00000000", -- 7154 - 0x1bf2  :    0 - 0x0
    "00001100", -- 7155 - 0x1bf3  :   12 - 0xc
    "11101100", -- 7156 - 0x1bf4  :  236 - 0xec
    "01100100", -- 7157 - 0x1bf5  :  100 - 0x64
    "11101100", -- 7158 - 0x1bf6  :  236 - 0xec
    "11101101", -- 7159 - 0x1bf7  :  237 - 0xed
    "00000000", -- 7160 - 0x1bf8  :    0 - 0x0
    "00000000", -- 7161 - 0x1bf9  :    0 - 0x0
    "00000000", -- 7162 - 0x1bfa  :    0 - 0x0
    "00000000", -- 7163 - 0x1bfb  :    0 - 0x0
    "00000000", -- 7164 - 0x1bfc  :    0 - 0x0
    "10001000", -- 7165 - 0x1bfd  :  136 - 0x88
    "00001000", -- 7166 - 0x1bfe  :    8 - 0x8
    "00001011", -- 7167 - 0x1bff  :   11 - 0xb
    "11100000", -- 7168 - 0x1c00  :  224 - 0xe0 -- Background 0xc0
    "11000000", -- 7169 - 0x1c01  :  192 - 0xc0
    "00000000", -- 7170 - 0x1c02  :    0 - 0x0
    "00110000", -- 7171 - 0x1c03  :   48 - 0x30
    "00110111", -- 7172 - 0x1c04  :   55 - 0x37
    "00010011", -- 7173 - 0x1c05  :   19 - 0x13
    "00110111", -- 7174 - 0x1c06  :   55 - 0x37
    "01110111", -- 7175 - 0x1c07  :  119 - 0x77
    "00000000", -- 7176 - 0x1c08  :    0 - 0x0
    "00000000", -- 7177 - 0x1c09  :    0 - 0x0
    "00000000", -- 7178 - 0x1c0a  :    0 - 0x0
    "00000000", -- 7179 - 0x1c0b  :    0 - 0x0
    "00000000", -- 7180 - 0x1c0c  :    0 - 0x0
    "00100100", -- 7181 - 0x1c0d  :   36 - 0x24
    "00100000", -- 7182 - 0x1c0e  :   32 - 0x20
    "10100000", -- 7183 - 0x1c0f  :  160 - 0xa0
    "00001111", -- 7184 - 0x1c10  :   15 - 0xf -- Background 0xc1
    "00001100", -- 7185 - 0x1c11  :   12 - 0xc
    "00000000", -- 7186 - 0x1c12  :    0 - 0x0
    "00000000", -- 7187 - 0x1c13  :    0 - 0x0
    "00000000", -- 7188 - 0x1c14  :    0 - 0x0
    "00000000", -- 7189 - 0x1c15  :    0 - 0x0
    "00000000", -- 7190 - 0x1c16  :    0 - 0x0
    "00000000", -- 7191 - 0x1c17  :    0 - 0x0
    "00000000", -- 7192 - 0x1c18  :    0 - 0x0
    "00000000", -- 7193 - 0x1c19  :    0 - 0x0
    "00000000", -- 7194 - 0x1c1a  :    0 - 0x0
    "00000000", -- 7195 - 0x1c1b  :    0 - 0x0
    "00000000", -- 7196 - 0x1c1c  :    0 - 0x0
    "00000000", -- 7197 - 0x1c1d  :    0 - 0x0
    "00000000", -- 7198 - 0x1c1e  :    0 - 0x0
    "00000000", -- 7199 - 0x1c1f  :    0 - 0x0
    "11110000", -- 7200 - 0x1c20  :  240 - 0xf0 -- Background 0xc2
    "00110000", -- 7201 - 0x1c21  :   48 - 0x30
    "00000000", -- 7202 - 0x1c22  :    0 - 0x0
    "00000000", -- 7203 - 0x1c23  :    0 - 0x0
    "00000000", -- 7204 - 0x1c24  :    0 - 0x0
    "00000000", -- 7205 - 0x1c25  :    0 - 0x0
    "00000000", -- 7206 - 0x1c26  :    0 - 0x0
    "00000000", -- 7207 - 0x1c27  :    0 - 0x0
    "00000000", -- 7208 - 0x1c28  :    0 - 0x0
    "00000000", -- 7209 - 0x1c29  :    0 - 0x0
    "00000000", -- 7210 - 0x1c2a  :    0 - 0x0
    "00000000", -- 7211 - 0x1c2b  :    0 - 0x0
    "00000000", -- 7212 - 0x1c2c  :    0 - 0x0
    "00000000", -- 7213 - 0x1c2d  :    0 - 0x0
    "00000000", -- 7214 - 0x1c2e  :    0 - 0x0
    "00000000", -- 7215 - 0x1c2f  :    0 - 0x0
    "00000000", -- 7216 - 0x1c30  :    0 - 0x0 -- Background 0xc3
    "00000000", -- 7217 - 0x1c31  :    0 - 0x0
    "00000000", -- 7218 - 0x1c32  :    0 - 0x0
    "00000100", -- 7219 - 0x1c33  :    4 - 0x4
    "00001101", -- 7220 - 0x1c34  :   13 - 0xd
    "00001111", -- 7221 - 0x1c35  :   15 - 0xf
    "00001100", -- 7222 - 0x1c36  :   12 - 0xc
    "00001100", -- 7223 - 0x1c37  :   12 - 0xc
    "00000000", -- 7224 - 0x1c38  :    0 - 0x0
    "00000000", -- 7225 - 0x1c39  :    0 - 0x0
    "00000000", -- 7226 - 0x1c3a  :    0 - 0x0
    "00001000", -- 7227 - 0x1c3b  :    8 - 0x8
    "00001011", -- 7228 - 0x1c3c  :   11 - 0xb
    "00001000", -- 7229 - 0x1c3d  :    8 - 0x8
    "00001000", -- 7230 - 0x1c3e  :    8 - 0x8
    "00001000", -- 7231 - 0x1c3f  :    8 - 0x8
    "00000000", -- 7232 - 0x1c40  :    0 - 0x0 -- Background 0xc4
    "00000000", -- 7233 - 0x1c41  :    0 - 0x0
    "00000000", -- 7234 - 0x1c42  :    0 - 0x0
    "00010000", -- 7235 - 0x1c43  :   16 - 0x10
    "01110000", -- 7236 - 0x1c44  :  112 - 0x70
    "11110000", -- 7237 - 0x1c45  :  240 - 0xf0
    "00110000", -- 7238 - 0x1c46  :   48 - 0x30
    "00110000", -- 7239 - 0x1c47  :   48 - 0x30
    "00000000", -- 7240 - 0x1c48  :    0 - 0x0
    "00000000", -- 7241 - 0x1c49  :    0 - 0x0
    "00000000", -- 7242 - 0x1c4a  :    0 - 0x0
    "00100000", -- 7243 - 0x1c4b  :   32 - 0x20
    "10100000", -- 7244 - 0x1c4c  :  160 - 0xa0
    "00100000", -- 7245 - 0x1c4d  :   32 - 0x20
    "00100000", -- 7246 - 0x1c4e  :   32 - 0x20
    "00100000", -- 7247 - 0x1c4f  :   32 - 0x20
    "11100100", -- 7248 - 0x1c50  :  228 - 0xe4 -- Background 0xc5
    "00100100", -- 7249 - 0x1c51  :   36 - 0x24
    "11100100", -- 7250 - 0x1c52  :  228 - 0xe4
    "11101111", -- 7251 - 0x1c53  :  239 - 0xef
    "00000111", -- 7252 - 0x1c54  :    7 - 0x7
    "00000110", -- 7253 - 0x1c55  :    6 - 0x6
    "00000100", -- 7254 - 0x1c56  :    4 - 0x4
    "00000100", -- 7255 - 0x1c57  :    4 - 0x4
    "00001000", -- 7256 - 0x1c58  :    8 - 0x8
    "11001000", -- 7257 - 0x1c59  :  200 - 0xc8
    "00001000", -- 7258 - 0x1c5a  :    8 - 0x8
    "00000011", -- 7259 - 0x1c5b  :    3 - 0x3
    "00000111", -- 7260 - 0x1c5c  :    7 - 0x7
    "00000111", -- 7261 - 0x1c5d  :    7 - 0x7
    "00000111", -- 7262 - 0x1c5e  :    7 - 0x7
    "00000011", -- 7263 - 0x1c5f  :    3 - 0x3
    "00010111", -- 7264 - 0x1c60  :   23 - 0x17 -- Background 0xc6
    "00010001", -- 7265 - 0x1c61  :   17 - 0x11
    "00010111", -- 7266 - 0x1c62  :   23 - 0x17
    "10110111", -- 7267 - 0x1c63  :  183 - 0xb7
    "11000000", -- 7268 - 0x1c64  :  192 - 0xc0
    "00100000", -- 7269 - 0x1c65  :   32 - 0x20
    "00100000", -- 7270 - 0x1c66  :   32 - 0x20
    "01100000", -- 7271 - 0x1c67  :   96 - 0x60
    "00100000", -- 7272 - 0x1c68  :   32 - 0x20
    "00100110", -- 7273 - 0x1c69  :   38 - 0x26
    "00100000", -- 7274 - 0x1c6a  :   32 - 0x20
    "11000000", -- 7275 - 0x1c6b  :  192 - 0xc0
    "11100000", -- 7276 - 0x1c6c  :  224 - 0xe0
    "11000000", -- 7277 - 0x1c6d  :  192 - 0xc0
    "11000000", -- 7278 - 0x1c6e  :  192 - 0xc0
    "10000000", -- 7279 - 0x1c6f  :  128 - 0x80
    "00000111", -- 7280 - 0x1c70  :    7 - 0x7 -- Background 0xc7
    "00000111", -- 7281 - 0x1c71  :    7 - 0x7
    "00000011", -- 7282 - 0x1c72  :    3 - 0x3
    "00000000", -- 7283 - 0x1c73  :    0 - 0x0
    "11100000", -- 7284 - 0x1c74  :  224 - 0xe0
    "00100000", -- 7285 - 0x1c75  :   32 - 0x20
    "11100000", -- 7286 - 0x1c76  :  224 - 0xe0
    "11100000", -- 7287 - 0x1c77  :  224 - 0xe0
    "00000000", -- 7288 - 0x1c78  :    0 - 0x0
    "00000000", -- 7289 - 0x1c79  :    0 - 0x0
    "00000000", -- 7290 - 0x1c7a  :    0 - 0x0
    "00000000", -- 7291 - 0x1c7b  :    0 - 0x0
    "00000000", -- 7292 - 0x1c7c  :    0 - 0x0
    "11000000", -- 7293 - 0x1c7d  :  192 - 0xc0
    "00000000", -- 7294 - 0x1c7e  :    0 - 0x0
    "00000000", -- 7295 - 0x1c7f  :    0 - 0x0
    "11100000", -- 7296 - 0x1c80  :  224 - 0xe0 -- Background 0xc8
    "11100000", -- 7297 - 0x1c81  :  224 - 0xe0
    "11000000", -- 7298 - 0x1c82  :  192 - 0xc0
    "00000000", -- 7299 - 0x1c83  :    0 - 0x0
    "00000111", -- 7300 - 0x1c84  :    7 - 0x7
    "00000001", -- 7301 - 0x1c85  :    1 - 0x1
    "00000111", -- 7302 - 0x1c86  :    7 - 0x7
    "00000111", -- 7303 - 0x1c87  :    7 - 0x7
    "00000000", -- 7304 - 0x1c88  :    0 - 0x0
    "00000000", -- 7305 - 0x1c89  :    0 - 0x0
    "00000000", -- 7306 - 0x1c8a  :    0 - 0x0
    "00000000", -- 7307 - 0x1c8b  :    0 - 0x0
    "00000000", -- 7308 - 0x1c8c  :    0 - 0x0
    "00000110", -- 7309 - 0x1c8d  :    6 - 0x6
    "00000000", -- 7310 - 0x1c8e  :    0 - 0x0
    "00000000", -- 7311 - 0x1c8f  :    0 - 0x0
    "00000001", -- 7312 - 0x1c90  :    1 - 0x1 -- Background 0xc9
    "00010011", -- 7313 - 0x1c91  :   19 - 0x13
    "00011111", -- 7314 - 0x1c92  :   31 - 0x1f
    "00001101", -- 7315 - 0x1c93  :   13 - 0xd
    "00000100", -- 7316 - 0x1c94  :    4 - 0x4
    "00001100", -- 7317 - 0x1c95  :   12 - 0xc
    "00010011", -- 7318 - 0x1c96  :   19 - 0x13
    "00011111", -- 7319 - 0x1c97  :   31 - 0x1f
    "00000000", -- 7320 - 0x1c98  :    0 - 0x0
    "00001111", -- 7321 - 0x1c99  :   15 - 0xf
    "00000000", -- 7322 - 0x1c9a  :    0 - 0x0
    "00001000", -- 7323 - 0x1c9b  :    8 - 0x8
    "00001000", -- 7324 - 0x1c9c  :    8 - 0x8
    "00000000", -- 7325 - 0x1c9d  :    0 - 0x0
    "00001111", -- 7326 - 0x1c9e  :   15 - 0xf
    "00000000", -- 7327 - 0x1c9f  :    0 - 0x0
    "01100000", -- 7328 - 0x1ca0  :   96 - 0x60 -- Background 0xca
    "01110000", -- 7329 - 0x1ca1  :  112 - 0x70
    "10100011", -- 7330 - 0x1ca2  :  163 - 0xa3
    "10000111", -- 7331 - 0x1ca3  :  135 - 0x87
    "11000110", -- 7332 - 0x1ca4  :  198 - 0xc6
    "01110100", -- 7333 - 0x1ca5  :  116 - 0x74
    "00000100", -- 7334 - 0x1ca6  :    4 - 0x4
    "10000111", -- 7335 - 0x1ca7  :  135 - 0x87
    "00000000", -- 7336 - 0x1ca8  :    0 - 0x0
    "00000000", -- 7337 - 0x1ca9  :    0 - 0x0
    "10000011", -- 7338 - 0x1caa  :  131 - 0x83
    "01000111", -- 7339 - 0x1cab  :   71 - 0x47
    "00110111", -- 7340 - 0x1cac  :   55 - 0x37
    "00000111", -- 7341 - 0x1cad  :    7 - 0x7
    "00000011", -- 7342 - 0x1cae  :    3 - 0x3
    "10000000", -- 7343 - 0x1caf  :  128 - 0x80
    "00000110", -- 7344 - 0x1cb0  :    6 - 0x6 -- Background 0xcb
    "00001111", -- 7345 - 0x1cb1  :   15 - 0xf
    "10000011", -- 7346 - 0x1cb2  :  131 - 0x83
    "11000001", -- 7347 - 0x1cb3  :  193 - 0xc1
    "00100000", -- 7348 - 0x1cb4  :   32 - 0x20
    "00100000", -- 7349 - 0x1cb5  :   32 - 0x20
    "01100000", -- 7350 - 0x1cb6  :   96 - 0x60
    "11100000", -- 7351 - 0x1cb7  :  224 - 0xe0
    "00000000", -- 7352 - 0x1cb8  :    0 - 0x0
    "00000000", -- 7353 - 0x1cb9  :    0 - 0x0
    "11000000", -- 7354 - 0x1cba  :  192 - 0xc0
    "11100000", -- 7355 - 0x1cbb  :  224 - 0xe0
    "11000000", -- 7356 - 0x1cbc  :  192 - 0xc0
    "11000000", -- 7357 - 0x1cbd  :  192 - 0xc0
    "10000000", -- 7358 - 0x1cbe  :  128 - 0x80
    "00000000", -- 7359 - 0x1cbf  :    0 - 0x0
    "10000111", -- 7360 - 0x1cc0  :  135 - 0x87 -- Background 0xcc
    "01000011", -- 7361 - 0x1cc1  :   67 - 0x43
    "00110000", -- 7362 - 0x1cc2  :   48 - 0x30
    "01100000", -- 7363 - 0x1cc3  :   96 - 0x60
    "11110000", -- 7364 - 0x1cc4  :  240 - 0xf0
    "11010000", -- 7365 - 0x1cc5  :  208 - 0xd0
    "10010000", -- 7366 - 0x1cc6  :  144 - 0x90
    "01100000", -- 7367 - 0x1cc7  :   96 - 0x60
    "01000000", -- 7368 - 0x1cc8  :   64 - 0x40
    "00110000", -- 7369 - 0x1cc9  :   48 - 0x30
    "00000000", -- 7370 - 0x1cca  :    0 - 0x0
    "00000000", -- 7371 - 0x1ccb  :    0 - 0x0
    "00000000", -- 7372 - 0x1ccc  :    0 - 0x0
    "01100000", -- 7373 - 0x1ccd  :   96 - 0x60
    "01100000", -- 7374 - 0x1cce  :   96 - 0x60
    "00000000", -- 7375 - 0x1ccf  :    0 - 0x0
    "11100000", -- 7376 - 0x1cd0  :  224 - 0xe0 -- Background 0xcd
    "11000000", -- 7377 - 0x1cd1  :  192 - 0xc0
    "00000000", -- 7378 - 0x1cd2  :    0 - 0x0
    "00000110", -- 7379 - 0x1cd3  :    6 - 0x6
    "00001111", -- 7380 - 0x1cd4  :   15 - 0xf
    "00001101", -- 7381 - 0x1cd5  :   13 - 0xd
    "00001001", -- 7382 - 0x1cd6  :    9 - 0x9
    "00000110", -- 7383 - 0x1cd7  :    6 - 0x6
    "00000000", -- 7384 - 0x1cd8  :    0 - 0x0
    "00000000", -- 7385 - 0x1cd9  :    0 - 0x0
    "00000000", -- 7386 - 0x1cda  :    0 - 0x0
    "00000000", -- 7387 - 0x1cdb  :    0 - 0x0
    "00000000", -- 7388 - 0x1cdc  :    0 - 0x0
    "00000110", -- 7389 - 0x1cdd  :    6 - 0x6
    "00000110", -- 7390 - 0x1cde  :    6 - 0x6
    "00000000", -- 7391 - 0x1cdf  :    0 - 0x0
    "11111100", -- 7392 - 0x1ce0  :  252 - 0xfc -- Background 0xce
    "11000000", -- 7393 - 0x1ce1  :  192 - 0xc0
    "11010001", -- 7394 - 0x1ce2  :  209 - 0xd1
    "11000010", -- 7395 - 0x1ce3  :  194 - 0xc2
    "10011110", -- 7396 - 0x1ce4  :  158 - 0x9e
    "10111111", -- 7397 - 0x1ce5  :  191 - 0xbf
    "10110000", -- 7398 - 0x1ce6  :  176 - 0xb0
    "10110011", -- 7399 - 0x1ce7  :  179 - 0xb3
    "00000000", -- 7400 - 0x1ce8  :    0 - 0x0
    "00000001", -- 7401 - 0x1ce9  :    1 - 0x1
    "00011011", -- 7402 - 0x1cea  :   27 - 0x1b
    "00010011", -- 7403 - 0x1ceb  :   19 - 0x13
    "00011111", -- 7404 - 0x1cec  :   31 - 0x1f
    "00111111", -- 7405 - 0x1ced  :   63 - 0x3f
    "00111111", -- 7406 - 0x1cee  :   63 - 0x3f
    "00111111", -- 7407 - 0x1cef  :   63 - 0x3f
    "00000111", -- 7408 - 0x1cf0  :    7 - 0x7 -- Background 0xcf
    "11110011", -- 7409 - 0x1cf1  :  243 - 0xf3
    "00001011", -- 7410 - 0x1cf2  :   11 - 0xb
    "01111011", -- 7411 - 0x1cf3  :  123 - 0x7b
    "01111011", -- 7412 - 0x1cf4  :  123 - 0x7b
    "11111001", -- 7413 - 0x1cf5  :  249 - 0xf9
    "00001101", -- 7414 - 0x1cf6  :   13 - 0xd
    "11101101", -- 7415 - 0x1cf7  :  237 - 0xed
    "00000000", -- 7416 - 0x1cf8  :    0 - 0x0
    "11111000", -- 7417 - 0x1cf9  :  248 - 0xf8
    "00001000", -- 7418 - 0x1cfa  :    8 - 0x8
    "00001000", -- 7419 - 0x1cfb  :    8 - 0x8
    "00001000", -- 7420 - 0x1cfc  :    8 - 0x8
    "11111000", -- 7421 - 0x1cfd  :  248 - 0xf8
    "11110000", -- 7422 - 0x1cfe  :  240 - 0xf0
    "11010000", -- 7423 - 0x1cff  :  208 - 0xd0
    "11111111", -- 7424 - 0x1d00  :  255 - 0xff -- Background 0xd0
    "11111111", -- 7425 - 0x1d01  :  255 - 0xff
    "11111111", -- 7426 - 0x1d02  :  255 - 0xff
    "11111111", -- 7427 - 0x1d03  :  255 - 0xff
    "11101110", -- 7428 - 0x1d04  :  238 - 0xee
    "11101110", -- 7429 - 0x1d05  :  238 - 0xee
    "11101110", -- 7430 - 0x1d06  :  238 - 0xee
    "11101110", -- 7431 - 0x1d07  :  238 - 0xee
    "00000000", -- 7432 - 0x1d08  :    0 - 0x0
    "00000000", -- 7433 - 0x1d09  :    0 - 0x0
    "01111100", -- 7434 - 0x1d0a  :  124 - 0x7c
    "11111110", -- 7435 - 0x1d0b  :  254 - 0xfe
    "11101110", -- 7436 - 0x1d0c  :  238 - 0xee
    "11101110", -- 7437 - 0x1d0d  :  238 - 0xee
    "11101110", -- 7438 - 0x1d0e  :  238 - 0xee
    "11101110", -- 7439 - 0x1d0f  :  238 - 0xee
    "11111111", -- 7440 - 0x1d10  :  255 - 0xff -- Background 0xd1
    "11111111", -- 7441 - 0x1d11  :  255 - 0xff
    "11111111", -- 7442 - 0x1d12  :  255 - 0xff
    "11111011", -- 7443 - 0x1d13  :  251 - 0xfb
    "11111011", -- 7444 - 0x1d14  :  251 - 0xfb
    "11111011", -- 7445 - 0x1d15  :  251 - 0xfb
    "11111011", -- 7446 - 0x1d16  :  251 - 0xfb
    "11111011", -- 7447 - 0x1d17  :  251 - 0xfb
    "00000000", -- 7448 - 0x1d18  :    0 - 0x0
    "00000000", -- 7449 - 0x1d19  :    0 - 0x0
    "00111000", -- 7450 - 0x1d1a  :   56 - 0x38
    "01111000", -- 7451 - 0x1d1b  :  120 - 0x78
    "01111000", -- 7452 - 0x1d1c  :  120 - 0x78
    "00111000", -- 7453 - 0x1d1d  :   56 - 0x38
    "00111000", -- 7454 - 0x1d1e  :   56 - 0x38
    "00111000", -- 7455 - 0x1d1f  :   56 - 0x38
    "11111111", -- 7456 - 0x1d20  :  255 - 0xff -- Background 0xd2
    "11111111", -- 7457 - 0x1d21  :  255 - 0xff
    "11111111", -- 7458 - 0x1d22  :  255 - 0xff
    "11111111", -- 7459 - 0x1d23  :  255 - 0xff
    "11101110", -- 7460 - 0x1d24  :  238 - 0xee
    "10001110", -- 7461 - 0x1d25  :  142 - 0x8e
    "11111110", -- 7462 - 0x1d26  :  254 - 0xfe
    "11111110", -- 7463 - 0x1d27  :  254 - 0xfe
    "00000000", -- 7464 - 0x1d28  :    0 - 0x0
    "00000000", -- 7465 - 0x1d29  :    0 - 0x0
    "01111100", -- 7466 - 0x1d2a  :  124 - 0x7c
    "11111110", -- 7467 - 0x1d2b  :  254 - 0xfe
    "11101110", -- 7468 - 0x1d2c  :  238 - 0xee
    "00001110", -- 7469 - 0x1d2d  :   14 - 0xe
    "00001110", -- 7470 - 0x1d2e  :   14 - 0xe
    "01111110", -- 7471 - 0x1d2f  :  126 - 0x7e
    "11111111", -- 7472 - 0x1d30  :  255 - 0xff -- Background 0xd3
    "11111111", -- 7473 - 0x1d31  :  255 - 0xff
    "11111111", -- 7474 - 0x1d32  :  255 - 0xff
    "11111111", -- 7475 - 0x1d33  :  255 - 0xff
    "11101110", -- 7476 - 0x1d34  :  238 - 0xee
    "10001110", -- 7477 - 0x1d35  :  142 - 0x8e
    "11111100", -- 7478 - 0x1d36  :  252 - 0xfc
    "11111101", -- 7479 - 0x1d37  :  253 - 0xfd
    "00000000", -- 7480 - 0x1d38  :    0 - 0x0
    "00000000", -- 7481 - 0x1d39  :    0 - 0x0
    "01111100", -- 7482 - 0x1d3a  :  124 - 0x7c
    "11111110", -- 7483 - 0x1d3b  :  254 - 0xfe
    "11101110", -- 7484 - 0x1d3c  :  238 - 0xee
    "00001110", -- 7485 - 0x1d3d  :   14 - 0xe
    "00111100", -- 7486 - 0x1d3e  :   60 - 0x3c
    "00111100", -- 7487 - 0x1d3f  :   60 - 0x3c
    "11111111", -- 7488 - 0x1d40  :  255 - 0xff -- Background 0xd4
    "11111111", -- 7489 - 0x1d41  :  255 - 0xff
    "11111111", -- 7490 - 0x1d42  :  255 - 0xff
    "11111110", -- 7491 - 0x1d43  :  254 - 0xfe
    "11101110", -- 7492 - 0x1d44  :  238 - 0xee
    "11101110", -- 7493 - 0x1d45  :  238 - 0xee
    "11101110", -- 7494 - 0x1d46  :  238 - 0xee
    "11101110", -- 7495 - 0x1d47  :  238 - 0xee
    "00000000", -- 7496 - 0x1d48  :    0 - 0x0
    "00000000", -- 7497 - 0x1d49  :    0 - 0x0
    "00111110", -- 7498 - 0x1d4a  :   62 - 0x3e
    "01111110", -- 7499 - 0x1d4b  :  126 - 0x7e
    "11101110", -- 7500 - 0x1d4c  :  238 - 0xee
    "11101110", -- 7501 - 0x1d4d  :  238 - 0xee
    "11101110", -- 7502 - 0x1d4e  :  238 - 0xee
    "11101110", -- 7503 - 0x1d4f  :  238 - 0xee
    "11111111", -- 7504 - 0x1d50  :  255 - 0xff -- Background 0xd5
    "11111111", -- 7505 - 0x1d51  :  255 - 0xff
    "11111111", -- 7506 - 0x1d52  :  255 - 0xff
    "11111101", -- 7507 - 0x1d53  :  253 - 0xfd
    "11100001", -- 7508 - 0x1d54  :  225 - 0xe1
    "11101111", -- 7509 - 0x1d55  :  239 - 0xef
    "11111111", -- 7510 - 0x1d56  :  255 - 0xff
    "11111111", -- 7511 - 0x1d57  :  255 - 0xff
    "00000000", -- 7512 - 0x1d58  :    0 - 0x0
    "00000000", -- 7513 - 0x1d59  :    0 - 0x0
    "11111100", -- 7514 - 0x1d5a  :  252 - 0xfc
    "11111100", -- 7515 - 0x1d5b  :  252 - 0xfc
    "11100000", -- 7516 - 0x1d5c  :  224 - 0xe0
    "11100000", -- 7517 - 0x1d5d  :  224 - 0xe0
    "11111100", -- 7518 - 0x1d5e  :  252 - 0xfc
    "11111110", -- 7519 - 0x1d5f  :  254 - 0xfe
    "11111111", -- 7520 - 0x1d60  :  255 - 0xff -- Background 0xd6
    "11111111", -- 7521 - 0x1d61  :  255 - 0xff
    "11111111", -- 7522 - 0x1d62  :  255 - 0xff
    "11111101", -- 7523 - 0x1d63  :  253 - 0xfd
    "11100001", -- 7524 - 0x1d64  :  225 - 0xe1
    "11101111", -- 7525 - 0x1d65  :  239 - 0xef
    "11111111", -- 7526 - 0x1d66  :  255 - 0xff
    "11111111", -- 7527 - 0x1d67  :  255 - 0xff
    "00000000", -- 7528 - 0x1d68  :    0 - 0x0
    "00000000", -- 7529 - 0x1d69  :    0 - 0x0
    "01111100", -- 7530 - 0x1d6a  :  124 - 0x7c
    "11111100", -- 7531 - 0x1d6b  :  252 - 0xfc
    "11100000", -- 7532 - 0x1d6c  :  224 - 0xe0
    "11100000", -- 7533 - 0x1d6d  :  224 - 0xe0
    "11111100", -- 7534 - 0x1d6e  :  252 - 0xfc
    "11111110", -- 7535 - 0x1d6f  :  254 - 0xfe
    "11111111", -- 7536 - 0x1d70  :  255 - 0xff -- Background 0xd7
    "11111111", -- 7537 - 0x1d71  :  255 - 0xff
    "11111111", -- 7538 - 0x1d72  :  255 - 0xff
    "11111110", -- 7539 - 0x1d73  :  254 - 0xfe
    "11101110", -- 7540 - 0x1d74  :  238 - 0xee
    "10001110", -- 7541 - 0x1d75  :  142 - 0x8e
    "11111110", -- 7542 - 0x1d76  :  254 - 0xfe
    "11111100", -- 7543 - 0x1d77  :  252 - 0xfc
    "00000000", -- 7544 - 0x1d78  :    0 - 0x0
    "00000000", -- 7545 - 0x1d79  :    0 - 0x0
    "11111110", -- 7546 - 0x1d7a  :  254 - 0xfe
    "11111110", -- 7547 - 0x1d7b  :  254 - 0xfe
    "11101110", -- 7548 - 0x1d7c  :  238 - 0xee
    "00001110", -- 7549 - 0x1d7d  :   14 - 0xe
    "00001110", -- 7550 - 0x1d7e  :   14 - 0xe
    "00011100", -- 7551 - 0x1d7f  :   28 - 0x1c
    "11111111", -- 7552 - 0x1d80  :  255 - 0xff -- Background 0xd8
    "11111111", -- 7553 - 0x1d81  :  255 - 0xff
    "11111111", -- 7554 - 0x1d82  :  255 - 0xff
    "11111111", -- 7555 - 0x1d83  :  255 - 0xff
    "11101110", -- 7556 - 0x1d84  :  238 - 0xee
    "11101110", -- 7557 - 0x1d85  :  238 - 0xee
    "11111100", -- 7558 - 0x1d86  :  252 - 0xfc
    "11111111", -- 7559 - 0x1d87  :  255 - 0xff
    "00000000", -- 7560 - 0x1d88  :    0 - 0x0
    "00000000", -- 7561 - 0x1d89  :    0 - 0x0
    "01111100", -- 7562 - 0x1d8a  :  124 - 0x7c
    "11111110", -- 7563 - 0x1d8b  :  254 - 0xfe
    "11101110", -- 7564 - 0x1d8c  :  238 - 0xee
    "11101110", -- 7565 - 0x1d8d  :  238 - 0xee
    "01111100", -- 7566 - 0x1d8e  :  124 - 0x7c
    "11111110", -- 7567 - 0x1d8f  :  254 - 0xfe
    "11111111", -- 7568 - 0x1d90  :  255 - 0xff -- Background 0xd9
    "11111111", -- 7569 - 0x1d91  :  255 - 0xff
    "11111111", -- 7570 - 0x1d92  :  255 - 0xff
    "11111111", -- 7571 - 0x1d93  :  255 - 0xff
    "11101110", -- 7572 - 0x1d94  :  238 - 0xee
    "11101110", -- 7573 - 0x1d95  :  238 - 0xee
    "11101110", -- 7574 - 0x1d96  :  238 - 0xee
    "11101110", -- 7575 - 0x1d97  :  238 - 0xee
    "00000000", -- 7576 - 0x1d98  :    0 - 0x0
    "00000000", -- 7577 - 0x1d99  :    0 - 0x0
    "01111100", -- 7578 - 0x1d9a  :  124 - 0x7c
    "11111110", -- 7579 - 0x1d9b  :  254 - 0xfe
    "11101110", -- 7580 - 0x1d9c  :  238 - 0xee
    "11101110", -- 7581 - 0x1d9d  :  238 - 0xee
    "11101110", -- 7582 - 0x1d9e  :  238 - 0xee
    "11101110", -- 7583 - 0x1d9f  :  238 - 0xee
    "00000000", -- 7584 - 0x1da0  :    0 - 0x0 -- Background 0xda
    "00000000", -- 7585 - 0x1da1  :    0 - 0x0
    "00000000", -- 7586 - 0x1da2  :    0 - 0x0
    "10000000", -- 7587 - 0x1da3  :  128 - 0x80
    "00000000", -- 7588 - 0x1da4  :    0 - 0x0
    "00000000", -- 7589 - 0x1da5  :    0 - 0x0
    "00000100", -- 7590 - 0x1da6  :    4 - 0x4
    "00000000", -- 7591 - 0x1da7  :    0 - 0x0
    "00000000", -- 7592 - 0x1da8  :    0 - 0x0
    "00100000", -- 7593 - 0x1da9  :   32 - 0x20
    "00000000", -- 7594 - 0x1daa  :    0 - 0x0
    "00000010", -- 7595 - 0x1dab  :    2 - 0x2
    "00000000", -- 7596 - 0x1dac  :    0 - 0x0
    "00100000", -- 7597 - 0x1dad  :   32 - 0x20
    "00000000", -- 7598 - 0x1dae  :    0 - 0x0
    "00000000", -- 7599 - 0x1daf  :    0 - 0x0
    "00000000", -- 7600 - 0x1db0  :    0 - 0x0 -- Background 0xdb
    "00000100", -- 7601 - 0x1db1  :    4 - 0x4
    "00000000", -- 7602 - 0x1db2  :    0 - 0x0
    "00010001", -- 7603 - 0x1db3  :   17 - 0x11
    "00000000", -- 7604 - 0x1db4  :    0 - 0x0
    "00000000", -- 7605 - 0x1db5  :    0 - 0x0
    "00000000", -- 7606 - 0x1db6  :    0 - 0x0
    "00100000", -- 7607 - 0x1db7  :   32 - 0x20
    "00100000", -- 7608 - 0x1db8  :   32 - 0x20
    "00000000", -- 7609 - 0x1db9  :    0 - 0x0
    "00000000", -- 7610 - 0x1dba  :    0 - 0x0
    "00000000", -- 7611 - 0x1dbb  :    0 - 0x0
    "10000000", -- 7612 - 0x1dbc  :  128 - 0x80
    "00000000", -- 7613 - 0x1dbd  :    0 - 0x0
    "00000100", -- 7614 - 0x1dbe  :    4 - 0x4
    "00000000", -- 7615 - 0x1dbf  :    0 - 0x0
    "00000000", -- 7616 - 0x1dc0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 7617 - 0x1dc1  :    0 - 0x0
    "00000000", -- 7618 - 0x1dc2  :    0 - 0x0
    "00100000", -- 7619 - 0x1dc3  :   32 - 0x20
    "00000000", -- 7620 - 0x1dc4  :    0 - 0x0
    "00000000", -- 7621 - 0x1dc5  :    0 - 0x0
    "00000000", -- 7622 - 0x1dc6  :    0 - 0x0
    "00000100", -- 7623 - 0x1dc7  :    4 - 0x4
    "00000000", -- 7624 - 0x1dc8  :    0 - 0x0
    "00001000", -- 7625 - 0x1dc9  :    8 - 0x8
    "00000000", -- 7626 - 0x1dca  :    0 - 0x0
    "00000000", -- 7627 - 0x1dcb  :    0 - 0x0
    "00000010", -- 7628 - 0x1dcc  :    2 - 0x2
    "00000000", -- 7629 - 0x1dcd  :    0 - 0x0
    "01000000", -- 7630 - 0x1dce  :   64 - 0x40
    "00000000", -- 7631 - 0x1dcf  :    0 - 0x0
    "00000000", -- 7632 - 0x1dd0  :    0 - 0x0 -- Background 0xdd
    "00000000", -- 7633 - 0x1dd1  :    0 - 0x0
    "00010001", -- 7634 - 0x1dd2  :   17 - 0x11
    "00000000", -- 7635 - 0x1dd3  :    0 - 0x0
    "00000000", -- 7636 - 0x1dd4  :    0 - 0x0
    "10000000", -- 7637 - 0x1dd5  :  128 - 0x80
    "00000000", -- 7638 - 0x1dd6  :    0 - 0x0
    "00000000", -- 7639 - 0x1dd7  :    0 - 0x0
    "00000000", -- 7640 - 0x1dd8  :    0 - 0x0
    "01000000", -- 7641 - 0x1dd9  :   64 - 0x40
    "00000000", -- 7642 - 0x1dda  :    0 - 0x0
    "00000000", -- 7643 - 0x1ddb  :    0 - 0x0
    "00000000", -- 7644 - 0x1ddc  :    0 - 0x0
    "00000000", -- 7645 - 0x1ddd  :    0 - 0x0
    "00000010", -- 7646 - 0x1dde  :    2 - 0x2
    "00100000", -- 7647 - 0x1ddf  :   32 - 0x20
    "10110011", -- 7648 - 0x1de0  :  179 - 0xb3 -- Background 0xde
    "10110011", -- 7649 - 0x1de1  :  179 - 0xb3
    "10110011", -- 7650 - 0x1de2  :  179 - 0xb3
    "10110011", -- 7651 - 0x1de3  :  179 - 0xb3
    "10110000", -- 7652 - 0x1de4  :  176 - 0xb0
    "10101111", -- 7653 - 0x1de5  :  175 - 0xaf
    "10011111", -- 7654 - 0x1de6  :  159 - 0x9f
    "11000000", -- 7655 - 0x1de7  :  192 - 0xc0
    "00111110", -- 7656 - 0x1de8  :   62 - 0x3e
    "00111111", -- 7657 - 0x1de9  :   63 - 0x3f
    "00111110", -- 7658 - 0x1dea  :   62 - 0x3e
    "00111100", -- 7659 - 0x1deb  :   60 - 0x3c
    "00111111", -- 7660 - 0x1dec  :   63 - 0x3f
    "00110000", -- 7661 - 0x1ded  :   48 - 0x30
    "00000000", -- 7662 - 0x1dee  :    0 - 0x0
    "00000000", -- 7663 - 0x1def  :    0 - 0x0
    "11101101", -- 7664 - 0x1df0  :  237 - 0xed -- Background 0xdf
    "11001101", -- 7665 - 0x1df1  :  205 - 0xcd
    "11001101", -- 7666 - 0x1df2  :  205 - 0xcd
    "00001101", -- 7667 - 0x1df3  :   13 - 0xd
    "00001101", -- 7668 - 0x1df4  :   13 - 0xd
    "11111101", -- 7669 - 0x1df5  :  253 - 0xfd
    "11111101", -- 7670 - 0x1df6  :  253 - 0xfd
    "00000011", -- 7671 - 0x1df7  :    3 - 0x3
    "00010000", -- 7672 - 0x1df8  :   16 - 0x10
    "10110000", -- 7673 - 0x1df9  :  176 - 0xb0
    "00110000", -- 7674 - 0x1dfa  :   48 - 0x30
    "11110000", -- 7675 - 0x1dfb  :  240 - 0xf0
    "11110000", -- 7676 - 0x1dfc  :  240 - 0xf0
    "00000000", -- 7677 - 0x1dfd  :    0 - 0x0
    "00000000", -- 7678 - 0x1dfe  :    0 - 0x0
    "00000000", -- 7679 - 0x1dff  :    0 - 0x0
    "11101110", -- 7680 - 0x1e00  :  238 - 0xee -- Background 0xe0
    "11101110", -- 7681 - 0x1e01  :  238 - 0xee
    "11101110", -- 7682 - 0x1e02  :  238 - 0xee
    "11101110", -- 7683 - 0x1e03  :  238 - 0xee
    "11111110", -- 7684 - 0x1e04  :  254 - 0xfe
    "11111100", -- 7685 - 0x1e05  :  252 - 0xfc
    "11000001", -- 7686 - 0x1e06  :  193 - 0xc1
    "11111111", -- 7687 - 0x1e07  :  255 - 0xff
    "11101110", -- 7688 - 0x1e08  :  238 - 0xee
    "11101110", -- 7689 - 0x1e09  :  238 - 0xee
    "11101110", -- 7690 - 0x1e0a  :  238 - 0xee
    "11101110", -- 7691 - 0x1e0b  :  238 - 0xee
    "11111110", -- 7692 - 0x1e0c  :  254 - 0xfe
    "01111100", -- 7693 - 0x1e0d  :  124 - 0x7c
    "00000000", -- 7694 - 0x1e0e  :    0 - 0x0
    "00000000", -- 7695 - 0x1e0f  :    0 - 0x0
    "11111011", -- 7696 - 0x1e10  :  251 - 0xfb -- Background 0xe1
    "11111011", -- 7697 - 0x1e11  :  251 - 0xfb
    "11111011", -- 7698 - 0x1e12  :  251 - 0xfb
    "11111011", -- 7699 - 0x1e13  :  251 - 0xfb
    "11111111", -- 7700 - 0x1e14  :  255 - 0xff
    "11111101", -- 7701 - 0x1e15  :  253 - 0xfd
    "11000001", -- 7702 - 0x1e16  :  193 - 0xc1
    "11111111", -- 7703 - 0x1e17  :  255 - 0xff
    "00111000", -- 7704 - 0x1e18  :   56 - 0x38
    "00111000", -- 7705 - 0x1e19  :   56 - 0x38
    "00111000", -- 7706 - 0x1e1a  :   56 - 0x38
    "00111000", -- 7707 - 0x1e1b  :   56 - 0x38
    "01111100", -- 7708 - 0x1e1c  :  124 - 0x7c
    "01111100", -- 7709 - 0x1e1d  :  124 - 0x7c
    "00000000", -- 7710 - 0x1e1e  :    0 - 0x0
    "00000000", -- 7711 - 0x1e1f  :    0 - 0x0
    "11111100", -- 7712 - 0x1e20  :  252 - 0xfc -- Background 0xe2
    "11100001", -- 7713 - 0x1e21  :  225 - 0xe1
    "11101111", -- 7714 - 0x1e22  :  239 - 0xef
    "11101111", -- 7715 - 0x1e23  :  239 - 0xef
    "11111111", -- 7716 - 0x1e24  :  255 - 0xff
    "11111110", -- 7717 - 0x1e25  :  254 - 0xfe
    "10000000", -- 7718 - 0x1e26  :  128 - 0x80
    "11111111", -- 7719 - 0x1e27  :  255 - 0xff
    "11111100", -- 7720 - 0x1e28  :  252 - 0xfc
    "11100000", -- 7721 - 0x1e29  :  224 - 0xe0
    "11100000", -- 7722 - 0x1e2a  :  224 - 0xe0
    "11100000", -- 7723 - 0x1e2b  :  224 - 0xe0
    "11111110", -- 7724 - 0x1e2c  :  254 - 0xfe
    "11111110", -- 7725 - 0x1e2d  :  254 - 0xfe
    "00000000", -- 7726 - 0x1e2e  :    0 - 0x0
    "00000000", -- 7727 - 0x1e2f  :    0 - 0x0
    "11101110", -- 7728 - 0x1e30  :  238 - 0xee -- Background 0xe3
    "11111110", -- 7729 - 0x1e31  :  254 - 0xfe
    "11111110", -- 7730 - 0x1e32  :  254 - 0xfe
    "11111110", -- 7731 - 0x1e33  :  254 - 0xfe
    "11111110", -- 7732 - 0x1e34  :  254 - 0xfe
    "11111100", -- 7733 - 0x1e35  :  252 - 0xfc
    "11000001", -- 7734 - 0x1e36  :  193 - 0xc1
    "11111111", -- 7735 - 0x1e37  :  255 - 0xff
    "00001110", -- 7736 - 0x1e38  :   14 - 0xe
    "00001110", -- 7737 - 0x1e39  :   14 - 0xe
    "00001110", -- 7738 - 0x1e3a  :   14 - 0xe
    "11101110", -- 7739 - 0x1e3b  :  238 - 0xee
    "11111110", -- 7740 - 0x1e3c  :  254 - 0xfe
    "01111100", -- 7741 - 0x1e3d  :  124 - 0x7c
    "00000000", -- 7742 - 0x1e3e  :    0 - 0x0
    "00000000", -- 7743 - 0x1e3f  :    0 - 0x0
    "11101110", -- 7744 - 0x1e40  :  238 - 0xee -- Background 0xe4
    "11101110", -- 7745 - 0x1e41  :  238 - 0xee
    "11111110", -- 7746 - 0x1e42  :  254 - 0xfe
    "11111110", -- 7747 - 0x1e43  :  254 - 0xfe
    "10001110", -- 7748 - 0x1e44  :  142 - 0x8e
    "11111110", -- 7749 - 0x1e45  :  254 - 0xfe
    "11111000", -- 7750 - 0x1e46  :  248 - 0xf8
    "11111111", -- 7751 - 0x1e47  :  255 - 0xff
    "11101110", -- 7752 - 0x1e48  :  238 - 0xee
    "11101110", -- 7753 - 0x1e49  :  238 - 0xee
    "11111110", -- 7754 - 0x1e4a  :  254 - 0xfe
    "11111110", -- 7755 - 0x1e4b  :  254 - 0xfe
    "00001110", -- 7756 - 0x1e4c  :   14 - 0xe
    "00001110", -- 7757 - 0x1e4d  :   14 - 0xe
    "00000000", -- 7758 - 0x1e4e  :    0 - 0x0
    "00000000", -- 7759 - 0x1e4f  :    0 - 0x0
    "10001110", -- 7760 - 0x1e50  :  142 - 0x8e -- Background 0xe5
    "11111110", -- 7761 - 0x1e51  :  254 - 0xfe
    "11111110", -- 7762 - 0x1e52  :  254 - 0xfe
    "11111110", -- 7763 - 0x1e53  :  254 - 0xfe
    "11111110", -- 7764 - 0x1e54  :  254 - 0xfe
    "11111100", -- 7765 - 0x1e55  :  252 - 0xfc
    "11000001", -- 7766 - 0x1e56  :  193 - 0xc1
    "11111111", -- 7767 - 0x1e57  :  255 - 0xff
    "00001110", -- 7768 - 0x1e58  :   14 - 0xe
    "00001110", -- 7769 - 0x1e59  :   14 - 0xe
    "00001110", -- 7770 - 0x1e5a  :   14 - 0xe
    "11101110", -- 7771 - 0x1e5b  :  238 - 0xee
    "11111110", -- 7772 - 0x1e5c  :  254 - 0xfe
    "01111100", -- 7773 - 0x1e5d  :  124 - 0x7c
    "00000000", -- 7774 - 0x1e5e  :    0 - 0x0
    "00000000", -- 7775 - 0x1e5f  :    0 - 0x0
    "11101110", -- 7776 - 0x1e60  :  238 - 0xee -- Background 0xe6
    "11101110", -- 7777 - 0x1e61  :  238 - 0xee
    "11101110", -- 7778 - 0x1e62  :  238 - 0xee
    "11101110", -- 7779 - 0x1e63  :  238 - 0xee
    "11111110", -- 7780 - 0x1e64  :  254 - 0xfe
    "11111100", -- 7781 - 0x1e65  :  252 - 0xfc
    "11000001", -- 7782 - 0x1e66  :  193 - 0xc1
    "11111111", -- 7783 - 0x1e67  :  255 - 0xff
    "11101110", -- 7784 - 0x1e68  :  238 - 0xee
    "11101110", -- 7785 - 0x1e69  :  238 - 0xee
    "11101110", -- 7786 - 0x1e6a  :  238 - 0xee
    "11101110", -- 7787 - 0x1e6b  :  238 - 0xee
    "11111110", -- 7788 - 0x1e6c  :  254 - 0xfe
    "01111100", -- 7789 - 0x1e6d  :  124 - 0x7c
    "00000000", -- 7790 - 0x1e6e  :    0 - 0x0
    "00000000", -- 7791 - 0x1e6f  :    0 - 0x0
    "11111101", -- 7792 - 0x1e70  :  253 - 0xfd -- Background 0xe7
    "11111101", -- 7793 - 0x1e71  :  253 - 0xfd
    "11111001", -- 7794 - 0x1e72  :  249 - 0xf9
    "11111011", -- 7795 - 0x1e73  :  251 - 0xfb
    "11111011", -- 7796 - 0x1e74  :  251 - 0xfb
    "11111011", -- 7797 - 0x1e75  :  251 - 0xfb
    "11100011", -- 7798 - 0x1e76  :  227 - 0xe3
    "11111111", -- 7799 - 0x1e77  :  255 - 0xff
    "00011100", -- 7800 - 0x1e78  :   28 - 0x1c
    "00011100", -- 7801 - 0x1e79  :   28 - 0x1c
    "00111000", -- 7802 - 0x1e7a  :   56 - 0x38
    "00111000", -- 7803 - 0x1e7b  :   56 - 0x38
    "00111000", -- 7804 - 0x1e7c  :   56 - 0x38
    "00111000", -- 7805 - 0x1e7d  :   56 - 0x38
    "00000000", -- 7806 - 0x1e7e  :    0 - 0x0
    "00000000", -- 7807 - 0x1e7f  :    0 - 0x0
    "11101110", -- 7808 - 0x1e80  :  238 - 0xee -- Background 0xe8
    "11101110", -- 7809 - 0x1e81  :  238 - 0xee
    "11101110", -- 7810 - 0x1e82  :  238 - 0xee
    "11101110", -- 7811 - 0x1e83  :  238 - 0xee
    "11111110", -- 7812 - 0x1e84  :  254 - 0xfe
    "11111100", -- 7813 - 0x1e85  :  252 - 0xfc
    "11000001", -- 7814 - 0x1e86  :  193 - 0xc1
    "11111111", -- 7815 - 0x1e87  :  255 - 0xff
    "11101110", -- 7816 - 0x1e88  :  238 - 0xee
    "11101110", -- 7817 - 0x1e89  :  238 - 0xee
    "11101110", -- 7818 - 0x1e8a  :  238 - 0xee
    "11101110", -- 7819 - 0x1e8b  :  238 - 0xee
    "11111110", -- 7820 - 0x1e8c  :  254 - 0xfe
    "01111100", -- 7821 - 0x1e8d  :  124 - 0x7c
    "00000000", -- 7822 - 0x1e8e  :    0 - 0x0
    "00000000", -- 7823 - 0x1e8f  :    0 - 0x0
    "11111110", -- 7824 - 0x1e90  :  254 - 0xfe -- Background 0xe9
    "11111110", -- 7825 - 0x1e91  :  254 - 0xfe
    "11001110", -- 7826 - 0x1e92  :  206 - 0xce
    "11111110", -- 7827 - 0x1e93  :  254 - 0xfe
    "11111110", -- 7828 - 0x1e94  :  254 - 0xfe
    "11111100", -- 7829 - 0x1e95  :  252 - 0xfc
    "11000001", -- 7830 - 0x1e96  :  193 - 0xc1
    "11111111", -- 7831 - 0x1e97  :  255 - 0xff
    "11111110", -- 7832 - 0x1e98  :  254 - 0xfe
    "01111110", -- 7833 - 0x1e99  :  126 - 0x7e
    "00001110", -- 7834 - 0x1e9a  :   14 - 0xe
    "00001110", -- 7835 - 0x1e9b  :   14 - 0xe
    "01111110", -- 7836 - 0x1e9c  :  126 - 0x7e
    "01111100", -- 7837 - 0x1e9d  :  124 - 0x7c
    "00000000", -- 7838 - 0x1e9e  :    0 - 0x0
    "00000000", -- 7839 - 0x1e9f  :    0 - 0x0
    "00000000", -- 7840 - 0x1ea0  :    0 - 0x0 -- Background 0xea
    "01110000", -- 7841 - 0x1ea1  :  112 - 0x70
    "00111000", -- 7842 - 0x1ea2  :   56 - 0x38
    "00000000", -- 7843 - 0x1ea3  :    0 - 0x0
    "00000010", -- 7844 - 0x1ea4  :    2 - 0x2
    "00000111", -- 7845 - 0x1ea5  :    7 - 0x7
    "00000011", -- 7846 - 0x1ea6  :    3 - 0x3
    "00000000", -- 7847 - 0x1ea7  :    0 - 0x0
    "00000000", -- 7848 - 0x1ea8  :    0 - 0x0
    "01110000", -- 7849 - 0x1ea9  :  112 - 0x70
    "00111000", -- 7850 - 0x1eaa  :   56 - 0x38
    "00000000", -- 7851 - 0x1eab  :    0 - 0x0
    "00000010", -- 7852 - 0x1eac  :    2 - 0x2
    "00000111", -- 7853 - 0x1ead  :    7 - 0x7
    "00000011", -- 7854 - 0x1eae  :    3 - 0x3
    "00000000", -- 7855 - 0x1eaf  :    0 - 0x0
    "00000000", -- 7856 - 0x1eb0  :    0 - 0x0 -- Background 0xeb
    "00001100", -- 7857 - 0x1eb1  :   12 - 0xc
    "00000110", -- 7858 - 0x1eb2  :    6 - 0x6
    "00000110", -- 7859 - 0x1eb3  :    6 - 0x6
    "01100000", -- 7860 - 0x1eb4  :   96 - 0x60
    "01110000", -- 7861 - 0x1eb5  :  112 - 0x70
    "00110000", -- 7862 - 0x1eb6  :   48 - 0x30
    "00000000", -- 7863 - 0x1eb7  :    0 - 0x0
    "00000000", -- 7864 - 0x1eb8  :    0 - 0x0
    "00001100", -- 7865 - 0x1eb9  :   12 - 0xc
    "00000110", -- 7866 - 0x1eba  :    6 - 0x6
    "00000110", -- 7867 - 0x1ebb  :    6 - 0x6
    "01100000", -- 7868 - 0x1ebc  :   96 - 0x60
    "01110000", -- 7869 - 0x1ebd  :  112 - 0x70
    "00110000", -- 7870 - 0x1ebe  :   48 - 0x30
    "00000000", -- 7871 - 0x1ebf  :    0 - 0x0
    "00000000", -- 7872 - 0x1ec0  :    0 - 0x0 -- Background 0xec
    "11000000", -- 7873 - 0x1ec1  :  192 - 0xc0
    "11100000", -- 7874 - 0x1ec2  :  224 - 0xe0
    "01100000", -- 7875 - 0x1ec3  :   96 - 0x60
    "00000000", -- 7876 - 0x1ec4  :    0 - 0x0
    "00001100", -- 7877 - 0x1ec5  :   12 - 0xc
    "00001110", -- 7878 - 0x1ec6  :   14 - 0xe
    "00000110", -- 7879 - 0x1ec7  :    6 - 0x6
    "00000000", -- 7880 - 0x1ec8  :    0 - 0x0
    "11000000", -- 7881 - 0x1ec9  :  192 - 0xc0
    "11100000", -- 7882 - 0x1eca  :  224 - 0xe0
    "01100000", -- 7883 - 0x1ecb  :   96 - 0x60
    "00000000", -- 7884 - 0x1ecc  :    0 - 0x0
    "00001100", -- 7885 - 0x1ecd  :   12 - 0xc
    "00001110", -- 7886 - 0x1ece  :   14 - 0xe
    "00000110", -- 7887 - 0x1ecf  :    6 - 0x6
    "01100000", -- 7888 - 0x1ed0  :   96 - 0x60 -- Background 0xed
    "01110000", -- 7889 - 0x1ed1  :  112 - 0x70
    "00110000", -- 7890 - 0x1ed2  :   48 - 0x30
    "00000000", -- 7891 - 0x1ed3  :    0 - 0x0
    "00000000", -- 7892 - 0x1ed4  :    0 - 0x0
    "00001100", -- 7893 - 0x1ed5  :   12 - 0xc
    "00001110", -- 7894 - 0x1ed6  :   14 - 0xe
    "00000110", -- 7895 - 0x1ed7  :    6 - 0x6
    "01100000", -- 7896 - 0x1ed8  :   96 - 0x60
    "01110000", -- 7897 - 0x1ed9  :  112 - 0x70
    "00110000", -- 7898 - 0x1eda  :   48 - 0x30
    "00000000", -- 7899 - 0x1edb  :    0 - 0x0
    "00000000", -- 7900 - 0x1edc  :    0 - 0x0
    "00001100", -- 7901 - 0x1edd  :   12 - 0xc
    "00001110", -- 7902 - 0x1ede  :   14 - 0xe
    "00000110", -- 7903 - 0x1edf  :    6 - 0x6
    "11111111", -- 7904 - 0x1ee0  :  255 - 0xff -- Background 0xee
    "11111111", -- 7905 - 0x1ee1  :  255 - 0xff
    "10111101", -- 7906 - 0x1ee2  :  189 - 0xbd
    "11111111", -- 7907 - 0x1ee3  :  255 - 0xff
    "11111111", -- 7908 - 0x1ee4  :  255 - 0xff
    "11111011", -- 7909 - 0x1ee5  :  251 - 0xfb
    "11111111", -- 7910 - 0x1ee6  :  255 - 0xff
    "11111111", -- 7911 - 0x1ee7  :  255 - 0xff
    "00000000", -- 7912 - 0x1ee8  :    0 - 0x0
    "00000000", -- 7913 - 0x1ee9  :    0 - 0x0
    "01000010", -- 7914 - 0x1eea  :   66 - 0x42
    "00000000", -- 7915 - 0x1eeb  :    0 - 0x0
    "00000000", -- 7916 - 0x1eec  :    0 - 0x0
    "00000100", -- 7917 - 0x1eed  :    4 - 0x4
    "00000000", -- 7918 - 0x1eee  :    0 - 0x0
    "00000000", -- 7919 - 0x1eef  :    0 - 0x0
    "11111111", -- 7920 - 0x1ef0  :  255 - 0xff -- Background 0xef
    "11111111", -- 7921 - 0x1ef1  :  255 - 0xff
    "11111011", -- 7922 - 0x1ef2  :  251 - 0xfb
    "11111111", -- 7923 - 0x1ef3  :  255 - 0xff
    "11011111", -- 7924 - 0x1ef4  :  223 - 0xdf
    "11111111", -- 7925 - 0x1ef5  :  255 - 0xff
    "11111111", -- 7926 - 0x1ef6  :  255 - 0xff
    "11111111", -- 7927 - 0x1ef7  :  255 - 0xff
    "00000000", -- 7928 - 0x1ef8  :    0 - 0x0
    "00000000", -- 7929 - 0x1ef9  :    0 - 0x0
    "00000100", -- 7930 - 0x1efa  :    4 - 0x4
    "00000000", -- 7931 - 0x1efb  :    0 - 0x0
    "00100000", -- 7932 - 0x1efc  :   32 - 0x20
    "00000000", -- 7933 - 0x1efd  :    0 - 0x0
    "00000000", -- 7934 - 0x1efe  :    0 - 0x0
    "00000000", -- 7935 - 0x1eff  :    0 - 0x0
    "00000000", -- 7936 - 0x1f00  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 7937 - 0x1f01  :    0 - 0x0
    "00000000", -- 7938 - 0x1f02  :    0 - 0x0
    "00000000", -- 7939 - 0x1f03  :    0 - 0x0
    "00000000", -- 7940 - 0x1f04  :    0 - 0x0
    "00000000", -- 7941 - 0x1f05  :    0 - 0x0
    "00000000", -- 7942 - 0x1f06  :    0 - 0x0
    "00000000", -- 7943 - 0x1f07  :    0 - 0x0
    "00000000", -- 7944 - 0x1f08  :    0 - 0x0
    "00000000", -- 7945 - 0x1f09  :    0 - 0x0
    "00000000", -- 7946 - 0x1f0a  :    0 - 0x0
    "00000000", -- 7947 - 0x1f0b  :    0 - 0x0
    "00000000", -- 7948 - 0x1f0c  :    0 - 0x0
    "00000000", -- 7949 - 0x1f0d  :    0 - 0x0
    "00000000", -- 7950 - 0x1f0e  :    0 - 0x0
    "00000000", -- 7951 - 0x1f0f  :    0 - 0x0
    "00000000", -- 7952 - 0x1f10  :    0 - 0x0 -- Background 0xf1
    "10000000", -- 7953 - 0x1f11  :  128 - 0x80
    "00000000", -- 7954 - 0x1f12  :    0 - 0x0
    "00000000", -- 7955 - 0x1f13  :    0 - 0x0
    "00000000", -- 7956 - 0x1f14  :    0 - 0x0
    "00000000", -- 7957 - 0x1f15  :    0 - 0x0
    "00000000", -- 7958 - 0x1f16  :    0 - 0x0
    "00000000", -- 7959 - 0x1f17  :    0 - 0x0
    "10000000", -- 7960 - 0x1f18  :  128 - 0x80
    "10000000", -- 7961 - 0x1f19  :  128 - 0x80
    "10000000", -- 7962 - 0x1f1a  :  128 - 0x80
    "10000000", -- 7963 - 0x1f1b  :  128 - 0x80
    "00000000", -- 7964 - 0x1f1c  :    0 - 0x0
    "00000000", -- 7965 - 0x1f1d  :    0 - 0x0
    "00000000", -- 7966 - 0x1f1e  :    0 - 0x0
    "00000000", -- 7967 - 0x1f1f  :    0 - 0x0
    "00000000", -- 7968 - 0x1f20  :    0 - 0x0 -- Background 0xf2
    "11000000", -- 7969 - 0x1f21  :  192 - 0xc0
    "00000000", -- 7970 - 0x1f22  :    0 - 0x0
    "00000000", -- 7971 - 0x1f23  :    0 - 0x0
    "00000000", -- 7972 - 0x1f24  :    0 - 0x0
    "00000000", -- 7973 - 0x1f25  :    0 - 0x0
    "00000000", -- 7974 - 0x1f26  :    0 - 0x0
    "00000000", -- 7975 - 0x1f27  :    0 - 0x0
    "11000000", -- 7976 - 0x1f28  :  192 - 0xc0
    "11000000", -- 7977 - 0x1f29  :  192 - 0xc0
    "11000000", -- 7978 - 0x1f2a  :  192 - 0xc0
    "11000000", -- 7979 - 0x1f2b  :  192 - 0xc0
    "00000000", -- 7980 - 0x1f2c  :    0 - 0x0
    "00000000", -- 7981 - 0x1f2d  :    0 - 0x0
    "00000000", -- 7982 - 0x1f2e  :    0 - 0x0
    "00000000", -- 7983 - 0x1f2f  :    0 - 0x0
    "00000000", -- 7984 - 0x1f30  :    0 - 0x0 -- Background 0xf3
    "11100000", -- 7985 - 0x1f31  :  224 - 0xe0
    "00000000", -- 7986 - 0x1f32  :    0 - 0x0
    "00000000", -- 7987 - 0x1f33  :    0 - 0x0
    "00000000", -- 7988 - 0x1f34  :    0 - 0x0
    "00000000", -- 7989 - 0x1f35  :    0 - 0x0
    "00000000", -- 7990 - 0x1f36  :    0 - 0x0
    "00000000", -- 7991 - 0x1f37  :    0 - 0x0
    "11100000", -- 7992 - 0x1f38  :  224 - 0xe0
    "11100000", -- 7993 - 0x1f39  :  224 - 0xe0
    "11100000", -- 7994 - 0x1f3a  :  224 - 0xe0
    "11100000", -- 7995 - 0x1f3b  :  224 - 0xe0
    "00000000", -- 7996 - 0x1f3c  :    0 - 0x0
    "00000000", -- 7997 - 0x1f3d  :    0 - 0x0
    "00000000", -- 7998 - 0x1f3e  :    0 - 0x0
    "00000000", -- 7999 - 0x1f3f  :    0 - 0x0
    "00000000", -- 8000 - 0x1f40  :    0 - 0x0 -- Background 0xf4
    "11110000", -- 8001 - 0x1f41  :  240 - 0xf0
    "00000000", -- 8002 - 0x1f42  :    0 - 0x0
    "00000000", -- 8003 - 0x1f43  :    0 - 0x0
    "00000000", -- 8004 - 0x1f44  :    0 - 0x0
    "00000000", -- 8005 - 0x1f45  :    0 - 0x0
    "00000000", -- 8006 - 0x1f46  :    0 - 0x0
    "00000000", -- 8007 - 0x1f47  :    0 - 0x0
    "11110000", -- 8008 - 0x1f48  :  240 - 0xf0
    "11110000", -- 8009 - 0x1f49  :  240 - 0xf0
    "11110000", -- 8010 - 0x1f4a  :  240 - 0xf0
    "11110000", -- 8011 - 0x1f4b  :  240 - 0xf0
    "00000000", -- 8012 - 0x1f4c  :    0 - 0x0
    "00000000", -- 8013 - 0x1f4d  :    0 - 0x0
    "00000000", -- 8014 - 0x1f4e  :    0 - 0x0
    "00000000", -- 8015 - 0x1f4f  :    0 - 0x0
    "00000000", -- 8016 - 0x1f50  :    0 - 0x0 -- Background 0xf5
    "11111000", -- 8017 - 0x1f51  :  248 - 0xf8
    "00000000", -- 8018 - 0x1f52  :    0 - 0x0
    "00000000", -- 8019 - 0x1f53  :    0 - 0x0
    "00000000", -- 8020 - 0x1f54  :    0 - 0x0
    "00000000", -- 8021 - 0x1f55  :    0 - 0x0
    "00000000", -- 8022 - 0x1f56  :    0 - 0x0
    "00000000", -- 8023 - 0x1f57  :    0 - 0x0
    "11111000", -- 8024 - 0x1f58  :  248 - 0xf8
    "11111000", -- 8025 - 0x1f59  :  248 - 0xf8
    "11111000", -- 8026 - 0x1f5a  :  248 - 0xf8
    "11111000", -- 8027 - 0x1f5b  :  248 - 0xf8
    "00000000", -- 8028 - 0x1f5c  :    0 - 0x0
    "00000000", -- 8029 - 0x1f5d  :    0 - 0x0
    "00000000", -- 8030 - 0x1f5e  :    0 - 0x0
    "00000000", -- 8031 - 0x1f5f  :    0 - 0x0
    "00000000", -- 8032 - 0x1f60  :    0 - 0x0 -- Background 0xf6
    "11111100", -- 8033 - 0x1f61  :  252 - 0xfc
    "00000000", -- 8034 - 0x1f62  :    0 - 0x0
    "00000000", -- 8035 - 0x1f63  :    0 - 0x0
    "00000000", -- 8036 - 0x1f64  :    0 - 0x0
    "00000000", -- 8037 - 0x1f65  :    0 - 0x0
    "00000000", -- 8038 - 0x1f66  :    0 - 0x0
    "00000000", -- 8039 - 0x1f67  :    0 - 0x0
    "11111100", -- 8040 - 0x1f68  :  252 - 0xfc
    "11111100", -- 8041 - 0x1f69  :  252 - 0xfc
    "11111100", -- 8042 - 0x1f6a  :  252 - 0xfc
    "11111100", -- 8043 - 0x1f6b  :  252 - 0xfc
    "00000000", -- 8044 - 0x1f6c  :    0 - 0x0
    "00000000", -- 8045 - 0x1f6d  :    0 - 0x0
    "00000000", -- 8046 - 0x1f6e  :    0 - 0x0
    "00000000", -- 8047 - 0x1f6f  :    0 - 0x0
    "00000000", -- 8048 - 0x1f70  :    0 - 0x0 -- Background 0xf7
    "11111110", -- 8049 - 0x1f71  :  254 - 0xfe
    "00000000", -- 8050 - 0x1f72  :    0 - 0x0
    "00000000", -- 8051 - 0x1f73  :    0 - 0x0
    "00000000", -- 8052 - 0x1f74  :    0 - 0x0
    "00000000", -- 8053 - 0x1f75  :    0 - 0x0
    "00000000", -- 8054 - 0x1f76  :    0 - 0x0
    "00000000", -- 8055 - 0x1f77  :    0 - 0x0
    "11111110", -- 8056 - 0x1f78  :  254 - 0xfe
    "11111110", -- 8057 - 0x1f79  :  254 - 0xfe
    "11111110", -- 8058 - 0x1f7a  :  254 - 0xfe
    "11111110", -- 8059 - 0x1f7b  :  254 - 0xfe
    "00000000", -- 8060 - 0x1f7c  :    0 - 0x0
    "00000000", -- 8061 - 0x1f7d  :    0 - 0x0
    "00000000", -- 8062 - 0x1f7e  :    0 - 0x0
    "00000000", -- 8063 - 0x1f7f  :    0 - 0x0
    "00000000", -- 8064 - 0x1f80  :    0 - 0x0 -- Background 0xf8
    "11111111", -- 8065 - 0x1f81  :  255 - 0xff
    "00000000", -- 8066 - 0x1f82  :    0 - 0x0
    "00000000", -- 8067 - 0x1f83  :    0 - 0x0
    "00000000", -- 8068 - 0x1f84  :    0 - 0x0
    "00000000", -- 8069 - 0x1f85  :    0 - 0x0
    "00000000", -- 8070 - 0x1f86  :    0 - 0x0
    "00000000", -- 8071 - 0x1f87  :    0 - 0x0
    "11111111", -- 8072 - 0x1f88  :  255 - 0xff
    "11111111", -- 8073 - 0x1f89  :  255 - 0xff
    "11111111", -- 8074 - 0x1f8a  :  255 - 0xff
    "11111111", -- 8075 - 0x1f8b  :  255 - 0xff
    "00000000", -- 8076 - 0x1f8c  :    0 - 0x0
    "00000000", -- 8077 - 0x1f8d  :    0 - 0x0
    "00000000", -- 8078 - 0x1f8e  :    0 - 0x0
    "00000000", -- 8079 - 0x1f8f  :    0 - 0x0
    "11111111", -- 8080 - 0x1f90  :  255 - 0xff -- Background 0xf9
    "11111111", -- 8081 - 0x1f91  :  255 - 0xff
    "11111111", -- 8082 - 0x1f92  :  255 - 0xff
    "11111111", -- 8083 - 0x1f93  :  255 - 0xff
    "10000000", -- 8084 - 0x1f94  :  128 - 0x80
    "10000000", -- 8085 - 0x1f95  :  128 - 0x80
    "11000000", -- 8086 - 0x1f96  :  192 - 0xc0
    "11000000", -- 8087 - 0x1f97  :  192 - 0xc0
    "00000000", -- 8088 - 0x1f98  :    0 - 0x0
    "00000000", -- 8089 - 0x1f99  :    0 - 0x0
    "00000000", -- 8090 - 0x1f9a  :    0 - 0x0
    "00000000", -- 8091 - 0x1f9b  :    0 - 0x0
    "01111111", -- 8092 - 0x1f9c  :  127 - 0x7f
    "01000000", -- 8093 - 0x1f9d  :   64 - 0x40
    "01000000", -- 8094 - 0x1f9e  :   64 - 0x40
    "01000000", -- 8095 - 0x1f9f  :   64 - 0x40
    "11111111", -- 8096 - 0x1fa0  :  255 - 0xff -- Background 0xfa
    "11111111", -- 8097 - 0x1fa1  :  255 - 0xff
    "11111111", -- 8098 - 0x1fa2  :  255 - 0xff
    "11111111", -- 8099 - 0x1fa3  :  255 - 0xff
    "00000000", -- 8100 - 0x1fa4  :    0 - 0x0
    "00000000", -- 8101 - 0x1fa5  :    0 - 0x0
    "00000000", -- 8102 - 0x1fa6  :    0 - 0x0
    "00000000", -- 8103 - 0x1fa7  :    0 - 0x0
    "00000000", -- 8104 - 0x1fa8  :    0 - 0x0
    "00000000", -- 8105 - 0x1fa9  :    0 - 0x0
    "00000000", -- 8106 - 0x1faa  :    0 - 0x0
    "00000000", -- 8107 - 0x1fab  :    0 - 0x0
    "11111111", -- 8108 - 0x1fac  :  255 - 0xff
    "00000000", -- 8109 - 0x1fad  :    0 - 0x0
    "00000000", -- 8110 - 0x1fae  :    0 - 0x0
    "00000000", -- 8111 - 0x1faf  :    0 - 0x0
    "11111111", -- 8112 - 0x1fb0  :  255 - 0xff -- Background 0xfb
    "11111111", -- 8113 - 0x1fb1  :  255 - 0xff
    "11111111", -- 8114 - 0x1fb2  :  255 - 0xff
    "11111111", -- 8115 - 0x1fb3  :  255 - 0xff
    "00000001", -- 8116 - 0x1fb4  :    1 - 0x1
    "00000000", -- 8117 - 0x1fb5  :    0 - 0x0
    "00000010", -- 8118 - 0x1fb6  :    2 - 0x2
    "00000010", -- 8119 - 0x1fb7  :    2 - 0x2
    "00000000", -- 8120 - 0x1fb8  :    0 - 0x0
    "00000000", -- 8121 - 0x1fb9  :    0 - 0x0
    "00000000", -- 8122 - 0x1fba  :    0 - 0x0
    "00000000", -- 8123 - 0x1fbb  :    0 - 0x0
    "11111110", -- 8124 - 0x1fbc  :  254 - 0xfe
    "00000010", -- 8125 - 0x1fbd  :    2 - 0x2
    "00000010", -- 8126 - 0x1fbe  :    2 - 0x2
    "00000010", -- 8127 - 0x1fbf  :    2 - 0x2
    "11000000", -- 8128 - 0x1fc0  :  192 - 0xc0 -- Background 0xfc
    "11000000", -- 8129 - 0x1fc1  :  192 - 0xc0
    "10000000", -- 8130 - 0x1fc2  :  128 - 0x80
    "10000000", -- 8131 - 0x1fc3  :  128 - 0x80
    "11000000", -- 8132 - 0x1fc4  :  192 - 0xc0
    "11111111", -- 8133 - 0x1fc5  :  255 - 0xff
    "11111111", -- 8134 - 0x1fc6  :  255 - 0xff
    "11111111", -- 8135 - 0x1fc7  :  255 - 0xff
    "01000000", -- 8136 - 0x1fc8  :   64 - 0x40
    "01000000", -- 8137 - 0x1fc9  :   64 - 0x40
    "01000000", -- 8138 - 0x1fca  :   64 - 0x40
    "01111111", -- 8139 - 0x1fcb  :  127 - 0x7f
    "00000000", -- 8140 - 0x1fcc  :    0 - 0x0
    "00000000", -- 8141 - 0x1fcd  :    0 - 0x0
    "00000000", -- 8142 - 0x1fce  :    0 - 0x0
    "00000000", -- 8143 - 0x1fcf  :    0 - 0x0
    "00000000", -- 8144 - 0x1fd0  :    0 - 0x0 -- Background 0xfd
    "00000000", -- 8145 - 0x1fd1  :    0 - 0x0
    "00000000", -- 8146 - 0x1fd2  :    0 - 0x0
    "00000000", -- 8147 - 0x1fd3  :    0 - 0x0
    "00000000", -- 8148 - 0x1fd4  :    0 - 0x0
    "11111111", -- 8149 - 0x1fd5  :  255 - 0xff
    "11111111", -- 8150 - 0x1fd6  :  255 - 0xff
    "11111111", -- 8151 - 0x1fd7  :  255 - 0xff
    "00000000", -- 8152 - 0x1fd8  :    0 - 0x0
    "00000000", -- 8153 - 0x1fd9  :    0 - 0x0
    "00000000", -- 8154 - 0x1fda  :    0 - 0x0
    "11111111", -- 8155 - 0x1fdb  :  255 - 0xff
    "00000000", -- 8156 - 0x1fdc  :    0 - 0x0
    "00000000", -- 8157 - 0x1fdd  :    0 - 0x0
    "00000000", -- 8158 - 0x1fde  :    0 - 0x0
    "00000000", -- 8159 - 0x1fdf  :    0 - 0x0
    "00000010", -- 8160 - 0x1fe0  :    2 - 0x2 -- Background 0xfe
    "00000010", -- 8161 - 0x1fe1  :    2 - 0x2
    "00000000", -- 8162 - 0x1fe2  :    0 - 0x0
    "00000000", -- 8163 - 0x1fe3  :    0 - 0x0
    "00000000", -- 8164 - 0x1fe4  :    0 - 0x0
    "11111111", -- 8165 - 0x1fe5  :  255 - 0xff
    "11111111", -- 8166 - 0x1fe6  :  255 - 0xff
    "11111111", -- 8167 - 0x1fe7  :  255 - 0xff
    "00000010", -- 8168 - 0x1fe8  :    2 - 0x2
    "00000010", -- 8169 - 0x1fe9  :    2 - 0x2
    "00000010", -- 8170 - 0x1fea  :    2 - 0x2
    "11111110", -- 8171 - 0x1feb  :  254 - 0xfe
    "00000000", -- 8172 - 0x1fec  :    0 - 0x0
    "00000000", -- 8173 - 0x1fed  :    0 - 0x0
    "00000000", -- 8174 - 0x1fee  :    0 - 0x0
    "00000000", -- 8175 - 0x1fef  :    0 - 0x0
    "11111111", -- 8176 - 0x1ff0  :  255 - 0xff -- Background 0xff
    "11111111", -- 8177 - 0x1ff1  :  255 - 0xff
    "11111111", -- 8178 - 0x1ff2  :  255 - 0xff
    "11111111", -- 8179 - 0x1ff3  :  255 - 0xff
    "11111111", -- 8180 - 0x1ff4  :  255 - 0xff
    "11111111", -- 8181 - 0x1ff5  :  255 - 0xff
    "11111111", -- 8182 - 0x1ff6  :  255 - 0xff
    "11111111", -- 8183 - 0x1ff7  :  255 - 0xff
    "00000000", -- 8184 - 0x1ff8  :    0 - 0x0
    "00000000", -- 8185 - 0x1ff9  :    0 - 0x0
    "00000000", -- 8186 - 0x1ffa  :    0 - 0x0
    "00000000", -- 8187 - 0x1ffb  :    0 - 0x0
    "00000000", -- 8188 - 0x1ffc  :    0 - 0x0
    "00000000", -- 8189 - 0x1ffd  :    0 - 0x0
    "00000000", -- 8190 - 0x1ffe  :    0 - 0x0
    "00000000"  -- 8191 - 0x1fff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
