--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables


---  Original memory dump file name: sprilo_ntable_00.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_SPRILO_00 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_SPRILO_00;

architecture BEHAVIORAL of ROM_NTABLE_SPRILO_00 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "11111010", --    0 -  0x0  :  250 - 0xfa
    "11111010", --    1 -  0x1  :  250 - 0xfa
    "11111010", --    2 -  0x2  :  250 - 0xfa
    "11101010", --    3 -  0x3  :  234 - 0xea
    "11111010", --    4 -  0x4  :  250 - 0xfa
    "11111010", --    5 -  0x5  :  250 - 0xfa
    "11111010", --    6 -  0x6  :  250 - 0xfa
    "11111010", --    7 -  0x7  :  250 - 0xfa
    "11111010", --    8 -  0x8  :  250 - 0xfa
    "11111010", --    9 -  0x9  :  250 - 0xfa
    "11111010", --   10 -  0xa  :  250 - 0xfa
    "11111010", --   11 -  0xb  :  250 - 0xfa
    "11111010", --   12 -  0xc  :  250 - 0xfa
    "11111010", --   13 -  0xd  :  250 - 0xfa
    "11101010", --   14 -  0xe  :  234 - 0xea
    "11111010", --   15 -  0xf  :  250 - 0xfa
    "11111010", --   16 - 0x10  :  250 - 0xfa
    "11111010", --   17 - 0x11  :  250 - 0xfa
    "11111010", --   18 - 0x12  :  250 - 0xfa
    "11111010", --   19 - 0x13  :  250 - 0xfa
    "11111010", --   20 - 0x14  :  250 - 0xfa
    "11111010", --   21 - 0x15  :  250 - 0xfa
    "11111010", --   22 - 0x16  :  250 - 0xfa
    "11111010", --   23 - 0x17  :  250 - 0xfa
    "11111010", --   24 - 0x18  :  250 - 0xfa
    "11111010", --   25 - 0x19  :  250 - 0xfa
    "11111010", --   26 - 0x1a  :  250 - 0xfa
    "11111010", --   27 - 0x1b  :  250 - 0xfa
    "11111010", --   28 - 0x1c  :  250 - 0xfa
    "11111010", --   29 - 0x1d  :  250 - 0xfa
    "11111010", --   30 - 0x1e  :  250 - 0xfa
    "11111010", --   31 - 0x1f  :  250 - 0xfa
    "11111010", --   32 - 0x20  :  250 - 0xfa
    "11100111", --   33 - 0x21  :  231 - 0xe7
    "11111011", --   34 - 0x22  :  251 - 0xfb
    "11111011", --   35 - 0x23  :  251 - 0xfb
    "11111011", --   36 - 0x24  :  251 - 0xfb
    "11111011", --   37 - 0x25  :  251 - 0xfb
    "11111011", --   38 - 0x26  :  251 - 0xfb
    "11111011", --   39 - 0x27  :  251 - 0xfb
    "11111011", --   40 - 0x28  :  251 - 0xfb
    "11111011", --   41 - 0x29  :  251 - 0xfb
    "11111011", --   42 - 0x2a  :  251 - 0xfb
    "11111011", --   43 - 0x2b  :  251 - 0xfb
    "11111011", --   44 - 0x2c  :  251 - 0xfb
    "11111011", --   45 - 0x2d  :  251 - 0xfb
    "11111011", --   46 - 0x2e  :  251 - 0xfb
    "11111011", --   47 - 0x2f  :  251 - 0xfb
    "11111011", --   48 - 0x30  :  251 - 0xfb
    "11111011", --   49 - 0x31  :  251 - 0xfb
    "11111011", --   50 - 0x32  :  251 - 0xfb
    "11111011", --   51 - 0x33  :  251 - 0xfb
    "11111011", --   52 - 0x34  :  251 - 0xfb
    "11111011", --   53 - 0x35  :  251 - 0xfb
    "11101000", --   54 - 0x36  :  232 - 0xe8
    "11111010", --   55 - 0x37  :  250 - 0xfa
    "11111010", --   56 - 0x38  :  250 - 0xfa
    "11101001", --   57 - 0x39  :  233 - 0xe9
    "11111001", --   58 - 0x3a  :  249 - 0xf9
    "11101001", --   59 - 0x3b  :  233 - 0xe9
    "11111010", --   60 - 0x3c  :  250 - 0xfa
    "11111010", --   61 - 0x3d  :  250 - 0xfa
    "11101001", --   62 - 0x3e  :  233 - 0xe9
    "11111010", --   63 - 0x3f  :  250 - 0xfa
    "11101010", --   64 - 0x40  :  234 - 0xea
    "11111100", --   65 - 0x41  :  252 - 0xfc
    "11111111", --   66 - 0x42  :  255 - 0xff
    "11111111", --   67 - 0x43  :  255 - 0xff
    "11111111", --   68 - 0x44  :  255 - 0xff
    "11111111", --   69 - 0x45  :  255 - 0xff
    "11111111", --   70 - 0x46  :  255 - 0xff
    "11111111", --   71 - 0x47  :  255 - 0xff
    "11111111", --   72 - 0x48  :  255 - 0xff
    "11111111", --   73 - 0x49  :  255 - 0xff
    "11111111", --   74 - 0x4a  :  255 - 0xff
    "11111111", --   75 - 0x4b  :  255 - 0xff
    "11111111", --   76 - 0x4c  :  255 - 0xff
    "11111111", --   77 - 0x4d  :  255 - 0xff
    "11111111", --   78 - 0x4e  :  255 - 0xff
    "11111111", --   79 - 0x4f  :  255 - 0xff
    "11111111", --   80 - 0x50  :  255 - 0xff
    "11111111", --   81 - 0x51  :  255 - 0xff
    "11111111", --   82 - 0x52  :  255 - 0xff
    "11111111", --   83 - 0x53  :  255 - 0xff
    "11111111", --   84 - 0x54  :  255 - 0xff
    "11111111", --   85 - 0x55  :  255 - 0xff
    "11101100", --   86 - 0x56  :  236 - 0xec
    "11111010", --   87 - 0x57  :  250 - 0xfa
    "11111010", --   88 - 0x58  :  250 - 0xfa
    "11111010", --   89 - 0x59  :  250 - 0xfa
    "11111010", --   90 - 0x5a  :  250 - 0xfa
    "11111010", --   91 - 0x5b  :  250 - 0xfa
    "11111010", --   92 - 0x5c  :  250 - 0xfa
    "11101001", --   93 - 0x5d  :  233 - 0xe9
    "11111010", --   94 - 0x5e  :  250 - 0xfa
    "11111010", --   95 - 0x5f  :  250 - 0xfa
    "11111010", --   96 - 0x60  :  250 - 0xfa
    "11111100", --   97 - 0x61  :  252 - 0xfc
    "11111111", --   98 - 0x62  :  255 - 0xff
    "11111111", --   99 - 0x63  :  255 - 0xff
    "11111111", --  100 - 0x64  :  255 - 0xff
    "11111111", --  101 - 0x65  :  255 - 0xff
    "11111101", --  102 - 0x66  :  253 - 0xfd
    "11111111", --  103 - 0x67  :  255 - 0xff
    "11111101", --  104 - 0x68  :  253 - 0xfd
    "11111111", --  105 - 0x69  :  255 - 0xff
    "11111101", --  106 - 0x6a  :  253 - 0xfd
    "11111111", --  107 - 0x6b  :  255 - 0xff
    "11111101", --  108 - 0x6c  :  253 - 0xfd
    "11111111", --  109 - 0x6d  :  255 - 0xff
    "11111101", --  110 - 0x6e  :  253 - 0xfd
    "11111111", --  111 - 0x6f  :  255 - 0xff
    "11111101", --  112 - 0x70  :  253 - 0xfd
    "11111111", --  113 - 0x71  :  255 - 0xff
    "11111101", --  114 - 0x72  :  253 - 0xfd
    "11111111", --  115 - 0x73  :  255 - 0xff
    "11111111", --  116 - 0x74  :  255 - 0xff
    "11111111", --  117 - 0x75  :  255 - 0xff
    "11101100", --  118 - 0x76  :  236 - 0xec
    "11111010", --  119 - 0x77  :  250 - 0xfa
    "11111010", --  120 - 0x78  :  250 - 0xfa
    "11111010", --  121 - 0x79  :  250 - 0xfa
    "11111010", --  122 - 0x7a  :  250 - 0xfa
    "11111010", --  123 - 0x7b  :  250 - 0xfa
    "11111010", --  124 - 0x7c  :  250 - 0xfa
    "11111010", --  125 - 0x7d  :  250 - 0xfa
    "11111010", --  126 - 0x7e  :  250 - 0xfa
    "11111010", --  127 - 0x7f  :  250 - 0xfa
    "11101001", --  128 - 0x80  :  233 - 0xe9
    "11111100", --  129 - 0x81  :  252 - 0xfc
    "11111111", --  130 - 0x82  :  255 - 0xff
    "11111111", --  131 - 0x83  :  255 - 0xff
    "11111111", --  132 - 0x84  :  255 - 0xff
    "11111111", --  133 - 0x85  :  255 - 0xff
    "11111101", --  134 - 0x86  :  253 - 0xfd
    "11111111", --  135 - 0x87  :  255 - 0xff
    "11111101", --  136 - 0x88  :  253 - 0xfd
    "11111111", --  137 - 0x89  :  255 - 0xff
    "11111101", --  138 - 0x8a  :  253 - 0xfd
    "11111111", --  139 - 0x8b  :  255 - 0xff
    "11111101", --  140 - 0x8c  :  253 - 0xfd
    "11111111", --  141 - 0x8d  :  255 - 0xff
    "11111101", --  142 - 0x8e  :  253 - 0xfd
    "11111111", --  143 - 0x8f  :  255 - 0xff
    "11111101", --  144 - 0x90  :  253 - 0xfd
    "11111111", --  145 - 0x91  :  255 - 0xff
    "11111101", --  146 - 0x92  :  253 - 0xfd
    "11111111", --  147 - 0x93  :  255 - 0xff
    "11111111", --  148 - 0x94  :  255 - 0xff
    "11111111", --  149 - 0x95  :  255 - 0xff
    "11101100", --  150 - 0x96  :  236 - 0xec
    "11101001", --  151 - 0x97  :  233 - 0xe9
    "11111010", --  152 - 0x98  :  250 - 0xfa
    "11111010", --  153 - 0x99  :  250 - 0xfa
    "11101010", --  154 - 0x9a  :  234 - 0xea
    "11111010", --  155 - 0x9b  :  250 - 0xfa
    "11111001", --  156 - 0x9c  :  249 - 0xf9
    "11111010", --  157 - 0x9d  :  250 - 0xfa
    "11111010", --  158 - 0x9e  :  250 - 0xfa
    "11111010", --  159 - 0x9f  :  250 - 0xfa
    "11111010", --  160 - 0xa0  :  250 - 0xfa
    "11111100", --  161 - 0xa1  :  252 - 0xfc
    "11111111", --  162 - 0xa2  :  255 - 0xff
    "11111111", --  163 - 0xa3  :  255 - 0xff
    "11111111", --  164 - 0xa4  :  255 - 0xff
    "11111111", --  165 - 0xa5  :  255 - 0xff
    "11111111", --  166 - 0xa6  :  255 - 0xff
    "11111111", --  167 - 0xa7  :  255 - 0xff
    "11111111", --  168 - 0xa8  :  255 - 0xff
    "11111111", --  169 - 0xa9  :  255 - 0xff
    "11111111", --  170 - 0xaa  :  255 - 0xff
    "11111111", --  171 - 0xab  :  255 - 0xff
    "11111111", --  172 - 0xac  :  255 - 0xff
    "11111111", --  173 - 0xad  :  255 - 0xff
    "11111111", --  174 - 0xae  :  255 - 0xff
    "11111111", --  175 - 0xaf  :  255 - 0xff
    "11111111", --  176 - 0xb0  :  255 - 0xff
    "11111111", --  177 - 0xb1  :  255 - 0xff
    "11111111", --  178 - 0xb2  :  255 - 0xff
    "11111111", --  179 - 0xb3  :  255 - 0xff
    "11111111", --  180 - 0xb4  :  255 - 0xff
    "11111111", --  181 - 0xb5  :  255 - 0xff
    "11110101", --  182 - 0xb6  :  245 - 0xf5
    "11111011", --  183 - 0xb7  :  251 - 0xfb
    "11111011", --  184 - 0xb8  :  251 - 0xfb
    "11111011", --  185 - 0xb9  :  251 - 0xfb
    "11111011", --  186 - 0xba  :  251 - 0xfb
    "11111011", --  187 - 0xbb  :  251 - 0xfb
    "11111011", --  188 - 0xbc  :  251 - 0xfb
    "11111011", --  189 - 0xbd  :  251 - 0xfb
    "11101000", --  190 - 0xbe  :  232 - 0xe8
    "11111010", --  191 - 0xbf  :  250 - 0xfa
    "11111010", --  192 - 0xc0  :  250 - 0xfa
    "11111100", --  193 - 0xc1  :  252 - 0xfc
    "11111111", --  194 - 0xc2  :  255 - 0xff
    "11111111", --  195 - 0xc3  :  255 - 0xff
    "11111111", --  196 - 0xc4  :  255 - 0xff
    "11111111", --  197 - 0xc5  :  255 - 0xff
    "11100101", --  198 - 0xc6  :  229 - 0xe5
    "11101011", --  199 - 0xc7  :  235 - 0xeb
    "11101011", --  200 - 0xc8  :  235 - 0xeb
    "11101011", --  201 - 0xc9  :  235 - 0xeb
    "11101011", --  202 - 0xca  :  235 - 0xeb
    "11101011", --  203 - 0xcb  :  235 - 0xeb
    "11101011", --  204 - 0xcc  :  235 - 0xeb
    "11101011", --  205 - 0xcd  :  235 - 0xeb
    "11101011", --  206 - 0xce  :  235 - 0xeb
    "11101011", --  207 - 0xcf  :  235 - 0xeb
    "11101011", --  208 - 0xd0  :  235 - 0xeb
    "11100110", --  209 - 0xd1  :  230 - 0xe6
    "11111111", --  210 - 0xd2  :  255 - 0xff
    "11111110", --  211 - 0xd3  :  254 - 0xfe
    "11111110", --  212 - 0xd4  :  254 - 0xfe
    "11111111", --  213 - 0xd5  :  255 - 0xff
    "11111111", --  214 - 0xd6  :  255 - 0xff
    "11111111", --  215 - 0xd7  :  255 - 0xff
    "11111111", --  216 - 0xd8  :  255 - 0xff
    "11111111", --  217 - 0xd9  :  255 - 0xff
    "11111111", --  218 - 0xda  :  255 - 0xff
    "11111111", --  219 - 0xdb  :  255 - 0xff
    "11111111", --  220 - 0xdc  :  255 - 0xff
    "11111111", --  221 - 0xdd  :  255 - 0xff
    "11101100", --  222 - 0xde  :  236 - 0xec
    "11111010", --  223 - 0xdf  :  250 - 0xfa
    "11111010", --  224 - 0xe0  :  250 - 0xfa
    "11111100", --  225 - 0xe1  :  252 - 0xfc
    "11111111", --  226 - 0xe2  :  255 - 0xff
    "11111110", --  227 - 0xe3  :  254 - 0xfe
    "11111110", --  228 - 0xe4  :  254 - 0xfe
    "11111111", --  229 - 0xe5  :  255 - 0xff
    "11101100", --  230 - 0xe6  :  236 - 0xec
    "11111010", --  231 - 0xe7  :  250 - 0xfa
    "11111010", --  232 - 0xe8  :  250 - 0xfa
    "11111001", --  233 - 0xe9  :  249 - 0xf9
    "11111010", --  234 - 0xea  :  250 - 0xfa
    "11111010", --  235 - 0xeb  :  250 - 0xfa
    "11111010", --  236 - 0xec  :  250 - 0xfa
    "11111010", --  237 - 0xed  :  250 - 0xfa
    "11111010", --  238 - 0xee  :  250 - 0xfa
    "11111010", --  239 - 0xef  :  250 - 0xfa
    "11111010", --  240 - 0xf0  :  250 - 0xfa
    "11111100", --  241 - 0xf1  :  252 - 0xfc
    "11111111", --  242 - 0xf2  :  255 - 0xff
    "11111111", --  243 - 0xf3  :  255 - 0xff
    "11111111", --  244 - 0xf4  :  255 - 0xff
    "11111111", --  245 - 0xf5  :  255 - 0xff
    "11111101", --  246 - 0xf6  :  253 - 0xfd
    "11111111", --  247 - 0xf7  :  255 - 0xff
    "11111101", --  248 - 0xf8  :  253 - 0xfd
    "11111111", --  249 - 0xf9  :  255 - 0xff
    "11111101", --  250 - 0xfa  :  253 - 0xfd
    "11111111", --  251 - 0xfb  :  255 - 0xff
    "11111111", --  252 - 0xfc  :  255 - 0xff
    "11111111", --  253 - 0xfd  :  255 - 0xff
    "11101100", --  254 - 0xfe  :  236 - 0xec
    "11111010", --  255 - 0xff  :  250 - 0xfa
    "11111010", --  256 - 0x100  :  250 - 0xfa
    "11111100", --  257 - 0x101  :  252 - 0xfc
    "11111111", --  258 - 0x102  :  255 - 0xff
    "11111111", --  259 - 0x103  :  255 - 0xff
    "11111111", --  260 - 0x104  :  255 - 0xff
    "11111111", --  261 - 0x105  :  255 - 0xff
    "11101100", --  262 - 0x106  :  236 - 0xec
    "11111010", --  263 - 0x107  :  250 - 0xfa
    "11111010", --  264 - 0x108  :  250 - 0xfa
    "11111010", --  265 - 0x109  :  250 - 0xfa
    "11111010", --  266 - 0x10a  :  250 - 0xfa
    "11111010", --  267 - 0x10b  :  250 - 0xfa
    "11111010", --  268 - 0x10c  :  250 - 0xfa
    "11111010", --  269 - 0x10d  :  250 - 0xfa
    "11111010", --  270 - 0x10e  :  250 - 0xfa
    "11111010", --  271 - 0x10f  :  250 - 0xfa
    "11111010", --  272 - 0x110  :  250 - 0xfa
    "11111100", --  273 - 0x111  :  252 - 0xfc
    "11111111", --  274 - 0x112  :  255 - 0xff
    "11111111", --  275 - 0x113  :  255 - 0xff
    "11111111", --  276 - 0x114  :  255 - 0xff
    "11111111", --  277 - 0x115  :  255 - 0xff
    "11111101", --  278 - 0x116  :  253 - 0xfd
    "11111111", --  279 - 0x117  :  255 - 0xff
    "11111101", --  280 - 0x118  :  253 - 0xfd
    "11111111", --  281 - 0x119  :  255 - 0xff
    "11111101", --  282 - 0x11a  :  253 - 0xfd
    "11111111", --  283 - 0x11b  :  255 - 0xff
    "11111111", --  284 - 0x11c  :  255 - 0xff
    "11111111", --  285 - 0x11d  :  255 - 0xff
    "11101100", --  286 - 0x11e  :  236 - 0xec
    "11111010", --  287 - 0x11f  :  250 - 0xfa
    "11111010", --  288 - 0x120  :  250 - 0xfa
    "11111100", --  289 - 0x121  :  252 - 0xfc
    "11111111", --  290 - 0x122  :  255 - 0xff
    "11111110", --  291 - 0x123  :  254 - 0xfe
    "11111110", --  292 - 0x124  :  254 - 0xfe
    "11111111", --  293 - 0x125  :  255 - 0xff
    "11101100", --  294 - 0x126  :  236 - 0xec
    "11111010", --  295 - 0x127  :  250 - 0xfa
    "11111010", --  296 - 0x128  :  250 - 0xfa
    "11101001", --  297 - 0x129  :  233 - 0xe9
    "11111010", --  298 - 0x12a  :  250 - 0xfa
    "11101001", --  299 - 0x12b  :  233 - 0xe9
    "11111010", --  300 - 0x12c  :  250 - 0xfa
    "11111010", --  301 - 0x12d  :  250 - 0xfa
    "11101001", --  302 - 0x12e  :  233 - 0xe9
    "11111010", --  303 - 0x12f  :  250 - 0xfa
    "11111010", --  304 - 0x130  :  250 - 0xfa
    "11111100", --  305 - 0x131  :  252 - 0xfc
    "11111111", --  306 - 0x132  :  255 - 0xff
    "11111111", --  307 - 0x133  :  255 - 0xff
    "11111111", --  308 - 0x134  :  255 - 0xff
    "11111111", --  309 - 0x135  :  255 - 0xff
    "11111111", --  310 - 0x136  :  255 - 0xff
    "11111111", --  311 - 0x137  :  255 - 0xff
    "11111111", --  312 - 0x138  :  255 - 0xff
    "11111111", --  313 - 0x139  :  255 - 0xff
    "11111111", --  314 - 0x13a  :  255 - 0xff
    "11111111", --  315 - 0x13b  :  255 - 0xff
    "11111111", --  316 - 0x13c  :  255 - 0xff
    "11111111", --  317 - 0x13d  :  255 - 0xff
    "11101100", --  318 - 0x13e  :  236 - 0xec
    "11111010", --  319 - 0x13f  :  250 - 0xfa
    "11111010", --  320 - 0x140  :  250 - 0xfa
    "11111100", --  321 - 0x141  :  252 - 0xfc
    "11111111", --  322 - 0x142  :  255 - 0xff
    "11111111", --  323 - 0x143  :  255 - 0xff
    "11111111", --  324 - 0x144  :  255 - 0xff
    "11111111", --  325 - 0x145  :  255 - 0xff
    "11101100", --  326 - 0x146  :  236 - 0xec
    "11111010", --  327 - 0x147  :  250 - 0xfa
    "11111010", --  328 - 0x148  :  250 - 0xfa
    "11111010", --  329 - 0x149  :  250 - 0xfa
    "11111010", --  330 - 0x14a  :  250 - 0xfa
    "11101001", --  331 - 0x14b  :  233 - 0xe9
    "11111010", --  332 - 0x14c  :  250 - 0xfa
    "11111010", --  333 - 0x14d  :  250 - 0xfa
    "11111010", --  334 - 0x14e  :  250 - 0xfa
    "11111010", --  335 - 0x14f  :  250 - 0xfa
    "11111010", --  336 - 0x150  :  250 - 0xfa
    "11110111", --  337 - 0x151  :  247 - 0xf7
    "11101011", --  338 - 0x152  :  235 - 0xeb
    "11101011", --  339 - 0x153  :  235 - 0xeb
    "11101011", --  340 - 0x154  :  235 - 0xeb
    "11101011", --  341 - 0x155  :  235 - 0xeb
    "11101011", --  342 - 0x156  :  235 - 0xeb
    "11101011", --  343 - 0x157  :  235 - 0xeb
    "11101011", --  344 - 0x158  :  235 - 0xeb
    "11100110", --  345 - 0x159  :  230 - 0xe6
    "11111111", --  346 - 0x15a  :  255 - 0xff
    "11111111", --  347 - 0x15b  :  255 - 0xff
    "11111111", --  348 - 0x15c  :  255 - 0xff
    "11111111", --  349 - 0x15d  :  255 - 0xff
    "11101100", --  350 - 0x15e  :  236 - 0xec
    "11111010", --  351 - 0x15f  :  250 - 0xfa
    "11111010", --  352 - 0x160  :  250 - 0xfa
    "11111100", --  353 - 0x161  :  252 - 0xfc
    "11111111", --  354 - 0x162  :  255 - 0xff
    "11111110", --  355 - 0x163  :  254 - 0xfe
    "11111110", --  356 - 0x164  :  254 - 0xfe
    "11111111", --  357 - 0x165  :  255 - 0xff
    "11101100", --  358 - 0x166  :  236 - 0xec
    "11111010", --  359 - 0x167  :  250 - 0xfa
    "11111010", --  360 - 0x168  :  250 - 0xfa
    "11111010", --  361 - 0x169  :  250 - 0xfa
    "11111010", --  362 - 0x16a  :  250 - 0xfa
    "11111010", --  363 - 0x16b  :  250 - 0xfa
    "11111010", --  364 - 0x16c  :  250 - 0xfa
    "11111010", --  365 - 0x16d  :  250 - 0xfa
    "11111010", --  366 - 0x16e  :  250 - 0xfa
    "11111010", --  367 - 0x16f  :  250 - 0xfa
    "11111010", --  368 - 0x170  :  250 - 0xfa
    "11111010", --  369 - 0x171  :  250 - 0xfa
    "11111010", --  370 - 0x172  :  250 - 0xfa
    "11111010", --  371 - 0x173  :  250 - 0xfa
    "11111010", --  372 - 0x174  :  250 - 0xfa
    "11111010", --  373 - 0x175  :  250 - 0xfa
    "11111010", --  374 - 0x176  :  250 - 0xfa
    "11101001", --  375 - 0x177  :  233 - 0xe9
    "11111010", --  376 - 0x178  :  250 - 0xfa
    "11111100", --  377 - 0x179  :  252 - 0xfc
    "11111111", --  378 - 0x17a  :  255 - 0xff
    "11111110", --  379 - 0x17b  :  254 - 0xfe
    "11111110", --  380 - 0x17c  :  254 - 0xfe
    "11111111", --  381 - 0x17d  :  255 - 0xff
    "11101100", --  382 - 0x17e  :  236 - 0xec
    "11111010", --  383 - 0x17f  :  250 - 0xfa
    "11101001", --  384 - 0x180  :  233 - 0xe9
    "11111100", --  385 - 0x181  :  252 - 0xfc
    "11111111", --  386 - 0x182  :  255 - 0xff
    "11111111", --  387 - 0x183  :  255 - 0xff
    "11111111", --  388 - 0x184  :  255 - 0xff
    "11111111", --  389 - 0x185  :  255 - 0xff
    "11101100", --  390 - 0x186  :  236 - 0xec
    "11111010", --  391 - 0x187  :  250 - 0xfa
    "11111010", --  392 - 0x188  :  250 - 0xfa
    "11111010", --  393 - 0x189  :  250 - 0xfa
    "11111010", --  394 - 0x18a  :  250 - 0xfa
    "11111010", --  395 - 0x18b  :  250 - 0xfa
    "11111010", --  396 - 0x18c  :  250 - 0xfa
    "11111010", --  397 - 0x18d  :  250 - 0xfa
    "11111010", --  398 - 0x18e  :  250 - 0xfa
    "11101001", --  399 - 0x18f  :  233 - 0xe9
    "11111010", --  400 - 0x190  :  250 - 0xfa
    "11101001", --  401 - 0x191  :  233 - 0xe9
    "11111010", --  402 - 0x192  :  250 - 0xfa
    "11111010", --  403 - 0x193  :  250 - 0xfa
    "11111010", --  404 - 0x194  :  250 - 0xfa
    "11111010", --  405 - 0x195  :  250 - 0xfa
    "11111010", --  406 - 0x196  :  250 - 0xfa
    "11111010", --  407 - 0x197  :  250 - 0xfa
    "11111010", --  408 - 0x198  :  250 - 0xfa
    "11111100", --  409 - 0x199  :  252 - 0xfc
    "11111111", --  410 - 0x19a  :  255 - 0xff
    "11111111", --  411 - 0x19b  :  255 - 0xff
    "11111111", --  412 - 0x19c  :  255 - 0xff
    "11111111", --  413 - 0x19d  :  255 - 0xff
    "11101100", --  414 - 0x19e  :  236 - 0xec
    "11111010", --  415 - 0x19f  :  250 - 0xfa
    "11111010", --  416 - 0x1a0  :  250 - 0xfa
    "11111100", --  417 - 0x1a1  :  252 - 0xfc
    "11111111", --  418 - 0x1a2  :  255 - 0xff
    "11111110", --  419 - 0x1a3  :  254 - 0xfe
    "11111110", --  420 - 0x1a4  :  254 - 0xfe
    "11111111", --  421 - 0x1a5  :  255 - 0xff
    "11101100", --  422 - 0x1a6  :  236 - 0xec
    "11111010", --  423 - 0x1a7  :  250 - 0xfa
    "11111001", --  424 - 0x1a8  :  249 - 0xf9
    "11111010", --  425 - 0x1a9  :  250 - 0xfa
    "11111010", --  426 - 0x1aa  :  250 - 0xfa
    "11101001", --  427 - 0x1ab  :  233 - 0xe9
    "11111010", --  428 - 0x1ac  :  250 - 0xfa
    "11111010", --  429 - 0x1ad  :  250 - 0xfa
    "11111010", --  430 - 0x1ae  :  250 - 0xfa
    "11111010", --  431 - 0x1af  :  250 - 0xfa
    "11111010", --  432 - 0x1b0  :  250 - 0xfa
    "11111010", --  433 - 0x1b1  :  250 - 0xfa
    "11111010", --  434 - 0x1b2  :  250 - 0xfa
    "11100111", --  435 - 0x1b3  :  231 - 0xe7
    "11111011", --  436 - 0x1b4  :  251 - 0xfb
    "11111011", --  437 - 0x1b5  :  251 - 0xfb
    "11111011", --  438 - 0x1b6  :  251 - 0xfb
    "11111011", --  439 - 0x1b7  :  251 - 0xfb
    "11111011", --  440 - 0x1b8  :  251 - 0xfb
    "11110110", --  441 - 0x1b9  :  246 - 0xf6
    "11111111", --  442 - 0x1ba  :  255 - 0xff
    "11111110", --  443 - 0x1bb  :  254 - 0xfe
    "11111110", --  444 - 0x1bc  :  254 - 0xfe
    "11111111", --  445 - 0x1bd  :  255 - 0xff
    "11101100", --  446 - 0x1be  :  236 - 0xec
    "11101001", --  447 - 0x1bf  :  233 - 0xe9
    "11111010", --  448 - 0x1c0  :  250 - 0xfa
    "11111100", --  449 - 0x1c1  :  252 - 0xfc
    "11111111", --  450 - 0x1c2  :  255 - 0xff
    "11111111", --  451 - 0x1c3  :  255 - 0xff
    "11111111", --  452 - 0x1c4  :  255 - 0xff
    "11111111", --  453 - 0x1c5  :  255 - 0xff
    "11101100", --  454 - 0x1c6  :  236 - 0xec
    "11111010", --  455 - 0x1c7  :  250 - 0xfa
    "11111010", --  456 - 0x1c8  :  250 - 0xfa
    "11111010", --  457 - 0x1c9  :  250 - 0xfa
    "11101001", --  458 - 0x1ca  :  233 - 0xe9
    "11111010", --  459 - 0x1cb  :  250 - 0xfa
    "11111010", --  460 - 0x1cc  :  250 - 0xfa
    "11111010", --  461 - 0x1cd  :  250 - 0xfa
    "11111010", --  462 - 0x1ce  :  250 - 0xfa
    "11111010", --  463 - 0x1cf  :  250 - 0xfa
    "11111010", --  464 - 0x1d0  :  250 - 0xfa
    "11111010", --  465 - 0x1d1  :  250 - 0xfa
    "11111010", --  466 - 0x1d2  :  250 - 0xfa
    "11111100", --  467 - 0x1d3  :  252 - 0xfc
    "11111111", --  468 - 0x1d4  :  255 - 0xff
    "11111111", --  469 - 0x1d5  :  255 - 0xff
    "11111111", --  470 - 0x1d6  :  255 - 0xff
    "11111111", --  471 - 0x1d7  :  255 - 0xff
    "11111111", --  472 - 0x1d8  :  255 - 0xff
    "11111111", --  473 - 0x1d9  :  255 - 0xff
    "11111111", --  474 - 0x1da  :  255 - 0xff
    "11111111", --  475 - 0x1db  :  255 - 0xff
    "11111111", --  476 - 0x1dc  :  255 - 0xff
    "11111111", --  477 - 0x1dd  :  255 - 0xff
    "11101100", --  478 - 0x1de  :  236 - 0xec
    "11111010", --  479 - 0x1df  :  250 - 0xfa
    "11101010", --  480 - 0x1e0  :  234 - 0xea
    "11111100", --  481 - 0x1e1  :  252 - 0xfc
    "11111111", --  482 - 0x1e2  :  255 - 0xff
    "11111110", --  483 - 0x1e3  :  254 - 0xfe
    "11111110", --  484 - 0x1e4  :  254 - 0xfe
    "11111111", --  485 - 0x1e5  :  255 - 0xff
    "11110101", --  486 - 0x1e6  :  245 - 0xf5
    "11111011", --  487 - 0x1e7  :  251 - 0xfb
    "11111011", --  488 - 0x1e8  :  251 - 0xfb
    "11111011", --  489 - 0x1e9  :  251 - 0xfb
    "11111011", --  490 - 0x1ea  :  251 - 0xfb
    "11111011", --  491 - 0x1eb  :  251 - 0xfb
    "11101000", --  492 - 0x1ec  :  232 - 0xe8
    "11111010", --  493 - 0x1ed  :  250 - 0xfa
    "11111010", --  494 - 0x1ee  :  250 - 0xfa
    "11111010", --  495 - 0x1ef  :  250 - 0xfa
    "11101001", --  496 - 0x1f0  :  233 - 0xe9
    "11111010", --  497 - 0x1f1  :  250 - 0xfa
    "11111010", --  498 - 0x1f2  :  250 - 0xfa
    "11111100", --  499 - 0x1f3  :  252 - 0xfc
    "11111111", --  500 - 0x1f4  :  255 - 0xff
    "11111111", --  501 - 0x1f5  :  255 - 0xff
    "11111111", --  502 - 0x1f6  :  255 - 0xff
    "11111111", --  503 - 0x1f7  :  255 - 0xff
    "11111101", --  504 - 0x1f8  :  253 - 0xfd
    "11111111", --  505 - 0x1f9  :  255 - 0xff
    "11111101", --  506 - 0x1fa  :  253 - 0xfd
    "11111111", --  507 - 0x1fb  :  255 - 0xff
    "11111111", --  508 - 0x1fc  :  255 - 0xff
    "11111111", --  509 - 0x1fd  :  255 - 0xff
    "11101100", --  510 - 0x1fe  :  236 - 0xec
    "11111010", --  511 - 0x1ff  :  250 - 0xfa
    "11111010", --  512 - 0x200  :  250 - 0xfa
    "11111100", --  513 - 0x201  :  252 - 0xfc
    "11111111", --  514 - 0x202  :  255 - 0xff
    "11111111", --  515 - 0x203  :  255 - 0xff
    "11111111", --  516 - 0x204  :  255 - 0xff
    "11111111", --  517 - 0x205  :  255 - 0xff
    "11111111", --  518 - 0x206  :  255 - 0xff
    "11111111", --  519 - 0x207  :  255 - 0xff
    "11111111", --  520 - 0x208  :  255 - 0xff
    "11111111", --  521 - 0x209  :  255 - 0xff
    "11111111", --  522 - 0x20a  :  255 - 0xff
    "11111111", --  523 - 0x20b  :  255 - 0xff
    "11101100", --  524 - 0x20c  :  236 - 0xec
    "11111010", --  525 - 0x20d  :  250 - 0xfa
    "11111010", --  526 - 0x20e  :  250 - 0xfa
    "11111010", --  527 - 0x20f  :  250 - 0xfa
    "11111010", --  528 - 0x210  :  250 - 0xfa
    "11111010", --  529 - 0x211  :  250 - 0xfa
    "11111010", --  530 - 0x212  :  250 - 0xfa
    "11111100", --  531 - 0x213  :  252 - 0xfc
    "11111111", --  532 - 0x214  :  255 - 0xff
    "11111111", --  533 - 0x215  :  255 - 0xff
    "11111111", --  534 - 0x216  :  255 - 0xff
    "11111111", --  535 - 0x217  :  255 - 0xff
    "11111101", --  536 - 0x218  :  253 - 0xfd
    "11111111", --  537 - 0x219  :  255 - 0xff
    "11111101", --  538 - 0x21a  :  253 - 0xfd
    "11111111", --  539 - 0x21b  :  255 - 0xff
    "11111111", --  540 - 0x21c  :  255 - 0xff
    "11111111", --  541 - 0x21d  :  255 - 0xff
    "11101100", --  542 - 0x21e  :  236 - 0xec
    "11101010", --  543 - 0x21f  :  234 - 0xea
    "11111010", --  544 - 0x220  :  250 - 0xfa
    "11111100", --  545 - 0x221  :  252 - 0xfc
    "11111111", --  546 - 0x222  :  255 - 0xff
    "11111111", --  547 - 0x223  :  255 - 0xff
    "11111111", --  548 - 0x224  :  255 - 0xff
    "11111111", --  549 - 0x225  :  255 - 0xff
    "11111101", --  550 - 0x226  :  253 - 0xfd
    "11111111", --  551 - 0x227  :  255 - 0xff
    "11111101", --  552 - 0x228  :  253 - 0xfd
    "11111111", --  553 - 0x229  :  255 - 0xff
    "11111111", --  554 - 0x22a  :  255 - 0xff
    "11111111", --  555 - 0x22b  :  255 - 0xff
    "11101100", --  556 - 0x22c  :  236 - 0xec
    "11111010", --  557 - 0x22d  :  250 - 0xfa
    "11111010", --  558 - 0x22e  :  250 - 0xfa
    "11111010", --  559 - 0x22f  :  250 - 0xfa
    "11111010", --  560 - 0x230  :  250 - 0xfa
    "11111010", --  561 - 0x231  :  250 - 0xfa
    "11111010", --  562 - 0x232  :  250 - 0xfa
    "11111100", --  563 - 0x233  :  252 - 0xfc
    "11111111", --  564 - 0x234  :  255 - 0xff
    "11111110", --  565 - 0x235  :  254 - 0xfe
    "11111110", --  566 - 0x236  :  254 - 0xfe
    "11111111", --  567 - 0x237  :  255 - 0xff
    "11111111", --  568 - 0x238  :  255 - 0xff
    "11111111", --  569 - 0x239  :  255 - 0xff
    "11111111", --  570 - 0x23a  :  255 - 0xff
    "11111111", --  571 - 0x23b  :  255 - 0xff
    "11111111", --  572 - 0x23c  :  255 - 0xff
    "11111111", --  573 - 0x23d  :  255 - 0xff
    "11101100", --  574 - 0x23e  :  236 - 0xec
    "11111010", --  575 - 0x23f  :  250 - 0xfa
    "11111010", --  576 - 0x240  :  250 - 0xfa
    "11111100", --  577 - 0x241  :  252 - 0xfc
    "11111111", --  578 - 0x242  :  255 - 0xff
    "11111111", --  579 - 0x243  :  255 - 0xff
    "11111111", --  580 - 0x244  :  255 - 0xff
    "11111111", --  581 - 0x245  :  255 - 0xff
    "11111101", --  582 - 0x246  :  253 - 0xfd
    "11111111", --  583 - 0x247  :  255 - 0xff
    "11111101", --  584 - 0x248  :  253 - 0xfd
    "11111111", --  585 - 0x249  :  255 - 0xff
    "11111111", --  586 - 0x24a  :  255 - 0xff
    "11111111", --  587 - 0x24b  :  255 - 0xff
    "11101100", --  588 - 0x24c  :  236 - 0xec
    "11111010", --  589 - 0x24d  :  250 - 0xfa
    "11111010", --  590 - 0x24e  :  250 - 0xfa
    "11101001", --  591 - 0x24f  :  233 - 0xe9
    "11111010", --  592 - 0x250  :  250 - 0xfa
    "11111010", --  593 - 0x251  :  250 - 0xfa
    "11111010", --  594 - 0x252  :  250 - 0xfa
    "11111100", --  595 - 0x253  :  252 - 0xfc
    "11111111", --  596 - 0x254  :  255 - 0xff
    "11111111", --  597 - 0x255  :  255 - 0xff
    "11111111", --  598 - 0x256  :  255 - 0xff
    "11111111", --  599 - 0x257  :  255 - 0xff
    "11100101", --  600 - 0x258  :  229 - 0xe5
    "11101011", --  601 - 0x259  :  235 - 0xeb
    "11101011", --  602 - 0x25a  :  235 - 0xeb
    "11101011", --  603 - 0x25b  :  235 - 0xeb
    "11101011", --  604 - 0x25c  :  235 - 0xeb
    "11101011", --  605 - 0x25d  :  235 - 0xeb
    "11111000", --  606 - 0x25e  :  248 - 0xf8
    "11111010", --  607 - 0x25f  :  250 - 0xfa
    "11111010", --  608 - 0x260  :  250 - 0xfa
    "11111100", --  609 - 0x261  :  252 - 0xfc
    "11111111", --  610 - 0x262  :  255 - 0xff
    "11111111", --  611 - 0x263  :  255 - 0xff
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111111", --  613 - 0x265  :  255 - 0xff
    "11111111", --  614 - 0x266  :  255 - 0xff
    "11111111", --  615 - 0x267  :  255 - 0xff
    "11111111", --  616 - 0x268  :  255 - 0xff
    "11111111", --  617 - 0x269  :  255 - 0xff
    "11111111", --  618 - 0x26a  :  255 - 0xff
    "11111111", --  619 - 0x26b  :  255 - 0xff
    "11101100", --  620 - 0x26c  :  236 - 0xec
    "11111010", --  621 - 0x26d  :  250 - 0xfa
    "11111010", --  622 - 0x26e  :  250 - 0xfa
    "11111010", --  623 - 0x26f  :  250 - 0xfa
    "11111010", --  624 - 0x270  :  250 - 0xfa
    "11111010", --  625 - 0x271  :  250 - 0xfa
    "11111010", --  626 - 0x272  :  250 - 0xfa
    "11111100", --  627 - 0x273  :  252 - 0xfc
    "11111111", --  628 - 0x274  :  255 - 0xff
    "11111110", --  629 - 0x275  :  254 - 0xfe
    "11111110", --  630 - 0x276  :  254 - 0xfe
    "11111111", --  631 - 0x277  :  255 - 0xff
    "11110101", --  632 - 0x278  :  245 - 0xf5
    "11111011", --  633 - 0x279  :  251 - 0xfb
    "11111011", --  634 - 0x27a  :  251 - 0xfb
    "11111011", --  635 - 0x27b  :  251 - 0xfb
    "11111011", --  636 - 0x27c  :  251 - 0xfb
    "11111011", --  637 - 0x27d  :  251 - 0xfb
    "11101000", --  638 - 0x27e  :  232 - 0xe8
    "11111010", --  639 - 0x27f  :  250 - 0xfa
    "11111010", --  640 - 0x280  :  250 - 0xfa
    "11110111", --  641 - 0x281  :  247 - 0xf7
    "11101011", --  642 - 0x282  :  235 - 0xeb
    "11101011", --  643 - 0x283  :  235 - 0xeb
    "11101011", --  644 - 0x284  :  235 - 0xeb
    "11101011", --  645 - 0x285  :  235 - 0xeb
    "11101011", --  646 - 0x286  :  235 - 0xeb
    "11100110", --  647 - 0x287  :  230 - 0xe6
    "11111111", --  648 - 0x288  :  255 - 0xff
    "11111111", --  649 - 0x289  :  255 - 0xff
    "11111111", --  650 - 0x28a  :  255 - 0xff
    "11111111", --  651 - 0x28b  :  255 - 0xff
    "11101100", --  652 - 0x28c  :  236 - 0xec
    "11111010", --  653 - 0x28d  :  250 - 0xfa
    "11111010", --  654 - 0x28e  :  250 - 0xfa
    "11101001", --  655 - 0x28f  :  233 - 0xe9
    "11111010", --  656 - 0x290  :  250 - 0xfa
    "11111010", --  657 - 0x291  :  250 - 0xfa
    "11111010", --  658 - 0x292  :  250 - 0xfa
    "11111100", --  659 - 0x293  :  252 - 0xfc
    "11111111", --  660 - 0x294  :  255 - 0xff
    "11111111", --  661 - 0x295  :  255 - 0xff
    "11111111", --  662 - 0x296  :  255 - 0xff
    "11111111", --  663 - 0x297  :  255 - 0xff
    "11111111", --  664 - 0x298  :  255 - 0xff
    "11111111", --  665 - 0x299  :  255 - 0xff
    "11111111", --  666 - 0x29a  :  255 - 0xff
    "11111111", --  667 - 0x29b  :  255 - 0xff
    "11111111", --  668 - 0x29c  :  255 - 0xff
    "11111111", --  669 - 0x29d  :  255 - 0xff
    "11101100", --  670 - 0x29e  :  236 - 0xec
    "11111010", --  671 - 0x29f  :  250 - 0xfa
    "11111010", --  672 - 0x2a0  :  250 - 0xfa
    "11111010", --  673 - 0x2a1  :  250 - 0xfa
    "11101010", --  674 - 0x2a2  :  234 - 0xea
    "11101001", --  675 - 0x2a3  :  233 - 0xe9
    "11111010", --  676 - 0x2a4  :  250 - 0xfa
    "11111010", --  677 - 0x2a5  :  250 - 0xfa
    "11111010", --  678 - 0x2a6  :  250 - 0xfa
    "11111100", --  679 - 0x2a7  :  252 - 0xfc
    "11111111", --  680 - 0x2a8  :  255 - 0xff
    "11111110", --  681 - 0x2a9  :  254 - 0xfe
    "11111110", --  682 - 0x2aa  :  254 - 0xfe
    "11111111", --  683 - 0x2ab  :  255 - 0xff
    "11101100", --  684 - 0x2ac  :  236 - 0xec
    "11111010", --  685 - 0x2ad  :  250 - 0xfa
    "11111010", --  686 - 0x2ae  :  250 - 0xfa
    "11111010", --  687 - 0x2af  :  250 - 0xfa
    "11111010", --  688 - 0x2b0  :  250 - 0xfa
    "11101001", --  689 - 0x2b1  :  233 - 0xe9
    "11111010", --  690 - 0x2b2  :  250 - 0xfa
    "11111100", --  691 - 0x2b3  :  252 - 0xfc
    "11111111", --  692 - 0x2b4  :  255 - 0xff
    "11111111", --  693 - 0x2b5  :  255 - 0xff
    "11111111", --  694 - 0x2b6  :  255 - 0xff
    "11111111", --  695 - 0x2b7  :  255 - 0xff
    "11111111", --  696 - 0x2b8  :  255 - 0xff
    "11111111", --  697 - 0x2b9  :  255 - 0xff
    "11111111", --  698 - 0x2ba  :  255 - 0xff
    "11111111", --  699 - 0x2bb  :  255 - 0xff
    "11111111", --  700 - 0x2bc  :  255 - 0xff
    "11111111", --  701 - 0x2bd  :  255 - 0xff
    "11101100", --  702 - 0x2be  :  236 - 0xec
    "11111010", --  703 - 0x2bf  :  250 - 0xfa
    "11111010", --  704 - 0x2c0  :  250 - 0xfa
    "11111010", --  705 - 0x2c1  :  250 - 0xfa
    "11111010", --  706 - 0x2c2  :  250 - 0xfa
    "11111010", --  707 - 0x2c3  :  250 - 0xfa
    "11111010", --  708 - 0x2c4  :  250 - 0xfa
    "11111010", --  709 - 0x2c5  :  250 - 0xfa
    "11101001", --  710 - 0x2c6  :  233 - 0xe9
    "11111100", --  711 - 0x2c7  :  252 - 0xfc
    "11111111", --  712 - 0x2c8  :  255 - 0xff
    "11111111", --  713 - 0x2c9  :  255 - 0xff
    "11111111", --  714 - 0x2ca  :  255 - 0xff
    "11111111", --  715 - 0x2cb  :  255 - 0xff
    "11101100", --  716 - 0x2cc  :  236 - 0xec
    "11111010", --  717 - 0x2cd  :  250 - 0xfa
    "11111010", --  718 - 0x2ce  :  250 - 0xfa
    "11111010", --  719 - 0x2cf  :  250 - 0xfa
    "11111010", --  720 - 0x2d0  :  250 - 0xfa
    "11111010", --  721 - 0x2d1  :  250 - 0xfa
    "11111010", --  722 - 0x2d2  :  250 - 0xfa
    "11110111", --  723 - 0x2d3  :  247 - 0xf7
    "11101011", --  724 - 0x2d4  :  235 - 0xeb
    "11101011", --  725 - 0x2d5  :  235 - 0xeb
    "11101011", --  726 - 0x2d6  :  235 - 0xeb
    "11101011", --  727 - 0x2d7  :  235 - 0xeb
    "11101011", --  728 - 0x2d8  :  235 - 0xeb
    "11100110", --  729 - 0x2d9  :  230 - 0xe6
    "11111111", --  730 - 0x2da  :  255 - 0xff
    "11111111", --  731 - 0x2db  :  255 - 0xff
    "11111111", --  732 - 0x2dc  :  255 - 0xff
    "11111111", --  733 - 0x2dd  :  255 - 0xff
    "11101100", --  734 - 0x2de  :  236 - 0xec
    "11111010", --  735 - 0x2df  :  250 - 0xfa
    "11111010", --  736 - 0x2e0  :  250 - 0xfa
    "11111010", --  737 - 0x2e1  :  250 - 0xfa
    "11101001", --  738 - 0x2e2  :  233 - 0xe9
    "11111010", --  739 - 0x2e3  :  250 - 0xfa
    "11111010", --  740 - 0x2e4  :  250 - 0xfa
    "11111010", --  741 - 0x2e5  :  250 - 0xfa
    "11111010", --  742 - 0x2e6  :  250 - 0xfa
    "11111100", --  743 - 0x2e7  :  252 - 0xfc
    "11111111", --  744 - 0x2e8  :  255 - 0xff
    "11111110", --  745 - 0x2e9  :  254 - 0xfe
    "11111110", --  746 - 0x2ea  :  254 - 0xfe
    "11111111", --  747 - 0x2eb  :  255 - 0xff
    "11110101", --  748 - 0x2ec  :  245 - 0xf5
    "11111011", --  749 - 0x2ed  :  251 - 0xfb
    "11111011", --  750 - 0x2ee  :  251 - 0xfb
    "11111011", --  751 - 0x2ef  :  251 - 0xfb
    "11111011", --  752 - 0x2f0  :  251 - 0xfb
    "11111011", --  753 - 0x2f1  :  251 - 0xfb
    "11111011", --  754 - 0x2f2  :  251 - 0xfb
    "11111011", --  755 - 0x2f3  :  251 - 0xfb
    "11111011", --  756 - 0x2f4  :  251 - 0xfb
    "11111011", --  757 - 0x2f5  :  251 - 0xfb
    "11111011", --  758 - 0x2f6  :  251 - 0xfb
    "11111011", --  759 - 0x2f7  :  251 - 0xfb
    "11111011", --  760 - 0x2f8  :  251 - 0xfb
    "11110110", --  761 - 0x2f9  :  246 - 0xf6
    "11111111", --  762 - 0x2fa  :  255 - 0xff
    "11111110", --  763 - 0x2fb  :  254 - 0xfe
    "11111110", --  764 - 0x2fc  :  254 - 0xfe
    "11111111", --  765 - 0x2fd  :  255 - 0xff
    "11101100", --  766 - 0x2fe  :  236 - 0xec
    "11111010", --  767 - 0x2ff  :  250 - 0xfa
    "11111010", --  768 - 0x300  :  250 - 0xfa
    "11111010", --  769 - 0x301  :  250 - 0xfa
    "11111010", --  770 - 0x302  :  250 - 0xfa
    "11111010", --  771 - 0x303  :  250 - 0xfa
    "11111010", --  772 - 0x304  :  250 - 0xfa
    "11111010", --  773 - 0x305  :  250 - 0xfa
    "11111010", --  774 - 0x306  :  250 - 0xfa
    "11111100", --  775 - 0x307  :  252 - 0xfc
    "11111111", --  776 - 0x308  :  255 - 0xff
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11111111", --  778 - 0x30a  :  255 - 0xff
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "11111111", --  780 - 0x30c  :  255 - 0xff
    "11111111", --  781 - 0x30d  :  255 - 0xff
    "11111111", --  782 - 0x30e  :  255 - 0xff
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "11111111", --  784 - 0x310  :  255 - 0xff
    "11111111", --  785 - 0x311  :  255 - 0xff
    "11101111", --  786 - 0x312  :  239 - 0xef
    "11111111", --  787 - 0x313  :  255 - 0xff
    "11111111", --  788 - 0x314  :  255 - 0xff
    "11111111", --  789 - 0x315  :  255 - 0xff
    "11111111", --  790 - 0x316  :  255 - 0xff
    "11111111", --  791 - 0x317  :  255 - 0xff
    "11111111", --  792 - 0x318  :  255 - 0xff
    "11111111", --  793 - 0x319  :  255 - 0xff
    "11111111", --  794 - 0x31a  :  255 - 0xff
    "11111111", --  795 - 0x31b  :  255 - 0xff
    "11111111", --  796 - 0x31c  :  255 - 0xff
    "11111111", --  797 - 0x31d  :  255 - 0xff
    "11101100", --  798 - 0x31e  :  236 - 0xec
    "11101001", --  799 - 0x31f  :  233 - 0xe9
    "11101010", --  800 - 0x320  :  234 - 0xea
    "00001101", --  801 - 0x321  :   13 - 0xd
    "00000001", --  802 - 0x322  :    1 - 0x1
    "00000010", --  803 - 0x323  :    2 - 0x2
    "00000010", --  804 - 0x324  :    2 - 0x2
    "11111010", --  805 - 0x325  :  250 - 0xfa
    "11111010", --  806 - 0x326  :  250 - 0xfa
    "11111100", --  807 - 0x327  :  252 - 0xfc
    "11111111", --  808 - 0x328  :  255 - 0xff
    "11111111", --  809 - 0x329  :  255 - 0xff
    "11111111", --  810 - 0x32a  :  255 - 0xff
    "11111111", --  811 - 0x32b  :  255 - 0xff
    "11111101", --  812 - 0x32c  :  253 - 0xfd
    "11111111", --  813 - 0x32d  :  255 - 0xff
    "11111101", --  814 - 0x32e  :  253 - 0xfd
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "11111101", --  816 - 0x330  :  253 - 0xfd
    "11111111", --  817 - 0x331  :  255 - 0xff
    "11101111", --  818 - 0x332  :  239 - 0xef
    "11111111", --  819 - 0x333  :  255 - 0xff
    "11111101", --  820 - 0x334  :  253 - 0xfd
    "11111111", --  821 - 0x335  :  255 - 0xff
    "11111101", --  822 - 0x336  :  253 - 0xfd
    "11111111", --  823 - 0x337  :  255 - 0xff
    "11111101", --  824 - 0x338  :  253 - 0xfd
    "11111111", --  825 - 0x339  :  255 - 0xff
    "11111111", --  826 - 0x33a  :  255 - 0xff
    "11111111", --  827 - 0x33b  :  255 - 0xff
    "11111111", --  828 - 0x33c  :  255 - 0xff
    "11111111", --  829 - 0x33d  :  255 - 0xff
    "11101100", --  830 - 0x33e  :  236 - 0xec
    "11111010", --  831 - 0x33f  :  250 - 0xfa
    "11111010", --  832 - 0x340  :  250 - 0xfa
    "11111010", --  833 - 0x341  :  250 - 0xfa
    "11111010", --  834 - 0x342  :  250 - 0xfa
    "11111010", --  835 - 0x343  :  250 - 0xfa
    "11111010", --  836 - 0x344  :  250 - 0xfa
    "11111010", --  837 - 0x345  :  250 - 0xfa
    "11111010", --  838 - 0x346  :  250 - 0xfa
    "11111100", --  839 - 0x347  :  252 - 0xfc
    "11111111", --  840 - 0x348  :  255 - 0xff
    "11111111", --  841 - 0x349  :  255 - 0xff
    "11111111", --  842 - 0x34a  :  255 - 0xff
    "11111111", --  843 - 0x34b  :  255 - 0xff
    "11111101", --  844 - 0x34c  :  253 - 0xfd
    "11111111", --  845 - 0x34d  :  255 - 0xff
    "11111101", --  846 - 0x34e  :  253 - 0xfd
    "11111111", --  847 - 0x34f  :  255 - 0xff
    "11111101", --  848 - 0x350  :  253 - 0xfd
    "11111111", --  849 - 0x351  :  255 - 0xff
    "11101111", --  850 - 0x352  :  239 - 0xef
    "11111111", --  851 - 0x353  :  255 - 0xff
    "11111101", --  852 - 0x354  :  253 - 0xfd
    "11111111", --  853 - 0x355  :  255 - 0xff
    "11111101", --  854 - 0x356  :  253 - 0xfd
    "11111111", --  855 - 0x357  :  255 - 0xff
    "11111101", --  856 - 0x358  :  253 - 0xfd
    "11111111", --  857 - 0x359  :  255 - 0xff
    "11111111", --  858 - 0x35a  :  255 - 0xff
    "11111111", --  859 - 0x35b  :  255 - 0xff
    "11111111", --  860 - 0x35c  :  255 - 0xff
    "11111111", --  861 - 0x35d  :  255 - 0xff
    "11101100", --  862 - 0x35e  :  236 - 0xec
    "11111010", --  863 - 0x35f  :  250 - 0xfa
    "11111010", --  864 - 0x360  :  250 - 0xfa
    "00001111", --  865 - 0x361  :   15 - 0xf
    "00000001", --  866 - 0x362  :    1 - 0x1
    "00010000", --  867 - 0x363  :   16 - 0x10
    "00000011", --  868 - 0x364  :    3 - 0x3
    "11111010", --  869 - 0x365  :  250 - 0xfa
    "11111010", --  870 - 0x366  :  250 - 0xfa
    "11111100", --  871 - 0x367  :  252 - 0xfc
    "11111111", --  872 - 0x368  :  255 - 0xff
    "11111111", --  873 - 0x369  :  255 - 0xff
    "11111111", --  874 - 0x36a  :  255 - 0xff
    "11111111", --  875 - 0x36b  :  255 - 0xff
    "11111111", --  876 - 0x36c  :  255 - 0xff
    "11111111", --  877 - 0x36d  :  255 - 0xff
    "11111111", --  878 - 0x36e  :  255 - 0xff
    "11111111", --  879 - 0x36f  :  255 - 0xff
    "11111111", --  880 - 0x370  :  255 - 0xff
    "11111111", --  881 - 0x371  :  255 - 0xff
    "11101111", --  882 - 0x372  :  239 - 0xef
    "11111111", --  883 - 0x373  :  255 - 0xff
    "11111111", --  884 - 0x374  :  255 - 0xff
    "11111111", --  885 - 0x375  :  255 - 0xff
    "11111111", --  886 - 0x376  :  255 - 0xff
    "11111111", --  887 - 0x377  :  255 - 0xff
    "11111111", --  888 - 0x378  :  255 - 0xff
    "11111111", --  889 - 0x379  :  255 - 0xff
    "11111111", --  890 - 0x37a  :  255 - 0xff
    "11111111", --  891 - 0x37b  :  255 - 0xff
    "11111111", --  892 - 0x37c  :  255 - 0xff
    "11111111", --  893 - 0x37d  :  255 - 0xff
    "11101100", --  894 - 0x37e  :  236 - 0xec
    "11111010", --  895 - 0x37f  :  250 - 0xfa
    "11111010", --  896 - 0x380  :  250 - 0xfa
    "11111010", --  897 - 0x381  :  250 - 0xfa
    "11111001", --  898 - 0x382  :  249 - 0xf9
    "11111010", --  899 - 0x383  :  250 - 0xfa
    "11111010", --  900 - 0x384  :  250 - 0xfa
    "11101010", --  901 - 0x385  :  234 - 0xea
    "11111010", --  902 - 0x386  :  250 - 0xfa
    "11110111", --  903 - 0x387  :  247 - 0xf7
    "11101011", --  904 - 0x388  :  235 - 0xeb
    "11101011", --  905 - 0x389  :  235 - 0xeb
    "11101011", --  906 - 0x38a  :  235 - 0xeb
    "11101011", --  907 - 0x38b  :  235 - 0xeb
    "11101011", --  908 - 0x38c  :  235 - 0xeb
    "11101011", --  909 - 0x38d  :  235 - 0xeb
    "11101011", --  910 - 0x38e  :  235 - 0xeb
    "11101011", --  911 - 0x38f  :  235 - 0xeb
    "11101011", --  912 - 0x390  :  235 - 0xeb
    "11101011", --  913 - 0x391  :  235 - 0xeb
    "11101011", --  914 - 0x392  :  235 - 0xeb
    "11101011", --  915 - 0x393  :  235 - 0xeb
    "11101011", --  916 - 0x394  :  235 - 0xeb
    "11101011", --  917 - 0x395  :  235 - 0xeb
    "11101011", --  918 - 0x396  :  235 - 0xeb
    "11101011", --  919 - 0x397  :  235 - 0xeb
    "11101011", --  920 - 0x398  :  235 - 0xeb
    "11101011", --  921 - 0x399  :  235 - 0xeb
    "11101011", --  922 - 0x39a  :  235 - 0xeb
    "11101011", --  923 - 0x39b  :  235 - 0xeb
    "11101011", --  924 - 0x39c  :  235 - 0xeb
    "11101011", --  925 - 0x39d  :  235 - 0xeb
    "11111000", --  926 - 0x39e  :  248 - 0xf8
    "11111010", --  927 - 0x39f  :  250 - 0xfa
    "11111010", --  928 - 0x3a0  :  250 - 0xfa
    "11111001", --  929 - 0x3a1  :  249 - 0xf9
    "11111010", --  930 - 0x3a2  :  250 - 0xfa
    "11111010", --  931 - 0x3a3  :  250 - 0xfa
    "11111010", --  932 - 0x3a4  :  250 - 0xfa
    "11111010", --  933 - 0x3a5  :  250 - 0xfa
    "11111010", --  934 - 0x3a6  :  250 - 0xfa
    "11111010", --  935 - 0x3a7  :  250 - 0xfa
    "11111010", --  936 - 0x3a8  :  250 - 0xfa
    "11111010", --  937 - 0x3a9  :  250 - 0xfa
    "11111010", --  938 - 0x3aa  :  250 - 0xfa
    "11111010", --  939 - 0x3ab  :  250 - 0xfa
    "11111010", --  940 - 0x3ac  :  250 - 0xfa
    "11111010", --  941 - 0x3ad  :  250 - 0xfa
    "11111010", --  942 - 0x3ae  :  250 - 0xfa
    "11111010", --  943 - 0x3af  :  250 - 0xfa
    "11111010", --  944 - 0x3b0  :  250 - 0xfa
    "11111010", --  945 - 0x3b1  :  250 - 0xfa
    "11111010", --  946 - 0x3b2  :  250 - 0xfa
    "11111010", --  947 - 0x3b3  :  250 - 0xfa
    "11111010", --  948 - 0x3b4  :  250 - 0xfa
    "11101001", --  949 - 0x3b5  :  233 - 0xe9
    "11111010", --  950 - 0x3b6  :  250 - 0xfa
    "11111010", --  951 - 0x3b7  :  250 - 0xfa
    "11111010", --  952 - 0x3b8  :  250 - 0xfa
    "11111010", --  953 - 0x3b9  :  250 - 0xfa
    "11111010", --  954 - 0x3ba  :  250 - 0xfa
    "11111010", --  955 - 0x3bb  :  250 - 0xfa
    "11101010", --  956 - 0x3bc  :  234 - 0xea
    "11111010", --  957 - 0x3bd  :  250 - 0xfa
    "11111010", --  958 - 0x3be  :  250 - 0xfa
    "11111010", --  959 - 0x3bf  :  250 - 0xfa
        ---- Attribute Table 0----
    "00010101", --  960 - 0x3c0  :   21 - 0x15
    "00000101", --  961 - 0x3c1  :    5 - 0x5
    "00000101", --  962 - 0x3c2  :    5 - 0x5
    "00000101", --  963 - 0x3c3  :    5 - 0x5
    "00000101", --  964 - 0x3c4  :    5 - 0x5
    "01000101", --  965 - 0x3c5  :   69 - 0x45
    "01010101", --  966 - 0x3c6  :   85 - 0x55
    "01010101", --  967 - 0x3c7  :   85 - 0x55
    "00010001", --  968 - 0x3c8  :   17 - 0x11
    "01000000", --  969 - 0x3c9  :   64 - 0x40
    "01010000", --  970 - 0x3ca  :   80 - 0x50
    "01010000", --  971 - 0x3cb  :   80 - 0x50
    "00010000", --  972 - 0x3cc  :   16 - 0x10
    "00000100", --  973 - 0x3cd  :    4 - 0x4
    "00000101", --  974 - 0x3ce  :    5 - 0x5
    "01000101", --  975 - 0x3cf  :   69 - 0x45
    "00010001", --  976 - 0x3d0  :   17 - 0x11
    "01000100", --  977 - 0x3d1  :   68 - 0x44
    "01010101", --  978 - 0x3d2  :   85 - 0x55
    "01010101", --  979 - 0x3d3  :   85 - 0x55
    "01010001", --  980 - 0x3d4  :   81 - 0x51
    "01010000", --  981 - 0x3d5  :   80 - 0x50
    "00010000", --  982 - 0x3d6  :   16 - 0x10
    "01000100", --  983 - 0x3d7  :   68 - 0x44
    "00010001", --  984 - 0x3d8  :   17 - 0x11
    "01000100", --  985 - 0x3d9  :   68 - 0x44
    "01010101", --  986 - 0x3da  :   85 - 0x55
    "01010101", --  987 - 0x3db  :   85 - 0x55
    "01010101", --  988 - 0x3dc  :   85 - 0x55
    "00000101", --  989 - 0x3dd  :    5 - 0x5
    "00000001", --  990 - 0x3de  :    1 - 0x1
    "01000100", --  991 - 0x3df  :   68 - 0x44
    "00010001", --  992 - 0x3e0  :   17 - 0x11
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "01010101", --  995 - 0x3e3  :   85 - 0x55
    "01010101", --  996 - 0x3e4  :   85 - 0x55
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "01010000", --  998 - 0x3e6  :   80 - 0x50
    "01010100", --  999 - 0x3e7  :   84 - 0x54
    "01010101", -- 1000 - 0x3e8  :   85 - 0x55
    "01010101", -- 1001 - 0x3e9  :   85 - 0x55
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "01010101", -- 1003 - 0x3eb  :   85 - 0x55
    "01010101", -- 1004 - 0x3ec  :   85 - 0x55
    "01010000", -- 1005 - 0x3ed  :   80 - 0x50
    "00010000", -- 1006 - 0x3ee  :   16 - 0x10
    "01000100", -- 1007 - 0x3ef  :   68 - 0x44
    "01010101", -- 1008 - 0x3f0  :   85 - 0x55
    "01010101", -- 1009 - 0x3f1  :   85 - 0x55
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "01000100", -- 1015 - 0x3f7  :   68 - 0x44
    "00000101", -- 1016 - 0x3f8  :    5 - 0x5
    "00000101", -- 1017 - 0x3f9  :    5 - 0x5
    "00000101", -- 1018 - 0x3fa  :    5 - 0x5
    "00000101", -- 1019 - 0x3fb  :    5 - 0x5
    "00000101", -- 1020 - 0x3fc  :    5 - 0x5
    "00000101", -- 1021 - 0x3fd  :    5 - 0x5
    "00000101", -- 1022 - 0x3fe  :    5 - 0x5
    "00000101", -- 1023 - 0x3ff  :    5 - 0x5
     ------- Name Table 1---------
    "00000000", -- 1024 - 0x400  :    0 - 0x0
    "00000000", -- 1025 - 0x401  :    0 - 0x0
    "00000000", -- 1026 - 0x402  :    0 - 0x0
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00000000", -- 1029 - 0x405  :    0 - 0x0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00000000", -- 1032 - 0x408  :    0 - 0x0
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "00000000", -- 1045 - 0x415  :    0 - 0x0
    "00000000", -- 1046 - 0x416  :    0 - 0x0
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0
    "00000000", -- 1057 - 0x421  :    0 - 0x0
    "00000000", -- 1058 - 0x422  :    0 - 0x0
    "00000000", -- 1059 - 0x423  :    0 - 0x0
    "00000000", -- 1060 - 0x424  :    0 - 0x0
    "00000000", -- 1061 - 0x425  :    0 - 0x0
    "00000000", -- 1062 - 0x426  :    0 - 0x0
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0
    "00000000", -- 1089 - 0x441  :    0 - 0x0
    "00000000", -- 1090 - 0x442  :    0 - 0x0
    "00000000", -- 1091 - 0x443  :    0 - 0x0
    "00000000", -- 1092 - 0x444  :    0 - 0x0
    "00000000", -- 1093 - 0x445  :    0 - 0x0
    "00000000", -- 1094 - 0x446  :    0 - 0x0
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00000000", -- 1096 - 0x448  :    0 - 0x0
    "00000000", -- 1097 - 0x449  :    0 - 0x0
    "00000000", -- 1098 - 0x44a  :    0 - 0x0
    "00000000", -- 1099 - 0x44b  :    0 - 0x0
    "00000000", -- 1100 - 0x44c  :    0 - 0x0
    "00000000", -- 1101 - 0x44d  :    0 - 0x0
    "00000000", -- 1102 - 0x44e  :    0 - 0x0
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0
    "00000000", -- 1105 - 0x451  :    0 - 0x0
    "00000000", -- 1106 - 0x452  :    0 - 0x0
    "00000000", -- 1107 - 0x453  :    0 - 0x0
    "00000000", -- 1108 - 0x454  :    0 - 0x0
    "00000000", -- 1109 - 0x455  :    0 - 0x0
    "00000000", -- 1110 - 0x456  :    0 - 0x0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00000000", -- 1112 - 0x458  :    0 - 0x0
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "00000000", -- 1114 - 0x45a  :    0 - 0x0
    "00000000", -- 1115 - 0x45b  :    0 - 0x0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00000000", -- 1117 - 0x45d  :    0 - 0x0
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000000", -- 1120 - 0x460  :    0 - 0x0
    "00000000", -- 1121 - 0x461  :    0 - 0x0
    "00000000", -- 1122 - 0x462  :    0 - 0x0
    "00000000", -- 1123 - 0x463  :    0 - 0x0
    "00000000", -- 1124 - 0x464  :    0 - 0x0
    "00000000", -- 1125 - 0x465  :    0 - 0x0
    "00000000", -- 1126 - 0x466  :    0 - 0x0
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000000", -- 1128 - 0x468  :    0 - 0x0
    "00000000", -- 1129 - 0x469  :    0 - 0x0
    "00000000", -- 1130 - 0x46a  :    0 - 0x0
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0
    "00000000", -- 1137 - 0x471  :    0 - 0x0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "00000000", -- 1140 - 0x474  :    0 - 0x0
    "00000000", -- 1141 - 0x475  :    0 - 0x0
    "00000000", -- 1142 - 0x476  :    0 - 0x0
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000000", -- 1144 - 0x478  :    0 - 0x0
    "00000000", -- 1145 - 0x479  :    0 - 0x0
    "00000000", -- 1146 - 0x47a  :    0 - 0x0
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00000000", -- 1156 - 0x484  :    0 - 0x0
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "00000000", -- 1158 - 0x486  :    0 - 0x0
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0
    "00000000", -- 1169 - 0x491  :    0 - 0x0
    "00000000", -- 1170 - 0x492  :    0 - 0x0
    "00000000", -- 1171 - 0x493  :    0 - 0x0
    "00000000", -- 1172 - 0x494  :    0 - 0x0
    "00000000", -- 1173 - 0x495  :    0 - 0x0
    "00000000", -- 1174 - 0x496  :    0 - 0x0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "00000000", -- 1176 - 0x498  :    0 - 0x0
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000000", -- 1186 - 0x4a2  :    0 - 0x0
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00000000", -- 1188 - 0x4a4  :    0 - 0x0
    "00000000", -- 1189 - 0x4a5  :    0 - 0x0
    "00000000", -- 1190 - 0x4a6  :    0 - 0x0
    "00000000", -- 1191 - 0x4a7  :    0 - 0x0
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00000000", -- 1194 - 0x4aa  :    0 - 0x0
    "00000000", -- 1195 - 0x4ab  :    0 - 0x0
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0
    "00000000", -- 1201 - 0x4b1  :    0 - 0x0
    "00000000", -- 1202 - 0x4b2  :    0 - 0x0
    "00000000", -- 1203 - 0x4b3  :    0 - 0x0
    "00000000", -- 1204 - 0x4b4  :    0 - 0x0
    "00000000", -- 1205 - 0x4b5  :    0 - 0x0
    "00000000", -- 1206 - 0x4b6  :    0 - 0x0
    "00000000", -- 1207 - 0x4b7  :    0 - 0x0
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0
    "00000000", -- 1217 - 0x4c1  :    0 - 0x0
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000000", -- 1219 - 0x4c3  :    0 - 0x0
    "00000000", -- 1220 - 0x4c4  :    0 - 0x0
    "00000000", -- 1221 - 0x4c5  :    0 - 0x0
    "00000000", -- 1222 - 0x4c6  :    0 - 0x0
    "00000000", -- 1223 - 0x4c7  :    0 - 0x0
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "00000000", -- 1228 - 0x4cc  :    0 - 0x0
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00000000", -- 1235 - 0x4d3  :    0 - 0x0
    "00000000", -- 1236 - 0x4d4  :    0 - 0x0
    "00000000", -- 1237 - 0x4d5  :    0 - 0x0
    "00000000", -- 1238 - 0x4d6  :    0 - 0x0
    "00000000", -- 1239 - 0x4d7  :    0 - 0x0
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0
    "00000000", -- 1249 - 0x4e1  :    0 - 0x0
    "00000000", -- 1250 - 0x4e2  :    0 - 0x0
    "00000000", -- 1251 - 0x4e3  :    0 - 0x0
    "00000000", -- 1252 - 0x4e4  :    0 - 0x0
    "00000000", -- 1253 - 0x4e5  :    0 - 0x0
    "00000000", -- 1254 - 0x4e6  :    0 - 0x0
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0
    "00000000", -- 1257 - 0x4e9  :    0 - 0x0
    "00000000", -- 1258 - 0x4ea  :    0 - 0x0
    "00000000", -- 1259 - 0x4eb  :    0 - 0x0
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00000000", -- 1261 - 0x4ed  :    0 - 0x0
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0
    "00000000", -- 1265 - 0x4f1  :    0 - 0x0
    "00000000", -- 1266 - 0x4f2  :    0 - 0x0
    "00000000", -- 1267 - 0x4f3  :    0 - 0x0
    "00000000", -- 1268 - 0x4f4  :    0 - 0x0
    "00000000", -- 1269 - 0x4f5  :    0 - 0x0
    "00000000", -- 1270 - 0x4f6  :    0 - 0x0
    "00000000", -- 1271 - 0x4f7  :    0 - 0x0
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0
    "00000000", -- 1281 - 0x501  :    0 - 0x0
    "00000000", -- 1282 - 0x502  :    0 - 0x0
    "00000000", -- 1283 - 0x503  :    0 - 0x0
    "00000000", -- 1284 - 0x504  :    0 - 0x0
    "00000000", -- 1285 - 0x505  :    0 - 0x0
    "00000000", -- 1286 - 0x506  :    0 - 0x0
    "00000000", -- 1287 - 0x507  :    0 - 0x0
    "00000000", -- 1288 - 0x508  :    0 - 0x0
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00000000", -- 1290 - 0x50a  :    0 - 0x0
    "00000000", -- 1291 - 0x50b  :    0 - 0x0
    "00000000", -- 1292 - 0x50c  :    0 - 0x0
    "00000000", -- 1293 - 0x50d  :    0 - 0x0
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00000000", -- 1296 - 0x510  :    0 - 0x0
    "00000000", -- 1297 - 0x511  :    0 - 0x0
    "00000000", -- 1298 - 0x512  :    0 - 0x0
    "00000000", -- 1299 - 0x513  :    0 - 0x0
    "00000000", -- 1300 - 0x514  :    0 - 0x0
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "00000000", -- 1302 - 0x516  :    0 - 0x0
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "00000000", -- 1304 - 0x518  :    0 - 0x0
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "00000000", -- 1306 - 0x51a  :    0 - 0x0
    "00000000", -- 1307 - 0x51b  :    0 - 0x0
    "00000000", -- 1308 - 0x51c  :    0 - 0x0
    "00000000", -- 1309 - 0x51d  :    0 - 0x0
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00000000", -- 1312 - 0x520  :    0 - 0x0
    "00000000", -- 1313 - 0x521  :    0 - 0x0
    "00000000", -- 1314 - 0x522  :    0 - 0x0
    "00000000", -- 1315 - 0x523  :    0 - 0x0
    "00000000", -- 1316 - 0x524  :    0 - 0x0
    "00000000", -- 1317 - 0x525  :    0 - 0x0
    "00000000", -- 1318 - 0x526  :    0 - 0x0
    "00000000", -- 1319 - 0x527  :    0 - 0x0
    "00000000", -- 1320 - 0x528  :    0 - 0x0
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "00000000", -- 1324 - 0x52c  :    0 - 0x0
    "00000000", -- 1325 - 0x52d  :    0 - 0x0
    "00000000", -- 1326 - 0x52e  :    0 - 0x0
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00000000", -- 1328 - 0x530  :    0 - 0x0
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "00000000", -- 1331 - 0x533  :    0 - 0x0
    "00000000", -- 1332 - 0x534  :    0 - 0x0
    "00000000", -- 1333 - 0x535  :    0 - 0x0
    "00000000", -- 1334 - 0x536  :    0 - 0x0
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "00000000", -- 1336 - 0x538  :    0 - 0x0
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "00000000", -- 1338 - 0x53a  :    0 - 0x0
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00000000", -- 1344 - 0x540  :    0 - 0x0
    "00000000", -- 1345 - 0x541  :    0 - 0x0
    "00000000", -- 1346 - 0x542  :    0 - 0x0
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00000000", -- 1349 - 0x545  :    0 - 0x0
    "00000000", -- 1350 - 0x546  :    0 - 0x0
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "00000000", -- 1352 - 0x548  :    0 - 0x0
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "00000000", -- 1354 - 0x54a  :    0 - 0x0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "00000000", -- 1357 - 0x54d  :    0 - 0x0
    "00000000", -- 1358 - 0x54e  :    0 - 0x0
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "00000000", -- 1380 - 0x564  :    0 - 0x0
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "00000000", -- 1386 - 0x56a  :    0 - 0x0
    "00000000", -- 1387 - 0x56b  :    0 - 0x0
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000000", -- 1396 - 0x574  :    0 - 0x0
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "00000000", -- 1408 - 0x580  :    0 - 0x0
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "00000000", -- 1410 - 0x582  :    0 - 0x0
    "00000000", -- 1411 - 0x583  :    0 - 0x0
    "00000000", -- 1412 - 0x584  :    0 - 0x0
    "00000000", -- 1413 - 0x585  :    0 - 0x0
    "00000000", -- 1414 - 0x586  :    0 - 0x0
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00000000", -- 1416 - 0x588  :    0 - 0x0
    "00000000", -- 1417 - 0x589  :    0 - 0x0
    "00000000", -- 1418 - 0x58a  :    0 - 0x0
    "00000000", -- 1419 - 0x58b  :    0 - 0x0
    "00000000", -- 1420 - 0x58c  :    0 - 0x0
    "00000000", -- 1421 - 0x58d  :    0 - 0x0
    "00000000", -- 1422 - 0x58e  :    0 - 0x0
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "00000000", -- 1424 - 0x590  :    0 - 0x0
    "00000000", -- 1425 - 0x591  :    0 - 0x0
    "00000000", -- 1426 - 0x592  :    0 - 0x0
    "00000000", -- 1427 - 0x593  :    0 - 0x0
    "00000000", -- 1428 - 0x594  :    0 - 0x0
    "00000000", -- 1429 - 0x595  :    0 - 0x0
    "00000000", -- 1430 - 0x596  :    0 - 0x0
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00000000", -- 1432 - 0x598  :    0 - 0x0
    "00000000", -- 1433 - 0x599  :    0 - 0x0
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00000000", -- 1435 - 0x59b  :    0 - 0x0
    "00000000", -- 1436 - 0x59c  :    0 - 0x0
    "00000000", -- 1437 - 0x59d  :    0 - 0x0
    "00000000", -- 1438 - 0x59e  :    0 - 0x0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "00000000", -- 1442 - 0x5a2  :    0 - 0x0
    "00000000", -- 1443 - 0x5a3  :    0 - 0x0
    "00000000", -- 1444 - 0x5a4  :    0 - 0x0
    "00000000", -- 1445 - 0x5a5  :    0 - 0x0
    "00000000", -- 1446 - 0x5a6  :    0 - 0x0
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "00000000", -- 1450 - 0x5aa  :    0 - 0x0
    "00000000", -- 1451 - 0x5ab  :    0 - 0x0
    "00000000", -- 1452 - 0x5ac  :    0 - 0x0
    "00000000", -- 1453 - 0x5ad  :    0 - 0x0
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00000000", -- 1461 - 0x5b5  :    0 - 0x0
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "00000000", -- 1466 - 0x5ba  :    0 - 0x0
    "00000000", -- 1467 - 0x5bb  :    0 - 0x0
    "00000000", -- 1468 - 0x5bc  :    0 - 0x0
    "00000000", -- 1469 - 0x5bd  :    0 - 0x0
    "00000000", -- 1470 - 0x5be  :    0 - 0x0
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0
    "00000000", -- 1473 - 0x5c1  :    0 - 0x0
    "00000000", -- 1474 - 0x5c2  :    0 - 0x0
    "00000000", -- 1475 - 0x5c3  :    0 - 0x0
    "00000000", -- 1476 - 0x5c4  :    0 - 0x0
    "00000000", -- 1477 - 0x5c5  :    0 - 0x0
    "00000000", -- 1478 - 0x5c6  :    0 - 0x0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "00000000", -- 1482 - 0x5ca  :    0 - 0x0
    "00000000", -- 1483 - 0x5cb  :    0 - 0x0
    "00000000", -- 1484 - 0x5cc  :    0 - 0x0
    "00000000", -- 1485 - 0x5cd  :    0 - 0x0
    "00000000", -- 1486 - 0x5ce  :    0 - 0x0
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0
    "00000000", -- 1489 - 0x5d1  :    0 - 0x0
    "00000000", -- 1490 - 0x5d2  :    0 - 0x0
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "00000000", -- 1492 - 0x5d4  :    0 - 0x0
    "00000000", -- 1493 - 0x5d5  :    0 - 0x0
    "00000000", -- 1494 - 0x5d6  :    0 - 0x0
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0
    "00000000", -- 1505 - 0x5e1  :    0 - 0x0
    "00000000", -- 1506 - 0x5e2  :    0 - 0x0
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "00000000", -- 1508 - 0x5e4  :    0 - 0x0
    "00000000", -- 1509 - 0x5e5  :    0 - 0x0
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00000000", -- 1514 - 0x5ea  :    0 - 0x0
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "00000000", -- 1516 - 0x5ec  :    0 - 0x0
    "00000000", -- 1517 - 0x5ed  :    0 - 0x0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000000", -- 1542 - 0x606  :    0 - 0x0
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00000000", -- 1544 - 0x608  :    0 - 0x0
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000000", -- 1578 - 0x62a  :    0 - 0x0
    "00000000", -- 1579 - 0x62b  :    0 - 0x0
    "00000000", -- 1580 - 0x62c  :    0 - 0x0
    "00000000", -- 1581 - 0x62d  :    0 - 0x0
    "00000000", -- 1582 - 0x62e  :    0 - 0x0
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "00000000", -- 1584 - 0x630  :    0 - 0x0
    "00000000", -- 1585 - 0x631  :    0 - 0x0
    "00000000", -- 1586 - 0x632  :    0 - 0x0
    "00000000", -- 1587 - 0x633  :    0 - 0x0
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "00000000", -- 1589 - 0x635  :    0 - 0x0
    "00000000", -- 1590 - 0x636  :    0 - 0x0
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00000000", -- 1592 - 0x638  :    0 - 0x0
    "00000000", -- 1593 - 0x639  :    0 - 0x0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "00000000", -- 1596 - 0x63c  :    0 - 0x0
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00000000", -- 1608 - 0x648  :    0 - 0x0
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "00000000", -- 1622 - 0x656  :    0 - 0x0
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00000000", -- 1680 - 0x690  :    0 - 0x0
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00000000", -- 1685 - 0x695  :    0 - 0x0
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00000000", -- 1688 - 0x698  :    0 - 0x0
    "00000000", -- 1689 - 0x699  :    0 - 0x0
    "00000000", -- 1690 - 0x69a  :    0 - 0x0
    "00000000", -- 1691 - 0x69b  :    0 - 0x0
    "00000000", -- 1692 - 0x69c  :    0 - 0x0
    "00000000", -- 1693 - 0x69d  :    0 - 0x0
    "00000000", -- 1694 - 0x69e  :    0 - 0x0
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0
    "00000000", -- 1705 - 0x6a9  :    0 - 0x0
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "00000000", -- 1715 - 0x6b3  :    0 - 0x0
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "00000000", -- 1720 - 0x6b8  :    0 - 0x0
    "00000000", -- 1721 - 0x6b9  :    0 - 0x0
    "00000000", -- 1722 - 0x6ba  :    0 - 0x0
    "00000000", -- 1723 - 0x6bb  :    0 - 0x0
    "00000000", -- 1724 - 0x6bc  :    0 - 0x0
    "00000000", -- 1725 - 0x6bd  :    0 - 0x0
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000000", -- 1734 - 0x6c6  :    0 - 0x0
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "00000000", -- 1738 - 0x6ca  :    0 - 0x0
    "00000000", -- 1739 - 0x6cb  :    0 - 0x0
    "00000000", -- 1740 - 0x6cc  :    0 - 0x0
    "00000000", -- 1741 - 0x6cd  :    0 - 0x0
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0
    "00000000", -- 1753 - 0x6d9  :    0 - 0x0
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "00000000", -- 1755 - 0x6db  :    0 - 0x0
    "00000000", -- 1756 - 0x6dc  :    0 - 0x0
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00000000", -- 1773 - 0x6ed  :    0 - 0x0
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0
    "00000000", -- 1777 - 0x6f1  :    0 - 0x0
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00000000", -- 1779 - 0x6f3  :    0 - 0x0
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "00000000", -- 1781 - 0x6f5  :    0 - 0x0
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "00000000", -- 1784 - 0x6f8  :    0 - 0x0
    "00000000", -- 1785 - 0x6f9  :    0 - 0x0
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "00000000", -- 1787 - 0x6fb  :    0 - 0x0
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "00000000", -- 1789 - 0x6fd  :    0 - 0x0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00000000", -- 1792 - 0x700  :    0 - 0x0
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000000", -- 1816 - 0x718  :    0 - 0x0
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000000", -- 1828 - 0x724  :    0 - 0x0
    "00000000", -- 1829 - 0x725  :    0 - 0x0
    "00000000", -- 1830 - 0x726  :    0 - 0x0
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "00000000", -- 1840 - 0x730  :    0 - 0x0
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "00000000", -- 1845 - 0x735  :    0 - 0x0
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
        ---- Attribute Table 1----
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
