//-   Sprites Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_NOVA_SPR
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table both color planes
      12'h0: dout <= 8'b11111111; //    0 : 255 - 0xff -- Sprite 0x0
      12'h1: dout <= 8'b11111111; //    1 : 255 - 0xff
      12'h2: dout <= 8'b11000000; //    2 : 192 - 0xc0
      12'h3: dout <= 8'b11000000; //    3 : 192 - 0xc0
      12'h4: dout <= 8'b11000000; //    4 : 192 - 0xc0
      12'h5: dout <= 8'b11000000; //    5 : 192 - 0xc0
      12'h6: dout <= 8'b11010101; //    6 : 213 - 0xd5
      12'h7: dout <= 8'b11111111; //    7 : 255 - 0xff
      12'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- plane 1
      12'h9: dout <= 8'b01111111; //    9 : 127 - 0x7f
      12'hA: dout <= 8'b01111111; //   10 : 127 - 0x7f
      12'hB: dout <= 8'b01111111; //   11 : 127 - 0x7f
      12'hC: dout <= 8'b01111111; //   12 : 127 - 0x7f
      12'hD: dout <= 8'b01111111; //   13 : 127 - 0x7f
      12'hE: dout <= 8'b01101010; //   14 : 106 - 0x6a
      12'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      12'h10: dout <= 8'b11111111; //   16 : 255 - 0xff -- Sprite 0x1
      12'h11: dout <= 8'b11111111; //   17 : 255 - 0xff
      12'h12: dout <= 8'b11001110; //   18 : 206 - 0xce
      12'h13: dout <= 8'b11000110; //   19 : 198 - 0xc6
      12'h14: dout <= 8'b11001110; //   20 : 206 - 0xce
      12'h15: dout <= 8'b11000110; //   21 : 198 - 0xc6
      12'h16: dout <= 8'b11101110; //   22 : 238 - 0xee
      12'h17: dout <= 8'b11111111; //   23 : 255 - 0xff
      12'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- plane 1
      12'h19: dout <= 8'b01111011; //   25 : 123 - 0x7b
      12'h1A: dout <= 8'b01110011; //   26 : 115 - 0x73
      12'h1B: dout <= 8'b01111011; //   27 : 123 - 0x7b
      12'h1C: dout <= 8'b01110011; //   28 : 115 - 0x73
      12'h1D: dout <= 8'b01111011; //   29 : 123 - 0x7b
      12'h1E: dout <= 8'b01010011; //   30 :  83 - 0x53
      12'h1F: dout <= 8'b00000000; //   31 :   0 - 0x0
      12'h20: dout <= 8'b11111111; //   32 : 255 - 0xff -- Sprite 0x2
      12'h21: dout <= 8'b11111111; //   33 : 255 - 0xff
      12'h22: dout <= 8'b01110001; //   34 : 113 - 0x71
      12'h23: dout <= 8'b00110011; //   35 :  51 - 0x33
      12'h24: dout <= 8'b01110001; //   36 : 113 - 0x71
      12'h25: dout <= 8'b00110011; //   37 :  51 - 0x33
      12'h26: dout <= 8'b01110101; //   38 : 117 - 0x75
      12'h27: dout <= 8'b11111111; //   39 : 255 - 0xff
      12'h28: dout <= 8'b00000000; //   40 :   0 - 0x0 -- plane 1
      12'h29: dout <= 8'b11011110; //   41 : 222 - 0xde
      12'h2A: dout <= 8'b10011110; //   42 : 158 - 0x9e
      12'h2B: dout <= 8'b11011100; //   43 : 220 - 0xdc
      12'h2C: dout <= 8'b10011110; //   44 : 158 - 0x9e
      12'h2D: dout <= 8'b11011100; //   45 : 220 - 0xdc
      12'h2E: dout <= 8'b10011010; //   46 : 154 - 0x9a
      12'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout <= 8'b11111111; //   48 : 255 - 0xff -- Sprite 0x3
      12'h31: dout <= 8'b11111111; //   49 : 255 - 0xff
      12'h32: dout <= 8'b00000011; //   50 :   3 - 0x3
      12'h33: dout <= 8'b00000001; //   51 :   1 - 0x1
      12'h34: dout <= 8'b00000011; //   52 :   3 - 0x3
      12'h35: dout <= 8'b00000001; //   53 :   1 - 0x1
      12'h36: dout <= 8'b10101011; //   54 : 171 - 0xab
      12'h37: dout <= 8'b11111111; //   55 : 255 - 0xff
      12'h38: dout <= 8'b00000000; //   56 :   0 - 0x0 -- plane 1
      12'h39: dout <= 8'b11111110; //   57 : 254 - 0xfe
      12'h3A: dout <= 8'b11111100; //   58 : 252 - 0xfc
      12'h3B: dout <= 8'b11111110; //   59 : 254 - 0xfe
      12'h3C: dout <= 8'b11111100; //   60 : 252 - 0xfc
      12'h3D: dout <= 8'b11111110; //   61 : 254 - 0xfe
      12'h3E: dout <= 8'b01010100; //   62 :  84 - 0x54
      12'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout <= 8'b11111111; //   64 : 255 - 0xff -- Sprite 0x4
      12'h41: dout <= 8'b11111111; //   65 : 255 - 0xff
      12'h42: dout <= 8'b11100000; //   66 : 224 - 0xe0
      12'h43: dout <= 8'b11000110; //   67 : 198 - 0xc6
      12'h44: dout <= 8'b11000110; //   68 : 198 - 0xc6
      12'h45: dout <= 8'b11110110; //   69 : 246 - 0xf6
      12'h46: dout <= 8'b11110000; //   70 : 240 - 0xf0
      12'h47: dout <= 8'b11110001; //   71 : 241 - 0xf1
      12'h48: dout <= 8'b00000000; //   72 :   0 - 0x0 -- plane 1
      12'h49: dout <= 8'b01111111; //   73 : 127 - 0x7f
      12'h4A: dout <= 8'b01011111; //   74 :  95 - 0x5f
      12'h4B: dout <= 8'b01111001; //   75 : 121 - 0x79
      12'h4C: dout <= 8'b01111001; //   76 : 121 - 0x79
      12'h4D: dout <= 8'b01001001; //   77 :  73 - 0x49
      12'h4E: dout <= 8'b01001111; //   78 :  79 - 0x4f
      12'h4F: dout <= 8'b01001110; //   79 :  78 - 0x4e
      12'h50: dout <= 8'b11000111; //   80 : 199 - 0xc7 -- Sprite 0x5
      12'h51: dout <= 8'b11001111; //   81 : 207 - 0xcf
      12'h52: dout <= 8'b11011111; //   82 : 223 - 0xdf
      12'h53: dout <= 8'b11011111; //   83 : 223 - 0xdf
      12'h54: dout <= 8'b11001110; //   84 : 206 - 0xce
      12'h55: dout <= 8'b11100000; //   85 : 224 - 0xe0
      12'h56: dout <= 8'b11111111; //   86 : 255 - 0xff
      12'h57: dout <= 8'b11111111; //   87 : 255 - 0xff
      12'h58: dout <= 8'b01111000; //   88 : 120 - 0x78 -- plane 1
      12'h59: dout <= 8'b01110000; //   89 : 112 - 0x70
      12'h5A: dout <= 8'b01100000; //   90 :  96 - 0x60
      12'h5B: dout <= 8'b01100000; //   91 :  96 - 0x60
      12'h5C: dout <= 8'b01110001; //   92 : 113 - 0x71
      12'h5D: dout <= 8'b01011111; //   93 :  95 - 0x5f
      12'h5E: dout <= 8'b01111111; //   94 : 127 - 0x7f
      12'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout <= 8'b11111111; //   96 : 255 - 0xff -- Sprite 0x6
      12'h61: dout <= 8'b11111111; //   97 : 255 - 0xff
      12'h62: dout <= 8'b00000111; //   98 :   7 - 0x7
      12'h63: dout <= 8'b01100011; //   99 :  99 - 0x63
      12'h64: dout <= 8'b01100011; //  100 :  99 - 0x63
      12'h65: dout <= 8'b01101111; //  101 : 111 - 0x6f
      12'h66: dout <= 8'b00001111; //  102 :  15 - 0xf
      12'h67: dout <= 8'b10001111; //  103 : 143 - 0x8f
      12'h68: dout <= 8'b00000000; //  104 :   0 - 0x0 -- plane 1
      12'h69: dout <= 8'b11111110; //  105 : 254 - 0xfe
      12'h6A: dout <= 8'b11111010; //  106 : 250 - 0xfa
      12'h6B: dout <= 8'b10011110; //  107 : 158 - 0x9e
      12'h6C: dout <= 8'b10011110; //  108 : 158 - 0x9e
      12'h6D: dout <= 8'b10010010; //  109 : 146 - 0x92
      12'h6E: dout <= 8'b11110010; //  110 : 242 - 0xf2
      12'h6F: dout <= 8'b01110010; //  111 : 114 - 0x72
      12'h70: dout <= 8'b11100011; //  112 : 227 - 0xe3 -- Sprite 0x7
      12'h71: dout <= 8'b11110011; //  113 : 243 - 0xf3
      12'h72: dout <= 8'b11111011; //  114 : 251 - 0xfb
      12'h73: dout <= 8'b11111011; //  115 : 251 - 0xfb
      12'h74: dout <= 8'b01110011; //  116 : 115 - 0x73
      12'h75: dout <= 8'b00000111; //  117 :   7 - 0x7
      12'h76: dout <= 8'b11111111; //  118 : 255 - 0xff
      12'h77: dout <= 8'b11111111; //  119 : 255 - 0xff
      12'h78: dout <= 8'b00011110; //  120 :  30 - 0x1e -- plane 1
      12'h79: dout <= 8'b00001110; //  121 :  14 - 0xe
      12'h7A: dout <= 8'b00000110; //  122 :   6 - 0x6
      12'h7B: dout <= 8'b00000110; //  123 :   6 - 0x6
      12'h7C: dout <= 8'b10001110; //  124 : 142 - 0x8e
      12'h7D: dout <= 8'b11111010; //  125 : 250 - 0xfa
      12'h7E: dout <= 8'b11111110; //  126 : 254 - 0xfe
      12'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout <= 8'b11111111; //  128 : 255 - 0xff -- Sprite 0x8
      12'h81: dout <= 8'b11010101; //  129 : 213 - 0xd5
      12'h82: dout <= 8'b10101010; //  130 : 170 - 0xaa
      12'h83: dout <= 8'b11010101; //  131 : 213 - 0xd5
      12'h84: dout <= 8'b10101010; //  132 : 170 - 0xaa
      12'h85: dout <= 8'b11010101; //  133 : 213 - 0xd5
      12'h86: dout <= 8'b10101010; //  134 : 170 - 0xaa
      12'h87: dout <= 8'b11010101; //  135 : 213 - 0xd5
      12'h88: dout <= 8'b00000000; //  136 :   0 - 0x0 -- plane 1
      12'h89: dout <= 8'b01111111; //  137 : 127 - 0x7f
      12'h8A: dout <= 8'b01011111; //  138 :  95 - 0x5f
      12'h8B: dout <= 8'b01111111; //  139 : 127 - 0x7f
      12'h8C: dout <= 8'b01111111; //  140 : 127 - 0x7f
      12'h8D: dout <= 8'b01111111; //  141 : 127 - 0x7f
      12'h8E: dout <= 8'b01111111; //  142 : 127 - 0x7f
      12'h8F: dout <= 8'b01111111; //  143 : 127 - 0x7f
      12'h90: dout <= 8'b10101010; //  144 : 170 - 0xaa -- Sprite 0x9
      12'h91: dout <= 8'b11010101; //  145 : 213 - 0xd5
      12'h92: dout <= 8'b10101010; //  146 : 170 - 0xaa
      12'h93: dout <= 8'b11010101; //  147 : 213 - 0xd5
      12'h94: dout <= 8'b10101010; //  148 : 170 - 0xaa
      12'h95: dout <= 8'b11110101; //  149 : 245 - 0xf5
      12'h96: dout <= 8'b10101010; //  150 : 170 - 0xaa
      12'h97: dout <= 8'b11111111; //  151 : 255 - 0xff
      12'h98: dout <= 8'b01111111; //  152 : 127 - 0x7f -- plane 1
      12'h99: dout <= 8'b01111111; //  153 : 127 - 0x7f
      12'h9A: dout <= 8'b01111111; //  154 : 127 - 0x7f
      12'h9B: dout <= 8'b01111111; //  155 : 127 - 0x7f
      12'h9C: dout <= 8'b01111111; //  156 : 127 - 0x7f
      12'h9D: dout <= 8'b01011111; //  157 :  95 - 0x5f
      12'h9E: dout <= 8'b01111111; //  158 : 127 - 0x7f
      12'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      12'hA0: dout <= 8'b11111111; //  160 : 255 - 0xff -- Sprite 0xa
      12'hA1: dout <= 8'b01010101; //  161 :  85 - 0x55
      12'hA2: dout <= 8'b10101111; //  162 : 175 - 0xaf
      12'hA3: dout <= 8'b01010101; //  163 :  85 - 0x55
      12'hA4: dout <= 8'b10101011; //  164 : 171 - 0xab
      12'hA5: dout <= 8'b01010101; //  165 :  85 - 0x55
      12'hA6: dout <= 8'b10101011; //  166 : 171 - 0xab
      12'hA7: dout <= 8'b01010101; //  167 :  85 - 0x55
      12'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0 -- plane 1
      12'hA9: dout <= 8'b11111110; //  169 : 254 - 0xfe
      12'hAA: dout <= 8'b11111010; //  170 : 250 - 0xfa
      12'hAB: dout <= 8'b11111110; //  171 : 254 - 0xfe
      12'hAC: dout <= 8'b11111110; //  172 : 254 - 0xfe
      12'hAD: dout <= 8'b11111110; //  173 : 254 - 0xfe
      12'hAE: dout <= 8'b11111110; //  174 : 254 - 0xfe
      12'hAF: dout <= 8'b11111110; //  175 : 254 - 0xfe
      12'hB0: dout <= 8'b10101011; //  176 : 171 - 0xab -- Sprite 0xb
      12'hB1: dout <= 8'b01010101; //  177 :  85 - 0x55
      12'hB2: dout <= 8'b10101011; //  178 : 171 - 0xab
      12'hB3: dout <= 8'b01010101; //  179 :  85 - 0x55
      12'hB4: dout <= 8'b10101011; //  180 : 171 - 0xab
      12'hB5: dout <= 8'b01010101; //  181 :  85 - 0x55
      12'hB6: dout <= 8'b10101011; //  182 : 171 - 0xab
      12'hB7: dout <= 8'b11111111; //  183 : 255 - 0xff
      12'hB8: dout <= 8'b11111110; //  184 : 254 - 0xfe -- plane 1
      12'hB9: dout <= 8'b11111110; //  185 : 254 - 0xfe
      12'hBA: dout <= 8'b11111110; //  186 : 254 - 0xfe
      12'hBB: dout <= 8'b11111110; //  187 : 254 - 0xfe
      12'hBC: dout <= 8'b11111110; //  188 : 254 - 0xfe
      12'hBD: dout <= 8'b11111010; //  189 : 250 - 0xfa
      12'hBE: dout <= 8'b11111110; //  190 : 254 - 0xfe
      12'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout <= 8'b11111111; //  192 : 255 - 0xff -- Sprite 0xc
      12'hC1: dout <= 8'b11010101; //  193 : 213 - 0xd5
      12'hC2: dout <= 8'b10100000; //  194 : 160 - 0xa0
      12'hC3: dout <= 8'b11010000; //  195 : 208 - 0xd0
      12'hC4: dout <= 8'b10001111; //  196 : 143 - 0x8f
      12'hC5: dout <= 8'b11001000; //  197 : 200 - 0xc8
      12'hC6: dout <= 8'b10001000; //  198 : 136 - 0x88
      12'hC7: dout <= 8'b11001000; //  199 : 200 - 0xc8
      12'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0 -- plane 1
      12'hC9: dout <= 8'b00111111; //  201 :  63 - 0x3f
      12'hCA: dout <= 8'b01011111; //  202 :  95 - 0x5f
      12'hCB: dout <= 8'b01101111; //  203 : 111 - 0x6f
      12'hCC: dout <= 8'b01110000; //  204 : 112 - 0x70
      12'hCD: dout <= 8'b01110111; //  205 : 119 - 0x77
      12'hCE: dout <= 8'b01110111; //  206 : 119 - 0x77
      12'hCF: dout <= 8'b01110111; //  207 : 119 - 0x77
      12'hD0: dout <= 8'b10001000; //  208 : 136 - 0x88 -- Sprite 0xd
      12'hD1: dout <= 8'b11001000; //  209 : 200 - 0xc8
      12'hD2: dout <= 8'b10001000; //  210 : 136 - 0x88
      12'hD3: dout <= 8'b11001111; //  211 : 207 - 0xcf
      12'hD4: dout <= 8'b10010000; //  212 : 144 - 0x90
      12'hD5: dout <= 8'b11100000; //  213 : 224 - 0xe0
      12'hD6: dout <= 8'b11101010; //  214 : 234 - 0xea
      12'hD7: dout <= 8'b11111111; //  215 : 255 - 0xff
      12'hD8: dout <= 8'b01110111; //  216 : 119 - 0x77 -- plane 1
      12'hD9: dout <= 8'b01110111; //  217 : 119 - 0x77
      12'hDA: dout <= 8'b01110111; //  218 : 119 - 0x77
      12'hDB: dout <= 8'b01110000; //  219 : 112 - 0x70
      12'hDC: dout <= 8'b01101111; //  220 : 111 - 0x6f
      12'hDD: dout <= 8'b01011111; //  221 :  95 - 0x5f
      12'hDE: dout <= 8'b00010101; //  222 :  21 - 0x15
      12'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      12'hE0: dout <= 8'b11111111; //  224 : 255 - 0xff -- Sprite 0xe
      12'hE1: dout <= 8'b01011011; //  225 :  91 - 0x5b
      12'hE2: dout <= 8'b00000111; //  226 :   7 - 0x7
      12'hE3: dout <= 8'b00001001; //  227 :   9 - 0x9
      12'hE4: dout <= 8'b11110011; //  228 : 243 - 0xf3
      12'hE5: dout <= 8'b00010001; //  229 :  17 - 0x11
      12'hE6: dout <= 8'b00010011; //  230 :  19 - 0x13
      12'hE7: dout <= 8'b00010001; //  231 :  17 - 0x11
      12'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0 -- plane 1
      12'hE9: dout <= 8'b11111100; //  233 : 252 - 0xfc
      12'hEA: dout <= 8'b11111000; //  234 : 248 - 0xf8
      12'hEB: dout <= 8'b11110110; //  235 : 246 - 0xf6
      12'hEC: dout <= 8'b00001100; //  236 :  12 - 0xc
      12'hED: dout <= 8'b11101110; //  237 : 238 - 0xee
      12'hEE: dout <= 8'b11101100; //  238 : 236 - 0xec
      12'hEF: dout <= 8'b11101110; //  239 : 238 - 0xee
      12'hF0: dout <= 8'b00010011; //  240 :  19 - 0x13 -- Sprite 0xf
      12'hF1: dout <= 8'b00010001; //  241 :  17 - 0x11
      12'hF2: dout <= 8'b00010011; //  242 :  19 - 0x13
      12'hF3: dout <= 8'b11110001; //  243 : 241 - 0xf1
      12'hF4: dout <= 8'b00001011; //  244 :  11 - 0xb
      12'hF5: dout <= 8'b00000101; //  245 :   5 - 0x5
      12'hF6: dout <= 8'b10101011; //  246 : 171 - 0xab
      12'hF7: dout <= 8'b11111111; //  247 : 255 - 0xff
      12'hF8: dout <= 8'b11101100; //  248 : 236 - 0xec -- plane 1
      12'hF9: dout <= 8'b11101110; //  249 : 238 - 0xee
      12'hFA: dout <= 8'b11101100; //  250 : 236 - 0xec
      12'hFB: dout <= 8'b00001110; //  251 :  14 - 0xe
      12'hFC: dout <= 8'b11110100; //  252 : 244 - 0xf4
      12'hFD: dout <= 8'b11111010; //  253 : 250 - 0xfa
      12'hFE: dout <= 8'b01010100; //  254 :  84 - 0x54
      12'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout <= 8'b11010000; //  256 : 208 - 0xd0 -- Sprite 0x10
      12'h101: dout <= 8'b10010000; //  257 : 144 - 0x90
      12'h102: dout <= 8'b11011111; //  258 : 223 - 0xdf
      12'h103: dout <= 8'b10011010; //  259 : 154 - 0x9a
      12'h104: dout <= 8'b11010101; //  260 : 213 - 0xd5
      12'h105: dout <= 8'b10011111; //  261 : 159 - 0x9f
      12'h106: dout <= 8'b11010000; //  262 : 208 - 0xd0
      12'h107: dout <= 8'b10010000; //  263 : 144 - 0x90
      12'h108: dout <= 8'b01100000; //  264 :  96 - 0x60 -- plane 1
      12'h109: dout <= 8'b01100000; //  265 :  96 - 0x60
      12'h10A: dout <= 8'b01100000; //  266 :  96 - 0x60
      12'h10B: dout <= 8'b01101111; //  267 : 111 - 0x6f
      12'h10C: dout <= 8'b01101010; //  268 : 106 - 0x6a
      12'h10D: dout <= 8'b01100000; //  269 :  96 - 0x60
      12'h10E: dout <= 8'b01100000; //  270 :  96 - 0x60
      12'h10F: dout <= 8'b01100000; //  271 :  96 - 0x60
      12'h110: dout <= 8'b00001001; //  272 :   9 - 0x9 -- Sprite 0x11
      12'h111: dout <= 8'b00001011; //  273 :  11 - 0xb
      12'h112: dout <= 8'b11111001; //  274 : 249 - 0xf9
      12'h113: dout <= 8'b10101011; //  275 : 171 - 0xab
      12'h114: dout <= 8'b01011001; //  276 :  89 - 0x59
      12'h115: dout <= 8'b11111011; //  277 : 251 - 0xfb
      12'h116: dout <= 8'b00001001; //  278 :   9 - 0x9
      12'h117: dout <= 8'b00001011; //  279 :  11 - 0xb
      12'h118: dout <= 8'b00000110; //  280 :   6 - 0x6 -- plane 1
      12'h119: dout <= 8'b00000100; //  281 :   4 - 0x4
      12'h11A: dout <= 8'b00000110; //  282 :   6 - 0x6
      12'h11B: dout <= 8'b11110100; //  283 : 244 - 0xf4
      12'h11C: dout <= 8'b10100110; //  284 : 166 - 0xa6
      12'h11D: dout <= 8'b00000100; //  285 :   4 - 0x4
      12'h11E: dout <= 8'b00000110; //  286 :   6 - 0x6
      12'h11F: dout <= 8'b00000100; //  287 :   4 - 0x4
      12'h120: dout <= 8'b00011000; //  288 :  24 - 0x18 -- Sprite 0x12
      12'h121: dout <= 8'b00010100; //  289 :  20 - 0x14
      12'h122: dout <= 8'b00010100; //  290 :  20 - 0x14
      12'h123: dout <= 8'b00111010; //  291 :  58 - 0x3a
      12'h124: dout <= 8'b00111010; //  292 :  58 - 0x3a
      12'h125: dout <= 8'b01111010; //  293 : 122 - 0x7a
      12'h126: dout <= 8'b01111010; //  294 : 122 - 0x7a
      12'h127: dout <= 8'b01111010; //  295 : 122 - 0x7a
      12'h128: dout <= 8'b00000000; //  296 :   0 - 0x0 -- plane 1
      12'h129: dout <= 8'b00001000; //  297 :   8 - 0x8
      12'h12A: dout <= 8'b00001000; //  298 :   8 - 0x8
      12'h12B: dout <= 8'b00011100; //  299 :  28 - 0x1c
      12'h12C: dout <= 8'b00011100; //  300 :  28 - 0x1c
      12'h12D: dout <= 8'b00111100; //  301 :  60 - 0x3c
      12'h12E: dout <= 8'b00111100; //  302 :  60 - 0x3c
      12'h12F: dout <= 8'b00111100; //  303 :  60 - 0x3c
      12'h130: dout <= 8'b11111011; //  304 : 251 - 0xfb -- Sprite 0x13
      12'h131: dout <= 8'b11111101; //  305 : 253 - 0xfd
      12'h132: dout <= 8'b11111101; //  306 : 253 - 0xfd
      12'h133: dout <= 8'b11111101; //  307 : 253 - 0xfd
      12'h134: dout <= 8'b11111101; //  308 : 253 - 0xfd
      12'h135: dout <= 8'b11111101; //  309 : 253 - 0xfd
      12'h136: dout <= 8'b10000001; //  310 : 129 - 0x81
      12'h137: dout <= 8'b11111111; //  311 : 255 - 0xff
      12'h138: dout <= 8'b00111100; //  312 :  60 - 0x3c -- plane 1
      12'h139: dout <= 8'b01111110; //  313 : 126 - 0x7e
      12'h13A: dout <= 8'b01111110; //  314 : 126 - 0x7e
      12'h13B: dout <= 8'b01111110; //  315 : 126 - 0x7e
      12'h13C: dout <= 8'b01111110; //  316 : 126 - 0x7e
      12'h13D: dout <= 8'b01111110; //  317 : 126 - 0x7e
      12'h13E: dout <= 8'b01111110; //  318 : 126 - 0x7e
      12'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x14
      12'h141: dout <= 8'b00000111; //  321 :   7 - 0x7
      12'h142: dout <= 8'b00000010; //  322 :   2 - 0x2
      12'h143: dout <= 8'b00000100; //  323 :   4 - 0x4
      12'h144: dout <= 8'b00000011; //  324 :   3 - 0x3
      12'h145: dout <= 8'b00000011; //  325 :   3 - 0x3
      12'h146: dout <= 8'b00001101; //  326 :  13 - 0xd
      12'h147: dout <= 8'b00010111; //  327 :  23 - 0x17
      12'h148: dout <= 8'b00000000; //  328 :   0 - 0x0 -- plane 1
      12'h149: dout <= 8'b00000000; //  329 :   0 - 0x0
      12'h14A: dout <= 8'b00000101; //  330 :   5 - 0x5
      12'h14B: dout <= 8'b00000011; //  331 :   3 - 0x3
      12'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      12'h14D: dout <= 8'b00000000; //  333 :   0 - 0x0
      12'h14E: dout <= 8'b00000010; //  334 :   2 - 0x2
      12'h14F: dout <= 8'b00001111; //  335 :  15 - 0xf
      12'h150: dout <= 8'b00101111; //  336 :  47 - 0x2f -- Sprite 0x15
      12'h151: dout <= 8'b01001111; //  337 :  79 - 0x4f
      12'h152: dout <= 8'b01001111; //  338 :  79 - 0x4f
      12'h153: dout <= 8'b01001111; //  339 :  79 - 0x4f
      12'h154: dout <= 8'b01001111; //  340 :  79 - 0x4f
      12'h155: dout <= 8'b00100111; //  341 :  39 - 0x27
      12'h156: dout <= 8'b00010000; //  342 :  16 - 0x10
      12'h157: dout <= 8'b00001111; //  343 :  15 - 0xf
      12'h158: dout <= 8'b00011100; //  344 :  28 - 0x1c -- plane 1
      12'h159: dout <= 8'b00111010; //  345 :  58 - 0x3a
      12'h15A: dout <= 8'b00111100; //  346 :  60 - 0x3c
      12'h15B: dout <= 8'b00111111; //  347 :  63 - 0x3f
      12'h15C: dout <= 8'b00111000; //  348 :  56 - 0x38
      12'h15D: dout <= 8'b00011110; //  349 :  30 - 0x1e
      12'h15E: dout <= 8'b00001111; //  350 :  15 - 0xf
      12'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x16
      12'h161: dout <= 8'b11100000; //  353 : 224 - 0xe0
      12'h162: dout <= 8'b10100000; //  354 : 160 - 0xa0
      12'h163: dout <= 8'b00100000; //  355 :  32 - 0x20
      12'h164: dout <= 8'b11000000; //  356 : 192 - 0xc0
      12'h165: dout <= 8'b01000000; //  357 :  64 - 0x40
      12'h166: dout <= 8'b00110000; //  358 :  48 - 0x30
      12'h167: dout <= 8'b11101000; //  359 : 232 - 0xe8
      12'h168: dout <= 8'b00000000; //  360 :   0 - 0x0 -- plane 1
      12'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      12'h16A: dout <= 8'b01000000; //  362 :  64 - 0x40
      12'h16B: dout <= 8'b11000000; //  363 : 192 - 0xc0
      12'h16C: dout <= 8'b00000000; //  364 :   0 - 0x0
      12'h16D: dout <= 8'b10000000; //  365 : 128 - 0x80
      12'h16E: dout <= 8'b11000000; //  366 : 192 - 0xc0
      12'h16F: dout <= 8'b01110000; //  367 : 112 - 0x70
      12'h170: dout <= 8'b11110100; //  368 : 244 - 0xf4 -- Sprite 0x17
      12'h171: dout <= 8'b11110010; //  369 : 242 - 0xf2
      12'h172: dout <= 8'b11110010; //  370 : 242 - 0xf2
      12'h173: dout <= 8'b11110010; //  371 : 242 - 0xf2
      12'h174: dout <= 8'b11110010; //  372 : 242 - 0xf2
      12'h175: dout <= 8'b11100100; //  373 : 228 - 0xe4
      12'h176: dout <= 8'b00001000; //  374 :   8 - 0x8
      12'h177: dout <= 8'b11110000; //  375 : 240 - 0xf0
      12'h178: dout <= 8'b00011000; //  376 :  24 - 0x18 -- plane 1
      12'h179: dout <= 8'b11111100; //  377 : 252 - 0xfc
      12'h17A: dout <= 8'b00111100; //  378 :  60 - 0x3c
      12'h17B: dout <= 8'b01011100; //  379 :  92 - 0x5c
      12'h17C: dout <= 8'b00111100; //  380 :  60 - 0x3c
      12'h17D: dout <= 8'b11111000; //  381 : 248 - 0xf8
      12'h17E: dout <= 8'b11110000; //  382 : 240 - 0xf0
      12'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      12'h180: dout <= 8'b00111111; //  384 :  63 - 0x3f -- Sprite 0x18
      12'h181: dout <= 8'b01000000; //  385 :  64 - 0x40
      12'h182: dout <= 8'b01000000; //  386 :  64 - 0x40
      12'h183: dout <= 8'b10000000; //  387 : 128 - 0x80
      12'h184: dout <= 8'b10000000; //  388 : 128 - 0x80
      12'h185: dout <= 8'b01111111; //  389 : 127 - 0x7f
      12'h186: dout <= 8'b00000001; //  390 :   1 - 0x1
      12'h187: dout <= 8'b01111111; //  391 : 127 - 0x7f
      12'h188: dout <= 8'b00000000; //  392 :   0 - 0x0 -- plane 1
      12'h189: dout <= 8'b00111111; //  393 :  63 - 0x3f
      12'h18A: dout <= 8'b00111111; //  394 :  63 - 0x3f
      12'h18B: dout <= 8'b01111111; //  395 : 127 - 0x7f
      12'h18C: dout <= 8'b01111111; //  396 : 127 - 0x7f
      12'h18D: dout <= 8'b00000000; //  397 :   0 - 0x0
      12'h18E: dout <= 8'b00000000; //  398 :   0 - 0x0
      12'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      12'h190: dout <= 8'b11111100; //  400 : 252 - 0xfc -- Sprite 0x19
      12'h191: dout <= 8'b00000010; //  401 :   2 - 0x2
      12'h192: dout <= 8'b00000010; //  402 :   2 - 0x2
      12'h193: dout <= 8'b00000001; //  403 :   1 - 0x1
      12'h194: dout <= 8'b00000001; //  404 :   1 - 0x1
      12'h195: dout <= 8'b11111110; //  405 : 254 - 0xfe
      12'h196: dout <= 8'b10000000; //  406 : 128 - 0x80
      12'h197: dout <= 8'b11111110; //  407 : 254 - 0xfe
      12'h198: dout <= 8'b00000000; //  408 :   0 - 0x0 -- plane 1
      12'h199: dout <= 8'b11111100; //  409 : 252 - 0xfc
      12'h19A: dout <= 8'b11111100; //  410 : 252 - 0xfc
      12'h19B: dout <= 8'b11111110; //  411 : 254 - 0xfe
      12'h19C: dout <= 8'b11111110; //  412 : 254 - 0xfe
      12'h19D: dout <= 8'b00000000; //  413 :   0 - 0x0
      12'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      12'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout <= 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x1a
      12'h1A1: dout <= 8'b00000000; //  417 :   0 - 0x0
      12'h1A2: dout <= 8'b00111111; //  418 :  63 - 0x3f
      12'h1A3: dout <= 8'b01000000; //  419 :  64 - 0x40
      12'h1A4: dout <= 8'b01000000; //  420 :  64 - 0x40
      12'h1A5: dout <= 8'b10000000; //  421 : 128 - 0x80
      12'h1A6: dout <= 8'b10000000; //  422 : 128 - 0x80
      12'h1A7: dout <= 8'b01111111; //  423 : 127 - 0x7f
      12'h1A8: dout <= 8'b00000000; //  424 :   0 - 0x0 -- plane 1
      12'h1A9: dout <= 8'b00000000; //  425 :   0 - 0x0
      12'h1AA: dout <= 8'b00000000; //  426 :   0 - 0x0
      12'h1AB: dout <= 8'b00111111; //  427 :  63 - 0x3f
      12'h1AC: dout <= 8'b00111111; //  428 :  63 - 0x3f
      12'h1AD: dout <= 8'b01111111; //  429 : 127 - 0x7f
      12'h1AE: dout <= 8'b01111111; //  430 : 127 - 0x7f
      12'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      12'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x1b
      12'h1B1: dout <= 8'b00000000; //  433 :   0 - 0x0
      12'h1B2: dout <= 8'b11111100; //  434 : 252 - 0xfc
      12'h1B3: dout <= 8'b00000010; //  435 :   2 - 0x2
      12'h1B4: dout <= 8'b00000010; //  436 :   2 - 0x2
      12'h1B5: dout <= 8'b00000001; //  437 :   1 - 0x1
      12'h1B6: dout <= 8'b00000001; //  438 :   1 - 0x1
      12'h1B7: dout <= 8'b11111110; //  439 : 254 - 0xfe
      12'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0 -- plane 1
      12'h1B9: dout <= 8'b00000000; //  441 :   0 - 0x0
      12'h1BA: dout <= 8'b00000000; //  442 :   0 - 0x0
      12'h1BB: dout <= 8'b11111100; //  443 : 252 - 0xfc
      12'h1BC: dout <= 8'b11111100; //  444 : 252 - 0xfc
      12'h1BD: dout <= 8'b11111110; //  445 : 254 - 0xfe
      12'h1BE: dout <= 8'b11111110; //  446 : 254 - 0xfe
      12'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout <= 8'b01111111; //  448 : 127 - 0x7f -- Sprite 0x1c
      12'h1C1: dout <= 8'b10000000; //  449 : 128 - 0x80
      12'h1C2: dout <= 8'b10000000; //  450 : 128 - 0x80
      12'h1C3: dout <= 8'b10000000; //  451 : 128 - 0x80
      12'h1C4: dout <= 8'b10011011; //  452 : 155 - 0x9b
      12'h1C5: dout <= 8'b10100100; //  453 : 164 - 0xa4
      12'h1C6: dout <= 8'b10100110; //  454 : 166 - 0xa6
      12'h1C7: dout <= 8'b10000000; //  455 : 128 - 0x80
      12'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0 -- plane 1
      12'h1C9: dout <= 8'b01111111; //  457 : 127 - 0x7f
      12'h1CA: dout <= 8'b01111111; //  458 : 127 - 0x7f
      12'h1CB: dout <= 8'b01111111; //  459 : 127 - 0x7f
      12'h1CC: dout <= 8'b01100100; //  460 : 100 - 0x64
      12'h1CD: dout <= 8'b01011011; //  461 :  91 - 0x5b
      12'h1CE: dout <= 8'b01011001; //  462 :  89 - 0x59
      12'h1CF: dout <= 8'b01111111; //  463 : 127 - 0x7f
      12'h1D0: dout <= 8'b10000000; //  464 : 128 - 0x80 -- Sprite 0x1d
      12'h1D1: dout <= 8'b01111111; //  465 : 127 - 0x7f
      12'h1D2: dout <= 8'b00000010; //  466 :   2 - 0x2
      12'h1D3: dout <= 8'b00000010; //  467 :   2 - 0x2
      12'h1D4: dout <= 8'b00000010; //  468 :   2 - 0x2
      12'h1D5: dout <= 8'b00000010; //  469 :   2 - 0x2
      12'h1D6: dout <= 8'b00000010; //  470 :   2 - 0x2
      12'h1D7: dout <= 8'b00001111; //  471 :  15 - 0xf
      12'h1D8: dout <= 8'b01111111; //  472 : 127 - 0x7f -- plane 1
      12'h1D9: dout <= 8'b00000000; //  473 :   0 - 0x0
      12'h1DA: dout <= 8'b00000001; //  474 :   1 - 0x1
      12'h1DB: dout <= 8'b00000001; //  475 :   1 - 0x1
      12'h1DC: dout <= 8'b00000001; //  476 :   1 - 0x1
      12'h1DD: dout <= 8'b00000001; //  477 :   1 - 0x1
      12'h1DE: dout <= 8'b00000001; //  478 :   1 - 0x1
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b11111110; //  480 : 254 - 0xfe -- Sprite 0x1e
      12'h1E1: dout <= 8'b00000001; //  481 :   1 - 0x1
      12'h1E2: dout <= 8'b00000001; //  482 :   1 - 0x1
      12'h1E3: dout <= 8'b00000001; //  483 :   1 - 0x1
      12'h1E4: dout <= 8'b01000001; //  484 :  65 - 0x41
      12'h1E5: dout <= 8'b11110101; //  485 : 245 - 0xf5
      12'h1E6: dout <= 8'b00011101; //  486 :  29 - 0x1d
      12'h1E7: dout <= 8'b00000001; //  487 :   1 - 0x1
      12'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0 -- plane 1
      12'h1E9: dout <= 8'b11111110; //  489 : 254 - 0xfe
      12'h1EA: dout <= 8'b11111110; //  490 : 254 - 0xfe
      12'h1EB: dout <= 8'b11111110; //  491 : 254 - 0xfe
      12'h1EC: dout <= 8'b10111110; //  492 : 190 - 0xbe
      12'h1ED: dout <= 8'b00001010; //  493 :  10 - 0xa
      12'h1EE: dout <= 8'b11100010; //  494 : 226 - 0xe2
      12'h1EF: dout <= 8'b11111110; //  495 : 254 - 0xfe
      12'h1F0: dout <= 8'b00000001; //  496 :   1 - 0x1 -- Sprite 0x1f
      12'h1F1: dout <= 8'b11111110; //  497 : 254 - 0xfe
      12'h1F2: dout <= 8'b01000000; //  498 :  64 - 0x40
      12'h1F3: dout <= 8'b01000000; //  499 :  64 - 0x40
      12'h1F4: dout <= 8'b01000000; //  500 :  64 - 0x40
      12'h1F5: dout <= 8'b01000000; //  501 :  64 - 0x40
      12'h1F6: dout <= 8'b01000000; //  502 :  64 - 0x40
      12'h1F7: dout <= 8'b11110000; //  503 : 240 - 0xf0
      12'h1F8: dout <= 8'b11111110; //  504 : 254 - 0xfe -- plane 1
      12'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout <= 8'b10000000; //  506 : 128 - 0x80
      12'h1FB: dout <= 8'b10000000; //  507 : 128 - 0x80
      12'h1FC: dout <= 8'b10000000; //  508 : 128 - 0x80
      12'h1FD: dout <= 8'b10000000; //  509 : 128 - 0x80
      12'h1FE: dout <= 8'b10000000; //  510 : 128 - 0x80
      12'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout <= 8'b00000111; //  512 :   7 - 0x7 -- Sprite 0x20
      12'h201: dout <= 8'b00011111; //  513 :  31 - 0x1f
      12'h202: dout <= 8'b00111111; //  514 :  63 - 0x3f
      12'h203: dout <= 8'b01111111; //  515 : 127 - 0x7f
      12'h204: dout <= 8'b01111111; //  516 : 127 - 0x7f
      12'h205: dout <= 8'b11111111; //  517 : 255 - 0xff
      12'h206: dout <= 8'b11111111; //  518 : 255 - 0xff
      12'h207: dout <= 8'b11111111; //  519 : 255 - 0xff
      12'h208: dout <= 8'b00000000; //  520 :   0 - 0x0 -- plane 1
      12'h209: dout <= 8'b00000000; //  521 :   0 - 0x0
      12'h20A: dout <= 8'b00000000; //  522 :   0 - 0x0
      12'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      12'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      12'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      12'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      12'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout <= 8'b11100000; //  528 : 224 - 0xe0 -- Sprite 0x21
      12'h211: dout <= 8'b11111000; //  529 : 248 - 0xf8
      12'h212: dout <= 8'b11111100; //  530 : 252 - 0xfc
      12'h213: dout <= 8'b11111110; //  531 : 254 - 0xfe
      12'h214: dout <= 8'b11111110; //  532 : 254 - 0xfe
      12'h215: dout <= 8'b11111111; //  533 : 255 - 0xff
      12'h216: dout <= 8'b11111111; //  534 : 255 - 0xff
      12'h217: dout <= 8'b11111111; //  535 : 255 - 0xff
      12'h218: dout <= 8'b00000000; //  536 :   0 - 0x0 -- plane 1
      12'h219: dout <= 8'b00000000; //  537 :   0 - 0x0
      12'h21A: dout <= 8'b00000000; //  538 :   0 - 0x0
      12'h21B: dout <= 8'b00000000; //  539 :   0 - 0x0
      12'h21C: dout <= 8'b00000000; //  540 :   0 - 0x0
      12'h21D: dout <= 8'b00000000; //  541 :   0 - 0x0
      12'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      12'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout <= 8'b00000111; //  544 :   7 - 0x7 -- Sprite 0x22
      12'h221: dout <= 8'b00011111; //  545 :  31 - 0x1f
      12'h222: dout <= 8'b00111111; //  546 :  63 - 0x3f
      12'h223: dout <= 8'b01111111; //  547 : 127 - 0x7f
      12'h224: dout <= 8'b01111111; //  548 : 127 - 0x7f
      12'h225: dout <= 8'b11111111; //  549 : 255 - 0xff
      12'h226: dout <= 8'b11111111; //  550 : 255 - 0xff
      12'h227: dout <= 8'b11111111; //  551 : 255 - 0xff
      12'h228: dout <= 8'b00000000; //  552 :   0 - 0x0 -- plane 1
      12'h229: dout <= 8'b00000000; //  553 :   0 - 0x0
      12'h22A: dout <= 8'b00011000; //  554 :  24 - 0x18
      12'h22B: dout <= 8'b00010000; //  555 :  16 - 0x10
      12'h22C: dout <= 8'b00011010; //  556 :  26 - 0x1a
      12'h22D: dout <= 8'b00010001; //  557 :  17 - 0x11
      12'h22E: dout <= 8'b00011010; //  558 :  26 - 0x1a
      12'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout <= 8'b11100000; //  560 : 224 - 0xe0 -- Sprite 0x23
      12'h231: dout <= 8'b11111000; //  561 : 248 - 0xf8
      12'h232: dout <= 8'b11111100; //  562 : 252 - 0xfc
      12'h233: dout <= 8'b11111110; //  563 : 254 - 0xfe
      12'h234: dout <= 8'b11111110; //  564 : 254 - 0xfe
      12'h235: dout <= 8'b11111111; //  565 : 255 - 0xff
      12'h236: dout <= 8'b11111111; //  566 : 255 - 0xff
      12'h237: dout <= 8'b11111111; //  567 : 255 - 0xff
      12'h238: dout <= 8'b00000000; //  568 :   0 - 0x0 -- plane 1
      12'h239: dout <= 8'b00000000; //  569 :   0 - 0x0
      12'h23A: dout <= 8'b00000000; //  570 :   0 - 0x0
      12'h23B: dout <= 8'b00101000; //  571 :  40 - 0x28
      12'h23C: dout <= 8'b10001100; //  572 : 140 - 0x8c
      12'h23D: dout <= 8'b00101000; //  573 :  40 - 0x28
      12'h23E: dout <= 8'b10101100; //  574 : 172 - 0xac
      12'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x24
      12'h241: dout <= 8'b00000000; //  577 :   0 - 0x0
      12'h242: dout <= 8'b00000000; //  578 :   0 - 0x0
      12'h243: dout <= 8'b00000000; //  579 :   0 - 0x0
      12'h244: dout <= 8'b00000000; //  580 :   0 - 0x0
      12'h245: dout <= 8'b00000000; //  581 :   0 - 0x0
      12'h246: dout <= 8'b00000000; //  582 :   0 - 0x0
      12'h247: dout <= 8'b00000000; //  583 :   0 - 0x0
      12'h248: dout <= 8'b00000000; //  584 :   0 - 0x0 -- plane 1
      12'h249: dout <= 8'b00000000; //  585 :   0 - 0x0
      12'h24A: dout <= 8'b00000000; //  586 :   0 - 0x0
      12'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      12'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      12'h24D: dout <= 8'b00000000; //  589 :   0 - 0x0
      12'h24E: dout <= 8'b00000000; //  590 :   0 - 0x0
      12'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout <= 8'b00101111; //  592 :  47 - 0x2f -- Sprite 0x25
      12'h251: dout <= 8'b01001111; //  593 :  79 - 0x4f
      12'h252: dout <= 8'b01001111; //  594 :  79 - 0x4f
      12'h253: dout <= 8'b01001111; //  595 :  79 - 0x4f
      12'h254: dout <= 8'b01001111; //  596 :  79 - 0x4f
      12'h255: dout <= 8'b00100111; //  597 :  39 - 0x27
      12'h256: dout <= 8'b00010000; //  598 :  16 - 0x10
      12'h257: dout <= 8'b00001111; //  599 :  15 - 0xf
      12'h258: dout <= 8'b00011100; //  600 :  28 - 0x1c -- plane 1
      12'h259: dout <= 8'b00111001; //  601 :  57 - 0x39
      12'h25A: dout <= 8'b00111111; //  602 :  63 - 0x3f
      12'h25B: dout <= 8'b00111110; //  603 :  62 - 0x3e
      12'h25C: dout <= 8'b00111111; //  604 :  63 - 0x3f
      12'h25D: dout <= 8'b00011110; //  605 :  30 - 0x1e
      12'h25E: dout <= 8'b00001111; //  606 :  15 - 0xf
      12'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout <= 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x26
      12'h261: dout <= 8'b11100000; //  609 : 224 - 0xe0
      12'h262: dout <= 8'b10100000; //  610 : 160 - 0xa0
      12'h263: dout <= 8'b00100000; //  611 :  32 - 0x20
      12'h264: dout <= 8'b11000000; //  612 : 192 - 0xc0
      12'h265: dout <= 8'b01000000; //  613 :  64 - 0x40
      12'h266: dout <= 8'b00110000; //  614 :  48 - 0x30
      12'h267: dout <= 8'b11101000; //  615 : 232 - 0xe8
      12'h268: dout <= 8'b00000000; //  616 :   0 - 0x0 -- plane 1
      12'h269: dout <= 8'b00000000; //  617 :   0 - 0x0
      12'h26A: dout <= 8'b01000000; //  618 :  64 - 0x40
      12'h26B: dout <= 8'b11000000; //  619 : 192 - 0xc0
      12'h26C: dout <= 8'b00000000; //  620 :   0 - 0x0
      12'h26D: dout <= 8'b10000000; //  621 : 128 - 0x80
      12'h26E: dout <= 8'b11000000; //  622 : 192 - 0xc0
      12'h26F: dout <= 8'b11110000; //  623 : 240 - 0xf0
      12'h270: dout <= 8'b11110100; //  624 : 244 - 0xf4 -- Sprite 0x27
      12'h271: dout <= 8'b11110010; //  625 : 242 - 0xf2
      12'h272: dout <= 8'b11110010; //  626 : 242 - 0xf2
      12'h273: dout <= 8'b11110010; //  627 : 242 - 0xf2
      12'h274: dout <= 8'b11110010; //  628 : 242 - 0xf2
      12'h275: dout <= 8'b11100100; //  629 : 228 - 0xe4
      12'h276: dout <= 8'b00001000; //  630 :   8 - 0x8
      12'h277: dout <= 8'b11110000; //  631 : 240 - 0xf0
      12'h278: dout <= 8'b00111000; //  632 :  56 - 0x38 -- plane 1
      12'h279: dout <= 8'b10011100; //  633 : 156 - 0x9c
      12'h27A: dout <= 8'b10011100; //  634 : 156 - 0x9c
      12'h27B: dout <= 8'b00111100; //  635 :  60 - 0x3c
      12'h27C: dout <= 8'b11111100; //  636 : 252 - 0xfc
      12'h27D: dout <= 8'b01111000; //  637 : 120 - 0x78
      12'h27E: dout <= 8'b11110000; //  638 : 240 - 0xf0
      12'h27F: dout <= 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout <= 8'b11111111; //  640 : 255 - 0xff -- Sprite 0x28
      12'h281: dout <= 8'b11010101; //  641 : 213 - 0xd5
      12'h282: dout <= 8'b10100011; //  642 : 163 - 0xa3
      12'h283: dout <= 8'b11010111; //  643 : 215 - 0xd7
      12'h284: dout <= 8'b10001111; //  644 : 143 - 0x8f
      12'h285: dout <= 8'b11001111; //  645 : 207 - 0xcf
      12'h286: dout <= 8'b10001011; //  646 : 139 - 0x8b
      12'h287: dout <= 8'b11001011; //  647 : 203 - 0xcb
      12'h288: dout <= 8'b00000000; //  648 :   0 - 0x0 -- plane 1
      12'h289: dout <= 8'b00111110; //  649 :  62 - 0x3e
      12'h28A: dout <= 8'b01011101; //  650 :  93 - 0x5d
      12'h28B: dout <= 8'b01101011; //  651 : 107 - 0x6b
      12'h28C: dout <= 8'b01110101; //  652 : 117 - 0x75
      12'h28D: dout <= 8'b01110001; //  653 : 113 - 0x71
      12'h28E: dout <= 8'b01110101; //  654 : 117 - 0x75
      12'h28F: dout <= 8'b01110100; //  655 : 116 - 0x74
      12'h290: dout <= 8'b10001111; //  656 : 143 - 0x8f -- Sprite 0x29
      12'h291: dout <= 8'b11001111; //  657 : 207 - 0xcf
      12'h292: dout <= 8'b10001111; //  658 : 143 - 0x8f
      12'h293: dout <= 8'b11001111; //  659 : 207 - 0xcf
      12'h294: dout <= 8'b10010000; //  660 : 144 - 0x90
      12'h295: dout <= 8'b11100000; //  661 : 224 - 0xe0
      12'h296: dout <= 8'b11101010; //  662 : 234 - 0xea
      12'h297: dout <= 8'b11111111; //  663 : 255 - 0xff
      12'h298: dout <= 8'b01110000; //  664 : 112 - 0x70 -- plane 1
      12'h299: dout <= 8'b01110111; //  665 : 119 - 0x77
      12'h29A: dout <= 8'b01110111; //  666 : 119 - 0x77
      12'h29B: dout <= 8'b01110000; //  667 : 112 - 0x70
      12'h29C: dout <= 8'b01101111; //  668 : 111 - 0x6f
      12'h29D: dout <= 8'b01011111; //  669 :  95 - 0x5f
      12'h29E: dout <= 8'b00010101; //  670 :  21 - 0x15
      12'h29F: dout <= 8'b00000000; //  671 :   0 - 0x0
      12'h2A0: dout <= 8'b11111111; //  672 : 255 - 0xff -- Sprite 0x2a
      12'h2A1: dout <= 8'b11011011; //  673 : 219 - 0xdb
      12'h2A2: dout <= 8'b11000111; //  674 : 199 - 0xc7
      12'h2A3: dout <= 8'b11101001; //  675 : 233 - 0xe9
      12'h2A4: dout <= 8'b11110011; //  676 : 243 - 0xf3
      12'h2A5: dout <= 8'b11110001; //  677 : 241 - 0xf1
      12'h2A6: dout <= 8'b11010011; //  678 : 211 - 0xd3
      12'h2A7: dout <= 8'b11010001; //  679 : 209 - 0xd1
      12'h2A8: dout <= 8'b00000000; //  680 :   0 - 0x0 -- plane 1
      12'h2A9: dout <= 8'b01111100; //  681 : 124 - 0x7c
      12'h2AA: dout <= 8'b10111000; //  682 : 184 - 0xb8
      12'h2AB: dout <= 8'b11010110; //  683 : 214 - 0xd6
      12'h2AC: dout <= 8'b10101100; //  684 : 172 - 0xac
      12'h2AD: dout <= 8'b10001110; //  685 : 142 - 0x8e
      12'h2AE: dout <= 8'b10101100; //  686 : 172 - 0xac
      12'h2AF: dout <= 8'b00101110; //  687 :  46 - 0x2e
      12'h2B0: dout <= 8'b11110011; //  688 : 243 - 0xf3 -- Sprite 0x2b
      12'h2B1: dout <= 8'b11110001; //  689 : 241 - 0xf1
      12'h2B2: dout <= 8'b11110011; //  690 : 243 - 0xf3
      12'h2B3: dout <= 8'b11110001; //  691 : 241 - 0xf1
      12'h2B4: dout <= 8'b00001011; //  692 :  11 - 0xb
      12'h2B5: dout <= 8'b00000101; //  693 :   5 - 0x5
      12'h2B6: dout <= 8'b10101011; //  694 : 171 - 0xab
      12'h2B7: dout <= 8'b11111111; //  695 : 255 - 0xff
      12'h2B8: dout <= 8'b00001100; //  696 :  12 - 0xc -- plane 1
      12'h2B9: dout <= 8'b11101110; //  697 : 238 - 0xee
      12'h2BA: dout <= 8'b11101100; //  698 : 236 - 0xec
      12'h2BB: dout <= 8'b00001110; //  699 :  14 - 0xe
      12'h2BC: dout <= 8'b11110100; //  700 : 244 - 0xf4
      12'h2BD: dout <= 8'b11111010; //  701 : 250 - 0xfa
      12'h2BE: dout <= 8'b01010100; //  702 :  84 - 0x54
      12'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout <= 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x2c
      12'h2C1: dout <= 8'b00000000; //  705 :   0 - 0x0
      12'h2C2: dout <= 8'b00000000; //  706 :   0 - 0x0
      12'h2C3: dout <= 8'b00000000; //  707 :   0 - 0x0
      12'h2C4: dout <= 8'b00000000; //  708 :   0 - 0x0
      12'h2C5: dout <= 8'b00000000; //  709 :   0 - 0x0
      12'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      12'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0 -- plane 1
      12'h2C9: dout <= 8'b00000000; //  713 :   0 - 0x0
      12'h2CA: dout <= 8'b00000000; //  714 :   0 - 0x0
      12'h2CB: dout <= 8'b00000000; //  715 :   0 - 0x0
      12'h2CC: dout <= 8'b00000000; //  716 :   0 - 0x0
      12'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      12'h2CE: dout <= 8'b00000000; //  718 :   0 - 0x0
      12'h2CF: dout <= 8'b00000000; //  719 :   0 - 0x0
      12'h2D0: dout <= 8'b00101111; //  720 :  47 - 0x2f -- Sprite 0x2d
      12'h2D1: dout <= 8'b01001111; //  721 :  79 - 0x4f
      12'h2D2: dout <= 8'b01001111; //  722 :  79 - 0x4f
      12'h2D3: dout <= 8'b01001111; //  723 :  79 - 0x4f
      12'h2D4: dout <= 8'b01001111; //  724 :  79 - 0x4f
      12'h2D5: dout <= 8'b00100111; //  725 :  39 - 0x27
      12'h2D6: dout <= 8'b00010000; //  726 :  16 - 0x10
      12'h2D7: dout <= 8'b00001111; //  727 :  15 - 0xf
      12'h2D8: dout <= 8'b00011110; //  728 :  30 - 0x1e -- plane 1
      12'h2D9: dout <= 8'b00111110; //  729 :  62 - 0x3e
      12'h2DA: dout <= 8'b00111110; //  730 :  62 - 0x3e
      12'h2DB: dout <= 8'b00111110; //  731 :  62 - 0x3e
      12'h2DC: dout <= 8'b00111111; //  732 :  63 - 0x3f
      12'h2DD: dout <= 8'b00011110; //  733 :  30 - 0x1e
      12'h2DE: dout <= 8'b00001111; //  734 :  15 - 0xf
      12'h2DF: dout <= 8'b00000000; //  735 :   0 - 0x0
      12'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x2e
      12'h2E1: dout <= 8'b00000000; //  737 :   0 - 0x0
      12'h2E2: dout <= 8'b00000000; //  738 :   0 - 0x0
      12'h2E3: dout <= 8'b00000000; //  739 :   0 - 0x0
      12'h2E4: dout <= 8'b00000000; //  740 :   0 - 0x0
      12'h2E5: dout <= 8'b00000000; //  741 :   0 - 0x0
      12'h2E6: dout <= 8'b00000000; //  742 :   0 - 0x0
      12'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0 -- plane 1
      12'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      12'h2EA: dout <= 8'b00000000; //  746 :   0 - 0x0
      12'h2EB: dout <= 8'b00000000; //  747 :   0 - 0x0
      12'h2EC: dout <= 8'b00000000; //  748 :   0 - 0x0
      12'h2ED: dout <= 8'b00000000; //  749 :   0 - 0x0
      12'h2EE: dout <= 8'b00000000; //  750 :   0 - 0x0
      12'h2EF: dout <= 8'b00000000; //  751 :   0 - 0x0
      12'h2F0: dout <= 8'b11110100; //  752 : 244 - 0xf4 -- Sprite 0x2f
      12'h2F1: dout <= 8'b11110010; //  753 : 242 - 0xf2
      12'h2F2: dout <= 8'b11110010; //  754 : 242 - 0xf2
      12'h2F3: dout <= 8'b11110010; //  755 : 242 - 0xf2
      12'h2F4: dout <= 8'b11110010; //  756 : 242 - 0xf2
      12'h2F5: dout <= 8'b11100100; //  757 : 228 - 0xe4
      12'h2F6: dout <= 8'b00001000; //  758 :   8 - 0x8
      12'h2F7: dout <= 8'b11110000; //  759 : 240 - 0xf0
      12'h2F8: dout <= 8'b01111000; //  760 : 120 - 0x78 -- plane 1
      12'h2F9: dout <= 8'b01111100; //  761 : 124 - 0x7c
      12'h2FA: dout <= 8'b01111100; //  762 : 124 - 0x7c
      12'h2FB: dout <= 8'b01111100; //  763 : 124 - 0x7c
      12'h2FC: dout <= 8'b11111100; //  764 : 252 - 0xfc
      12'h2FD: dout <= 8'b01111000; //  765 : 120 - 0x78
      12'h2FE: dout <= 8'b11110000; //  766 : 240 - 0xf0
      12'h2FF: dout <= 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout <= 8'b00011000; //  768 :  24 - 0x18 -- Sprite 0x30
      12'h301: dout <= 8'b00100100; //  769 :  36 - 0x24
      12'h302: dout <= 8'b01000010; //  770 :  66 - 0x42
      12'h303: dout <= 8'b10100101; //  771 : 165 - 0xa5
      12'h304: dout <= 8'b11100111; //  772 : 231 - 0xe7
      12'h305: dout <= 8'b00100100; //  773 :  36 - 0x24
      12'h306: dout <= 8'b00100100; //  774 :  36 - 0x24
      12'h307: dout <= 8'b00111100; //  775 :  60 - 0x3c
      12'h308: dout <= 8'b00000000; //  776 :   0 - 0x0 -- plane 1
      12'h309: dout <= 8'b00011000; //  777 :  24 - 0x18
      12'h30A: dout <= 8'b00111100; //  778 :  60 - 0x3c
      12'h30B: dout <= 8'b01011010; //  779 :  90 - 0x5a
      12'h30C: dout <= 8'b00011000; //  780 :  24 - 0x18
      12'h30D: dout <= 8'b00011000; //  781 :  24 - 0x18
      12'h30E: dout <= 8'b00011000; //  782 :  24 - 0x18
      12'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      12'h310: dout <= 8'b00111100; //  784 :  60 - 0x3c -- Sprite 0x31
      12'h311: dout <= 8'b00100100; //  785 :  36 - 0x24
      12'h312: dout <= 8'b00100100; //  786 :  36 - 0x24
      12'h313: dout <= 8'b01100110; //  787 : 102 - 0x66
      12'h314: dout <= 8'b10100101; //  788 : 165 - 0xa5
      12'h315: dout <= 8'b01000010; //  789 :  66 - 0x42
      12'h316: dout <= 8'b00100100; //  790 :  36 - 0x24
      12'h317: dout <= 8'b00011000; //  791 :  24 - 0x18
      12'h318: dout <= 8'b00000000; //  792 :   0 - 0x0 -- plane 1
      12'h319: dout <= 8'b00011000; //  793 :  24 - 0x18
      12'h31A: dout <= 8'b00011000; //  794 :  24 - 0x18
      12'h31B: dout <= 8'b00011000; //  795 :  24 - 0x18
      12'h31C: dout <= 8'b01011010; //  796 :  90 - 0x5a
      12'h31D: dout <= 8'b00111100; //  797 :  60 - 0x3c
      12'h31E: dout <= 8'b00011000; //  798 :  24 - 0x18
      12'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout <= 8'b00000010; //  800 :   2 - 0x2 -- Sprite 0x32
      12'h321: dout <= 8'b00000010; //  801 :   2 - 0x2
      12'h322: dout <= 8'b00000011; //  802 :   3 - 0x3
      12'h323: dout <= 8'b00000010; //  803 :   2 - 0x2
      12'h324: dout <= 8'b00000010; //  804 :   2 - 0x2
      12'h325: dout <= 8'b00000010; //  805 :   2 - 0x2
      12'h326: dout <= 8'b00000011; //  806 :   3 - 0x3
      12'h327: dout <= 8'b00000010; //  807 :   2 - 0x2
      12'h328: dout <= 8'b00000001; //  808 :   1 - 0x1 -- plane 1
      12'h329: dout <= 8'b00000001; //  809 :   1 - 0x1
      12'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      12'h32B: dout <= 8'b00000001; //  811 :   1 - 0x1
      12'h32C: dout <= 8'b00000001; //  812 :   1 - 0x1
      12'h32D: dout <= 8'b00000001; //  813 :   1 - 0x1
      12'h32E: dout <= 8'b00000000; //  814 :   0 - 0x0
      12'h32F: dout <= 8'b00000001; //  815 :   1 - 0x1
      12'h330: dout <= 8'b01000000; //  816 :  64 - 0x40 -- Sprite 0x33
      12'h331: dout <= 8'b11000000; //  817 : 192 - 0xc0
      12'h332: dout <= 8'b01000000; //  818 :  64 - 0x40
      12'h333: dout <= 8'b01000000; //  819 :  64 - 0x40
      12'h334: dout <= 8'b01000000; //  820 :  64 - 0x40
      12'h335: dout <= 8'b11000000; //  821 : 192 - 0xc0
      12'h336: dout <= 8'b01000000; //  822 :  64 - 0x40
      12'h337: dout <= 8'b01000000; //  823 :  64 - 0x40
      12'h338: dout <= 8'b10000000; //  824 : 128 - 0x80 -- plane 1
      12'h339: dout <= 8'b00000000; //  825 :   0 - 0x0
      12'h33A: dout <= 8'b10000000; //  826 : 128 - 0x80
      12'h33B: dout <= 8'b10000000; //  827 : 128 - 0x80
      12'h33C: dout <= 8'b10000000; //  828 : 128 - 0x80
      12'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      12'h33E: dout <= 8'b10000000; //  830 : 128 - 0x80
      12'h33F: dout <= 8'b10000000; //  831 : 128 - 0x80
      12'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x34
      12'h341: dout <= 8'b00011000; //  833 :  24 - 0x18
      12'h342: dout <= 8'b00111100; //  834 :  60 - 0x3c
      12'h343: dout <= 8'b01100010; //  835 :  98 - 0x62
      12'h344: dout <= 8'b01100001; //  836 :  97 - 0x61
      12'h345: dout <= 8'b11000000; //  837 : 192 - 0xc0
      12'h346: dout <= 8'b11000000; //  838 : 192 - 0xc0
      12'h347: dout <= 8'b11000000; //  839 : 192 - 0xc0
      12'h348: dout <= 8'b00000000; //  840 :   0 - 0x0 -- plane 1
      12'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout <= 8'b00011000; //  842 :  24 - 0x18
      12'h34B: dout <= 8'b00111100; //  843 :  60 - 0x3c
      12'h34C: dout <= 8'b00111110; //  844 :  62 - 0x3e
      12'h34D: dout <= 8'b01111111; //  845 : 127 - 0x7f
      12'h34E: dout <= 8'b01111111; //  846 : 127 - 0x7f
      12'h34F: dout <= 8'b01111111; //  847 : 127 - 0x7f
      12'h350: dout <= 8'b01100000; //  848 :  96 - 0x60 -- Sprite 0x35
      12'h351: dout <= 8'b01100000; //  849 :  96 - 0x60
      12'h352: dout <= 8'b00110000; //  850 :  48 - 0x30
      12'h353: dout <= 8'b00011000; //  851 :  24 - 0x18
      12'h354: dout <= 8'b00001100; //  852 :  12 - 0xc
      12'h355: dout <= 8'b00000110; //  853 :   6 - 0x6
      12'h356: dout <= 8'b00000010; //  854 :   2 - 0x2
      12'h357: dout <= 8'b00000001; //  855 :   1 - 0x1
      12'h358: dout <= 8'b00111111; //  856 :  63 - 0x3f -- plane 1
      12'h359: dout <= 8'b00111111; //  857 :  63 - 0x3f
      12'h35A: dout <= 8'b00011111; //  858 :  31 - 0x1f
      12'h35B: dout <= 8'b00001111; //  859 :  15 - 0xf
      12'h35C: dout <= 8'b00000111; //  860 :   7 - 0x7
      12'h35D: dout <= 8'b00000011; //  861 :   3 - 0x3
      12'h35E: dout <= 8'b00000001; //  862 :   1 - 0x1
      12'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout <= 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x36
      12'h361: dout <= 8'b00011000; //  865 :  24 - 0x18
      12'h362: dout <= 8'b00100100; //  866 :  36 - 0x24
      12'h363: dout <= 8'b01000010; //  867 :  66 - 0x42
      12'h364: dout <= 8'b10000010; //  868 : 130 - 0x82
      12'h365: dout <= 8'b00000001; //  869 :   1 - 0x1
      12'h366: dout <= 8'b00000001; //  870 :   1 - 0x1
      12'h367: dout <= 8'b00000001; //  871 :   1 - 0x1
      12'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- plane 1
      12'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout <= 8'b00011000; //  874 :  24 - 0x18
      12'h36B: dout <= 8'b00111100; //  875 :  60 - 0x3c
      12'h36C: dout <= 8'b01111100; //  876 : 124 - 0x7c
      12'h36D: dout <= 8'b11111110; //  877 : 254 - 0xfe
      12'h36E: dout <= 8'b11111110; //  878 : 254 - 0xfe
      12'h36F: dout <= 8'b11111110; //  879 : 254 - 0xfe
      12'h370: dout <= 8'b00000010; //  880 :   2 - 0x2 -- Sprite 0x37
      12'h371: dout <= 8'b00000010; //  881 :   2 - 0x2
      12'h372: dout <= 8'b00000100; //  882 :   4 - 0x4
      12'h373: dout <= 8'b00001000; //  883 :   8 - 0x8
      12'h374: dout <= 8'b00010000; //  884 :  16 - 0x10
      12'h375: dout <= 8'b00100000; //  885 :  32 - 0x20
      12'h376: dout <= 8'b01000000; //  886 :  64 - 0x40
      12'h377: dout <= 8'b10000000; //  887 : 128 - 0x80
      12'h378: dout <= 8'b11111100; //  888 : 252 - 0xfc -- plane 1
      12'h379: dout <= 8'b11111100; //  889 : 252 - 0xfc
      12'h37A: dout <= 8'b11111000; //  890 : 248 - 0xf8
      12'h37B: dout <= 8'b11110000; //  891 : 240 - 0xf0
      12'h37C: dout <= 8'b11100000; //  892 : 224 - 0xe0
      12'h37D: dout <= 8'b11000000; //  893 : 192 - 0xc0
      12'h37E: dout <= 8'b10000000; //  894 : 128 - 0x80
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x38
      12'h381: dout <= 8'b00000110; //  897 :   6 - 0x6
      12'h382: dout <= 8'b00001101; //  898 :  13 - 0xd
      12'h383: dout <= 8'b00001100; //  899 :  12 - 0xc
      12'h384: dout <= 8'b00001100; //  900 :  12 - 0xc
      12'h385: dout <= 8'b00000110; //  901 :   6 - 0x6
      12'h386: dout <= 8'b00000010; //  902 :   2 - 0x2
      12'h387: dout <= 8'b00000001; //  903 :   1 - 0x1
      12'h388: dout <= 8'b00000000; //  904 :   0 - 0x0 -- plane 1
      12'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout <= 8'b00000110; //  906 :   6 - 0x6
      12'h38B: dout <= 8'b00000111; //  907 :   7 - 0x7
      12'h38C: dout <= 8'b00000111; //  908 :   7 - 0x7
      12'h38D: dout <= 8'b00000011; //  909 :   3 - 0x3
      12'h38E: dout <= 8'b00000001; //  910 :   1 - 0x1
      12'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      12'h390: dout <= 8'b11111111; //  912 : 255 - 0xff -- Sprite 0x39
      12'h391: dout <= 8'b00000000; //  913 :   0 - 0x0
      12'h392: dout <= 8'b00000000; //  914 :   0 - 0x0
      12'h393: dout <= 8'b00000000; //  915 :   0 - 0x0
      12'h394: dout <= 8'b00000000; //  916 :   0 - 0x0
      12'h395: dout <= 8'b00000000; //  917 :   0 - 0x0
      12'h396: dout <= 8'b00000000; //  918 :   0 - 0x0
      12'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout <= 8'b00000000; //  920 :   0 - 0x0 -- plane 1
      12'h399: dout <= 8'b00000000; //  921 :   0 - 0x0
      12'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      12'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      12'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      12'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      12'h39E: dout <= 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x3a
      12'h3A1: dout <= 8'b01100000; //  929 :  96 - 0x60
      12'h3A2: dout <= 8'b10010000; //  930 : 144 - 0x90
      12'h3A3: dout <= 8'b00010000; //  931 :  16 - 0x10
      12'h3A4: dout <= 8'b00010000; //  932 :  16 - 0x10
      12'h3A5: dout <= 8'b00100000; //  933 :  32 - 0x20
      12'h3A6: dout <= 8'b01000000; //  934 :  64 - 0x40
      12'h3A7: dout <= 8'b10000000; //  935 : 128 - 0x80
      12'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0 -- plane 1
      12'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout <= 8'b01100000; //  938 :  96 - 0x60
      12'h3AB: dout <= 8'b11100000; //  939 : 224 - 0xe0
      12'h3AC: dout <= 8'b11100000; //  940 : 224 - 0xe0
      12'h3AD: dout <= 8'b11000000; //  941 : 192 - 0xc0
      12'h3AE: dout <= 8'b10000000; //  942 : 128 - 0x80
      12'h3AF: dout <= 8'b00000000; //  943 :   0 - 0x0
      12'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x3b
      12'h3B1: dout <= 8'b01010100; //  945 :  84 - 0x54
      12'h3B2: dout <= 8'b00000010; //  946 :   2 - 0x2
      12'h3B3: dout <= 8'b01000000; //  947 :  64 - 0x40
      12'h3B4: dout <= 8'b00000010; //  948 :   2 - 0x2
      12'h3B5: dout <= 8'b01000000; //  949 :  64 - 0x40
      12'h3B6: dout <= 8'b00101010; //  950 :  42 - 0x2a
      12'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout <= 8'b00000000; //  952 :   0 - 0x0 -- plane 1
      12'h3B9: dout <= 8'b00101010; //  953 :  42 - 0x2a
      12'h3BA: dout <= 8'b01000000; //  954 :  64 - 0x40
      12'h3BB: dout <= 8'b00000010; //  955 :   2 - 0x2
      12'h3BC: dout <= 8'b01000000; //  956 :  64 - 0x40
      12'h3BD: dout <= 8'b00000010; //  957 :   2 - 0x2
      12'h3BE: dout <= 8'b01010100; //  958 :  84 - 0x54
      12'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout <= 8'b11111111; //  960 : 255 - 0xff -- Sprite 0x3c
      12'h3C1: dout <= 8'b11111111; //  961 : 255 - 0xff
      12'h3C2: dout <= 8'b11111111; //  962 : 255 - 0xff
      12'h3C3: dout <= 8'b11111111; //  963 : 255 - 0xff
      12'h3C4: dout <= 8'b11111111; //  964 : 255 - 0xff
      12'h3C5: dout <= 8'b11111111; //  965 : 255 - 0xff
      12'h3C6: dout <= 8'b11111111; //  966 : 255 - 0xff
      12'h3C7: dout <= 8'b11111111; //  967 : 255 - 0xff
      12'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- plane 1
      12'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x3d
      12'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      12'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      12'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout <= 8'b11111111; //  984 : 255 - 0xff -- plane 1
      12'h3D9: dout <= 8'b11111111; //  985 : 255 - 0xff
      12'h3DA: dout <= 8'b11111111; //  986 : 255 - 0xff
      12'h3DB: dout <= 8'b11111111; //  987 : 255 - 0xff
      12'h3DC: dout <= 8'b11111111; //  988 : 255 - 0xff
      12'h3DD: dout <= 8'b11111111; //  989 : 255 - 0xff
      12'h3DE: dout <= 8'b11111111; //  990 : 255 - 0xff
      12'h3DF: dout <= 8'b11111111; //  991 : 255 - 0xff
      12'h3E0: dout <= 8'b11111111; //  992 : 255 - 0xff -- Sprite 0x3e
      12'h3E1: dout <= 8'b11111111; //  993 : 255 - 0xff
      12'h3E2: dout <= 8'b11111111; //  994 : 255 - 0xff
      12'h3E3: dout <= 8'b11111111; //  995 : 255 - 0xff
      12'h3E4: dout <= 8'b11111111; //  996 : 255 - 0xff
      12'h3E5: dout <= 8'b11111111; //  997 : 255 - 0xff
      12'h3E6: dout <= 8'b11111111; //  998 : 255 - 0xff
      12'h3E7: dout <= 8'b11111111; //  999 : 255 - 0xff
      12'h3E8: dout <= 8'b11111111; // 1000 : 255 - 0xff -- plane 1
      12'h3E9: dout <= 8'b11111111; // 1001 : 255 - 0xff
      12'h3EA: dout <= 8'b11111111; // 1002 : 255 - 0xff
      12'h3EB: dout <= 8'b11111111; // 1003 : 255 - 0xff
      12'h3EC: dout <= 8'b11111111; // 1004 : 255 - 0xff
      12'h3ED: dout <= 8'b11111111; // 1005 : 255 - 0xff
      12'h3EE: dout <= 8'b11111111; // 1006 : 255 - 0xff
      12'h3EF: dout <= 8'b11111111; // 1007 : 255 - 0xff
      12'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x3f
      12'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout <= 8'b00000000; // 1012 :   0 - 0x0
      12'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0 -- plane 1
      12'h3F9: dout <= 8'b00000000; // 1017 :   0 - 0x0
      12'h3FA: dout <= 8'b00000000; // 1018 :   0 - 0x0
      12'h3FB: dout <= 8'b00000000; // 1019 :   0 - 0x0
      12'h3FC: dout <= 8'b00000000; // 1020 :   0 - 0x0
      12'h3FD: dout <= 8'b00000000; // 1021 :   0 - 0x0
      12'h3FE: dout <= 8'b00000000; // 1022 :   0 - 0x0
      12'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout <= 8'b00111100; // 1024 :  60 - 0x3c -- Sprite 0x40
      12'h401: dout <= 8'b01000010; // 1025 :  66 - 0x42
      12'h402: dout <= 8'b10011001; // 1026 : 153 - 0x99
      12'h403: dout <= 8'b10100101; // 1027 : 165 - 0xa5
      12'h404: dout <= 8'b10100101; // 1028 : 165 - 0xa5
      12'h405: dout <= 8'b10011010; // 1029 : 154 - 0x9a
      12'h406: dout <= 8'b01000000; // 1030 :  64 - 0x40
      12'h407: dout <= 8'b00111100; // 1031 :  60 - 0x3c
      12'h408: dout <= 8'b00000000; // 1032 :   0 - 0x0 -- plane 1
      12'h409: dout <= 8'b00000000; // 1033 :   0 - 0x0
      12'h40A: dout <= 8'b00000000; // 1034 :   0 - 0x0
      12'h40B: dout <= 8'b00000000; // 1035 :   0 - 0x0
      12'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      12'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      12'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout <= 8'b00001100; // 1040 :  12 - 0xc -- Sprite 0x41
      12'h411: dout <= 8'b00010010; // 1041 :  18 - 0x12
      12'h412: dout <= 8'b00100010; // 1042 :  34 - 0x22
      12'h413: dout <= 8'b00100010; // 1043 :  34 - 0x22
      12'h414: dout <= 8'b01111110; // 1044 : 126 - 0x7e
      12'h415: dout <= 8'b00100010; // 1045 :  34 - 0x22
      12'h416: dout <= 8'b00100100; // 1046 :  36 - 0x24
      12'h417: dout <= 8'b00000000; // 1047 :   0 - 0x0
      12'h418: dout <= 8'b00000000; // 1048 :   0 - 0x0 -- plane 1
      12'h419: dout <= 8'b00000000; // 1049 :   0 - 0x0
      12'h41A: dout <= 8'b00000000; // 1050 :   0 - 0x0
      12'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      12'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout <= 8'b00111100; // 1056 :  60 - 0x3c -- Sprite 0x42
      12'h421: dout <= 8'b01000010; // 1057 :  66 - 0x42
      12'h422: dout <= 8'b01010010; // 1058 :  82 - 0x52
      12'h423: dout <= 8'b00011100; // 1059 :  28 - 0x1c
      12'h424: dout <= 8'b00010010; // 1060 :  18 - 0x12
      12'h425: dout <= 8'b00110010; // 1061 :  50 - 0x32
      12'h426: dout <= 8'b00011100; // 1062 :  28 - 0x1c
      12'h427: dout <= 8'b00000000; // 1063 :   0 - 0x0
      12'h428: dout <= 8'b00000000; // 1064 :   0 - 0x0 -- plane 1
      12'h429: dout <= 8'b00000000; // 1065 :   0 - 0x0
      12'h42A: dout <= 8'b00000000; // 1066 :   0 - 0x0
      12'h42B: dout <= 8'b00000000; // 1067 :   0 - 0x0
      12'h42C: dout <= 8'b00000000; // 1068 :   0 - 0x0
      12'h42D: dout <= 8'b00000000; // 1069 :   0 - 0x0
      12'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      12'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout <= 8'b00011000; // 1072 :  24 - 0x18 -- Sprite 0x43
      12'h431: dout <= 8'b00100100; // 1073 :  36 - 0x24
      12'h432: dout <= 8'b01010100; // 1074 :  84 - 0x54
      12'h433: dout <= 8'b01001000; // 1075 :  72 - 0x48
      12'h434: dout <= 8'b01000010; // 1076 :  66 - 0x42
      12'h435: dout <= 8'b00100100; // 1077 :  36 - 0x24
      12'h436: dout <= 8'b00011000; // 1078 :  24 - 0x18
      12'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout <= 8'b00000000; // 1080 :   0 - 0x0 -- plane 1
      12'h439: dout <= 8'b00000000; // 1081 :   0 - 0x0
      12'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      12'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      12'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      12'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout <= 8'b01011000; // 1088 :  88 - 0x58 -- Sprite 0x44
      12'h441: dout <= 8'b11100100; // 1089 : 228 - 0xe4
      12'h442: dout <= 8'b01000010; // 1090 :  66 - 0x42
      12'h443: dout <= 8'b01000010; // 1091 :  66 - 0x42
      12'h444: dout <= 8'b00100010; // 1092 :  34 - 0x22
      12'h445: dout <= 8'b01100100; // 1093 : 100 - 0x64
      12'h446: dout <= 8'b00111000; // 1094 :  56 - 0x38
      12'h447: dout <= 8'b00000000; // 1095 :   0 - 0x0
      12'h448: dout <= 8'b00000000; // 1096 :   0 - 0x0 -- plane 1
      12'h449: dout <= 8'b00000000; // 1097 :   0 - 0x0
      12'h44A: dout <= 8'b00000000; // 1098 :   0 - 0x0
      12'h44B: dout <= 8'b00000000; // 1099 :   0 - 0x0
      12'h44C: dout <= 8'b00000000; // 1100 :   0 - 0x0
      12'h44D: dout <= 8'b00000000; // 1101 :   0 - 0x0
      12'h44E: dout <= 8'b00000000; // 1102 :   0 - 0x0
      12'h44F: dout <= 8'b00000000; // 1103 :   0 - 0x0
      12'h450: dout <= 8'b00011100; // 1104 :  28 - 0x1c -- Sprite 0x45
      12'h451: dout <= 8'b00100000; // 1105 :  32 - 0x20
      12'h452: dout <= 8'b00100000; // 1106 :  32 - 0x20
      12'h453: dout <= 8'b00101100; // 1107 :  44 - 0x2c
      12'h454: dout <= 8'b01110000; // 1108 : 112 - 0x70
      12'h455: dout <= 8'b00100010; // 1109 :  34 - 0x22
      12'h456: dout <= 8'b00011100; // 1110 :  28 - 0x1c
      12'h457: dout <= 8'b00000000; // 1111 :   0 - 0x0
      12'h458: dout <= 8'b00000000; // 1112 :   0 - 0x0 -- plane 1
      12'h459: dout <= 8'b00000000; // 1113 :   0 - 0x0
      12'h45A: dout <= 8'b00000000; // 1114 :   0 - 0x0
      12'h45B: dout <= 8'b00000000; // 1115 :   0 - 0x0
      12'h45C: dout <= 8'b00000000; // 1116 :   0 - 0x0
      12'h45D: dout <= 8'b00000000; // 1117 :   0 - 0x0
      12'h45E: dout <= 8'b00000000; // 1118 :   0 - 0x0
      12'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout <= 8'b00011100; // 1120 :  28 - 0x1c -- Sprite 0x46
      12'h461: dout <= 8'b00100000; // 1121 :  32 - 0x20
      12'h462: dout <= 8'b00100000; // 1122 :  32 - 0x20
      12'h463: dout <= 8'b00101100; // 1123 :  44 - 0x2c
      12'h464: dout <= 8'b01110000; // 1124 : 112 - 0x70
      12'h465: dout <= 8'b00010000; // 1125 :  16 - 0x10
      12'h466: dout <= 8'b00010000; // 1126 :  16 - 0x10
      12'h467: dout <= 8'b00000000; // 1127 :   0 - 0x0
      12'h468: dout <= 8'b00000000; // 1128 :   0 - 0x0 -- plane 1
      12'h469: dout <= 8'b00000000; // 1129 :   0 - 0x0
      12'h46A: dout <= 8'b00000000; // 1130 :   0 - 0x0
      12'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      12'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      12'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      12'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      12'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      12'h470: dout <= 8'b00011000; // 1136 :  24 - 0x18 -- Sprite 0x47
      12'h471: dout <= 8'b00100100; // 1137 :  36 - 0x24
      12'h472: dout <= 8'b01000000; // 1138 :  64 - 0x40
      12'h473: dout <= 8'b01001110; // 1139 :  78 - 0x4e
      12'h474: dout <= 8'b01000010; // 1140 :  66 - 0x42
      12'h475: dout <= 8'b00100100; // 1141 :  36 - 0x24
      12'h476: dout <= 8'b00011000; // 1142 :  24 - 0x18
      12'h477: dout <= 8'b00000000; // 1143 :   0 - 0x0
      12'h478: dout <= 8'b00000000; // 1144 :   0 - 0x0 -- plane 1
      12'h479: dout <= 8'b00000000; // 1145 :   0 - 0x0
      12'h47A: dout <= 8'b00000000; // 1146 :   0 - 0x0
      12'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      12'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      12'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      12'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      12'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout <= 8'b00100000; // 1152 :  32 - 0x20 -- Sprite 0x48
      12'h481: dout <= 8'b01000100; // 1153 :  68 - 0x44
      12'h482: dout <= 8'b01000100; // 1154 :  68 - 0x44
      12'h483: dout <= 8'b01000100; // 1155 :  68 - 0x44
      12'h484: dout <= 8'b11111100; // 1156 : 252 - 0xfc
      12'h485: dout <= 8'b01000100; // 1157 :  68 - 0x44
      12'h486: dout <= 8'b01001000; // 1158 :  72 - 0x48
      12'h487: dout <= 8'b00000000; // 1159 :   0 - 0x0
      12'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0 -- plane 1
      12'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      12'h48A: dout <= 8'b00000000; // 1162 :   0 - 0x0
      12'h48B: dout <= 8'b00000000; // 1163 :   0 - 0x0
      12'h48C: dout <= 8'b00000000; // 1164 :   0 - 0x0
      12'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      12'h48E: dout <= 8'b00000000; // 1166 :   0 - 0x0
      12'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout <= 8'b00010000; // 1168 :  16 - 0x10 -- Sprite 0x49
      12'h491: dout <= 8'b00010000; // 1169 :  16 - 0x10
      12'h492: dout <= 8'b00010000; // 1170 :  16 - 0x10
      12'h493: dout <= 8'b00010000; // 1171 :  16 - 0x10
      12'h494: dout <= 8'b00010000; // 1172 :  16 - 0x10
      12'h495: dout <= 8'b00001000; // 1173 :   8 - 0x8
      12'h496: dout <= 8'b00001000; // 1174 :   8 - 0x8
      12'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      12'h498: dout <= 8'b00000000; // 1176 :   0 - 0x0 -- plane 1
      12'h499: dout <= 8'b00000000; // 1177 :   0 - 0x0
      12'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      12'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      12'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      12'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      12'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      12'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      12'h4A0: dout <= 8'b00001000; // 1184 :   8 - 0x8 -- Sprite 0x4a
      12'h4A1: dout <= 8'b00001000; // 1185 :   8 - 0x8
      12'h4A2: dout <= 8'b00000100; // 1186 :   4 - 0x4
      12'h4A3: dout <= 8'b00000100; // 1187 :   4 - 0x4
      12'h4A4: dout <= 8'b01000100; // 1188 :  68 - 0x44
      12'h4A5: dout <= 8'b01001000; // 1189 :  72 - 0x48
      12'h4A6: dout <= 8'b00110000; // 1190 :  48 - 0x30
      12'h4A7: dout <= 8'b00000000; // 1191 :   0 - 0x0
      12'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0 -- plane 1
      12'h4A9: dout <= 8'b00000000; // 1193 :   0 - 0x0
      12'h4AA: dout <= 8'b00000000; // 1194 :   0 - 0x0
      12'h4AB: dout <= 8'b00000000; // 1195 :   0 - 0x0
      12'h4AC: dout <= 8'b00000000; // 1196 :   0 - 0x0
      12'h4AD: dout <= 8'b00000000; // 1197 :   0 - 0x0
      12'h4AE: dout <= 8'b00000000; // 1198 :   0 - 0x0
      12'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      12'h4B0: dout <= 8'b01000100; // 1200 :  68 - 0x44 -- Sprite 0x4b
      12'h4B1: dout <= 8'b01000100; // 1201 :  68 - 0x44
      12'h4B2: dout <= 8'b01001000; // 1202 :  72 - 0x48
      12'h4B3: dout <= 8'b01110000; // 1203 : 112 - 0x70
      12'h4B4: dout <= 8'b01001000; // 1204 :  72 - 0x48
      12'h4B5: dout <= 8'b00100100; // 1205 :  36 - 0x24
      12'h4B6: dout <= 8'b00100010; // 1206 :  34 - 0x22
      12'h4B7: dout <= 8'b00000000; // 1207 :   0 - 0x0
      12'h4B8: dout <= 8'b00000000; // 1208 :   0 - 0x0 -- plane 1
      12'h4B9: dout <= 8'b00000000; // 1209 :   0 - 0x0
      12'h4BA: dout <= 8'b00000000; // 1210 :   0 - 0x0
      12'h4BB: dout <= 8'b00000000; // 1211 :   0 - 0x0
      12'h4BC: dout <= 8'b00000000; // 1212 :   0 - 0x0
      12'h4BD: dout <= 8'b00000000; // 1213 :   0 - 0x0
      12'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      12'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      12'h4C0: dout <= 8'b00010000; // 1216 :  16 - 0x10 -- Sprite 0x4c
      12'h4C1: dout <= 8'b00100000; // 1217 :  32 - 0x20
      12'h4C2: dout <= 8'b00100000; // 1218 :  32 - 0x20
      12'h4C3: dout <= 8'b00100000; // 1219 :  32 - 0x20
      12'h4C4: dout <= 8'b01000000; // 1220 :  64 - 0x40
      12'h4C5: dout <= 8'b01000000; // 1221 :  64 - 0x40
      12'h4C6: dout <= 8'b01000110; // 1222 :  70 - 0x46
      12'h4C7: dout <= 8'b00111000; // 1223 :  56 - 0x38
      12'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0 -- plane 1
      12'h4C9: dout <= 8'b00000000; // 1225 :   0 - 0x0
      12'h4CA: dout <= 8'b00000000; // 1226 :   0 - 0x0
      12'h4CB: dout <= 8'b00000000; // 1227 :   0 - 0x0
      12'h4CC: dout <= 8'b00000000; // 1228 :   0 - 0x0
      12'h4CD: dout <= 8'b00000000; // 1229 :   0 - 0x0
      12'h4CE: dout <= 8'b00000000; // 1230 :   0 - 0x0
      12'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      12'h4D0: dout <= 8'b00100100; // 1232 :  36 - 0x24 -- Sprite 0x4d
      12'h4D1: dout <= 8'b01011010; // 1233 :  90 - 0x5a
      12'h4D2: dout <= 8'b01011010; // 1234 :  90 - 0x5a
      12'h4D3: dout <= 8'b01011010; // 1235 :  90 - 0x5a
      12'h4D4: dout <= 8'b01000010; // 1236 :  66 - 0x42
      12'h4D5: dout <= 8'b01000010; // 1237 :  66 - 0x42
      12'h4D6: dout <= 8'b00100010; // 1238 :  34 - 0x22
      12'h4D7: dout <= 8'b00000000; // 1239 :   0 - 0x0
      12'h4D8: dout <= 8'b00000000; // 1240 :   0 - 0x0 -- plane 1
      12'h4D9: dout <= 8'b00000000; // 1241 :   0 - 0x0
      12'h4DA: dout <= 8'b00000000; // 1242 :   0 - 0x0
      12'h4DB: dout <= 8'b00000000; // 1243 :   0 - 0x0
      12'h4DC: dout <= 8'b00000000; // 1244 :   0 - 0x0
      12'h4DD: dout <= 8'b00000000; // 1245 :   0 - 0x0
      12'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      12'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout <= 8'b00100100; // 1248 :  36 - 0x24 -- Sprite 0x4e
      12'h4E1: dout <= 8'b01010010; // 1249 :  82 - 0x52
      12'h4E2: dout <= 8'b01010010; // 1250 :  82 - 0x52
      12'h4E3: dout <= 8'b01010010; // 1251 :  82 - 0x52
      12'h4E4: dout <= 8'b01010010; // 1252 :  82 - 0x52
      12'h4E5: dout <= 8'b01010010; // 1253 :  82 - 0x52
      12'h4E6: dout <= 8'b01001100; // 1254 :  76 - 0x4c
      12'h4E7: dout <= 8'b00000000; // 1255 :   0 - 0x0
      12'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0 -- plane 1
      12'h4E9: dout <= 8'b00000000; // 1257 :   0 - 0x0
      12'h4EA: dout <= 8'b00000000; // 1258 :   0 - 0x0
      12'h4EB: dout <= 8'b00000000; // 1259 :   0 - 0x0
      12'h4EC: dout <= 8'b00000000; // 1260 :   0 - 0x0
      12'h4ED: dout <= 8'b00000000; // 1261 :   0 - 0x0
      12'h4EE: dout <= 8'b00000000; // 1262 :   0 - 0x0
      12'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout <= 8'b00111000; // 1264 :  56 - 0x38 -- Sprite 0x4f
      12'h4F1: dout <= 8'b01000100; // 1265 :  68 - 0x44
      12'h4F2: dout <= 8'b10000010; // 1266 : 130 - 0x82
      12'h4F3: dout <= 8'b10000010; // 1267 : 130 - 0x82
      12'h4F4: dout <= 8'b10000010; // 1268 : 130 - 0x82
      12'h4F5: dout <= 8'b01000100; // 1269 :  68 - 0x44
      12'h4F6: dout <= 8'b00111000; // 1270 :  56 - 0x38
      12'h4F7: dout <= 8'b00000000; // 1271 :   0 - 0x0
      12'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0 -- plane 1
      12'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      12'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      12'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      12'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      12'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout <= 8'b01111111; // 1280 : 127 - 0x7f -- Sprite 0x50
      12'h501: dout <= 8'b11000000; // 1281 : 192 - 0xc0
      12'h502: dout <= 8'b10000000; // 1282 : 128 - 0x80
      12'h503: dout <= 8'b10000000; // 1283 : 128 - 0x80
      12'h504: dout <= 8'b10000000; // 1284 : 128 - 0x80
      12'h505: dout <= 8'b11000011; // 1285 : 195 - 0xc3
      12'h506: dout <= 8'b11111111; // 1286 : 255 - 0xff
      12'h507: dout <= 8'b11111111; // 1287 : 255 - 0xff
      12'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0 -- plane 1
      12'h509: dout <= 8'b00111111; // 1289 :  63 - 0x3f
      12'h50A: dout <= 8'b01111111; // 1290 : 127 - 0x7f
      12'h50B: dout <= 8'b01111111; // 1291 : 127 - 0x7f
      12'h50C: dout <= 8'b01111111; // 1292 : 127 - 0x7f
      12'h50D: dout <= 8'b00111100; // 1293 :  60 - 0x3c
      12'h50E: dout <= 8'b00000000; // 1294 :   0 - 0x0
      12'h50F: dout <= 8'b01000000; // 1295 :  64 - 0x40
      12'h510: dout <= 8'b11111110; // 1296 : 254 - 0xfe -- Sprite 0x51
      12'h511: dout <= 8'b00000011; // 1297 :   3 - 0x3
      12'h512: dout <= 8'b00000001; // 1298 :   1 - 0x1
      12'h513: dout <= 8'b00000001; // 1299 :   1 - 0x1
      12'h514: dout <= 8'b00000001; // 1300 :   1 - 0x1
      12'h515: dout <= 8'b11000011; // 1301 : 195 - 0xc3
      12'h516: dout <= 8'b11111111; // 1302 : 255 - 0xff
      12'h517: dout <= 8'b11111111; // 1303 : 255 - 0xff
      12'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0 -- plane 1
      12'h519: dout <= 8'b11111100; // 1305 : 252 - 0xfc
      12'h51A: dout <= 8'b11111110; // 1306 : 254 - 0xfe
      12'h51B: dout <= 8'b11111110; // 1307 : 254 - 0xfe
      12'h51C: dout <= 8'b11111110; // 1308 : 254 - 0xfe
      12'h51D: dout <= 8'b00111100; // 1309 :  60 - 0x3c
      12'h51E: dout <= 8'b00000000; // 1310 :   0 - 0x0
      12'h51F: dout <= 8'b00000010; // 1311 :   2 - 0x2
      12'h520: dout <= 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0x52
      12'h521: dout <= 8'b00000111; // 1313 :   7 - 0x7
      12'h522: dout <= 8'b00001100; // 1314 :  12 - 0xc
      12'h523: dout <= 8'b00011000; // 1315 :  24 - 0x18
      12'h524: dout <= 8'b00110000; // 1316 :  48 - 0x30
      12'h525: dout <= 8'b01100000; // 1317 :  96 - 0x60
      12'h526: dout <= 8'b01000000; // 1318 :  64 - 0x40
      12'h527: dout <= 8'b01001111; // 1319 :  79 - 0x4f
      12'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0 -- plane 1
      12'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      12'h52A: dout <= 8'b00000011; // 1322 :   3 - 0x3
      12'h52B: dout <= 8'b00000111; // 1323 :   7 - 0x7
      12'h52C: dout <= 8'b00001111; // 1324 :  15 - 0xf
      12'h52D: dout <= 8'b00011111; // 1325 :  31 - 0x1f
      12'h52E: dout <= 8'b00111111; // 1326 :  63 - 0x3f
      12'h52F: dout <= 8'b00110000; // 1327 :  48 - 0x30
      12'h530: dout <= 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0x53
      12'h531: dout <= 8'b11110000; // 1329 : 240 - 0xf0
      12'h532: dout <= 8'b01010000; // 1330 :  80 - 0x50
      12'h533: dout <= 8'b01001000; // 1331 :  72 - 0x48
      12'h534: dout <= 8'b01001100; // 1332 :  76 - 0x4c
      12'h535: dout <= 8'b01000100; // 1333 :  68 - 0x44
      12'h536: dout <= 8'b10000010; // 1334 : 130 - 0x82
      12'h537: dout <= 8'b10000011; // 1335 : 131 - 0x83
      12'h538: dout <= 8'b00000000; // 1336 :   0 - 0x0 -- plane 1
      12'h539: dout <= 8'b00000000; // 1337 :   0 - 0x0
      12'h53A: dout <= 8'b10100000; // 1338 : 160 - 0xa0
      12'h53B: dout <= 8'b10110000; // 1339 : 176 - 0xb0
      12'h53C: dout <= 8'b10110000; // 1340 : 176 - 0xb0
      12'h53D: dout <= 8'b10111000; // 1341 : 184 - 0xb8
      12'h53E: dout <= 8'b01111100; // 1342 : 124 - 0x7c
      12'h53F: dout <= 8'b01111100; // 1343 : 124 - 0x7c
      12'h540: dout <= 8'b01111111; // 1344 : 127 - 0x7f -- Sprite 0x54
      12'h541: dout <= 8'b11011110; // 1345 : 222 - 0xde
      12'h542: dout <= 8'b10001110; // 1346 : 142 - 0x8e
      12'h543: dout <= 8'b11000101; // 1347 : 197 - 0xc5
      12'h544: dout <= 8'b10010010; // 1348 : 146 - 0x92
      12'h545: dout <= 8'b11000111; // 1349 : 199 - 0xc7
      12'h546: dout <= 8'b11100010; // 1350 : 226 - 0xe2
      12'h547: dout <= 8'b11010000; // 1351 : 208 - 0xd0
      12'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0 -- plane 1
      12'h549: dout <= 8'b00100001; // 1353 :  33 - 0x21
      12'h54A: dout <= 8'b01110001; // 1354 : 113 - 0x71
      12'h54B: dout <= 8'b00111010; // 1355 :  58 - 0x3a
      12'h54C: dout <= 8'b01101101; // 1356 : 109 - 0x6d
      12'h54D: dout <= 8'b00111000; // 1357 :  56 - 0x38
      12'h54E: dout <= 8'b00011101; // 1358 :  29 - 0x1d
      12'h54F: dout <= 8'b00101111; // 1359 :  47 - 0x2f
      12'h550: dout <= 8'b11111111; // 1360 : 255 - 0xff -- Sprite 0x55
      12'h551: dout <= 8'b11011110; // 1361 : 222 - 0xde
      12'h552: dout <= 8'b10001110; // 1362 : 142 - 0x8e
      12'h553: dout <= 8'b11000101; // 1363 : 197 - 0xc5
      12'h554: dout <= 8'b10010010; // 1364 : 146 - 0x92
      12'h555: dout <= 8'b01000111; // 1365 :  71 - 0x47
      12'h556: dout <= 8'b11100010; // 1366 : 226 - 0xe2
      12'h557: dout <= 8'b01010000; // 1367 :  80 - 0x50
      12'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0 -- plane 1
      12'h559: dout <= 8'b00100001; // 1369 :  33 - 0x21
      12'h55A: dout <= 8'b01110001; // 1370 : 113 - 0x71
      12'h55B: dout <= 8'b00111010; // 1371 :  58 - 0x3a
      12'h55C: dout <= 8'b01101101; // 1372 : 109 - 0x6d
      12'h55D: dout <= 8'b10111000; // 1373 : 184 - 0xb8
      12'h55E: dout <= 8'b00011101; // 1374 :  29 - 0x1d
      12'h55F: dout <= 8'b10101111; // 1375 : 175 - 0xaf
      12'h560: dout <= 8'b11111110; // 1376 : 254 - 0xfe -- Sprite 0x56
      12'h561: dout <= 8'b11011111; // 1377 : 223 - 0xdf
      12'h562: dout <= 8'b10001111; // 1378 : 143 - 0x8f
      12'h563: dout <= 8'b11000101; // 1379 : 197 - 0xc5
      12'h564: dout <= 8'b10010011; // 1380 : 147 - 0x93
      12'h565: dout <= 8'b01000111; // 1381 :  71 - 0x47
      12'h566: dout <= 8'b11100011; // 1382 : 227 - 0xe3
      12'h567: dout <= 8'b01010001; // 1383 :  81 - 0x51
      12'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0 -- plane 1
      12'h569: dout <= 8'b00100000; // 1385 :  32 - 0x20
      12'h56A: dout <= 8'b01110000; // 1386 : 112 - 0x70
      12'h56B: dout <= 8'b00111010; // 1387 :  58 - 0x3a
      12'h56C: dout <= 8'b01101100; // 1388 : 108 - 0x6c
      12'h56D: dout <= 8'b10111000; // 1389 : 184 - 0xb8
      12'h56E: dout <= 8'b00011100; // 1390 :  28 - 0x1c
      12'h56F: dout <= 8'b10101110; // 1391 : 174 - 0xae
      12'h570: dout <= 8'b01111111; // 1392 : 127 - 0x7f -- Sprite 0x57
      12'h571: dout <= 8'b10000000; // 1393 : 128 - 0x80
      12'h572: dout <= 8'b10110011; // 1394 : 179 - 0xb3
      12'h573: dout <= 8'b01001100; // 1395 :  76 - 0x4c
      12'h574: dout <= 8'b00111111; // 1396 :  63 - 0x3f
      12'h575: dout <= 8'b00000011; // 1397 :   3 - 0x3
      12'h576: dout <= 8'b00000000; // 1398 :   0 - 0x0
      12'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0 -- plane 1
      12'h579: dout <= 8'b01111111; // 1401 : 127 - 0x7f
      12'h57A: dout <= 8'b01001100; // 1402 :  76 - 0x4c
      12'h57B: dout <= 8'b00110011; // 1403 :  51 - 0x33
      12'h57C: dout <= 8'b00000000; // 1404 :   0 - 0x0
      12'h57D: dout <= 8'b00000000; // 1405 :   0 - 0x0
      12'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      12'h57F: dout <= 8'b00000000; // 1407 :   0 - 0x0
      12'h580: dout <= 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0x58
      12'h581: dout <= 8'b00000000; // 1409 :   0 - 0x0
      12'h582: dout <= 8'b00110011; // 1410 :  51 - 0x33
      12'h583: dout <= 8'b11001100; // 1411 : 204 - 0xcc
      12'h584: dout <= 8'b00110011; // 1412 :  51 - 0x33
      12'h585: dout <= 8'b11111111; // 1413 : 255 - 0xff
      12'h586: dout <= 8'b00000000; // 1414 :   0 - 0x0
      12'h587: dout <= 8'b00000000; // 1415 :   0 - 0x0
      12'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0 -- plane 1
      12'h589: dout <= 8'b11111111; // 1417 : 255 - 0xff
      12'h58A: dout <= 8'b11001100; // 1418 : 204 - 0xcc
      12'h58B: dout <= 8'b00110011; // 1419 :  51 - 0x33
      12'h58C: dout <= 8'b11001100; // 1420 : 204 - 0xcc
      12'h58D: dout <= 8'b00000000; // 1421 :   0 - 0x0
      12'h58E: dout <= 8'b00000000; // 1422 :   0 - 0x0
      12'h58F: dout <= 8'b00000000; // 1423 :   0 - 0x0
      12'h590: dout <= 8'b11111110; // 1424 : 254 - 0xfe -- Sprite 0x59
      12'h591: dout <= 8'b00000001; // 1425 :   1 - 0x1
      12'h592: dout <= 8'b00110011; // 1426 :  51 - 0x33
      12'h593: dout <= 8'b11001110; // 1427 : 206 - 0xce
      12'h594: dout <= 8'b00111100; // 1428 :  60 - 0x3c
      12'h595: dout <= 8'b11000000; // 1429 : 192 - 0xc0
      12'h596: dout <= 8'b00000000; // 1430 :   0 - 0x0
      12'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      12'h598: dout <= 8'b00000000; // 1432 :   0 - 0x0 -- plane 1
      12'h599: dout <= 8'b11111110; // 1433 : 254 - 0xfe
      12'h59A: dout <= 8'b11001100; // 1434 : 204 - 0xcc
      12'h59B: dout <= 8'b00110000; // 1435 :  48 - 0x30
      12'h59C: dout <= 8'b11000000; // 1436 : 192 - 0xc0
      12'h59D: dout <= 8'b00000000; // 1437 :   0 - 0x0
      12'h59E: dout <= 8'b00000000; // 1438 :   0 - 0x0
      12'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout <= 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0x5a
      12'h5A1: dout <= 8'b00000000; // 1441 :   0 - 0x0
      12'h5A2: dout <= 8'b00000000; // 1442 :   0 - 0x0
      12'h5A3: dout <= 8'b00000000; // 1443 :   0 - 0x0
      12'h5A4: dout <= 8'b00000000; // 1444 :   0 - 0x0
      12'h5A5: dout <= 8'b00000000; // 1445 :   0 - 0x0
      12'h5A6: dout <= 8'b00000000; // 1446 :   0 - 0x0
      12'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      12'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0 -- plane 1
      12'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      12'h5AA: dout <= 8'b00000000; // 1450 :   0 - 0x0
      12'h5AB: dout <= 8'b00000000; // 1451 :   0 - 0x0
      12'h5AC: dout <= 8'b00000000; // 1452 :   0 - 0x0
      12'h5AD: dout <= 8'b00000000; // 1453 :   0 - 0x0
      12'h5AE: dout <= 8'b00000000; // 1454 :   0 - 0x0
      12'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      12'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0x5b
      12'h5B1: dout <= 8'b00000000; // 1457 :   0 - 0x0
      12'h5B2: dout <= 8'b00000000; // 1458 :   0 - 0x0
      12'h5B3: dout <= 8'b00000001; // 1459 :   1 - 0x1
      12'h5B4: dout <= 8'b00000011; // 1460 :   3 - 0x3
      12'h5B5: dout <= 8'b00000011; // 1461 :   3 - 0x3
      12'h5B6: dout <= 8'b00000111; // 1462 :   7 - 0x7
      12'h5B7: dout <= 8'b00111111; // 1463 :  63 - 0x3f
      12'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0 -- plane 1
      12'h5B9: dout <= 8'b00000000; // 1465 :   0 - 0x0
      12'h5BA: dout <= 8'b00000000; // 1466 :   0 - 0x0
      12'h5BB: dout <= 8'b00000000; // 1467 :   0 - 0x0
      12'h5BC: dout <= 8'b00000001; // 1468 :   1 - 0x1
      12'h5BD: dout <= 8'b00000001; // 1469 :   1 - 0x1
      12'h5BE: dout <= 8'b00000011; // 1470 :   3 - 0x3
      12'h5BF: dout <= 8'b00000011; // 1471 :   3 - 0x3
      12'h5C0: dout <= 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0x5c
      12'h5C1: dout <= 8'b00000001; // 1473 :   1 - 0x1
      12'h5C2: dout <= 8'b01111111; // 1474 : 127 - 0x7f
      12'h5C3: dout <= 8'b11111111; // 1475 : 255 - 0xff
      12'h5C4: dout <= 8'b11111111; // 1476 : 255 - 0xff
      12'h5C5: dout <= 8'b11111111; // 1477 : 255 - 0xff
      12'h5C6: dout <= 8'b11111111; // 1478 : 255 - 0xff
      12'h5C7: dout <= 8'b11111111; // 1479 : 255 - 0xff
      12'h5C8: dout <= 8'b00000000; // 1480 :   0 - 0x0 -- plane 1
      12'h5C9: dout <= 8'b00000000; // 1481 :   0 - 0x0
      12'h5CA: dout <= 8'b00000001; // 1482 :   1 - 0x1
      12'h5CB: dout <= 8'b01111110; // 1483 : 126 - 0x7e
      12'h5CC: dout <= 8'b11111111; // 1484 : 255 - 0xff
      12'h5CD: dout <= 8'b11111111; // 1485 : 255 - 0xff
      12'h5CE: dout <= 8'b11111111; // 1486 : 255 - 0xff
      12'h5CF: dout <= 8'b11111111; // 1487 : 255 - 0xff
      12'h5D0: dout <= 8'b11111111; // 1488 : 255 - 0xff -- Sprite 0x5d
      12'h5D1: dout <= 8'b11111111; // 1489 : 255 - 0xff
      12'h5D2: dout <= 8'b11111111; // 1490 : 255 - 0xff
      12'h5D3: dout <= 8'b11111111; // 1491 : 255 - 0xff
      12'h5D4: dout <= 8'b11111111; // 1492 : 255 - 0xff
      12'h5D5: dout <= 8'b11111111; // 1493 : 255 - 0xff
      12'h5D6: dout <= 8'b11111111; // 1494 : 255 - 0xff
      12'h5D7: dout <= 8'b11111111; // 1495 : 255 - 0xff
      12'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0 -- plane 1
      12'h5D9: dout <= 8'b11111111; // 1497 : 255 - 0xff
      12'h5DA: dout <= 8'b11111111; // 1498 : 255 - 0xff
      12'h5DB: dout <= 8'b11111111; // 1499 : 255 - 0xff
      12'h5DC: dout <= 8'b01111111; // 1500 : 127 - 0x7f
      12'h5DD: dout <= 8'b11111111; // 1501 : 255 - 0xff
      12'h5DE: dout <= 8'b11111111; // 1502 : 255 - 0xff
      12'h5DF: dout <= 8'b11111111; // 1503 : 255 - 0xff
      12'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0x5e
      12'h5E1: dout <= 8'b10000000; // 1505 : 128 - 0x80
      12'h5E2: dout <= 8'b11111110; // 1506 : 254 - 0xfe
      12'h5E3: dout <= 8'b11111111; // 1507 : 255 - 0xff
      12'h5E4: dout <= 8'b11111111; // 1508 : 255 - 0xff
      12'h5E5: dout <= 8'b11111111; // 1509 : 255 - 0xff
      12'h5E6: dout <= 8'b11111111; // 1510 : 255 - 0xff
      12'h5E7: dout <= 8'b11111111; // 1511 : 255 - 0xff
      12'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0 -- plane 1
      12'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      12'h5EA: dout <= 8'b10000000; // 1514 : 128 - 0x80
      12'h5EB: dout <= 8'b01111110; // 1515 : 126 - 0x7e
      12'h5EC: dout <= 8'b10111111; // 1516 : 191 - 0xbf
      12'h5ED: dout <= 8'b11111111; // 1517 : 255 - 0xff
      12'h5EE: dout <= 8'b11111111; // 1518 : 255 - 0xff
      12'h5EF: dout <= 8'b11111111; // 1519 : 255 - 0xff
      12'h5F0: dout <= 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0x5f
      12'h5F1: dout <= 8'b00000000; // 1521 :   0 - 0x0
      12'h5F2: dout <= 8'b00000000; // 1522 :   0 - 0x0
      12'h5F3: dout <= 8'b10000000; // 1523 : 128 - 0x80
      12'h5F4: dout <= 8'b11000000; // 1524 : 192 - 0xc0
      12'h5F5: dout <= 8'b11000000; // 1525 : 192 - 0xc0
      12'h5F6: dout <= 8'b11100000; // 1526 : 224 - 0xe0
      12'h5F7: dout <= 8'b11111000; // 1527 : 248 - 0xf8
      12'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- plane 1
      12'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      12'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      12'h5FC: dout <= 8'b10000000; // 1532 : 128 - 0x80
      12'h5FD: dout <= 8'b10000000; // 1533 : 128 - 0x80
      12'h5FE: dout <= 8'b11000000; // 1534 : 192 - 0xc0
      12'h5FF: dout <= 8'b11000000; // 1535 : 192 - 0xc0
      12'h600: dout <= 8'b11111111; // 1536 : 255 - 0xff -- Sprite 0x60
      12'h601: dout <= 8'b11111111; // 1537 : 255 - 0xff
      12'h602: dout <= 8'b11111111; // 1538 : 255 - 0xff
      12'h603: dout <= 8'b11111111; // 1539 : 255 - 0xff
      12'h604: dout <= 8'b11111111; // 1540 : 255 - 0xff
      12'h605: dout <= 8'b11111111; // 1541 : 255 - 0xff
      12'h606: dout <= 8'b11111111; // 1542 : 255 - 0xff
      12'h607: dout <= 8'b11111111; // 1543 : 255 - 0xff
      12'h608: dout <= 8'b01111111; // 1544 : 127 - 0x7f -- plane 1
      12'h609: dout <= 8'b01111111; // 1545 : 127 - 0x7f
      12'h60A: dout <= 8'b01111101; // 1546 : 125 - 0x7d
      12'h60B: dout <= 8'b01111111; // 1547 : 127 - 0x7f
      12'h60C: dout <= 8'b00111111; // 1548 :  63 - 0x3f
      12'h60D: dout <= 8'b01111111; // 1549 : 127 - 0x7f
      12'h60E: dout <= 8'b01111111; // 1550 : 127 - 0x7f
      12'h60F: dout <= 8'b01110111; // 1551 : 119 - 0x77
      12'h610: dout <= 8'b11111111; // 1552 : 255 - 0xff -- Sprite 0x61
      12'h611: dout <= 8'b11111111; // 1553 : 255 - 0xff
      12'h612: dout <= 8'b11111111; // 1554 : 255 - 0xff
      12'h613: dout <= 8'b11111111; // 1555 : 255 - 0xff
      12'h614: dout <= 8'b11111111; // 1556 : 255 - 0xff
      12'h615: dout <= 8'b11111111; // 1557 : 255 - 0xff
      12'h616: dout <= 8'b11111111; // 1558 : 255 - 0xff
      12'h617: dout <= 8'b11111111; // 1559 : 255 - 0xff
      12'h618: dout <= 8'b11111110; // 1560 : 254 - 0xfe -- plane 1
      12'h619: dout <= 8'b11111110; // 1561 : 254 - 0xfe
      12'h61A: dout <= 8'b11111100; // 1562 : 252 - 0xfc
      12'h61B: dout <= 8'b11111110; // 1563 : 254 - 0xfe
      12'h61C: dout <= 8'b10111110; // 1564 : 190 - 0xbe
      12'h61D: dout <= 8'b11111110; // 1565 : 254 - 0xfe
      12'h61E: dout <= 8'b11111110; // 1566 : 254 - 0xfe
      12'h61F: dout <= 8'b11110110; // 1567 : 246 - 0xf6
      12'h620: dout <= 8'b01111000; // 1568 : 120 - 0x78 -- Sprite 0x62
      12'h621: dout <= 8'b01100000; // 1569 :  96 - 0x60
      12'h622: dout <= 8'b01000000; // 1570 :  64 - 0x40
      12'h623: dout <= 8'b01000000; // 1571 :  64 - 0x40
      12'h624: dout <= 8'b01000000; // 1572 :  64 - 0x40
      12'h625: dout <= 8'b01100000; // 1573 :  96 - 0x60
      12'h626: dout <= 8'b00110000; // 1574 :  48 - 0x30
      12'h627: dout <= 8'b00011111; // 1575 :  31 - 0x1f
      12'h628: dout <= 8'b00000111; // 1576 :   7 - 0x7 -- plane 1
      12'h629: dout <= 8'b00011111; // 1577 :  31 - 0x1f
      12'h62A: dout <= 8'b00111111; // 1578 :  63 - 0x3f
      12'h62B: dout <= 8'b00111111; // 1579 :  63 - 0x3f
      12'h62C: dout <= 8'b00111111; // 1580 :  63 - 0x3f
      12'h62D: dout <= 8'b00011111; // 1581 :  31 - 0x1f
      12'h62E: dout <= 8'b00001111; // 1582 :  15 - 0xf
      12'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout <= 8'b10000001; // 1584 : 129 - 0x81 -- Sprite 0x63
      12'h631: dout <= 8'b10000011; // 1585 : 131 - 0x83
      12'h632: dout <= 8'b11000001; // 1586 : 193 - 0xc1
      12'h633: dout <= 8'b01000011; // 1587 :  67 - 0x43
      12'h634: dout <= 8'b01000001; // 1588 :  65 - 0x41
      12'h635: dout <= 8'b01100011; // 1589 :  99 - 0x63
      12'h636: dout <= 8'b00100110; // 1590 :  38 - 0x26
      12'h637: dout <= 8'b11111000; // 1591 : 248 - 0xf8
      12'h638: dout <= 8'b01111110; // 1592 : 126 - 0x7e -- plane 1
      12'h639: dout <= 8'b01111100; // 1593 : 124 - 0x7c
      12'h63A: dout <= 8'b00111110; // 1594 :  62 - 0x3e
      12'h63B: dout <= 8'b10111100; // 1595 : 188 - 0xbc
      12'h63C: dout <= 8'b10111110; // 1596 : 190 - 0xbe
      12'h63D: dout <= 8'b10011100; // 1597 : 156 - 0x9c
      12'h63E: dout <= 8'b11011000; // 1598 : 216 - 0xd8
      12'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout <= 8'b10111001; // 1600 : 185 - 0xb9 -- Sprite 0x64
      12'h641: dout <= 8'b10010100; // 1601 : 148 - 0x94
      12'h642: dout <= 8'b10001110; // 1602 : 142 - 0x8e
      12'h643: dout <= 8'b11000101; // 1603 : 197 - 0xc5
      12'h644: dout <= 8'b10010010; // 1604 : 146 - 0x92
      12'h645: dout <= 8'b11000111; // 1605 : 199 - 0xc7
      12'h646: dout <= 8'b11100010; // 1606 : 226 - 0xe2
      12'h647: dout <= 8'b11010000; // 1607 : 208 - 0xd0
      12'h648: dout <= 8'b01000110; // 1608 :  70 - 0x46 -- plane 1
      12'h649: dout <= 8'b01101011; // 1609 : 107 - 0x6b
      12'h64A: dout <= 8'b01110001; // 1610 : 113 - 0x71
      12'h64B: dout <= 8'b00111010; // 1611 :  58 - 0x3a
      12'h64C: dout <= 8'b01101101; // 1612 : 109 - 0x6d
      12'h64D: dout <= 8'b00111000; // 1613 :  56 - 0x38
      12'h64E: dout <= 8'b00011101; // 1614 :  29 - 0x1d
      12'h64F: dout <= 8'b00101111; // 1615 :  47 - 0x2f
      12'h650: dout <= 8'b10111001; // 1616 : 185 - 0xb9 -- Sprite 0x65
      12'h651: dout <= 8'b00010100; // 1617 :  20 - 0x14
      12'h652: dout <= 8'b10001110; // 1618 : 142 - 0x8e
      12'h653: dout <= 8'b11000101; // 1619 : 197 - 0xc5
      12'h654: dout <= 8'b10010010; // 1620 : 146 - 0x92
      12'h655: dout <= 8'b01000111; // 1621 :  71 - 0x47
      12'h656: dout <= 8'b11100010; // 1622 : 226 - 0xe2
      12'h657: dout <= 8'b01010000; // 1623 :  80 - 0x50
      12'h658: dout <= 8'b01000110; // 1624 :  70 - 0x46 -- plane 1
      12'h659: dout <= 8'b11101011; // 1625 : 235 - 0xeb
      12'h65A: dout <= 8'b01110001; // 1626 : 113 - 0x71
      12'h65B: dout <= 8'b00111010; // 1627 :  58 - 0x3a
      12'h65C: dout <= 8'b01101101; // 1628 : 109 - 0x6d
      12'h65D: dout <= 8'b10111000; // 1629 : 184 - 0xb8
      12'h65E: dout <= 8'b00011101; // 1630 :  29 - 0x1d
      12'h65F: dout <= 8'b10101111; // 1631 : 175 - 0xaf
      12'h660: dout <= 8'b10111001; // 1632 : 185 - 0xb9 -- Sprite 0x66
      12'h661: dout <= 8'b00010101; // 1633 :  21 - 0x15
      12'h662: dout <= 8'b10001111; // 1634 : 143 - 0x8f
      12'h663: dout <= 8'b11000101; // 1635 : 197 - 0xc5
      12'h664: dout <= 8'b10010011; // 1636 : 147 - 0x93
      12'h665: dout <= 8'b01000111; // 1637 :  71 - 0x47
      12'h666: dout <= 8'b11100011; // 1638 : 227 - 0xe3
      12'h667: dout <= 8'b01010001; // 1639 :  81 - 0x51
      12'h668: dout <= 8'b01000110; // 1640 :  70 - 0x46 -- plane 1
      12'h669: dout <= 8'b11101010; // 1641 : 234 - 0xea
      12'h66A: dout <= 8'b01110000; // 1642 : 112 - 0x70
      12'h66B: dout <= 8'b00111010; // 1643 :  58 - 0x3a
      12'h66C: dout <= 8'b01101100; // 1644 : 108 - 0x6c
      12'h66D: dout <= 8'b10111000; // 1645 : 184 - 0xb8
      12'h66E: dout <= 8'b00011100; // 1646 :  28 - 0x1c
      12'h66F: dout <= 8'b10101110; // 1647 : 174 - 0xae
      12'h670: dout <= 8'b01111111; // 1648 : 127 - 0x7f -- Sprite 0x67
      12'h671: dout <= 8'b10000000; // 1649 : 128 - 0x80
      12'h672: dout <= 8'b11001100; // 1650 : 204 - 0xcc
      12'h673: dout <= 8'b01111111; // 1651 : 127 - 0x7f
      12'h674: dout <= 8'b00111111; // 1652 :  63 - 0x3f
      12'h675: dout <= 8'b00000011; // 1653 :   3 - 0x3
      12'h676: dout <= 8'b00000000; // 1654 :   0 - 0x0
      12'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      12'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- plane 1
      12'h679: dout <= 8'b01111111; // 1657 : 127 - 0x7f
      12'h67A: dout <= 8'b01111111; // 1658 : 127 - 0x7f
      12'h67B: dout <= 8'b00110011; // 1659 :  51 - 0x33
      12'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      12'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      12'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout <= 8'b11111111; // 1664 : 255 - 0xff -- Sprite 0x68
      12'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout <= 8'b11001100; // 1666 : 204 - 0xcc
      12'h683: dout <= 8'b00110011; // 1667 :  51 - 0x33
      12'h684: dout <= 8'b11111111; // 1668 : 255 - 0xff
      12'h685: dout <= 8'b11111111; // 1669 : 255 - 0xff
      12'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      12'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      12'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- plane 1
      12'h689: dout <= 8'b11111111; // 1673 : 255 - 0xff
      12'h68A: dout <= 8'b11111111; // 1674 : 255 - 0xff
      12'h68B: dout <= 8'b11111111; // 1675 : 255 - 0xff
      12'h68C: dout <= 8'b11001100; // 1676 : 204 - 0xcc
      12'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      12'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      12'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout <= 8'b11111110; // 1680 : 254 - 0xfe -- Sprite 0x69
      12'h691: dout <= 8'b00000001; // 1681 :   1 - 0x1
      12'h692: dout <= 8'b11001101; // 1682 : 205 - 0xcd
      12'h693: dout <= 8'b00111110; // 1683 :  62 - 0x3e
      12'h694: dout <= 8'b11111100; // 1684 : 252 - 0xfc
      12'h695: dout <= 8'b11000000; // 1685 : 192 - 0xc0
      12'h696: dout <= 8'b00000000; // 1686 :   0 - 0x0
      12'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      12'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0 -- plane 1
      12'h699: dout <= 8'b11111110; // 1689 : 254 - 0xfe
      12'h69A: dout <= 8'b11111110; // 1690 : 254 - 0xfe
      12'h69B: dout <= 8'b11110000; // 1691 : 240 - 0xf0
      12'h69C: dout <= 8'b11000000; // 1692 : 192 - 0xc0
      12'h69D: dout <= 8'b00000000; // 1693 :   0 - 0x0
      12'h69E: dout <= 8'b00000000; // 1694 :   0 - 0x0
      12'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      12'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0x6a
      12'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      12'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      12'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      12'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      12'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      12'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      12'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0 -- plane 1
      12'h6A9: dout <= 8'b00000000; // 1705 :   0 - 0x0
      12'h6AA: dout <= 8'b00000000; // 1706 :   0 - 0x0
      12'h6AB: dout <= 8'b00000000; // 1707 :   0 - 0x0
      12'h6AC: dout <= 8'b00000000; // 1708 :   0 - 0x0
      12'h6AD: dout <= 8'b00000000; // 1709 :   0 - 0x0
      12'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      12'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout <= 8'b01111111; // 1712 : 127 - 0x7f -- Sprite 0x6b
      12'h6B1: dout <= 8'b11111111; // 1713 : 255 - 0xff
      12'h6B2: dout <= 8'b11111111; // 1714 : 255 - 0xff
      12'h6B3: dout <= 8'b11111111; // 1715 : 255 - 0xff
      12'h6B4: dout <= 8'b01111111; // 1716 : 127 - 0x7f
      12'h6B5: dout <= 8'b00110000; // 1717 :  48 - 0x30
      12'h6B6: dout <= 8'b00001111; // 1718 :  15 - 0xf
      12'h6B7: dout <= 8'b00000000; // 1719 :   0 - 0x0
      12'h6B8: dout <= 8'b00111101; // 1720 :  61 - 0x3d -- plane 1
      12'h6B9: dout <= 8'b01111111; // 1721 : 127 - 0x7f
      12'h6BA: dout <= 8'b01111111; // 1722 : 127 - 0x7f
      12'h6BB: dout <= 8'b01111111; // 1723 : 127 - 0x7f
      12'h6BC: dout <= 8'b00111111; // 1724 :  63 - 0x3f
      12'h6BD: dout <= 8'b00001111; // 1725 :  15 - 0xf
      12'h6BE: dout <= 8'b00000000; // 1726 :   0 - 0x0
      12'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout <= 8'b11111111; // 1728 : 255 - 0xff -- Sprite 0x6c
      12'h6C1: dout <= 8'b11111111; // 1729 : 255 - 0xff
      12'h6C2: dout <= 8'b11111111; // 1730 : 255 - 0xff
      12'h6C3: dout <= 8'b11111111; // 1731 : 255 - 0xff
      12'h6C4: dout <= 8'b11111111; // 1732 : 255 - 0xff
      12'h6C5: dout <= 8'b11111110; // 1733 : 254 - 0xfe
      12'h6C6: dout <= 8'b00000001; // 1734 :   1 - 0x1
      12'h6C7: dout <= 8'b11111110; // 1735 : 254 - 0xfe
      12'h6C8: dout <= 8'b11111111; // 1736 : 255 - 0xff -- plane 1
      12'h6C9: dout <= 8'b11111111; // 1737 : 255 - 0xff
      12'h6CA: dout <= 8'b11111111; // 1738 : 255 - 0xff
      12'h6CB: dout <= 8'b11111111; // 1739 : 255 - 0xff
      12'h6CC: dout <= 8'b11111111; // 1740 : 255 - 0xff
      12'h6CD: dout <= 8'b11111111; // 1741 : 255 - 0xff
      12'h6CE: dout <= 8'b11111110; // 1742 : 254 - 0xfe
      12'h6CF: dout <= 8'b00000000; // 1743 :   0 - 0x0
      12'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0x6d
      12'h6D1: dout <= 8'b00000000; // 1745 :   0 - 0x0
      12'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      12'h6D3: dout <= 8'b00000000; // 1747 :   0 - 0x0
      12'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      12'h6D5: dout <= 8'b00000000; // 1749 :   0 - 0x0
      12'h6D6: dout <= 8'b00000000; // 1750 :   0 - 0x0
      12'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      12'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0 -- plane 1
      12'h6D9: dout <= 8'b00000000; // 1753 :   0 - 0x0
      12'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      12'h6DB: dout <= 8'b00000000; // 1755 :   0 - 0x0
      12'h6DC: dout <= 8'b00000000; // 1756 :   0 - 0x0
      12'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      12'h6DE: dout <= 8'b00000000; // 1758 :   0 - 0x0
      12'h6DF: dout <= 8'b00000000; // 1759 :   0 - 0x0
      12'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0x6e
      12'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      12'h6E5: dout <= 8'b00000000; // 1765 :   0 - 0x0
      12'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      12'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      12'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- plane 1
      12'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      12'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      12'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      12'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      12'h6ED: dout <= 8'b00000000; // 1773 :   0 - 0x0
      12'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      12'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      12'h6F0: dout <= 8'b11111100; // 1776 : 252 - 0xfc -- Sprite 0x6f
      12'h6F1: dout <= 8'b11111110; // 1777 : 254 - 0xfe
      12'h6F2: dout <= 8'b11111111; // 1778 : 255 - 0xff
      12'h6F3: dout <= 8'b11111111; // 1779 : 255 - 0xff
      12'h6F4: dout <= 8'b11110010; // 1780 : 242 - 0xf2
      12'h6F5: dout <= 8'b00001100; // 1781 :  12 - 0xc
      12'h6F6: dout <= 8'b11110000; // 1782 : 240 - 0xf0
      12'h6F7: dout <= 8'b00000000; // 1783 :   0 - 0x0
      12'h6F8: dout <= 8'b10111000; // 1784 : 184 - 0xb8 -- plane 1
      12'h6F9: dout <= 8'b11111100; // 1785 : 252 - 0xfc
      12'h6FA: dout <= 8'b11111110; // 1786 : 254 - 0xfe
      12'h6FB: dout <= 8'b11111110; // 1787 : 254 - 0xfe
      12'h6FC: dout <= 8'b11111100; // 1788 : 252 - 0xfc
      12'h6FD: dout <= 8'b11110000; // 1789 : 240 - 0xf0
      12'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      12'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout <= 8'b01111111; // 1792 : 127 - 0x7f -- Sprite 0x70
      12'h701: dout <= 8'b11000000; // 1793 : 192 - 0xc0
      12'h702: dout <= 8'b10000000; // 1794 : 128 - 0x80
      12'h703: dout <= 8'b10000000; // 1795 : 128 - 0x80
      12'h704: dout <= 8'b11100011; // 1796 : 227 - 0xe3
      12'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      12'h706: dout <= 8'b11111111; // 1798 : 255 - 0xff
      12'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      12'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0 -- plane 1
      12'h709: dout <= 8'b00111111; // 1801 :  63 - 0x3f
      12'h70A: dout <= 8'b01111111; // 1802 : 127 - 0x7f
      12'h70B: dout <= 8'b01111111; // 1803 : 127 - 0x7f
      12'h70C: dout <= 8'b00011100; // 1804 :  28 - 0x1c
      12'h70D: dout <= 8'b00000000; // 1805 :   0 - 0x0
      12'h70E: dout <= 8'b00000000; // 1806 :   0 - 0x0
      12'h70F: dout <= 8'b00000000; // 1807 :   0 - 0x0
      12'h710: dout <= 8'b11111111; // 1808 : 255 - 0xff -- Sprite 0x71
      12'h711: dout <= 8'b00000000; // 1809 :   0 - 0x0
      12'h712: dout <= 8'b00000000; // 1810 :   0 - 0x0
      12'h713: dout <= 8'b00000000; // 1811 :   0 - 0x0
      12'h714: dout <= 8'b00000000; // 1812 :   0 - 0x0
      12'h715: dout <= 8'b11000011; // 1813 : 195 - 0xc3
      12'h716: dout <= 8'b11111111; // 1814 : 255 - 0xff
      12'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      12'h718: dout <= 8'b00000000; // 1816 :   0 - 0x0 -- plane 1
      12'h719: dout <= 8'b11111111; // 1817 : 255 - 0xff
      12'h71A: dout <= 8'b11111111; // 1818 : 255 - 0xff
      12'h71B: dout <= 8'b11111111; // 1819 : 255 - 0xff
      12'h71C: dout <= 8'b11111111; // 1820 : 255 - 0xff
      12'h71D: dout <= 8'b00111100; // 1821 :  60 - 0x3c
      12'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      12'h720: dout <= 8'b11111110; // 1824 : 254 - 0xfe -- Sprite 0x72
      12'h721: dout <= 8'b00000011; // 1825 :   3 - 0x3
      12'h722: dout <= 8'b00000001; // 1826 :   1 - 0x1
      12'h723: dout <= 8'b00000001; // 1827 :   1 - 0x1
      12'h724: dout <= 8'b11000111; // 1828 : 199 - 0xc7
      12'h725: dout <= 8'b11111111; // 1829 : 255 - 0xff
      12'h726: dout <= 8'b11111111; // 1830 : 255 - 0xff
      12'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      12'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0 -- plane 1
      12'h729: dout <= 8'b11111100; // 1833 : 252 - 0xfc
      12'h72A: dout <= 8'b11111110; // 1834 : 254 - 0xfe
      12'h72B: dout <= 8'b11111110; // 1835 : 254 - 0xfe
      12'h72C: dout <= 8'b00111000; // 1836 :  56 - 0x38
      12'h72D: dout <= 8'b00000000; // 1837 :   0 - 0x0
      12'h72E: dout <= 8'b00000000; // 1838 :   0 - 0x0
      12'h72F: dout <= 8'b00000000; // 1839 :   0 - 0x0
      12'h730: dout <= 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0x73
      12'h731: dout <= 8'b11111111; // 1841 : 255 - 0xff
      12'h732: dout <= 8'b11111111; // 1842 : 255 - 0xff
      12'h733: dout <= 8'b11111111; // 1843 : 255 - 0xff
      12'h734: dout <= 8'b11111111; // 1844 : 255 - 0xff
      12'h735: dout <= 8'b11111111; // 1845 : 255 - 0xff
      12'h736: dout <= 8'b11111111; // 1846 : 255 - 0xff
      12'h737: dout <= 8'b11111111; // 1847 : 255 - 0xff
      12'h738: dout <= 8'b11111111; // 1848 : 255 - 0xff -- plane 1
      12'h739: dout <= 8'b11111111; // 1849 : 255 - 0xff
      12'h73A: dout <= 8'b11111101; // 1850 : 253 - 0xfd
      12'h73B: dout <= 8'b11111111; // 1851 : 255 - 0xff
      12'h73C: dout <= 8'b10111111; // 1852 : 191 - 0xbf
      12'h73D: dout <= 8'b11111111; // 1853 : 255 - 0xff
      12'h73E: dout <= 8'b11111111; // 1854 : 255 - 0xff
      12'h73F: dout <= 8'b11110111; // 1855 : 247 - 0xf7
      12'h740: dout <= 8'b10111001; // 1856 : 185 - 0xb9 -- Sprite 0x74
      12'h741: dout <= 8'b10010100; // 1857 : 148 - 0x94
      12'h742: dout <= 8'b10001110; // 1858 : 142 - 0x8e
      12'h743: dout <= 8'b11000101; // 1859 : 197 - 0xc5
      12'h744: dout <= 8'b10010010; // 1860 : 146 - 0x92
      12'h745: dout <= 8'b11000111; // 1861 : 199 - 0xc7
      12'h746: dout <= 8'b11100010; // 1862 : 226 - 0xe2
      12'h747: dout <= 8'b01111111; // 1863 : 127 - 0x7f
      12'h748: dout <= 8'b01000110; // 1864 :  70 - 0x46 -- plane 1
      12'h749: dout <= 8'b01101011; // 1865 : 107 - 0x6b
      12'h74A: dout <= 8'b01110001; // 1866 : 113 - 0x71
      12'h74B: dout <= 8'b00111010; // 1867 :  58 - 0x3a
      12'h74C: dout <= 8'b01101101; // 1868 : 109 - 0x6d
      12'h74D: dout <= 8'b00111000; // 1869 :  56 - 0x38
      12'h74E: dout <= 8'b00011101; // 1870 :  29 - 0x1d
      12'h74F: dout <= 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout <= 8'b10111001; // 1872 : 185 - 0xb9 -- Sprite 0x75
      12'h751: dout <= 8'b00010100; // 1873 :  20 - 0x14
      12'h752: dout <= 8'b10001110; // 1874 : 142 - 0x8e
      12'h753: dout <= 8'b11000101; // 1875 : 197 - 0xc5
      12'h754: dout <= 8'b10010010; // 1876 : 146 - 0x92
      12'h755: dout <= 8'b01000111; // 1877 :  71 - 0x47
      12'h756: dout <= 8'b11100010; // 1878 : 226 - 0xe2
      12'h757: dout <= 8'b11111111; // 1879 : 255 - 0xff
      12'h758: dout <= 8'b01000110; // 1880 :  70 - 0x46 -- plane 1
      12'h759: dout <= 8'b11101011; // 1881 : 235 - 0xeb
      12'h75A: dout <= 8'b01110001; // 1882 : 113 - 0x71
      12'h75B: dout <= 8'b00111010; // 1883 :  58 - 0x3a
      12'h75C: dout <= 8'b01101101; // 1884 : 109 - 0x6d
      12'h75D: dout <= 8'b10111000; // 1885 : 184 - 0xb8
      12'h75E: dout <= 8'b00011101; // 1886 :  29 - 0x1d
      12'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      12'h760: dout <= 8'b10111001; // 1888 : 185 - 0xb9 -- Sprite 0x76
      12'h761: dout <= 8'b00010101; // 1889 :  21 - 0x15
      12'h762: dout <= 8'b10001111; // 1890 : 143 - 0x8f
      12'h763: dout <= 8'b11000101; // 1891 : 197 - 0xc5
      12'h764: dout <= 8'b10010011; // 1892 : 147 - 0x93
      12'h765: dout <= 8'b01000111; // 1893 :  71 - 0x47
      12'h766: dout <= 8'b11100011; // 1894 : 227 - 0xe3
      12'h767: dout <= 8'b11111110; // 1895 : 254 - 0xfe
      12'h768: dout <= 8'b01000110; // 1896 :  70 - 0x46 -- plane 1
      12'h769: dout <= 8'b11101010; // 1897 : 234 - 0xea
      12'h76A: dout <= 8'b01110000; // 1898 : 112 - 0x70
      12'h76B: dout <= 8'b00111010; // 1899 :  58 - 0x3a
      12'h76C: dout <= 8'b01101100; // 1900 : 108 - 0x6c
      12'h76D: dout <= 8'b10111000; // 1901 : 184 - 0xb8
      12'h76E: dout <= 8'b00011100; // 1902 :  28 - 0x1c
      12'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      12'h770: dout <= 8'b11111111; // 1904 : 255 - 0xff -- Sprite 0x77
      12'h771: dout <= 8'b11111111; // 1905 : 255 - 0xff
      12'h772: dout <= 8'b11111111; // 1906 : 255 - 0xff
      12'h773: dout <= 8'b11111111; // 1907 : 255 - 0xff
      12'h774: dout <= 8'b11111111; // 1908 : 255 - 0xff
      12'h775: dout <= 8'b11111111; // 1909 : 255 - 0xff
      12'h776: dout <= 8'b11111111; // 1910 : 255 - 0xff
      12'h777: dout <= 8'b11111111; // 1911 : 255 - 0xff
      12'h778: dout <= 8'b10000001; // 1912 : 129 - 0x81 -- plane 1
      12'h779: dout <= 8'b11111111; // 1913 : 255 - 0xff
      12'h77A: dout <= 8'b11111101; // 1914 : 253 - 0xfd
      12'h77B: dout <= 8'b11111111; // 1915 : 255 - 0xff
      12'h77C: dout <= 8'b10111111; // 1916 : 191 - 0xbf
      12'h77D: dout <= 8'b11111111; // 1917 : 255 - 0xff
      12'h77E: dout <= 8'b11111111; // 1918 : 255 - 0xff
      12'h77F: dout <= 8'b11110111; // 1919 : 247 - 0xf7
      12'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0x78
      12'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0 -- plane 1
      12'h789: dout <= 8'b00000000; // 1929 :   0 - 0x0
      12'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      12'h78B: dout <= 8'b00000000; // 1931 :   0 - 0x0
      12'h78C: dout <= 8'b00000000; // 1932 :   0 - 0x0
      12'h78D: dout <= 8'b00000000; // 1933 :   0 - 0x0
      12'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      12'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0x79
      12'h791: dout <= 8'b00000000; // 1937 :   0 - 0x0
      12'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0 -- plane 1
      12'h799: dout <= 8'b00000000; // 1945 :   0 - 0x0
      12'h79A: dout <= 8'b00000000; // 1946 :   0 - 0x0
      12'h79B: dout <= 8'b00000000; // 1947 :   0 - 0x0
      12'h79C: dout <= 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout <= 8'b00000000; // 1949 :   0 - 0x0
      12'h79E: dout <= 8'b00000000; // 1950 :   0 - 0x0
      12'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      12'h7A0: dout <= 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0x7a
      12'h7A1: dout <= 8'b00000000; // 1953 :   0 - 0x0
      12'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      12'h7A3: dout <= 8'b00000000; // 1955 :   0 - 0x0
      12'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      12'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      12'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout <= 8'b00000000; // 1960 :   0 - 0x0 -- plane 1
      12'h7A9: dout <= 8'b00000000; // 1961 :   0 - 0x0
      12'h7AA: dout <= 8'b00000000; // 1962 :   0 - 0x0
      12'h7AB: dout <= 8'b00000000; // 1963 :   0 - 0x0
      12'h7AC: dout <= 8'b00000000; // 1964 :   0 - 0x0
      12'h7AD: dout <= 8'b00000000; // 1965 :   0 - 0x0
      12'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      12'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0x7b
      12'h7B1: dout <= 8'b00000000; // 1969 :   0 - 0x0
      12'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      12'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      12'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      12'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      12'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout <= 8'b00000000; // 1976 :   0 - 0x0 -- plane 1
      12'h7B9: dout <= 8'b00000000; // 1977 :   0 - 0x0
      12'h7BA: dout <= 8'b00000000; // 1978 :   0 - 0x0
      12'h7BB: dout <= 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout <= 8'b00000000; // 1982 :   0 - 0x0
      12'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout <= 8'b00100010; // 1984 :  34 - 0x22 -- Sprite 0x7c
      12'h7C1: dout <= 8'b01010101; // 1985 :  85 - 0x55
      12'h7C2: dout <= 8'b10101010; // 1986 : 170 - 0xaa
      12'h7C3: dout <= 8'b00000101; // 1987 :   5 - 0x5
      12'h7C4: dout <= 8'b00000100; // 1988 :   4 - 0x4
      12'h7C5: dout <= 8'b00001010; // 1989 :  10 - 0xa
      12'h7C6: dout <= 8'b01010000; // 1990 :  80 - 0x50
      12'h7C7: dout <= 8'b00000010; // 1991 :   2 - 0x2
      12'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0 -- plane 1
      12'h7C9: dout <= 8'b00100010; // 1993 :  34 - 0x22
      12'h7CA: dout <= 8'b01110111; // 1994 : 119 - 0x77
      12'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      12'h7CC: dout <= 8'b11111011; // 1996 : 251 - 0xfb
      12'h7CD: dout <= 8'b11110101; // 1997 : 245 - 0xf5
      12'h7CE: dout <= 8'b11101111; // 1998 : 239 - 0xef
      12'h7CF: dout <= 8'b11111111; // 1999 : 255 - 0xff
      12'h7D0: dout <= 8'b01110011; // 2000 : 115 - 0x73 -- Sprite 0x7d
      12'h7D1: dout <= 8'b11111111; // 2001 : 255 - 0xff
      12'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      12'h7D3: dout <= 8'b10111101; // 2003 : 189 - 0xbd
      12'h7D4: dout <= 8'b01101110; // 2004 : 110 - 0x6e
      12'h7D5: dout <= 8'b00001010; // 2005 :  10 - 0xa
      12'h7D6: dout <= 8'b01010000; // 2006 :  80 - 0x50
      12'h7D7: dout <= 8'b00000010; // 2007 :   2 - 0x2
      12'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0 -- plane 1
      12'h7D9: dout <= 8'b01110011; // 2009 : 115 - 0x73
      12'h7DA: dout <= 8'b11111111; // 2010 : 255 - 0xff
      12'h7DB: dout <= 8'b11111111; // 2011 : 255 - 0xff
      12'h7DC: dout <= 8'b11111011; // 2012 : 251 - 0xfb
      12'h7DD: dout <= 8'b11111101; // 2013 : 253 - 0xfd
      12'h7DE: dout <= 8'b11101111; // 2014 : 239 - 0xef
      12'h7DF: dout <= 8'b11111111; // 2015 : 255 - 0xff
      12'h7E0: dout <= 8'b00100000; // 2016 :  32 - 0x20 -- Sprite 0x7e
      12'h7E1: dout <= 8'b01010000; // 2017 :  80 - 0x50
      12'h7E2: dout <= 8'b10000100; // 2018 : 132 - 0x84
      12'h7E3: dout <= 8'b00000000; // 2019 :   0 - 0x0
      12'h7E4: dout <= 8'b00100100; // 2020 :  36 - 0x24
      12'h7E5: dout <= 8'b01011010; // 2021 :  90 - 0x5a
      12'h7E6: dout <= 8'b00010000; // 2022 :  16 - 0x10
      12'h7E7: dout <= 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout <= 8'b11011111; // 2024 : 223 - 0xdf -- plane 1
      12'h7E9: dout <= 8'b10101111; // 2025 : 175 - 0xaf
      12'h7EA: dout <= 8'b01111111; // 2026 : 127 - 0x7f
      12'h7EB: dout <= 8'b11111111; // 2027 : 255 - 0xff
      12'h7EC: dout <= 8'b11111011; // 2028 : 251 - 0xfb
      12'h7ED: dout <= 8'b11110101; // 2029 : 245 - 0xf5
      12'h7EE: dout <= 8'b11101111; // 2030 : 239 - 0xef
      12'h7EF: dout <= 8'b11111111; // 2031 : 255 - 0xff
      12'h7F0: dout <= 8'b11111111; // 2032 : 255 - 0xff -- Sprite 0x7f
      12'h7F1: dout <= 8'b01010000; // 2033 :  80 - 0x50
      12'h7F2: dout <= 8'b10000100; // 2034 : 132 - 0x84
      12'h7F3: dout <= 8'b00000000; // 2035 :   0 - 0x0
      12'h7F4: dout <= 8'b00100100; // 2036 :  36 - 0x24
      12'h7F5: dout <= 8'b01011010; // 2037 :  90 - 0x5a
      12'h7F6: dout <= 8'b00010000; // 2038 :  16 - 0x10
      12'h7F7: dout <= 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0 -- plane 1
      12'h7F9: dout <= 8'b10101111; // 2041 : 175 - 0xaf
      12'h7FA: dout <= 8'b01111111; // 2042 : 127 - 0x7f
      12'h7FB: dout <= 8'b11111111; // 2043 : 255 - 0xff
      12'h7FC: dout <= 8'b11111011; // 2044 : 251 - 0xfb
      12'h7FD: dout <= 8'b11110101; // 2045 : 245 - 0xf5
      12'h7FE: dout <= 8'b11101111; // 2046 : 239 - 0xef
      12'h7FF: dout <= 8'b11111111; // 2047 : 255 - 0xff
      12'h800: dout <= 8'b11111111; // 2048 : 255 - 0xff -- Sprite 0x80
      12'h801: dout <= 8'b10000000; // 2049 : 128 - 0x80
      12'h802: dout <= 8'b11001111; // 2050 : 207 - 0xcf
      12'h803: dout <= 8'b01001000; // 2051 :  72 - 0x48
      12'h804: dout <= 8'b11001111; // 2052 : 207 - 0xcf
      12'h805: dout <= 8'b10000000; // 2053 : 128 - 0x80
      12'h806: dout <= 8'b11001111; // 2054 : 207 - 0xcf
      12'h807: dout <= 8'b01001000; // 2055 :  72 - 0x48
      12'h808: dout <= 8'b00000000; // 2056 :   0 - 0x0 -- plane 1
      12'h809: dout <= 8'b01111111; // 2057 : 127 - 0x7f
      12'h80A: dout <= 8'b00110000; // 2058 :  48 - 0x30
      12'h80B: dout <= 8'b00110000; // 2059 :  48 - 0x30
      12'h80C: dout <= 8'b00110000; // 2060 :  48 - 0x30
      12'h80D: dout <= 8'b01111111; // 2061 : 127 - 0x7f
      12'h80E: dout <= 8'b00110000; // 2062 :  48 - 0x30
      12'h80F: dout <= 8'b00110000; // 2063 :  48 - 0x30
      12'h810: dout <= 8'b11111111; // 2064 : 255 - 0xff -- Sprite 0x81
      12'h811: dout <= 8'b10000000; // 2065 : 128 - 0x80
      12'h812: dout <= 8'b11111111; // 2066 : 255 - 0xff
      12'h813: dout <= 8'b10000000; // 2067 : 128 - 0x80
      12'h814: dout <= 8'b10000000; // 2068 : 128 - 0x80
      12'h815: dout <= 8'b11011111; // 2069 : 223 - 0xdf
      12'h816: dout <= 8'b10110000; // 2070 : 176 - 0xb0
      12'h817: dout <= 8'b11000000; // 2071 : 192 - 0xc0
      12'h818: dout <= 8'b00000000; // 2072 :   0 - 0x0 -- plane 1
      12'h819: dout <= 8'b01111111; // 2073 : 127 - 0x7f
      12'h81A: dout <= 8'b00000000; // 2074 :   0 - 0x0
      12'h81B: dout <= 8'b01111111; // 2075 : 127 - 0x7f
      12'h81C: dout <= 8'b01111111; // 2076 : 127 - 0x7f
      12'h81D: dout <= 8'b00100000; // 2077 :  32 - 0x20
      12'h81E: dout <= 8'b01000000; // 2078 :  64 - 0x40
      12'h81F: dout <= 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout <= 8'b11111111; // 2080 : 255 - 0xff -- Sprite 0x82
      12'h821: dout <= 8'b00000001; // 2081 :   1 - 0x1
      12'h822: dout <= 8'b11110011; // 2082 : 243 - 0xf3
      12'h823: dout <= 8'b00010010; // 2083 :  18 - 0x12
      12'h824: dout <= 8'b11110011; // 2084 : 243 - 0xf3
      12'h825: dout <= 8'b00000001; // 2085 :   1 - 0x1
      12'h826: dout <= 8'b11110011; // 2086 : 243 - 0xf3
      12'h827: dout <= 8'b00010010; // 2087 :  18 - 0x12
      12'h828: dout <= 8'b00000000; // 2088 :   0 - 0x0 -- plane 1
      12'h829: dout <= 8'b11111110; // 2089 : 254 - 0xfe
      12'h82A: dout <= 8'b00001100; // 2090 :  12 - 0xc
      12'h82B: dout <= 8'b00001100; // 2091 :  12 - 0xc
      12'h82C: dout <= 8'b00001100; // 2092 :  12 - 0xc
      12'h82D: dout <= 8'b11111110; // 2093 : 254 - 0xfe
      12'h82E: dout <= 8'b00001100; // 2094 :  12 - 0xc
      12'h82F: dout <= 8'b00001100; // 2095 :  12 - 0xc
      12'h830: dout <= 8'b11111111; // 2096 : 255 - 0xff -- Sprite 0x83
      12'h831: dout <= 8'b00000000; // 2097 :   0 - 0x0
      12'h832: dout <= 8'b11111111; // 2098 : 255 - 0xff
      12'h833: dout <= 8'b00000000; // 2099 :   0 - 0x0
      12'h834: dout <= 8'b00000000; // 2100 :   0 - 0x0
      12'h835: dout <= 8'b11111111; // 2101 : 255 - 0xff
      12'h836: dout <= 8'b00000000; // 2102 :   0 - 0x0
      12'h837: dout <= 8'b00000000; // 2103 :   0 - 0x0
      12'h838: dout <= 8'b00000000; // 2104 :   0 - 0x0 -- plane 1
      12'h839: dout <= 8'b11111111; // 2105 : 255 - 0xff
      12'h83A: dout <= 8'b00000000; // 2106 :   0 - 0x0
      12'h83B: dout <= 8'b11111111; // 2107 : 255 - 0xff
      12'h83C: dout <= 8'b11111111; // 2108 : 255 - 0xff
      12'h83D: dout <= 8'b00000000; // 2109 :   0 - 0x0
      12'h83E: dout <= 8'b00000000; // 2110 :   0 - 0x0
      12'h83F: dout <= 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout <= 8'b11111111; // 2112 : 255 - 0xff -- Sprite 0x84
      12'h841: dout <= 8'b10000010; // 2113 : 130 - 0x82
      12'h842: dout <= 8'b00010000; // 2114 :  16 - 0x10
      12'h843: dout <= 8'b00000000; // 2115 :   0 - 0x0
      12'h844: dout <= 8'b00000000; // 2116 :   0 - 0x0
      12'h845: dout <= 8'b00010000; // 2117 :  16 - 0x10
      12'h846: dout <= 8'b01000100; // 2118 :  68 - 0x44
      12'h847: dout <= 8'b11111111; // 2119 : 255 - 0xff
      12'h848: dout <= 8'b00000000; // 2120 :   0 - 0x0 -- plane 1
      12'h849: dout <= 8'b11111111; // 2121 : 255 - 0xff
      12'h84A: dout <= 8'b11111111; // 2122 : 255 - 0xff
      12'h84B: dout <= 8'b11111111; // 2123 : 255 - 0xff
      12'h84C: dout <= 8'b11111111; // 2124 : 255 - 0xff
      12'h84D: dout <= 8'b11101111; // 2125 : 239 - 0xef
      12'h84E: dout <= 8'b10111011; // 2126 : 187 - 0xbb
      12'h84F: dout <= 8'b00000000; // 2127 :   0 - 0x0
      12'h850: dout <= 8'b11111111; // 2128 : 255 - 0xff -- Sprite 0x85
      12'h851: dout <= 8'b00000001; // 2129 :   1 - 0x1
      12'h852: dout <= 8'b11111111; // 2130 : 255 - 0xff
      12'h853: dout <= 8'b00000001; // 2131 :   1 - 0x1
      12'h854: dout <= 8'b00000001; // 2132 :   1 - 0x1
      12'h855: dout <= 8'b11110011; // 2133 : 243 - 0xf3
      12'h856: dout <= 8'b00001101; // 2134 :  13 - 0xd
      12'h857: dout <= 8'b00000011; // 2135 :   3 - 0x3
      12'h858: dout <= 8'b00000000; // 2136 :   0 - 0x0 -- plane 1
      12'h859: dout <= 8'b11111110; // 2137 : 254 - 0xfe
      12'h85A: dout <= 8'b00000000; // 2138 :   0 - 0x0
      12'h85B: dout <= 8'b11111110; // 2139 : 254 - 0xfe
      12'h85C: dout <= 8'b11111110; // 2140 : 254 - 0xfe
      12'h85D: dout <= 8'b00001100; // 2141 :  12 - 0xc
      12'h85E: dout <= 8'b00000010; // 2142 :   2 - 0x2
      12'h85F: dout <= 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout <= 8'b00000000; // 2144 :   0 - 0x0 -- Sprite 0x86
      12'h861: dout <= 8'b00000000; // 2145 :   0 - 0x0
      12'h862: dout <= 8'b00000000; // 2146 :   0 - 0x0
      12'h863: dout <= 8'b00000000; // 2147 :   0 - 0x0
      12'h864: dout <= 8'b00000000; // 2148 :   0 - 0x0
      12'h865: dout <= 8'b00000000; // 2149 :   0 - 0x0
      12'h866: dout <= 8'b00000000; // 2150 :   0 - 0x0
      12'h867: dout <= 8'b00000000; // 2151 :   0 - 0x0
      12'h868: dout <= 8'b00000000; // 2152 :   0 - 0x0 -- plane 1
      12'h869: dout <= 8'b00000000; // 2153 :   0 - 0x0
      12'h86A: dout <= 8'b00000000; // 2154 :   0 - 0x0
      12'h86B: dout <= 8'b00000000; // 2155 :   0 - 0x0
      12'h86C: dout <= 8'b00000000; // 2156 :   0 - 0x0
      12'h86D: dout <= 8'b00000000; // 2157 :   0 - 0x0
      12'h86E: dout <= 8'b00000000; // 2158 :   0 - 0x0
      12'h86F: dout <= 8'b00000000; // 2159 :   0 - 0x0
      12'h870: dout <= 8'b00000000; // 2160 :   0 - 0x0 -- Sprite 0x87
      12'h871: dout <= 8'b00000000; // 2161 :   0 - 0x0
      12'h872: dout <= 8'b00000000; // 2162 :   0 - 0x0
      12'h873: dout <= 8'b00000000; // 2163 :   0 - 0x0
      12'h874: dout <= 8'b00000000; // 2164 :   0 - 0x0
      12'h875: dout <= 8'b00000000; // 2165 :   0 - 0x0
      12'h876: dout <= 8'b00000000; // 2166 :   0 - 0x0
      12'h877: dout <= 8'b00000000; // 2167 :   0 - 0x0
      12'h878: dout <= 8'b00000000; // 2168 :   0 - 0x0 -- plane 1
      12'h879: dout <= 8'b00000000; // 2169 :   0 - 0x0
      12'h87A: dout <= 8'b00000000; // 2170 :   0 - 0x0
      12'h87B: dout <= 8'b00000000; // 2171 :   0 - 0x0
      12'h87C: dout <= 8'b00000000; // 2172 :   0 - 0x0
      12'h87D: dout <= 8'b00000000; // 2173 :   0 - 0x0
      12'h87E: dout <= 8'b00000000; // 2174 :   0 - 0x0
      12'h87F: dout <= 8'b00000000; // 2175 :   0 - 0x0
      12'h880: dout <= 8'b00000111; // 2176 :   7 - 0x7 -- Sprite 0x88
      12'h881: dout <= 8'b00011110; // 2177 :  30 - 0x1e
      12'h882: dout <= 8'b00101111; // 2178 :  47 - 0x2f
      12'h883: dout <= 8'b01010011; // 2179 :  83 - 0x53
      12'h884: dout <= 8'b01101110; // 2180 : 110 - 0x6e
      12'h885: dout <= 8'b11011011; // 2181 : 219 - 0xdb
      12'h886: dout <= 8'b11111010; // 2182 : 250 - 0xfa
      12'h887: dout <= 8'b11010101; // 2183 : 213 - 0xd5
      12'h888: dout <= 8'b00000000; // 2184 :   0 - 0x0 -- plane 1
      12'h889: dout <= 8'b00000111; // 2185 :   7 - 0x7
      12'h88A: dout <= 8'b00011111; // 2186 :  31 - 0x1f
      12'h88B: dout <= 8'b00111100; // 2187 :  60 - 0x3c
      12'h88C: dout <= 8'b00110001; // 2188 :  49 - 0x31
      12'h88D: dout <= 8'b01110100; // 2189 : 116 - 0x74
      12'h88E: dout <= 8'b01100101; // 2190 : 101 - 0x65
      12'h88F: dout <= 8'b01101010; // 2191 : 106 - 0x6a
      12'h890: dout <= 8'b10111011; // 2192 : 187 - 0xbb -- Sprite 0x89
      12'h891: dout <= 8'b11110010; // 2193 : 242 - 0xf2
      12'h892: dout <= 8'b11011101; // 2194 : 221 - 0xdd
      12'h893: dout <= 8'b01001111; // 2195 :  79 - 0x4f
      12'h894: dout <= 8'b01111011; // 2196 : 123 - 0x7b
      12'h895: dout <= 8'b00110010; // 2197 :  50 - 0x32
      12'h896: dout <= 8'b00011111; // 2198 :  31 - 0x1f
      12'h897: dout <= 8'b00000111; // 2199 :   7 - 0x7
      12'h898: dout <= 8'b01100100; // 2200 : 100 - 0x64 -- plane 1
      12'h899: dout <= 8'b01101101; // 2201 : 109 - 0x6d
      12'h89A: dout <= 8'b01110010; // 2202 : 114 - 0x72
      12'h89B: dout <= 8'b00110000; // 2203 :  48 - 0x30
      12'h89C: dout <= 8'b00111100; // 2204 :  60 - 0x3c
      12'h89D: dout <= 8'b00011111; // 2205 :  31 - 0x1f
      12'h89E: dout <= 8'b00000111; // 2206 :   7 - 0x7
      12'h89F: dout <= 8'b00000000; // 2207 :   0 - 0x0
      12'h8A0: dout <= 8'b11100000; // 2208 : 224 - 0xe0 -- Sprite 0x8a
      12'h8A1: dout <= 8'b11011000; // 2209 : 216 - 0xd8
      12'h8A2: dout <= 8'b01010100; // 2210 :  84 - 0x54
      12'h8A3: dout <= 8'b11101010; // 2211 : 234 - 0xea
      12'h8A4: dout <= 8'b10111010; // 2212 : 186 - 0xba
      12'h8A5: dout <= 8'b10010011; // 2213 : 147 - 0x93
      12'h8A6: dout <= 8'b11011111; // 2214 : 223 - 0xdf
      12'h8A7: dout <= 8'b10111101; // 2215 : 189 - 0xbd
      12'h8A8: dout <= 8'b00000000; // 2216 :   0 - 0x0 -- plane 1
      12'h8A9: dout <= 8'b11100000; // 2217 : 224 - 0xe0
      12'h8AA: dout <= 8'b11111000; // 2218 : 248 - 0xf8
      12'h8AB: dout <= 8'b00111100; // 2219 :  60 - 0x3c
      12'h8AC: dout <= 8'b01001100; // 2220 :  76 - 0x4c
      12'h8AD: dout <= 8'b01101110; // 2221 : 110 - 0x6e
      12'h8AE: dout <= 8'b00100110; // 2222 :  38 - 0x26
      12'h8AF: dout <= 8'b01000110; // 2223 :  70 - 0x46
      12'h8B0: dout <= 8'b01101011; // 2224 : 107 - 0x6b -- Sprite 0x8b
      12'h8B1: dout <= 8'b10011111; // 2225 : 159 - 0x9f
      12'h8B2: dout <= 8'b01011101; // 2226 :  93 - 0x5d
      12'h8B3: dout <= 8'b10110110; // 2227 : 182 - 0xb6
      12'h8B4: dout <= 8'b11101010; // 2228 : 234 - 0xea
      12'h8B5: dout <= 8'b11001100; // 2229 : 204 - 0xcc
      12'h8B6: dout <= 8'b01111000; // 2230 : 120 - 0x78
      12'h8B7: dout <= 8'b11100000; // 2231 : 224 - 0xe0
      12'h8B8: dout <= 8'b10010110; // 2232 : 150 - 0x96 -- plane 1
      12'h8B9: dout <= 8'b01100110; // 2233 : 102 - 0x66
      12'h8BA: dout <= 8'b10101110; // 2234 : 174 - 0xae
      12'h8BB: dout <= 8'b01001100; // 2235 :  76 - 0x4c
      12'h8BC: dout <= 8'b00111100; // 2236 :  60 - 0x3c
      12'h8BD: dout <= 8'b11111000; // 2237 : 248 - 0xf8
      12'h8BE: dout <= 8'b11100000; // 2238 : 224 - 0xe0
      12'h8BF: dout <= 8'b00000000; // 2239 :   0 - 0x0
      12'h8C0: dout <= 8'b00000111; // 2240 :   7 - 0x7 -- Sprite 0x8c
      12'h8C1: dout <= 8'b00011000; // 2241 :  24 - 0x18
      12'h8C2: dout <= 8'b00100011; // 2242 :  35 - 0x23
      12'h8C3: dout <= 8'b01001100; // 2243 :  76 - 0x4c
      12'h8C4: dout <= 8'b01110000; // 2244 : 112 - 0x70
      12'h8C5: dout <= 8'b10100001; // 2245 : 161 - 0xa1
      12'h8C6: dout <= 8'b10100110; // 2246 : 166 - 0xa6
      12'h8C7: dout <= 8'b10101000; // 2247 : 168 - 0xa8
      12'h8C8: dout <= 8'b00000000; // 2248 :   0 - 0x0 -- plane 1
      12'h8C9: dout <= 8'b00000111; // 2249 :   7 - 0x7
      12'h8CA: dout <= 8'b00011111; // 2250 :  31 - 0x1f
      12'h8CB: dout <= 8'b00111111; // 2251 :  63 - 0x3f
      12'h8CC: dout <= 8'b00111111; // 2252 :  63 - 0x3f
      12'h8CD: dout <= 8'b01111111; // 2253 : 127 - 0x7f
      12'h8CE: dout <= 8'b01111111; // 2254 : 127 - 0x7f
      12'h8CF: dout <= 8'b01111111; // 2255 : 127 - 0x7f
      12'h8D0: dout <= 8'b10100101; // 2256 : 165 - 0xa5 -- Sprite 0x8d
      12'h8D1: dout <= 8'b10100010; // 2257 : 162 - 0xa2
      12'h8D2: dout <= 8'b10010000; // 2258 : 144 - 0x90
      12'h8D3: dout <= 8'b01001000; // 2259 :  72 - 0x48
      12'h8D4: dout <= 8'b01000111; // 2260 :  71 - 0x47
      12'h8D5: dout <= 8'b00100000; // 2261 :  32 - 0x20
      12'h8D6: dout <= 8'b00011001; // 2262 :  25 - 0x19
      12'h8D7: dout <= 8'b00000111; // 2263 :   7 - 0x7
      12'h8D8: dout <= 8'b01111111; // 2264 : 127 - 0x7f -- plane 1
      12'h8D9: dout <= 8'b01111111; // 2265 : 127 - 0x7f
      12'h8DA: dout <= 8'b01111111; // 2266 : 127 - 0x7f
      12'h8DB: dout <= 8'b00111111; // 2267 :  63 - 0x3f
      12'h8DC: dout <= 8'b00111111; // 2268 :  63 - 0x3f
      12'h8DD: dout <= 8'b00011111; // 2269 :  31 - 0x1f
      12'h8DE: dout <= 8'b00000111; // 2270 :   7 - 0x7
      12'h8DF: dout <= 8'b00000000; // 2271 :   0 - 0x0
      12'h8E0: dout <= 8'b11100000; // 2272 : 224 - 0xe0 -- Sprite 0x8e
      12'h8E1: dout <= 8'b00011000; // 2273 :  24 - 0x18
      12'h8E2: dout <= 8'b00000100; // 2274 :   4 - 0x4
      12'h8E3: dout <= 8'b11000010; // 2275 : 194 - 0xc2
      12'h8E4: dout <= 8'b00110010; // 2276 :  50 - 0x32
      12'h8E5: dout <= 8'b00001001; // 2277 :   9 - 0x9
      12'h8E6: dout <= 8'b11000101; // 2278 : 197 - 0xc5
      12'h8E7: dout <= 8'b00100101; // 2279 :  37 - 0x25
      12'h8E8: dout <= 8'b00000000; // 2280 :   0 - 0x0 -- plane 1
      12'h8E9: dout <= 8'b11100000; // 2281 : 224 - 0xe0
      12'h8EA: dout <= 8'b11111000; // 2282 : 248 - 0xf8
      12'h8EB: dout <= 8'b11111100; // 2283 : 252 - 0xfc
      12'h8EC: dout <= 8'b11111100; // 2284 : 252 - 0xfc
      12'h8ED: dout <= 8'b11111110; // 2285 : 254 - 0xfe
      12'h8EE: dout <= 8'b11111110; // 2286 : 254 - 0xfe
      12'h8EF: dout <= 8'b11111110; // 2287 : 254 - 0xfe
      12'h8F0: dout <= 8'b10100101; // 2288 : 165 - 0xa5 -- Sprite 0x8f
      12'h8F1: dout <= 8'b01100101; // 2289 : 101 - 0x65
      12'h8F2: dout <= 8'b01000101; // 2290 :  69 - 0x45
      12'h8F3: dout <= 8'b10001010; // 2291 : 138 - 0x8a
      12'h8F4: dout <= 8'b10010010; // 2292 : 146 - 0x92
      12'h8F5: dout <= 8'b00100100; // 2293 :  36 - 0x24
      12'h8F6: dout <= 8'b11011000; // 2294 : 216 - 0xd8
      12'h8F7: dout <= 8'b11100000; // 2295 : 224 - 0xe0
      12'h8F8: dout <= 8'b11111110; // 2296 : 254 - 0xfe -- plane 1
      12'h8F9: dout <= 8'b11111110; // 2297 : 254 - 0xfe
      12'h8FA: dout <= 8'b11111110; // 2298 : 254 - 0xfe
      12'h8FB: dout <= 8'b11111100; // 2299 : 252 - 0xfc
      12'h8FC: dout <= 8'b11111100; // 2300 : 252 - 0xfc
      12'h8FD: dout <= 8'b11111000; // 2301 : 248 - 0xf8
      12'h8FE: dout <= 8'b11100000; // 2302 : 224 - 0xe0
      12'h8FF: dout <= 8'b00000000; // 2303 :   0 - 0x0
      12'h900: dout <= 8'b00000000; // 2304 :   0 - 0x0 -- Sprite 0x90
      12'h901: dout <= 8'b00000000; // 2305 :   0 - 0x0
      12'h902: dout <= 8'b00100000; // 2306 :  32 - 0x20
      12'h903: dout <= 8'b00110000; // 2307 :  48 - 0x30
      12'h904: dout <= 8'b00101100; // 2308 :  44 - 0x2c
      12'h905: dout <= 8'b00100010; // 2309 :  34 - 0x22
      12'h906: dout <= 8'b00010001; // 2310 :  17 - 0x11
      12'h907: dout <= 8'b00001000; // 2311 :   8 - 0x8
      12'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0 -- plane 1
      12'h909: dout <= 8'b00000000; // 2313 :   0 - 0x0
      12'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout <= 8'b00000000; // 2315 :   0 - 0x0
      12'h90C: dout <= 8'b00010000; // 2316 :  16 - 0x10
      12'h90D: dout <= 8'b00011100; // 2317 :  28 - 0x1c
      12'h90E: dout <= 8'b00001110; // 2318 :  14 - 0xe
      12'h90F: dout <= 8'b00000111; // 2319 :   7 - 0x7
      12'h910: dout <= 8'b00000100; // 2320 :   4 - 0x4 -- Sprite 0x91
      12'h911: dout <= 8'b11110010; // 2321 : 242 - 0xf2
      12'h912: dout <= 8'b11001111; // 2322 : 207 - 0xcf
      12'h913: dout <= 8'b00110000; // 2323 :  48 - 0x30
      12'h914: dout <= 8'b00001100; // 2324 :  12 - 0xc
      12'h915: dout <= 8'b11111111; // 2325 : 255 - 0xff
      12'h916: dout <= 8'b10000000; // 2326 : 128 - 0x80
      12'h917: dout <= 8'b11111111; // 2327 : 255 - 0xff
      12'h918: dout <= 8'b00000011; // 2328 :   3 - 0x3 -- plane 1
      12'h919: dout <= 8'b00000001; // 2329 :   1 - 0x1
      12'h91A: dout <= 8'b00110000; // 2330 :  48 - 0x30
      12'h91B: dout <= 8'b00001111; // 2331 :  15 - 0xf
      12'h91C: dout <= 8'b00000011; // 2332 :   3 - 0x3
      12'h91D: dout <= 8'b00000000; // 2333 :   0 - 0x0
      12'h91E: dout <= 8'b01111111; // 2334 : 127 - 0x7f
      12'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout <= 8'b01000010; // 2336 :  66 - 0x42 -- Sprite 0x92
      12'h921: dout <= 8'b10100101; // 2337 : 165 - 0xa5
      12'h922: dout <= 8'b10100101; // 2338 : 165 - 0xa5
      12'h923: dout <= 8'b10011001; // 2339 : 153 - 0x99
      12'h924: dout <= 8'b10011001; // 2340 : 153 - 0x99
      12'h925: dout <= 8'b10011001; // 2341 : 153 - 0x99
      12'h926: dout <= 8'b00000001; // 2342 :   1 - 0x1
      12'h927: dout <= 8'b00000000; // 2343 :   0 - 0x0
      12'h928: dout <= 8'b00000000; // 2344 :   0 - 0x0 -- plane 1
      12'h929: dout <= 8'b01000010; // 2345 :  66 - 0x42
      12'h92A: dout <= 8'b01000010; // 2346 :  66 - 0x42
      12'h92B: dout <= 8'b01100110; // 2347 : 102 - 0x66
      12'h92C: dout <= 8'b01100110; // 2348 : 102 - 0x66
      12'h92D: dout <= 8'b01100110; // 2349 : 102 - 0x66
      12'h92E: dout <= 8'b11111110; // 2350 : 254 - 0xfe
      12'h92F: dout <= 8'b11111111; // 2351 : 255 - 0xff
      12'h930: dout <= 8'b11111111; // 2352 : 255 - 0xff -- Sprite 0x93
      12'h931: dout <= 8'b11111111; // 2353 : 255 - 0xff
      12'h932: dout <= 8'b11111111; // 2354 : 255 - 0xff
      12'h933: dout <= 8'b10000001; // 2355 : 129 - 0x81
      12'h934: dout <= 8'b11111111; // 2356 : 255 - 0xff
      12'h935: dout <= 8'b11111111; // 2357 : 255 - 0xff
      12'h936: dout <= 8'b11111111; // 2358 : 255 - 0xff
      12'h937: dout <= 8'b10000001; // 2359 : 129 - 0x81
      12'h938: dout <= 8'b01111110; // 2360 : 126 - 0x7e -- plane 1
      12'h939: dout <= 8'b01111110; // 2361 : 126 - 0x7e
      12'h93A: dout <= 8'b01111110; // 2362 : 126 - 0x7e
      12'h93B: dout <= 8'b01111110; // 2363 : 126 - 0x7e
      12'h93C: dout <= 8'b01111110; // 2364 : 126 - 0x7e
      12'h93D: dout <= 8'b01111110; // 2365 : 126 - 0x7e
      12'h93E: dout <= 8'b01111110; // 2366 : 126 - 0x7e
      12'h93F: dout <= 8'b01111110; // 2367 : 126 - 0x7e
      12'h940: dout <= 8'b00000000; // 2368 :   0 - 0x0 -- Sprite 0x94
      12'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout <= 8'b00000100; // 2370 :   4 - 0x4
      12'h943: dout <= 8'b00001100; // 2371 :  12 - 0xc
      12'h944: dout <= 8'b00110100; // 2372 :  52 - 0x34
      12'h945: dout <= 8'b01000100; // 2373 :  68 - 0x44
      12'h946: dout <= 8'b10001000; // 2374 : 136 - 0x88
      12'h947: dout <= 8'b00010000; // 2375 :  16 - 0x10
      12'h948: dout <= 8'b00000000; // 2376 :   0 - 0x0 -- plane 1
      12'h949: dout <= 8'b00000000; // 2377 :   0 - 0x0
      12'h94A: dout <= 8'b00000000; // 2378 :   0 - 0x0
      12'h94B: dout <= 8'b00000000; // 2379 :   0 - 0x0
      12'h94C: dout <= 8'b00001000; // 2380 :   8 - 0x8
      12'h94D: dout <= 8'b00111000; // 2381 :  56 - 0x38
      12'h94E: dout <= 8'b01110000; // 2382 : 112 - 0x70
      12'h94F: dout <= 8'b11100000; // 2383 : 224 - 0xe0
      12'h950: dout <= 8'b00100000; // 2384 :  32 - 0x20 -- Sprite 0x95
      12'h951: dout <= 8'b01001111; // 2385 :  79 - 0x4f
      12'h952: dout <= 8'b11110011; // 2386 : 243 - 0xf3
      12'h953: dout <= 8'b00001100; // 2387 :  12 - 0xc
      12'h954: dout <= 8'b00110000; // 2388 :  48 - 0x30
      12'h955: dout <= 8'b11111111; // 2389 : 255 - 0xff
      12'h956: dout <= 8'b00000001; // 2390 :   1 - 0x1
      12'h957: dout <= 8'b11111111; // 2391 : 255 - 0xff
      12'h958: dout <= 8'b11000000; // 2392 : 192 - 0xc0 -- plane 1
      12'h959: dout <= 8'b10000000; // 2393 : 128 - 0x80
      12'h95A: dout <= 8'b00001100; // 2394 :  12 - 0xc
      12'h95B: dout <= 8'b11110000; // 2395 : 240 - 0xf0
      12'h95C: dout <= 8'b11000000; // 2396 : 192 - 0xc0
      12'h95D: dout <= 8'b00000000; // 2397 :   0 - 0x0
      12'h95E: dout <= 8'b11111110; // 2398 : 254 - 0xfe
      12'h95F: dout <= 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout <= 8'b01111111; // 2400 : 127 - 0x7f -- Sprite 0x96
      12'h961: dout <= 8'b11111111; // 2401 : 255 - 0xff
      12'h962: dout <= 8'b11111111; // 2402 : 255 - 0xff
      12'h963: dout <= 8'b11111111; // 2403 : 255 - 0xff
      12'h964: dout <= 8'b11111011; // 2404 : 251 - 0xfb
      12'h965: dout <= 8'b11111111; // 2405 : 255 - 0xff
      12'h966: dout <= 8'b11111111; // 2406 : 255 - 0xff
      12'h967: dout <= 8'b11111111; // 2407 : 255 - 0xff
      12'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0 -- plane 1
      12'h969: dout <= 8'b00111111; // 2409 :  63 - 0x3f
      12'h96A: dout <= 8'b01111111; // 2410 : 127 - 0x7f
      12'h96B: dout <= 8'b01111111; // 2411 : 127 - 0x7f
      12'h96C: dout <= 8'b01111111; // 2412 : 127 - 0x7f
      12'h96D: dout <= 8'b01111111; // 2413 : 127 - 0x7f
      12'h96E: dout <= 8'b01111111; // 2414 : 127 - 0x7f
      12'h96F: dout <= 8'b01111111; // 2415 : 127 - 0x7f
      12'h970: dout <= 8'b11111111; // 2416 : 255 - 0xff -- Sprite 0x97
      12'h971: dout <= 8'b11111111; // 2417 : 255 - 0xff
      12'h972: dout <= 8'b11111111; // 2418 : 255 - 0xff
      12'h973: dout <= 8'b11111111; // 2419 : 255 - 0xff
      12'h974: dout <= 8'b11111111; // 2420 : 255 - 0xff
      12'h975: dout <= 8'b11111111; // 2421 : 255 - 0xff
      12'h976: dout <= 8'b11111110; // 2422 : 254 - 0xfe
      12'h977: dout <= 8'b11111111; // 2423 : 255 - 0xff
      12'h978: dout <= 8'b01111111; // 2424 : 127 - 0x7f -- plane 1
      12'h979: dout <= 8'b01111111; // 2425 : 127 - 0x7f
      12'h97A: dout <= 8'b00111111; // 2426 :  63 - 0x3f
      12'h97B: dout <= 8'b01111111; // 2427 : 127 - 0x7f
      12'h97C: dout <= 8'b01111111; // 2428 : 127 - 0x7f
      12'h97D: dout <= 8'b01111111; // 2429 : 127 - 0x7f
      12'h97E: dout <= 8'b01111111; // 2430 : 127 - 0x7f
      12'h97F: dout <= 8'b01111111; // 2431 : 127 - 0x7f
      12'h980: dout <= 8'b11111111; // 2432 : 255 - 0xff -- Sprite 0x98
      12'h981: dout <= 8'b10111111; // 2433 : 191 - 0xbf
      12'h982: dout <= 8'b11111111; // 2434 : 255 - 0xff
      12'h983: dout <= 8'b11111111; // 2435 : 255 - 0xff
      12'h984: dout <= 8'b11111011; // 2436 : 251 - 0xfb
      12'h985: dout <= 8'b11111111; // 2437 : 255 - 0xff
      12'h986: dout <= 8'b11111111; // 2438 : 255 - 0xff
      12'h987: dout <= 8'b11111111; // 2439 : 255 - 0xff
      12'h988: dout <= 8'b00000000; // 2440 :   0 - 0x0 -- plane 1
      12'h989: dout <= 8'b11011111; // 2441 : 223 - 0xdf
      12'h98A: dout <= 8'b11111111; // 2442 : 255 - 0xff
      12'h98B: dout <= 8'b11111111; // 2443 : 255 - 0xff
      12'h98C: dout <= 8'b11111111; // 2444 : 255 - 0xff
      12'h98D: dout <= 8'b11111111; // 2445 : 255 - 0xff
      12'h98E: dout <= 8'b11111111; // 2446 : 255 - 0xff
      12'h98F: dout <= 8'b11111111; // 2447 : 255 - 0xff
      12'h990: dout <= 8'b11111111; // 2448 : 255 - 0xff -- Sprite 0x99
      12'h991: dout <= 8'b11111111; // 2449 : 255 - 0xff
      12'h992: dout <= 8'b11111111; // 2450 : 255 - 0xff
      12'h993: dout <= 8'b11111111; // 2451 : 255 - 0xff
      12'h994: dout <= 8'b11111111; // 2452 : 255 - 0xff
      12'h995: dout <= 8'b11111111; // 2453 : 255 - 0xff
      12'h996: dout <= 8'b11111110; // 2454 : 254 - 0xfe
      12'h997: dout <= 8'b11111111; // 2455 : 255 - 0xff
      12'h998: dout <= 8'b11111111; // 2456 : 255 - 0xff -- plane 1
      12'h999: dout <= 8'b11111111; // 2457 : 255 - 0xff
      12'h99A: dout <= 8'b10111111; // 2458 : 191 - 0xbf
      12'h99B: dout <= 8'b11111111; // 2459 : 255 - 0xff
      12'h99C: dout <= 8'b11111111; // 2460 : 255 - 0xff
      12'h99D: dout <= 8'b11111111; // 2461 : 255 - 0xff
      12'h99E: dout <= 8'b11111111; // 2462 : 255 - 0xff
      12'h99F: dout <= 8'b11111111; // 2463 : 255 - 0xff
      12'h9A0: dout <= 8'b11111110; // 2464 : 254 - 0xfe -- Sprite 0x9a
      12'h9A1: dout <= 8'b11111111; // 2465 : 255 - 0xff
      12'h9A2: dout <= 8'b11111111; // 2466 : 255 - 0xff
      12'h9A3: dout <= 8'b11111111; // 2467 : 255 - 0xff
      12'h9A4: dout <= 8'b11111011; // 2468 : 251 - 0xfb
      12'h9A5: dout <= 8'b11111111; // 2469 : 255 - 0xff
      12'h9A6: dout <= 8'b11111111; // 2470 : 255 - 0xff
      12'h9A7: dout <= 8'b11111111; // 2471 : 255 - 0xff
      12'h9A8: dout <= 8'b00000000; // 2472 :   0 - 0x0 -- plane 1
      12'h9A9: dout <= 8'b10111100; // 2473 : 188 - 0xbc
      12'h9AA: dout <= 8'b11111110; // 2474 : 254 - 0xfe
      12'h9AB: dout <= 8'b11111110; // 2475 : 254 - 0xfe
      12'h9AC: dout <= 8'b11111110; // 2476 : 254 - 0xfe
      12'h9AD: dout <= 8'b11111110; // 2477 : 254 - 0xfe
      12'h9AE: dout <= 8'b11111110; // 2478 : 254 - 0xfe
      12'h9AF: dout <= 8'b11111110; // 2479 : 254 - 0xfe
      12'h9B0: dout <= 8'b11111111; // 2480 : 255 - 0xff -- Sprite 0x9b
      12'h9B1: dout <= 8'b11111111; // 2481 : 255 - 0xff
      12'h9B2: dout <= 8'b11111111; // 2482 : 255 - 0xff
      12'h9B3: dout <= 8'b11111111; // 2483 : 255 - 0xff
      12'h9B4: dout <= 8'b11111111; // 2484 : 255 - 0xff
      12'h9B5: dout <= 8'b11111111; // 2485 : 255 - 0xff
      12'h9B6: dout <= 8'b11111111; // 2486 : 255 - 0xff
      12'h9B7: dout <= 8'b11111111; // 2487 : 255 - 0xff
      12'h9B8: dout <= 8'b11111110; // 2488 : 254 - 0xfe -- plane 1
      12'h9B9: dout <= 8'b11111110; // 2489 : 254 - 0xfe
      12'h9BA: dout <= 8'b10111110; // 2490 : 190 - 0xbe
      12'h9BB: dout <= 8'b11111110; // 2491 : 254 - 0xfe
      12'h9BC: dout <= 8'b11111110; // 2492 : 254 - 0xfe
      12'h9BD: dout <= 8'b11111110; // 2493 : 254 - 0xfe
      12'h9BE: dout <= 8'b11111110; // 2494 : 254 - 0xfe
      12'h9BF: dout <= 8'b11111110; // 2495 : 254 - 0xfe
      12'h9C0: dout <= 8'b11111111; // 2496 : 255 - 0xff -- Sprite 0x9c
      12'h9C1: dout <= 8'b11111111; // 2497 : 255 - 0xff
      12'h9C2: dout <= 8'b10100000; // 2498 : 160 - 0xa0
      12'h9C3: dout <= 8'b10010000; // 2499 : 144 - 0x90
      12'h9C4: dout <= 8'b10001000; // 2500 : 136 - 0x88
      12'h9C5: dout <= 8'b10000100; // 2501 : 132 - 0x84
      12'h9C6: dout <= 8'b01101010; // 2502 : 106 - 0x6a
      12'h9C7: dout <= 8'b00111111; // 2503 :  63 - 0x3f
      12'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0 -- plane 1
      12'h9C9: dout <= 8'b00111111; // 2505 :  63 - 0x3f
      12'h9CA: dout <= 8'b01011111; // 2506 :  95 - 0x5f
      12'h9CB: dout <= 8'b01101111; // 2507 : 111 - 0x6f
      12'h9CC: dout <= 8'b01110111; // 2508 : 119 - 0x77
      12'h9CD: dout <= 8'b01111011; // 2509 : 123 - 0x7b
      12'h9CE: dout <= 8'b00010101; // 2510 :  21 - 0x15
      12'h9CF: dout <= 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout <= 8'b11111111; // 2512 : 255 - 0xff -- Sprite 0x9d
      12'h9D1: dout <= 8'b11111111; // 2513 : 255 - 0xff
      12'h9D2: dout <= 8'b00100001; // 2514 :  33 - 0x21
      12'h9D3: dout <= 8'b00010001; // 2515 :  17 - 0x11
      12'h9D4: dout <= 8'b00001001; // 2516 :   9 - 0x9
      12'h9D5: dout <= 8'b00000101; // 2517 :   5 - 0x5
      12'h9D6: dout <= 8'b10101010; // 2518 : 170 - 0xaa
      12'h9D7: dout <= 8'b11111100; // 2519 : 252 - 0xfc
      12'h9D8: dout <= 8'b00000000; // 2520 :   0 - 0x0 -- plane 1
      12'h9D9: dout <= 8'b10111110; // 2521 : 190 - 0xbe
      12'h9DA: dout <= 8'b11011110; // 2522 : 222 - 0xde
      12'h9DB: dout <= 8'b11101110; // 2523 : 238 - 0xee
      12'h9DC: dout <= 8'b11110110; // 2524 : 246 - 0xf6
      12'h9DD: dout <= 8'b11111010; // 2525 : 250 - 0xfa
      12'h9DE: dout <= 8'b01010100; // 2526 :  84 - 0x54
      12'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout <= 8'b11111111; // 2528 : 255 - 0xff -- Sprite 0x9e
      12'h9E1: dout <= 8'b11111111; // 2529 : 255 - 0xff
      12'h9E2: dout <= 8'b00100000; // 2530 :  32 - 0x20
      12'h9E3: dout <= 8'b00010000; // 2531 :  16 - 0x10
      12'h9E4: dout <= 8'b00001000; // 2532 :   8 - 0x8
      12'h9E5: dout <= 8'b00000100; // 2533 :   4 - 0x4
      12'h9E6: dout <= 8'b10101010; // 2534 : 170 - 0xaa
      12'h9E7: dout <= 8'b11111111; // 2535 : 255 - 0xff
      12'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0 -- plane 1
      12'h9E9: dout <= 8'b10111111; // 2537 : 191 - 0xbf
      12'h9EA: dout <= 8'b11011111; // 2538 : 223 - 0xdf
      12'h9EB: dout <= 8'b11101111; // 2539 : 239 - 0xef
      12'h9EC: dout <= 8'b11110111; // 2540 : 247 - 0xf7
      12'h9ED: dout <= 8'b11111011; // 2541 : 251 - 0xfb
      12'h9EE: dout <= 8'b01010101; // 2542 :  85 - 0x55
      12'h9EF: dout <= 8'b00000000; // 2543 :   0 - 0x0
      12'h9F0: dout <= 8'b00000000; // 2544 :   0 - 0x0 -- Sprite 0x9f
      12'h9F1: dout <= 8'b00000000; // 2545 :   0 - 0x0
      12'h9F2: dout <= 8'b00000000; // 2546 :   0 - 0x0
      12'h9F3: dout <= 8'b00000000; // 2547 :   0 - 0x0
      12'h9F4: dout <= 8'b00000000; // 2548 :   0 - 0x0
      12'h9F5: dout <= 8'b00000000; // 2549 :   0 - 0x0
      12'h9F6: dout <= 8'b00000000; // 2550 :   0 - 0x0
      12'h9F7: dout <= 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- plane 1
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout <= 8'b11111111; // 2560 : 255 - 0xff -- Sprite 0xa0
      12'hA01: dout <= 8'b11010101; // 2561 : 213 - 0xd5
      12'hA02: dout <= 8'b11111111; // 2562 : 255 - 0xff
      12'hA03: dout <= 8'b00000010; // 2563 :   2 - 0x2
      12'hA04: dout <= 8'b00000010; // 2564 :   2 - 0x2
      12'hA05: dout <= 8'b00000010; // 2565 :   2 - 0x2
      12'hA06: dout <= 8'b00000010; // 2566 :   2 - 0x2
      12'hA07: dout <= 8'b00000010; // 2567 :   2 - 0x2
      12'hA08: dout <= 8'b00000000; // 2568 :   0 - 0x0 -- plane 1
      12'hA09: dout <= 8'b01111111; // 2569 : 127 - 0x7f
      12'hA0A: dout <= 8'b00000000; // 2570 :   0 - 0x0
      12'hA0B: dout <= 8'b00000001; // 2571 :   1 - 0x1
      12'hA0C: dout <= 8'b00000001; // 2572 :   1 - 0x1
      12'hA0D: dout <= 8'b00000001; // 2573 :   1 - 0x1
      12'hA0E: dout <= 8'b00000001; // 2574 :   1 - 0x1
      12'hA0F: dout <= 8'b00000001; // 2575 :   1 - 0x1
      12'hA10: dout <= 8'b00000010; // 2576 :   2 - 0x2 -- Sprite 0xa1
      12'hA11: dout <= 8'b00000010; // 2577 :   2 - 0x2
      12'hA12: dout <= 8'b00000010; // 2578 :   2 - 0x2
      12'hA13: dout <= 8'b00000010; // 2579 :   2 - 0x2
      12'hA14: dout <= 8'b00000010; // 2580 :   2 - 0x2
      12'hA15: dout <= 8'b00000010; // 2581 :   2 - 0x2
      12'hA16: dout <= 8'b00000010; // 2582 :   2 - 0x2
      12'hA17: dout <= 8'b00000010; // 2583 :   2 - 0x2
      12'hA18: dout <= 8'b00000001; // 2584 :   1 - 0x1 -- plane 1
      12'hA19: dout <= 8'b00000001; // 2585 :   1 - 0x1
      12'hA1A: dout <= 8'b00000001; // 2586 :   1 - 0x1
      12'hA1B: dout <= 8'b00000001; // 2587 :   1 - 0x1
      12'hA1C: dout <= 8'b00000001; // 2588 :   1 - 0x1
      12'hA1D: dout <= 8'b00000001; // 2589 :   1 - 0x1
      12'hA1E: dout <= 8'b00000001; // 2590 :   1 - 0x1
      12'hA1F: dout <= 8'b00000001; // 2591 :   1 - 0x1
      12'hA20: dout <= 8'b11111111; // 2592 : 255 - 0xff -- Sprite 0xa2
      12'hA21: dout <= 8'b01010101; // 2593 :  85 - 0x55
      12'hA22: dout <= 8'b11111111; // 2594 : 255 - 0xff
      12'hA23: dout <= 8'b01000000; // 2595 :  64 - 0x40
      12'hA24: dout <= 8'b01000000; // 2596 :  64 - 0x40
      12'hA25: dout <= 8'b01000000; // 2597 :  64 - 0x40
      12'hA26: dout <= 8'b01000000; // 2598 :  64 - 0x40
      12'hA27: dout <= 8'b01000000; // 2599 :  64 - 0x40
      12'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0 -- plane 1
      12'hA29: dout <= 8'b11111110; // 2601 : 254 - 0xfe
      12'hA2A: dout <= 8'b00000000; // 2602 :   0 - 0x0
      12'hA2B: dout <= 8'b10000000; // 2603 : 128 - 0x80
      12'hA2C: dout <= 8'b10000000; // 2604 : 128 - 0x80
      12'hA2D: dout <= 8'b10000000; // 2605 : 128 - 0x80
      12'hA2E: dout <= 8'b10000000; // 2606 : 128 - 0x80
      12'hA2F: dout <= 8'b10000000; // 2607 : 128 - 0x80
      12'hA30: dout <= 8'b01000000; // 2608 :  64 - 0x40 -- Sprite 0xa3
      12'hA31: dout <= 8'b01000000; // 2609 :  64 - 0x40
      12'hA32: dout <= 8'b01000000; // 2610 :  64 - 0x40
      12'hA33: dout <= 8'b01000000; // 2611 :  64 - 0x40
      12'hA34: dout <= 8'b01000000; // 2612 :  64 - 0x40
      12'hA35: dout <= 8'b01000000; // 2613 :  64 - 0x40
      12'hA36: dout <= 8'b01000000; // 2614 :  64 - 0x40
      12'hA37: dout <= 8'b01000000; // 2615 :  64 - 0x40
      12'hA38: dout <= 8'b10000000; // 2616 : 128 - 0x80 -- plane 1
      12'hA39: dout <= 8'b10000000; // 2617 : 128 - 0x80
      12'hA3A: dout <= 8'b10000000; // 2618 : 128 - 0x80
      12'hA3B: dout <= 8'b10000000; // 2619 : 128 - 0x80
      12'hA3C: dout <= 8'b10000000; // 2620 : 128 - 0x80
      12'hA3D: dout <= 8'b10000000; // 2621 : 128 - 0x80
      12'hA3E: dout <= 8'b10000000; // 2622 : 128 - 0x80
      12'hA3F: dout <= 8'b10000000; // 2623 : 128 - 0x80
      12'hA40: dout <= 8'b00110001; // 2624 :  49 - 0x31 -- Sprite 0xa4
      12'hA41: dout <= 8'b01001000; // 2625 :  72 - 0x48
      12'hA42: dout <= 8'b01000101; // 2626 :  69 - 0x45
      12'hA43: dout <= 8'b10000101; // 2627 : 133 - 0x85
      12'hA44: dout <= 8'b10000011; // 2628 : 131 - 0x83
      12'hA45: dout <= 8'b10000010; // 2629 : 130 - 0x82
      12'hA46: dout <= 8'b01100010; // 2630 :  98 - 0x62
      12'hA47: dout <= 8'b00010010; // 2631 :  18 - 0x12
      12'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0 -- plane 1
      12'hA49: dout <= 8'b00110000; // 2633 :  48 - 0x30
      12'hA4A: dout <= 8'b00111000; // 2634 :  56 - 0x38
      12'hA4B: dout <= 8'b01111000; // 2635 : 120 - 0x78
      12'hA4C: dout <= 8'b01111100; // 2636 : 124 - 0x7c
      12'hA4D: dout <= 8'b01111101; // 2637 : 125 - 0x7d
      12'hA4E: dout <= 8'b00011101; // 2638 :  29 - 0x1d
      12'hA4F: dout <= 8'b00001101; // 2639 :  13 - 0xd
      12'hA50: dout <= 8'b00110010; // 2640 :  50 - 0x32 -- Sprite 0xa5
      12'hA51: dout <= 8'b00100010; // 2641 :  34 - 0x22
      12'hA52: dout <= 8'b01000010; // 2642 :  66 - 0x42
      12'hA53: dout <= 8'b01000000; // 2643 :  64 - 0x40
      12'hA54: dout <= 8'b01000000; // 2644 :  64 - 0x40
      12'hA55: dout <= 8'b00100000; // 2645 :  32 - 0x20
      12'hA56: dout <= 8'b00011110; // 2646 :  30 - 0x1e
      12'hA57: dout <= 8'b00000111; // 2647 :   7 - 0x7
      12'hA58: dout <= 8'b00001101; // 2648 :  13 - 0xd -- plane 1
      12'hA59: dout <= 8'b00011101; // 2649 :  29 - 0x1d
      12'hA5A: dout <= 8'b00111101; // 2650 :  61 - 0x3d
      12'hA5B: dout <= 8'b00111111; // 2651 :  63 - 0x3f
      12'hA5C: dout <= 8'b00111111; // 2652 :  63 - 0x3f
      12'hA5D: dout <= 8'b00011111; // 2653 :  31 - 0x1f
      12'hA5E: dout <= 8'b00000001; // 2654 :   1 - 0x1
      12'hA5F: dout <= 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout <= 8'b10000000; // 2656 : 128 - 0x80 -- Sprite 0xa6
      12'hA61: dout <= 8'b11100000; // 2657 : 224 - 0xe0
      12'hA62: dout <= 8'b00111000; // 2658 :  56 - 0x38
      12'hA63: dout <= 8'b00100100; // 2659 :  36 - 0x24
      12'hA64: dout <= 8'b00000100; // 2660 :   4 - 0x4
      12'hA65: dout <= 8'b00001000; // 2661 :   8 - 0x8
      12'hA66: dout <= 8'b00110000; // 2662 :  48 - 0x30
      12'hA67: dout <= 8'b00100000; // 2663 :  32 - 0x20
      12'hA68: dout <= 8'b00000000; // 2664 :   0 - 0x0 -- plane 1
      12'hA69: dout <= 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout <= 8'b11100000; // 2666 : 224 - 0xe0
      12'hA6B: dout <= 8'b11111000; // 2667 : 248 - 0xf8
      12'hA6C: dout <= 8'b11111000; // 2668 : 248 - 0xf8
      12'hA6D: dout <= 8'b11110000; // 2669 : 240 - 0xf0
      12'hA6E: dout <= 8'b11000000; // 2670 : 192 - 0xc0
      12'hA6F: dout <= 8'b11000000; // 2671 : 192 - 0xc0
      12'hA70: dout <= 8'b00110000; // 2672 :  48 - 0x30 -- Sprite 0xa7
      12'hA71: dout <= 8'b00001000; // 2673 :   8 - 0x8
      12'hA72: dout <= 8'b00001000; // 2674 :   8 - 0x8
      12'hA73: dout <= 8'b00110000; // 2675 :  48 - 0x30
      12'hA74: dout <= 8'b00100000; // 2676 :  32 - 0x20
      12'hA75: dout <= 8'b00100000; // 2677 :  32 - 0x20
      12'hA76: dout <= 8'b00110000; // 2678 :  48 - 0x30
      12'hA77: dout <= 8'b11110000; // 2679 : 240 - 0xf0
      12'hA78: dout <= 8'b11000000; // 2680 : 192 - 0xc0 -- plane 1
      12'hA79: dout <= 8'b11110000; // 2681 : 240 - 0xf0
      12'hA7A: dout <= 8'b11110000; // 2682 : 240 - 0xf0
      12'hA7B: dout <= 8'b11000000; // 2683 : 192 - 0xc0
      12'hA7C: dout <= 8'b11000000; // 2684 : 192 - 0xc0
      12'hA7D: dout <= 8'b11000000; // 2685 : 192 - 0xc0
      12'hA7E: dout <= 8'b11000000; // 2686 : 192 - 0xc0
      12'hA7F: dout <= 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout <= 8'b11111111; // 2688 : 255 - 0xff -- Sprite 0xa8
      12'hA81: dout <= 8'b11010010; // 2689 : 210 - 0xd2
      12'hA82: dout <= 8'b11110100; // 2690 : 244 - 0xf4
      12'hA83: dout <= 8'b11011000; // 2691 : 216 - 0xd8
      12'hA84: dout <= 8'b11111000; // 2692 : 248 - 0xf8
      12'hA85: dout <= 8'b11010100; // 2693 : 212 - 0xd4
      12'hA86: dout <= 8'b11110010; // 2694 : 242 - 0xf2
      12'hA87: dout <= 8'b11010001; // 2695 : 209 - 0xd1
      12'hA88: dout <= 8'b00000000; // 2696 :   0 - 0x0 -- plane 1
      12'hA89: dout <= 8'b01100000; // 2697 :  96 - 0x60
      12'hA8A: dout <= 8'b01100000; // 2698 :  96 - 0x60
      12'hA8B: dout <= 8'b01100000; // 2699 :  96 - 0x60
      12'hA8C: dout <= 8'b01100000; // 2700 :  96 - 0x60
      12'hA8D: dout <= 8'b01100000; // 2701 :  96 - 0x60
      12'hA8E: dout <= 8'b01100000; // 2702 :  96 - 0x60
      12'hA8F: dout <= 8'b01100000; // 2703 :  96 - 0x60
      12'hA90: dout <= 8'b11110001; // 2704 : 241 - 0xf1 -- Sprite 0xa9
      12'hA91: dout <= 8'b11010010; // 2705 : 210 - 0xd2
      12'hA92: dout <= 8'b11110100; // 2706 : 244 - 0xf4
      12'hA93: dout <= 8'b11011000; // 2707 : 216 - 0xd8
      12'hA94: dout <= 8'b11111000; // 2708 : 248 - 0xf8
      12'hA95: dout <= 8'b11010100; // 2709 : 212 - 0xd4
      12'hA96: dout <= 8'b11110010; // 2710 : 242 - 0xf2
      12'hA97: dout <= 8'b11111111; // 2711 : 255 - 0xff
      12'hA98: dout <= 8'b01100000; // 2712 :  96 - 0x60 -- plane 1
      12'hA99: dout <= 8'b01100000; // 2713 :  96 - 0x60
      12'hA9A: dout <= 8'b01100000; // 2714 :  96 - 0x60
      12'hA9B: dout <= 8'b01100000; // 2715 :  96 - 0x60
      12'hA9C: dout <= 8'b01100000; // 2716 :  96 - 0x60
      12'hA9D: dout <= 8'b01100000; // 2717 :  96 - 0x60
      12'hA9E: dout <= 8'b01100000; // 2718 :  96 - 0x60
      12'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout <= 8'b11111111; // 2720 : 255 - 0xff -- Sprite 0xaa
      12'hAA1: dout <= 8'b01000010; // 2721 :  66 - 0x42
      12'hAA2: dout <= 8'b00100100; // 2722 :  36 - 0x24
      12'hAA3: dout <= 8'b00011000; // 2723 :  24 - 0x18
      12'hAA4: dout <= 8'b00011000; // 2724 :  24 - 0x18
      12'hAA5: dout <= 8'b00100100; // 2725 :  36 - 0x24
      12'hAA6: dout <= 8'b01000010; // 2726 :  66 - 0x42
      12'hAA7: dout <= 8'b10000001; // 2727 : 129 - 0x81
      12'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0 -- plane 1
      12'hAA9: dout <= 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout <= 8'b00000000; // 2730 :   0 - 0x0
      12'hAAB: dout <= 8'b00000000; // 2731 :   0 - 0x0
      12'hAAC: dout <= 8'b00000000; // 2732 :   0 - 0x0
      12'hAAD: dout <= 8'b00000000; // 2733 :   0 - 0x0
      12'hAAE: dout <= 8'b00000000; // 2734 :   0 - 0x0
      12'hAAF: dout <= 8'b00000000; // 2735 :   0 - 0x0
      12'hAB0: dout <= 8'b10000001; // 2736 : 129 - 0x81 -- Sprite 0xab
      12'hAB1: dout <= 8'b01000010; // 2737 :  66 - 0x42
      12'hAB2: dout <= 8'b00100100; // 2738 :  36 - 0x24
      12'hAB3: dout <= 8'b00011000; // 2739 :  24 - 0x18
      12'hAB4: dout <= 8'b00011000; // 2740 :  24 - 0x18
      12'hAB5: dout <= 8'b00100100; // 2741 :  36 - 0x24
      12'hAB6: dout <= 8'b01000010; // 2742 :  66 - 0x42
      12'hAB7: dout <= 8'b11111111; // 2743 : 255 - 0xff
      12'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0 -- plane 1
      12'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout <= 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout <= 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout <= 8'b11111111; // 2752 : 255 - 0xff -- Sprite 0xac
      12'hAC1: dout <= 8'b01001101; // 2753 :  77 - 0x4d
      12'hAC2: dout <= 8'b00101111; // 2754 :  47 - 0x2f
      12'hAC3: dout <= 8'b00011101; // 2755 :  29 - 0x1d
      12'hAC4: dout <= 8'b00011111; // 2756 :  31 - 0x1f
      12'hAC5: dout <= 8'b00101101; // 2757 :  45 - 0x2d
      12'hAC6: dout <= 8'b01001111; // 2758 :  79 - 0x4f
      12'hAC7: dout <= 8'b10001101; // 2759 : 141 - 0x8d
      12'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0 -- plane 1
      12'hAC9: dout <= 8'b00000110; // 2761 :   6 - 0x6
      12'hACA: dout <= 8'b00000110; // 2762 :   6 - 0x6
      12'hACB: dout <= 8'b00000110; // 2763 :   6 - 0x6
      12'hACC: dout <= 8'b00000110; // 2764 :   6 - 0x6
      12'hACD: dout <= 8'b00000110; // 2765 :   6 - 0x6
      12'hACE: dout <= 8'b00000110; // 2766 :   6 - 0x6
      12'hACF: dout <= 8'b00000110; // 2767 :   6 - 0x6
      12'hAD0: dout <= 8'b10001111; // 2768 : 143 - 0x8f -- Sprite 0xad
      12'hAD1: dout <= 8'b01001101; // 2769 :  77 - 0x4d
      12'hAD2: dout <= 8'b00101111; // 2770 :  47 - 0x2f
      12'hAD3: dout <= 8'b00011101; // 2771 :  29 - 0x1d
      12'hAD4: dout <= 8'b00011111; // 2772 :  31 - 0x1f
      12'hAD5: dout <= 8'b00101101; // 2773 :  45 - 0x2d
      12'hAD6: dout <= 8'b01001111; // 2774 :  79 - 0x4f
      12'hAD7: dout <= 8'b11111111; // 2775 : 255 - 0xff
      12'hAD8: dout <= 8'b00000110; // 2776 :   6 - 0x6 -- plane 1
      12'hAD9: dout <= 8'b00000110; // 2777 :   6 - 0x6
      12'hADA: dout <= 8'b00000110; // 2778 :   6 - 0x6
      12'hADB: dout <= 8'b00000110; // 2779 :   6 - 0x6
      12'hADC: dout <= 8'b00000110; // 2780 :   6 - 0x6
      12'hADD: dout <= 8'b00000110; // 2781 :   6 - 0x6
      12'hADE: dout <= 8'b00000110; // 2782 :   6 - 0x6
      12'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout <= 8'b00000001; // 2784 :   1 - 0x1 -- Sprite 0xae
      12'hAE1: dout <= 8'b00000011; // 2785 :   3 - 0x3
      12'hAE2: dout <= 8'b00000110; // 2786 :   6 - 0x6
      12'hAE3: dout <= 8'b00000111; // 2787 :   7 - 0x7
      12'hAE4: dout <= 8'b00000111; // 2788 :   7 - 0x7
      12'hAE5: dout <= 8'b00000111; // 2789 :   7 - 0x7
      12'hAE6: dout <= 8'b00000110; // 2790 :   6 - 0x6
      12'hAE7: dout <= 8'b00000111; // 2791 :   7 - 0x7
      12'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0 -- plane 1
      12'hAE9: dout <= 8'b00000001; // 2793 :   1 - 0x1
      12'hAEA: dout <= 8'b00000011; // 2794 :   3 - 0x3
      12'hAEB: dout <= 8'b00000010; // 2795 :   2 - 0x2
      12'hAEC: dout <= 8'b00000010; // 2796 :   2 - 0x2
      12'hAED: dout <= 8'b00000000; // 2797 :   0 - 0x0
      12'hAEE: dout <= 8'b00000011; // 2798 :   3 - 0x3
      12'hAEF: dout <= 8'b00000010; // 2799 :   2 - 0x2
      12'hAF0: dout <= 8'b00000110; // 2800 :   6 - 0x6 -- Sprite 0xaf
      12'hAF1: dout <= 8'b00000110; // 2801 :   6 - 0x6
      12'hAF2: dout <= 8'b00001110; // 2802 :  14 - 0xe
      12'hAF3: dout <= 8'b00001111; // 2803 :  15 - 0xf
      12'hAF4: dout <= 8'b00001110; // 2804 :  14 - 0xe
      12'hAF5: dout <= 8'b00011010; // 2805 :  26 - 0x1a
      12'hAF6: dout <= 8'b00011011; // 2806 :  27 - 0x1b
      12'hAF7: dout <= 8'b00001111; // 2807 :  15 - 0xf
      12'hAF8: dout <= 8'b00000001; // 2808 :   1 - 0x1 -- plane 1
      12'hAF9: dout <= 8'b00000011; // 2809 :   3 - 0x3
      12'hAFA: dout <= 8'b00000101; // 2810 :   5 - 0x5
      12'hAFB: dout <= 8'b00000100; // 2811 :   4 - 0x4
      12'hAFC: dout <= 8'b00000101; // 2812 :   5 - 0x5
      12'hAFD: dout <= 8'b00001101; // 2813 :  13 - 0xd
      12'hAFE: dout <= 8'b00001100; // 2814 :  12 - 0xc
      12'hAFF: dout <= 8'b00000001; // 2815 :   1 - 0x1
      12'hB00: dout <= 8'b00000000; // 2816 :   0 - 0x0 -- Sprite 0xb0
      12'hB01: dout <= 8'b11000000; // 2817 : 192 - 0xc0
      12'hB02: dout <= 8'b11110000; // 2818 : 240 - 0xf0
      12'hB03: dout <= 8'b10001000; // 2819 : 136 - 0x88
      12'hB04: dout <= 8'b00010100; // 2820 :  20 - 0x14
      12'hB05: dout <= 8'b01101000; // 2821 : 104 - 0x68
      12'hB06: dout <= 8'b10101000; // 2822 : 168 - 0xa8
      12'hB07: dout <= 8'b00101100; // 2823 :  44 - 0x2c
      12'hB08: dout <= 8'b00000000; // 2824 :   0 - 0x0 -- plane 1
      12'hB09: dout <= 8'b00000000; // 2825 :   0 - 0x0
      12'hB0A: dout <= 8'b01000000; // 2826 :  64 - 0x40
      12'hB0B: dout <= 8'b11110000; // 2827 : 240 - 0xf0
      12'hB0C: dout <= 8'b11101000; // 2828 : 232 - 0xe8
      12'hB0D: dout <= 8'b10010000; // 2829 : 144 - 0x90
      12'hB0E: dout <= 8'b01010000; // 2830 :  80 - 0x50
      12'hB0F: dout <= 8'b11010000; // 2831 : 208 - 0xd0
      12'hB10: dout <= 8'b00000100; // 2832 :   4 - 0x4 -- Sprite 0xb1
      12'hB11: dout <= 8'b00111000; // 2833 :  56 - 0x38
      12'hB12: dout <= 8'b00010000; // 2834 :  16 - 0x10
      12'hB13: dout <= 8'b10100000; // 2835 : 160 - 0xa0
      12'hB14: dout <= 8'b01100000; // 2836 :  96 - 0x60
      12'hB15: dout <= 8'b00100000; // 2837 :  32 - 0x20
      12'hB16: dout <= 8'b00010000; // 2838 :  16 - 0x10
      12'hB17: dout <= 8'b10001000; // 2839 : 136 - 0x88
      12'hB18: dout <= 8'b11111000; // 2840 : 248 - 0xf8 -- plane 1
      12'hB19: dout <= 8'b11000000; // 2841 : 192 - 0xc0
      12'hB1A: dout <= 8'b11100000; // 2842 : 224 - 0xe0
      12'hB1B: dout <= 8'b01000000; // 2843 :  64 - 0x40
      12'hB1C: dout <= 8'b10000000; // 2844 : 128 - 0x80
      12'hB1D: dout <= 8'b11000000; // 2845 : 192 - 0xc0
      12'hB1E: dout <= 8'b11100000; // 2846 : 224 - 0xe0
      12'hB1F: dout <= 8'b01110000; // 2847 : 112 - 0x70
      12'hB20: dout <= 8'b00001111; // 2848 :  15 - 0xf -- Sprite 0xb2
      12'hB21: dout <= 8'b00011011; // 2849 :  27 - 0x1b
      12'hB22: dout <= 8'b00011011; // 2850 :  27 - 0x1b
      12'hB23: dout <= 8'b00001110; // 2851 :  14 - 0xe
      12'hB24: dout <= 8'b00000110; // 2852 :   6 - 0x6
      12'hB25: dout <= 8'b00001100; // 2853 :  12 - 0xc
      12'hB26: dout <= 8'b00001100; // 2854 :  12 - 0xc
      12'hB27: dout <= 8'b00111111; // 2855 :  63 - 0x3f
      12'hB28: dout <= 8'b00000001; // 2856 :   1 - 0x1 -- plane 1
      12'hB29: dout <= 8'b00001101; // 2857 :  13 - 0xd
      12'hB2A: dout <= 8'b00001101; // 2858 :  13 - 0xd
      12'hB2B: dout <= 8'b00000011; // 2859 :   3 - 0x3
      12'hB2C: dout <= 8'b00000011; // 2860 :   3 - 0x3
      12'hB2D: dout <= 8'b00000111; // 2861 :   7 - 0x7
      12'hB2E: dout <= 8'b00000111; // 2862 :   7 - 0x7
      12'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout <= 8'b01111111; // 2864 : 127 - 0x7f -- Sprite 0xb3
      12'hB31: dout <= 8'b01100000; // 2865 :  96 - 0x60
      12'hB32: dout <= 8'b01100000; // 2866 :  96 - 0x60
      12'hB33: dout <= 8'b01100000; // 2867 :  96 - 0x60
      12'hB34: dout <= 8'b01100000; // 2868 :  96 - 0x60
      12'hB35: dout <= 8'b01100000; // 2869 :  96 - 0x60
      12'hB36: dout <= 8'b01101010; // 2870 : 106 - 0x6a
      12'hB37: dout <= 8'b01111111; // 2871 : 127 - 0x7f
      12'hB38: dout <= 8'b00111111; // 2872 :  63 - 0x3f -- plane 1
      12'hB39: dout <= 8'b00111111; // 2873 :  63 - 0x3f
      12'hB3A: dout <= 8'b00111111; // 2874 :  63 - 0x3f
      12'hB3B: dout <= 8'b00111111; // 2875 :  63 - 0x3f
      12'hB3C: dout <= 8'b00111111; // 2876 :  63 - 0x3f
      12'hB3D: dout <= 8'b00111111; // 2877 :  63 - 0x3f
      12'hB3E: dout <= 8'b00110101; // 2878 :  53 - 0x35
      12'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout <= 8'b01001000; // 2880 :  72 - 0x48 -- Sprite 0xb4
      12'hB41: dout <= 8'b00110000; // 2881 :  48 - 0x30
      12'hB42: dout <= 8'b00010000; // 2882 :  16 - 0x10
      12'hB43: dout <= 8'b00010000; // 2883 :  16 - 0x10
      12'hB44: dout <= 8'b00001000; // 2884 :   8 - 0x8
      12'hB45: dout <= 8'b00001000; // 2885 :   8 - 0x8
      12'hB46: dout <= 8'b00001000; // 2886 :   8 - 0x8
      12'hB47: dout <= 8'b11111100; // 2887 : 252 - 0xfc
      12'hB48: dout <= 8'b10110000; // 2888 : 176 - 0xb0 -- plane 1
      12'hB49: dout <= 8'b11000000; // 2889 : 192 - 0xc0
      12'hB4A: dout <= 8'b11100000; // 2890 : 224 - 0xe0
      12'hB4B: dout <= 8'b11100000; // 2891 : 224 - 0xe0
      12'hB4C: dout <= 8'b11110000; // 2892 : 240 - 0xf0
      12'hB4D: dout <= 8'b11110000; // 2893 : 240 - 0xf0
      12'hB4E: dout <= 8'b11110000; // 2894 : 240 - 0xf0
      12'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout <= 8'b11111110; // 2896 : 254 - 0xfe -- Sprite 0xb5
      12'hB51: dout <= 8'b00000110; // 2897 :   6 - 0x6
      12'hB52: dout <= 8'b00000010; // 2898 :   2 - 0x2
      12'hB53: dout <= 8'b00000110; // 2899 :   6 - 0x6
      12'hB54: dout <= 8'b00000010; // 2900 :   2 - 0x2
      12'hB55: dout <= 8'b00000110; // 2901 :   6 - 0x6
      12'hB56: dout <= 8'b10101010; // 2902 : 170 - 0xaa
      12'hB57: dout <= 8'b11111110; // 2903 : 254 - 0xfe
      12'hB58: dout <= 8'b11111100; // 2904 : 252 - 0xfc -- plane 1
      12'hB59: dout <= 8'b11111000; // 2905 : 248 - 0xf8
      12'hB5A: dout <= 8'b11111100; // 2906 : 252 - 0xfc
      12'hB5B: dout <= 8'b11111000; // 2907 : 248 - 0xf8
      12'hB5C: dout <= 8'b11111100; // 2908 : 252 - 0xfc
      12'hB5D: dout <= 8'b11111000; // 2909 : 248 - 0xf8
      12'hB5E: dout <= 8'b01010100; // 2910 :  84 - 0x54
      12'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout <= 8'b11111111; // 2912 : 255 - 0xff -- Sprite 0xb6
      12'hB61: dout <= 8'b10000000; // 2913 : 128 - 0x80
      12'hB62: dout <= 8'b10000000; // 2914 : 128 - 0x80
      12'hB63: dout <= 8'b10000000; // 2915 : 128 - 0x80
      12'hB64: dout <= 8'b10000000; // 2916 : 128 - 0x80
      12'hB65: dout <= 8'b10000000; // 2917 : 128 - 0x80
      12'hB66: dout <= 8'b10010101; // 2918 : 149 - 0x95
      12'hB67: dout <= 8'b11111111; // 2919 : 255 - 0xff
      12'hB68: dout <= 8'b00000000; // 2920 :   0 - 0x0 -- plane 1
      12'hB69: dout <= 8'b01111111; // 2921 : 127 - 0x7f
      12'hB6A: dout <= 8'b01111111; // 2922 : 127 - 0x7f
      12'hB6B: dout <= 8'b01111111; // 2923 : 127 - 0x7f
      12'hB6C: dout <= 8'b01111111; // 2924 : 127 - 0x7f
      12'hB6D: dout <= 8'b01111111; // 2925 : 127 - 0x7f
      12'hB6E: dout <= 8'b01101010; // 2926 : 106 - 0x6a
      12'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout <= 8'b11111111; // 2928 : 255 - 0xff -- Sprite 0xb7
      12'hB71: dout <= 8'b10000100; // 2929 : 132 - 0x84
      12'hB72: dout <= 8'b10001100; // 2930 : 140 - 0x8c
      12'hB73: dout <= 8'b10000100; // 2931 : 132 - 0x84
      12'hB74: dout <= 8'b10001100; // 2932 : 140 - 0x8c
      12'hB75: dout <= 8'b10000100; // 2933 : 132 - 0x84
      12'hB76: dout <= 8'b10101100; // 2934 : 172 - 0xac
      12'hB77: dout <= 8'b11111111; // 2935 : 255 - 0xff
      12'hB78: dout <= 8'b00000000; // 2936 :   0 - 0x0 -- plane 1
      12'hB79: dout <= 8'b01111011; // 2937 : 123 - 0x7b
      12'hB7A: dout <= 8'b01110011; // 2938 : 115 - 0x73
      12'hB7B: dout <= 8'b01111011; // 2939 : 123 - 0x7b
      12'hB7C: dout <= 8'b01110011; // 2940 : 115 - 0x73
      12'hB7D: dout <= 8'b01111011; // 2941 : 123 - 0x7b
      12'hB7E: dout <= 8'b01010011; // 2942 :  83 - 0x53
      12'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout <= 8'b11111111; // 2944 : 255 - 0xff -- Sprite 0xb8
      12'hB81: dout <= 8'b00100001; // 2945 :  33 - 0x21
      12'hB82: dout <= 8'b01100001; // 2946 :  97 - 0x61
      12'hB83: dout <= 8'b00100011; // 2947 :  35 - 0x23
      12'hB84: dout <= 8'b01100001; // 2948 :  97 - 0x61
      12'hB85: dout <= 8'b00100011; // 2949 :  35 - 0x23
      12'hB86: dout <= 8'b01100101; // 2950 : 101 - 0x65
      12'hB87: dout <= 8'b11111111; // 2951 : 255 - 0xff
      12'hB88: dout <= 8'b00000000; // 2952 :   0 - 0x0 -- plane 1
      12'hB89: dout <= 8'b11011110; // 2953 : 222 - 0xde
      12'hB8A: dout <= 8'b10011110; // 2954 : 158 - 0x9e
      12'hB8B: dout <= 8'b11011100; // 2955 : 220 - 0xdc
      12'hB8C: dout <= 8'b10011110; // 2956 : 158 - 0x9e
      12'hB8D: dout <= 8'b11011100; // 2957 : 220 - 0xdc
      12'hB8E: dout <= 8'b10011010; // 2958 : 154 - 0x9a
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b11111111; // 2960 : 255 - 0xff -- Sprite 0xb9
      12'hB91: dout <= 8'b00000001; // 2961 :   1 - 0x1
      12'hB92: dout <= 8'b00000011; // 2962 :   3 - 0x3
      12'hB93: dout <= 8'b00000001; // 2963 :   1 - 0x1
      12'hB94: dout <= 8'b00000011; // 2964 :   3 - 0x3
      12'hB95: dout <= 8'b00000001; // 2965 :   1 - 0x1
      12'hB96: dout <= 8'b10101011; // 2966 : 171 - 0xab
      12'hB97: dout <= 8'b11111111; // 2967 : 255 - 0xff
      12'hB98: dout <= 8'b00000000; // 2968 :   0 - 0x0 -- plane 1
      12'hB99: dout <= 8'b11111110; // 2969 : 254 - 0xfe
      12'hB9A: dout <= 8'b11111100; // 2970 : 252 - 0xfc
      12'hB9B: dout <= 8'b11111110; // 2971 : 254 - 0xfe
      12'hB9C: dout <= 8'b11111100; // 2972 : 252 - 0xfc
      12'hB9D: dout <= 8'b11111110; // 2973 : 254 - 0xfe
      12'hB9E: dout <= 8'b01010100; // 2974 :  84 - 0x54
      12'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout <= 8'b11111111; // 2976 : 255 - 0xff -- Sprite 0xba
      12'hBA1: dout <= 8'b11010101; // 2977 : 213 - 0xd5
      12'hBA2: dout <= 8'b10101010; // 2978 : 170 - 0xaa
      12'hBA3: dout <= 8'b11111111; // 2979 : 255 - 0xff
      12'hBA4: dout <= 8'b10000000; // 2980 : 128 - 0x80
      12'hBA5: dout <= 8'b10000000; // 2981 : 128 - 0x80
      12'hBA6: dout <= 8'b10010101; // 2982 : 149 - 0x95
      12'hBA7: dout <= 8'b11111111; // 2983 : 255 - 0xff
      12'hBA8: dout <= 8'b00000000; // 2984 :   0 - 0x0 -- plane 1
      12'hBA9: dout <= 8'b01111111; // 2985 : 127 - 0x7f
      12'hBAA: dout <= 8'b01111111; // 2986 : 127 - 0x7f
      12'hBAB: dout <= 8'b00000000; // 2987 :   0 - 0x0
      12'hBAC: dout <= 8'b01111111; // 2988 : 127 - 0x7f
      12'hBAD: dout <= 8'b01111111; // 2989 : 127 - 0x7f
      12'hBAE: dout <= 8'b01101010; // 2990 : 106 - 0x6a
      12'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout <= 8'b00000000; // 2992 :   0 - 0x0 -- Sprite 0xbb
      12'hBB1: dout <= 8'b00000000; // 2993 :   0 - 0x0
      12'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      12'hBB3: dout <= 8'b00000000; // 2995 :   0 - 0x0
      12'hBB4: dout <= 8'b00000000; // 2996 :   0 - 0x0
      12'hBB5: dout <= 8'b00000000; // 2997 :   0 - 0x0
      12'hBB6: dout <= 8'b00000000; // 2998 :   0 - 0x0
      12'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0 -- plane 1
      12'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      12'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      12'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      12'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      12'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b11111111; // 3008 : 255 - 0xff -- Sprite 0xbc
      12'hBC1: dout <= 8'b01010101; // 3009 :  85 - 0x55
      12'hBC2: dout <= 8'b10101011; // 3010 : 171 - 0xab
      12'hBC3: dout <= 8'b11111111; // 3011 : 255 - 0xff
      12'hBC4: dout <= 8'b01100001; // 3012 :  97 - 0x61
      12'hBC5: dout <= 8'b00100011; // 3013 :  35 - 0x23
      12'hBC6: dout <= 8'b01100101; // 3014 : 101 - 0x65
      12'hBC7: dout <= 8'b11111111; // 3015 : 255 - 0xff
      12'hBC8: dout <= 8'b00000000; // 3016 :   0 - 0x0 -- plane 1
      12'hBC9: dout <= 8'b11111110; // 3017 : 254 - 0xfe
      12'hBCA: dout <= 8'b11111110; // 3018 : 254 - 0xfe
      12'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout <= 8'b10011110; // 3020 : 158 - 0x9e
      12'hBCD: dout <= 8'b11011100; // 3021 : 220 - 0xdc
      12'hBCE: dout <= 8'b10011010; // 3022 : 154 - 0x9a
      12'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout <= 8'b00000000; // 3024 :   0 - 0x0 -- Sprite 0xbd
      12'hBD1: dout <= 8'b00000000; // 3025 :   0 - 0x0
      12'hBD2: dout <= 8'b00000000; // 3026 :   0 - 0x0
      12'hBD3: dout <= 8'b00000000; // 3027 :   0 - 0x0
      12'hBD4: dout <= 8'b00000000; // 3028 :   0 - 0x0
      12'hBD5: dout <= 8'b00000000; // 3029 :   0 - 0x0
      12'hBD6: dout <= 8'b00000000; // 3030 :   0 - 0x0
      12'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0 -- plane 1
      12'hBD9: dout <= 8'b00000000; // 3033 :   0 - 0x0
      12'hBDA: dout <= 8'b00000000; // 3034 :   0 - 0x0
      12'hBDB: dout <= 8'b00000000; // 3035 :   0 - 0x0
      12'hBDC: dout <= 8'b00000000; // 3036 :   0 - 0x0
      12'hBDD: dout <= 8'b00000000; // 3037 :   0 - 0x0
      12'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout <= 8'b00000000; // 3040 :   0 - 0x0 -- Sprite 0xbe
      12'hBE1: dout <= 8'b00000000; // 3041 :   0 - 0x0
      12'hBE2: dout <= 8'b00000000; // 3042 :   0 - 0x0
      12'hBE3: dout <= 8'b00000000; // 3043 :   0 - 0x0
      12'hBE4: dout <= 8'b00000000; // 3044 :   0 - 0x0
      12'hBE5: dout <= 8'b00000000; // 3045 :   0 - 0x0
      12'hBE6: dout <= 8'b00000000; // 3046 :   0 - 0x0
      12'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      12'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0 -- plane 1
      12'hBE9: dout <= 8'b00000000; // 3049 :   0 - 0x0
      12'hBEA: dout <= 8'b00000000; // 3050 :   0 - 0x0
      12'hBEB: dout <= 8'b00000000; // 3051 :   0 - 0x0
      12'hBEC: dout <= 8'b00000000; // 3052 :   0 - 0x0
      12'hBED: dout <= 8'b00000000; // 3053 :   0 - 0x0
      12'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      12'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Sprite 0xbf
      12'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      12'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      12'hBF4: dout <= 8'b00000000; // 3060 :   0 - 0x0
      12'hBF5: dout <= 8'b00000000; // 3061 :   0 - 0x0
      12'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      12'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0 -- plane 1
      12'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      12'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      12'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      12'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout <= 8'b00000000; // 3072 :   0 - 0x0 -- Sprite 0xc0
      12'hC01: dout <= 8'b00000000; // 3073 :   0 - 0x0
      12'hC02: dout <= 8'b00000000; // 3074 :   0 - 0x0
      12'hC03: dout <= 8'b00000000; // 3075 :   0 - 0x0
      12'hC04: dout <= 8'b00000000; // 3076 :   0 - 0x0
      12'hC05: dout <= 8'b00000000; // 3077 :   0 - 0x0
      12'hC06: dout <= 8'b00000000; // 3078 :   0 - 0x0
      12'hC07: dout <= 8'b00000000; // 3079 :   0 - 0x0
      12'hC08: dout <= 8'b00000000; // 3080 :   0 - 0x0 -- plane 1
      12'hC09: dout <= 8'b00000000; // 3081 :   0 - 0x0
      12'hC0A: dout <= 8'b00000000; // 3082 :   0 - 0x0
      12'hC0B: dout <= 8'b00000000; // 3083 :   0 - 0x0
      12'hC0C: dout <= 8'b00000000; // 3084 :   0 - 0x0
      12'hC0D: dout <= 8'b00000000; // 3085 :   0 - 0x0
      12'hC0E: dout <= 8'b00000000; // 3086 :   0 - 0x0
      12'hC0F: dout <= 8'b00000000; // 3087 :   0 - 0x0
      12'hC10: dout <= 8'b00000000; // 3088 :   0 - 0x0 -- Sprite 0xc1
      12'hC11: dout <= 8'b00000000; // 3089 :   0 - 0x0
      12'hC12: dout <= 8'b00000000; // 3090 :   0 - 0x0
      12'hC13: dout <= 8'b00000000; // 3091 :   0 - 0x0
      12'hC14: dout <= 8'b00000000; // 3092 :   0 - 0x0
      12'hC15: dout <= 8'b00000000; // 3093 :   0 - 0x0
      12'hC16: dout <= 8'b00000000; // 3094 :   0 - 0x0
      12'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      12'hC18: dout <= 8'b00000000; // 3096 :   0 - 0x0 -- plane 1
      12'hC19: dout <= 8'b00000000; // 3097 :   0 - 0x0
      12'hC1A: dout <= 8'b00000000; // 3098 :   0 - 0x0
      12'hC1B: dout <= 8'b00000000; // 3099 :   0 - 0x0
      12'hC1C: dout <= 8'b00000000; // 3100 :   0 - 0x0
      12'hC1D: dout <= 8'b00000000; // 3101 :   0 - 0x0
      12'hC1E: dout <= 8'b00000000; // 3102 :   0 - 0x0
      12'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout <= 8'b00000000; // 3104 :   0 - 0x0 -- Sprite 0xc2
      12'hC21: dout <= 8'b00000000; // 3105 :   0 - 0x0
      12'hC22: dout <= 8'b00000000; // 3106 :   0 - 0x0
      12'hC23: dout <= 8'b00000000; // 3107 :   0 - 0x0
      12'hC24: dout <= 8'b00000000; // 3108 :   0 - 0x0
      12'hC25: dout <= 8'b00000000; // 3109 :   0 - 0x0
      12'hC26: dout <= 8'b00000000; // 3110 :   0 - 0x0
      12'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      12'hC28: dout <= 8'b00000000; // 3112 :   0 - 0x0 -- plane 1
      12'hC29: dout <= 8'b00000000; // 3113 :   0 - 0x0
      12'hC2A: dout <= 8'b00000000; // 3114 :   0 - 0x0
      12'hC2B: dout <= 8'b00000000; // 3115 :   0 - 0x0
      12'hC2C: dout <= 8'b00000000; // 3116 :   0 - 0x0
      12'hC2D: dout <= 8'b00000000; // 3117 :   0 - 0x0
      12'hC2E: dout <= 8'b00000000; // 3118 :   0 - 0x0
      12'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      12'hC30: dout <= 8'b00000000; // 3120 :   0 - 0x0 -- Sprite 0xc3
      12'hC31: dout <= 8'b00000000; // 3121 :   0 - 0x0
      12'hC32: dout <= 8'b00000000; // 3122 :   0 - 0x0
      12'hC33: dout <= 8'b00000000; // 3123 :   0 - 0x0
      12'hC34: dout <= 8'b00000000; // 3124 :   0 - 0x0
      12'hC35: dout <= 8'b00000000; // 3125 :   0 - 0x0
      12'hC36: dout <= 8'b00000000; // 3126 :   0 - 0x0
      12'hC37: dout <= 8'b00000000; // 3127 :   0 - 0x0
      12'hC38: dout <= 8'b00000000; // 3128 :   0 - 0x0 -- plane 1
      12'hC39: dout <= 8'b00000000; // 3129 :   0 - 0x0
      12'hC3A: dout <= 8'b00000000; // 3130 :   0 - 0x0
      12'hC3B: dout <= 8'b00000000; // 3131 :   0 - 0x0
      12'hC3C: dout <= 8'b00000000; // 3132 :   0 - 0x0
      12'hC3D: dout <= 8'b00000000; // 3133 :   0 - 0x0
      12'hC3E: dout <= 8'b00000000; // 3134 :   0 - 0x0
      12'hC3F: dout <= 8'b00000000; // 3135 :   0 - 0x0
      12'hC40: dout <= 8'b00000000; // 3136 :   0 - 0x0 -- Sprite 0xc4
      12'hC41: dout <= 8'b00000000; // 3137 :   0 - 0x0
      12'hC42: dout <= 8'b00000000; // 3138 :   0 - 0x0
      12'hC43: dout <= 8'b00000000; // 3139 :   0 - 0x0
      12'hC44: dout <= 8'b00000000; // 3140 :   0 - 0x0
      12'hC45: dout <= 8'b00000000; // 3141 :   0 - 0x0
      12'hC46: dout <= 8'b00000000; // 3142 :   0 - 0x0
      12'hC47: dout <= 8'b00000000; // 3143 :   0 - 0x0
      12'hC48: dout <= 8'b00000000; // 3144 :   0 - 0x0 -- plane 1
      12'hC49: dout <= 8'b00000000; // 3145 :   0 - 0x0
      12'hC4A: dout <= 8'b00000000; // 3146 :   0 - 0x0
      12'hC4B: dout <= 8'b00000000; // 3147 :   0 - 0x0
      12'hC4C: dout <= 8'b00000000; // 3148 :   0 - 0x0
      12'hC4D: dout <= 8'b00000000; // 3149 :   0 - 0x0
      12'hC4E: dout <= 8'b00000000; // 3150 :   0 - 0x0
      12'hC4F: dout <= 8'b00000000; // 3151 :   0 - 0x0
      12'hC50: dout <= 8'b00000000; // 3152 :   0 - 0x0 -- Sprite 0xc5
      12'hC51: dout <= 8'b00000000; // 3153 :   0 - 0x0
      12'hC52: dout <= 8'b00000001; // 3154 :   1 - 0x1
      12'hC53: dout <= 8'b00000110; // 3155 :   6 - 0x6
      12'hC54: dout <= 8'b00001010; // 3156 :  10 - 0xa
      12'hC55: dout <= 8'b00010100; // 3157 :  20 - 0x14
      12'hC56: dout <= 8'b00010000; // 3158 :  16 - 0x10
      12'hC57: dout <= 8'b00101000; // 3159 :  40 - 0x28
      12'hC58: dout <= 8'b00000000; // 3160 :   0 - 0x0 -- plane 1
      12'hC59: dout <= 8'b00000000; // 3161 :   0 - 0x0
      12'hC5A: dout <= 8'b00000000; // 3162 :   0 - 0x0
      12'hC5B: dout <= 8'b00000001; // 3163 :   1 - 0x1
      12'hC5C: dout <= 8'b00000111; // 3164 :   7 - 0x7
      12'hC5D: dout <= 8'b00001111; // 3165 :  15 - 0xf
      12'hC5E: dout <= 8'b00001111; // 3166 :  15 - 0xf
      12'hC5F: dout <= 8'b00011111; // 3167 :  31 - 0x1f
      12'hC60: dout <= 8'b00011111; // 3168 :  31 - 0x1f -- Sprite 0xc6
      12'hC61: dout <= 8'b01100000; // 3169 :  96 - 0x60
      12'hC62: dout <= 8'b10100000; // 3170 : 160 - 0xa0
      12'hC63: dout <= 8'b01000000; // 3171 :  64 - 0x40
      12'hC64: dout <= 8'b00000000; // 3172 :   0 - 0x0
      12'hC65: dout <= 8'b00000000; // 3173 :   0 - 0x0
      12'hC66: dout <= 8'b00000000; // 3174 :   0 - 0x0
      12'hC67: dout <= 8'b00000000; // 3175 :   0 - 0x0
      12'hC68: dout <= 8'b00000000; // 3176 :   0 - 0x0 -- plane 1
      12'hC69: dout <= 8'b00011111; // 3177 :  31 - 0x1f
      12'hC6A: dout <= 8'b01111111; // 3178 : 127 - 0x7f
      12'hC6B: dout <= 8'b11111111; // 3179 : 255 - 0xff
      12'hC6C: dout <= 8'b11111111; // 3180 : 255 - 0xff
      12'hC6D: dout <= 8'b11111111; // 3181 : 255 - 0xff
      12'hC6E: dout <= 8'b11111111; // 3182 : 255 - 0xff
      12'hC6F: dout <= 8'b11111111; // 3183 : 255 - 0xff
      12'hC70: dout <= 8'b00110000; // 3184 :  48 - 0x30 -- Sprite 0xc7
      12'hC71: dout <= 8'b01000000; // 3185 :  64 - 0x40
      12'hC72: dout <= 8'b01100000; // 3186 :  96 - 0x60
      12'hC73: dout <= 8'b11000000; // 3187 : 192 - 0xc0
      12'hC74: dout <= 8'b10000000; // 3188 : 128 - 0x80
      12'hC75: dout <= 8'b10100000; // 3189 : 160 - 0xa0
      12'hC76: dout <= 8'b11000000; // 3190 : 192 - 0xc0
      12'hC77: dout <= 8'b10000000; // 3191 : 128 - 0x80
      12'hC78: dout <= 8'b00011111; // 3192 :  31 - 0x1f -- plane 1
      12'hC79: dout <= 8'b00111111; // 3193 :  63 - 0x3f
      12'hC7A: dout <= 8'b00111111; // 3194 :  63 - 0x3f
      12'hC7B: dout <= 8'b01111111; // 3195 : 127 - 0x7f
      12'hC7C: dout <= 8'b01111111; // 3196 : 127 - 0x7f
      12'hC7D: dout <= 8'b01111111; // 3197 : 127 - 0x7f
      12'hC7E: dout <= 8'b01111111; // 3198 : 127 - 0x7f
      12'hC7F: dout <= 8'b01111111; // 3199 : 127 - 0x7f
      12'hC80: dout <= 8'b11111111; // 3200 : 255 - 0xff -- Sprite 0xc8
      12'hC81: dout <= 8'b00000000; // 3201 :   0 - 0x0
      12'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      12'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      12'hC84: dout <= 8'b00000000; // 3204 :   0 - 0x0
      12'hC85: dout <= 8'b00000000; // 3205 :   0 - 0x0
      12'hC86: dout <= 8'b00000000; // 3206 :   0 - 0x0
      12'hC87: dout <= 8'b00000000; // 3207 :   0 - 0x0
      12'hC88: dout <= 8'b00000000; // 3208 :   0 - 0x0 -- plane 1
      12'hC89: dout <= 8'b11111111; // 3209 : 255 - 0xff
      12'hC8A: dout <= 8'b11111111; // 3210 : 255 - 0xff
      12'hC8B: dout <= 8'b11111111; // 3211 : 255 - 0xff
      12'hC8C: dout <= 8'b11111111; // 3212 : 255 - 0xff
      12'hC8D: dout <= 8'b11111111; // 3213 : 255 - 0xff
      12'hC8E: dout <= 8'b11111111; // 3214 : 255 - 0xff
      12'hC8F: dout <= 8'b11111111; // 3215 : 255 - 0xff
      12'hC90: dout <= 8'b00010100; // 3216 :  20 - 0x14 -- Sprite 0xc9
      12'hC91: dout <= 8'b00101010; // 3217 :  42 - 0x2a
      12'hC92: dout <= 8'b00010110; // 3218 :  22 - 0x16
      12'hC93: dout <= 8'b00101011; // 3219 :  43 - 0x2b
      12'hC94: dout <= 8'b00010101; // 3220 :  21 - 0x15
      12'hC95: dout <= 8'b00101011; // 3221 :  43 - 0x2b
      12'hC96: dout <= 8'b00010101; // 3222 :  21 - 0x15
      12'hC97: dout <= 8'b00101011; // 3223 :  43 - 0x2b
      12'hC98: dout <= 8'b11101000; // 3224 : 232 - 0xe8 -- plane 1
      12'hC99: dout <= 8'b11010100; // 3225 : 212 - 0xd4
      12'hC9A: dout <= 8'b11101000; // 3226 : 232 - 0xe8
      12'hC9B: dout <= 8'b11010100; // 3227 : 212 - 0xd4
      12'hC9C: dout <= 8'b11101010; // 3228 : 234 - 0xea
      12'hC9D: dout <= 8'b11010100; // 3229 : 212 - 0xd4
      12'hC9E: dout <= 8'b11101010; // 3230 : 234 - 0xea
      12'hC9F: dout <= 8'b11010100; // 3231 : 212 - 0xd4
      12'hCA0: dout <= 8'b00000000; // 3232 :   0 - 0x0 -- Sprite 0xca
      12'hCA1: dout <= 8'b00000100; // 3233 :   4 - 0x4
      12'hCA2: dout <= 8'b00000100; // 3234 :   4 - 0x4
      12'hCA3: dout <= 8'b00000101; // 3235 :   5 - 0x5
      12'hCA4: dout <= 8'b00010101; // 3236 :  21 - 0x15
      12'hCA5: dout <= 8'b00010101; // 3237 :  21 - 0x15
      12'hCA6: dout <= 8'b01010101; // 3238 :  85 - 0x55
      12'hCA7: dout <= 8'b01010101; // 3239 :  85 - 0x55
      12'hCA8: dout <= 8'b00000000; // 3240 :   0 - 0x0 -- plane 1
      12'hCA9: dout <= 8'b00000000; // 3241 :   0 - 0x0
      12'hCAA: dout <= 8'b00000000; // 3242 :   0 - 0x0
      12'hCAB: dout <= 8'b00000000; // 3243 :   0 - 0x0
      12'hCAC: dout <= 8'b00000000; // 3244 :   0 - 0x0
      12'hCAD: dout <= 8'b00000000; // 3245 :   0 - 0x0
      12'hCAE: dout <= 8'b00000000; // 3246 :   0 - 0x0
      12'hCAF: dout <= 8'b00000000; // 3247 :   0 - 0x0
      12'hCB0: dout <= 8'b00000000; // 3248 :   0 - 0x0 -- Sprite 0xcb
      12'hCB1: dout <= 8'b00000000; // 3249 :   0 - 0x0
      12'hCB2: dout <= 8'b00010000; // 3250 :  16 - 0x10
      12'hCB3: dout <= 8'b00010000; // 3251 :  16 - 0x10
      12'hCB4: dout <= 8'b01010001; // 3252 :  81 - 0x51
      12'hCB5: dout <= 8'b01010101; // 3253 :  85 - 0x55
      12'hCB6: dout <= 8'b01010101; // 3254 :  85 - 0x55
      12'hCB7: dout <= 8'b01010101; // 3255 :  85 - 0x55
      12'hCB8: dout <= 8'b00000000; // 3256 :   0 - 0x0 -- plane 1
      12'hCB9: dout <= 8'b00000000; // 3257 :   0 - 0x0
      12'hCBA: dout <= 8'b00000000; // 3258 :   0 - 0x0
      12'hCBB: dout <= 8'b00000000; // 3259 :   0 - 0x0
      12'hCBC: dout <= 8'b00000000; // 3260 :   0 - 0x0
      12'hCBD: dout <= 8'b00000000; // 3261 :   0 - 0x0
      12'hCBE: dout <= 8'b00000000; // 3262 :   0 - 0x0
      12'hCBF: dout <= 8'b00000000; // 3263 :   0 - 0x0
      12'hCC0: dout <= 8'b00000000; // 3264 :   0 - 0x0 -- Sprite 0xcc
      12'hCC1: dout <= 8'b00000000; // 3265 :   0 - 0x0
      12'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      12'hCC3: dout <= 8'b00000101; // 3267 :   5 - 0x5
      12'hCC4: dout <= 8'b00001111; // 3268 :  15 - 0xf
      12'hCC5: dout <= 8'b00000111; // 3269 :   7 - 0x7
      12'hCC6: dout <= 8'b00000011; // 3270 :   3 - 0x3
      12'hCC7: dout <= 8'b00000001; // 3271 :   1 - 0x1
      12'hCC8: dout <= 8'b00000000; // 3272 :   0 - 0x0 -- plane 1
      12'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      12'hCCA: dout <= 8'b00000000; // 3274 :   0 - 0x0
      12'hCCB: dout <= 8'b00000000; // 3275 :   0 - 0x0
      12'hCCC: dout <= 8'b00000101; // 3276 :   5 - 0x5
      12'hCCD: dout <= 8'b00000010; // 3277 :   2 - 0x2
      12'hCCE: dout <= 8'b00000001; // 3278 :   1 - 0x1
      12'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout <= 8'b00000000; // 3280 :   0 - 0x0 -- Sprite 0xcd
      12'hCD1: dout <= 8'b00000000; // 3281 :   0 - 0x0
      12'hCD2: dout <= 8'b10000000; // 3282 : 128 - 0x80
      12'hCD3: dout <= 8'b11010000; // 3283 : 208 - 0xd0
      12'hCD4: dout <= 8'b11111000; // 3284 : 248 - 0xf8
      12'hCD5: dout <= 8'b11110000; // 3285 : 240 - 0xf0
      12'hCD6: dout <= 8'b11100000; // 3286 : 224 - 0xe0
      12'hCD7: dout <= 8'b11000000; // 3287 : 192 - 0xc0
      12'hCD8: dout <= 8'b00000000; // 3288 :   0 - 0x0 -- plane 1
      12'hCD9: dout <= 8'b00000000; // 3289 :   0 - 0x0
      12'hCDA: dout <= 8'b00000000; // 3290 :   0 - 0x0
      12'hCDB: dout <= 8'b10000000; // 3291 : 128 - 0x80
      12'hCDC: dout <= 8'b01010000; // 3292 :  80 - 0x50
      12'hCDD: dout <= 8'b10100000; // 3293 : 160 - 0xa0
      12'hCDE: dout <= 8'b01000000; // 3294 :  64 - 0x40
      12'hCDF: dout <= 8'b10000000; // 3295 : 128 - 0x80
      12'hCE0: dout <= 8'b00000000; // 3296 :   0 - 0x0 -- Sprite 0xce
      12'hCE1: dout <= 8'b00000000; // 3297 :   0 - 0x0
      12'hCE2: dout <= 8'b00000000; // 3298 :   0 - 0x0
      12'hCE3: dout <= 8'b01111000; // 3299 : 120 - 0x78
      12'hCE4: dout <= 8'b11001111; // 3300 : 207 - 0xcf
      12'hCE5: dout <= 8'b10000000; // 3301 : 128 - 0x80
      12'hCE6: dout <= 8'b11001111; // 3302 : 207 - 0xcf
      12'hCE7: dout <= 8'b01001000; // 3303 :  72 - 0x48
      12'hCE8: dout <= 8'b00000000; // 3304 :   0 - 0x0 -- plane 1
      12'hCE9: dout <= 8'b00000000; // 3305 :   0 - 0x0
      12'hCEA: dout <= 8'b00000000; // 3306 :   0 - 0x0
      12'hCEB: dout <= 8'b00000000; // 3307 :   0 - 0x0
      12'hCEC: dout <= 8'b00110000; // 3308 :  48 - 0x30
      12'hCED: dout <= 8'b01111111; // 3309 : 127 - 0x7f
      12'hCEE: dout <= 8'b00110000; // 3310 :  48 - 0x30
      12'hCEF: dout <= 8'b00110000; // 3311 :  48 - 0x30
      12'hCF0: dout <= 8'b00000000; // 3312 :   0 - 0x0 -- Sprite 0xcf
      12'hCF1: dout <= 8'b00000000; // 3313 :   0 - 0x0
      12'hCF2: dout <= 8'b00000000; // 3314 :   0 - 0x0
      12'hCF3: dout <= 8'b00011110; // 3315 :  30 - 0x1e
      12'hCF4: dout <= 8'b11110011; // 3316 : 243 - 0xf3
      12'hCF5: dout <= 8'b00000001; // 3317 :   1 - 0x1
      12'hCF6: dout <= 8'b11110011; // 3318 : 243 - 0xf3
      12'hCF7: dout <= 8'b00010010; // 3319 :  18 - 0x12
      12'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0 -- plane 1
      12'hCF9: dout <= 8'b00000000; // 3321 :   0 - 0x0
      12'hCFA: dout <= 8'b00000000; // 3322 :   0 - 0x0
      12'hCFB: dout <= 8'b00000000; // 3323 :   0 - 0x0
      12'hCFC: dout <= 8'b00001100; // 3324 :  12 - 0xc
      12'hCFD: dout <= 8'b11111110; // 3325 : 254 - 0xfe
      12'hCFE: dout <= 8'b00001100; // 3326 :  12 - 0xc
      12'hCFF: dout <= 8'b00001100; // 3327 :  12 - 0xc
      12'hD00: dout <= 8'b00000000; // 3328 :   0 - 0x0 -- Sprite 0xd0
      12'hD01: dout <= 8'b00000000; // 3329 :   0 - 0x0
      12'hD02: dout <= 8'b00000000; // 3330 :   0 - 0x0
      12'hD03: dout <= 8'b00000000; // 3331 :   0 - 0x0
      12'hD04: dout <= 8'b00000000; // 3332 :   0 - 0x0
      12'hD05: dout <= 8'b00000000; // 3333 :   0 - 0x0
      12'hD06: dout <= 8'b00000000; // 3334 :   0 - 0x0
      12'hD07: dout <= 8'b00000000; // 3335 :   0 - 0x0
      12'hD08: dout <= 8'b00000000; // 3336 :   0 - 0x0 -- plane 1
      12'hD09: dout <= 8'b00000000; // 3337 :   0 - 0x0
      12'hD0A: dout <= 8'b00000000; // 3338 :   0 - 0x0
      12'hD0B: dout <= 8'b00000000; // 3339 :   0 - 0x0
      12'hD0C: dout <= 8'b00000000; // 3340 :   0 - 0x0
      12'hD0D: dout <= 8'b00000000; // 3341 :   0 - 0x0
      12'hD0E: dout <= 8'b00000000; // 3342 :   0 - 0x0
      12'hD0F: dout <= 8'b00000000; // 3343 :   0 - 0x0
      12'hD10: dout <= 8'b00000000; // 3344 :   0 - 0x0 -- Sprite 0xd1
      12'hD11: dout <= 8'b00000000; // 3345 :   0 - 0x0
      12'hD12: dout <= 8'b00000000; // 3346 :   0 - 0x0
      12'hD13: dout <= 8'b00000000; // 3347 :   0 - 0x0
      12'hD14: dout <= 8'b00000000; // 3348 :   0 - 0x0
      12'hD15: dout <= 8'b00000000; // 3349 :   0 - 0x0
      12'hD16: dout <= 8'b00000000; // 3350 :   0 - 0x0
      12'hD17: dout <= 8'b00000000; // 3351 :   0 - 0x0
      12'hD18: dout <= 8'b00000000; // 3352 :   0 - 0x0 -- plane 1
      12'hD19: dout <= 8'b00000000; // 3353 :   0 - 0x0
      12'hD1A: dout <= 8'b00000000; // 3354 :   0 - 0x0
      12'hD1B: dout <= 8'b00000000; // 3355 :   0 - 0x0
      12'hD1C: dout <= 8'b00000000; // 3356 :   0 - 0x0
      12'hD1D: dout <= 8'b00000000; // 3357 :   0 - 0x0
      12'hD1E: dout <= 8'b00000000; // 3358 :   0 - 0x0
      12'hD1F: dout <= 8'b00000000; // 3359 :   0 - 0x0
      12'hD20: dout <= 8'b00001000; // 3360 :   8 - 0x8 -- Sprite 0xd2
      12'hD21: dout <= 8'b00001100; // 3361 :  12 - 0xc
      12'hD22: dout <= 8'b00001000; // 3362 :   8 - 0x8
      12'hD23: dout <= 8'b00001000; // 3363 :   8 - 0x8
      12'hD24: dout <= 8'b00001010; // 3364 :  10 - 0xa
      12'hD25: dout <= 8'b00001000; // 3365 :   8 - 0x8
      12'hD26: dout <= 8'b00001000; // 3366 :   8 - 0x8
      12'hD27: dout <= 8'b00001100; // 3367 :  12 - 0xc
      12'hD28: dout <= 8'b00000111; // 3368 :   7 - 0x7 -- plane 1
      12'hD29: dout <= 8'b00000111; // 3369 :   7 - 0x7
      12'hD2A: dout <= 8'b00000111; // 3370 :   7 - 0x7
      12'hD2B: dout <= 8'b00000111; // 3371 :   7 - 0x7
      12'hD2C: dout <= 8'b00000111; // 3372 :   7 - 0x7
      12'hD2D: dout <= 8'b00000111; // 3373 :   7 - 0x7
      12'hD2E: dout <= 8'b00000111; // 3374 :   7 - 0x7
      12'hD2F: dout <= 8'b00000111; // 3375 :   7 - 0x7
      12'hD30: dout <= 8'b00010000; // 3376 :  16 - 0x10 -- Sprite 0xd3
      12'hD31: dout <= 8'b00010000; // 3377 :  16 - 0x10
      12'hD32: dout <= 8'b00110000; // 3378 :  48 - 0x30
      12'hD33: dout <= 8'b00010000; // 3379 :  16 - 0x10
      12'hD34: dout <= 8'b01010000; // 3380 :  80 - 0x50
      12'hD35: dout <= 8'b00010000; // 3381 :  16 - 0x10
      12'hD36: dout <= 8'b00110000; // 3382 :  48 - 0x30
      12'hD37: dout <= 8'b00010000; // 3383 :  16 - 0x10
      12'hD38: dout <= 8'b11100000; // 3384 : 224 - 0xe0 -- plane 1
      12'hD39: dout <= 8'b11100000; // 3385 : 224 - 0xe0
      12'hD3A: dout <= 8'b11000000; // 3386 : 192 - 0xc0
      12'hD3B: dout <= 8'b11100000; // 3387 : 224 - 0xe0
      12'hD3C: dout <= 8'b10100000; // 3388 : 160 - 0xa0
      12'hD3D: dout <= 8'b11100000; // 3389 : 224 - 0xe0
      12'hD3E: dout <= 8'b11000000; // 3390 : 192 - 0xc0
      12'hD3F: dout <= 8'b11100000; // 3391 : 224 - 0xe0
      12'hD40: dout <= 8'b00000000; // 3392 :   0 - 0x0 -- Sprite 0xd4
      12'hD41: dout <= 8'b00000000; // 3393 :   0 - 0x0
      12'hD42: dout <= 8'b00000000; // 3394 :   0 - 0x0
      12'hD43: dout <= 8'b00000000; // 3395 :   0 - 0x0
      12'hD44: dout <= 8'b00000000; // 3396 :   0 - 0x0
      12'hD45: dout <= 8'b00000000; // 3397 :   0 - 0x0
      12'hD46: dout <= 8'b00000000; // 3398 :   0 - 0x0
      12'hD47: dout <= 8'b00000000; // 3399 :   0 - 0x0
      12'hD48: dout <= 8'b00000000; // 3400 :   0 - 0x0 -- plane 1
      12'hD49: dout <= 8'b00000000; // 3401 :   0 - 0x0
      12'hD4A: dout <= 8'b00000000; // 3402 :   0 - 0x0
      12'hD4B: dout <= 8'b00000000; // 3403 :   0 - 0x0
      12'hD4C: dout <= 8'b00000000; // 3404 :   0 - 0x0
      12'hD4D: dout <= 8'b00000000; // 3405 :   0 - 0x0
      12'hD4E: dout <= 8'b00000000; // 3406 :   0 - 0x0
      12'hD4F: dout <= 8'b00000000; // 3407 :   0 - 0x0
      12'hD50: dout <= 8'b11111000; // 3408 : 248 - 0xf8 -- Sprite 0xd5
      12'hD51: dout <= 8'b00000110; // 3409 :   6 - 0x6
      12'hD52: dout <= 8'b00000001; // 3410 :   1 - 0x1
      12'hD53: dout <= 8'b00000000; // 3411 :   0 - 0x0
      12'hD54: dout <= 8'b00000000; // 3412 :   0 - 0x0
      12'hD55: dout <= 8'b00000000; // 3413 :   0 - 0x0
      12'hD56: dout <= 8'b00000000; // 3414 :   0 - 0x0
      12'hD57: dout <= 8'b00000000; // 3415 :   0 - 0x0
      12'hD58: dout <= 8'b00000000; // 3416 :   0 - 0x0 -- plane 1
      12'hD59: dout <= 8'b11111000; // 3417 : 248 - 0xf8
      12'hD5A: dout <= 8'b11111110; // 3418 : 254 - 0xfe
      12'hD5B: dout <= 8'b11111111; // 3419 : 255 - 0xff
      12'hD5C: dout <= 8'b11111111; // 3420 : 255 - 0xff
      12'hD5D: dout <= 8'b11111111; // 3421 : 255 - 0xff
      12'hD5E: dout <= 8'b11111111; // 3422 : 255 - 0xff
      12'hD5F: dout <= 8'b11111111; // 3423 : 255 - 0xff
      12'hD60: dout <= 8'b00000000; // 3424 :   0 - 0x0 -- Sprite 0xd6
      12'hD61: dout <= 8'b00000000; // 3425 :   0 - 0x0
      12'hD62: dout <= 8'b10000000; // 3426 : 128 - 0x80
      12'hD63: dout <= 8'b01100000; // 3427 :  96 - 0x60
      12'hD64: dout <= 8'b01010000; // 3428 :  80 - 0x50
      12'hD65: dout <= 8'b10101000; // 3429 : 168 - 0xa8
      12'hD66: dout <= 8'b01011000; // 3430 :  88 - 0x58
      12'hD67: dout <= 8'b00101100; // 3431 :  44 - 0x2c
      12'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0 -- plane 1
      12'hD69: dout <= 8'b00000000; // 3433 :   0 - 0x0
      12'hD6A: dout <= 8'b00000000; // 3434 :   0 - 0x0
      12'hD6B: dout <= 8'b10000000; // 3435 : 128 - 0x80
      12'hD6C: dout <= 8'b10100000; // 3436 : 160 - 0xa0
      12'hD6D: dout <= 8'b01010000; // 3437 :  80 - 0x50
      12'hD6E: dout <= 8'b10100000; // 3438 : 160 - 0xa0
      12'hD6F: dout <= 8'b11010000; // 3439 : 208 - 0xd0
      12'hD70: dout <= 8'b10100000; // 3440 : 160 - 0xa0 -- Sprite 0xd7
      12'hD71: dout <= 8'b11000000; // 3441 : 192 - 0xc0
      12'hD72: dout <= 8'b10000000; // 3442 : 128 - 0x80
      12'hD73: dout <= 8'b01010000; // 3443 :  80 - 0x50
      12'hD74: dout <= 8'b01100000; // 3444 :  96 - 0x60
      12'hD75: dout <= 8'b00111000; // 3445 :  56 - 0x38
      12'hD76: dout <= 8'b00001000; // 3446 :   8 - 0x8
      12'hD77: dout <= 8'b00000111; // 3447 :   7 - 0x7
      12'hD78: dout <= 8'b01111111; // 3448 : 127 - 0x7f -- plane 1
      12'hD79: dout <= 8'b01111111; // 3449 : 127 - 0x7f
      12'hD7A: dout <= 8'b01111111; // 3450 : 127 - 0x7f
      12'hD7B: dout <= 8'b00111111; // 3451 :  63 - 0x3f
      12'hD7C: dout <= 8'b00111111; // 3452 :  63 - 0x3f
      12'hD7D: dout <= 8'b00001111; // 3453 :  15 - 0xf
      12'hD7E: dout <= 8'b00000111; // 3454 :   7 - 0x7
      12'hD7F: dout <= 8'b00000000; // 3455 :   0 - 0x0
      12'hD80: dout <= 8'b00000000; // 3456 :   0 - 0x0 -- Sprite 0xd8
      12'hD81: dout <= 8'b00000000; // 3457 :   0 - 0x0
      12'hD82: dout <= 8'b00000000; // 3458 :   0 - 0x0
      12'hD83: dout <= 8'b00000000; // 3459 :   0 - 0x0
      12'hD84: dout <= 8'b00000000; // 3460 :   0 - 0x0
      12'hD85: dout <= 8'b00000000; // 3461 :   0 - 0x0
      12'hD86: dout <= 8'b00000000; // 3462 :   0 - 0x0
      12'hD87: dout <= 8'b11111111; // 3463 : 255 - 0xff
      12'hD88: dout <= 8'b11111111; // 3464 : 255 - 0xff -- plane 1
      12'hD89: dout <= 8'b11111111; // 3465 : 255 - 0xff
      12'hD8A: dout <= 8'b11111111; // 3466 : 255 - 0xff
      12'hD8B: dout <= 8'b11111111; // 3467 : 255 - 0xff
      12'hD8C: dout <= 8'b11111111; // 3468 : 255 - 0xff
      12'hD8D: dout <= 8'b11111111; // 3469 : 255 - 0xff
      12'hD8E: dout <= 8'b11111111; // 3470 : 255 - 0xff
      12'hD8F: dout <= 8'b00000000; // 3471 :   0 - 0x0
      12'hD90: dout <= 8'b00010101; // 3472 :  21 - 0x15 -- Sprite 0xd9
      12'hD91: dout <= 8'b00101011; // 3473 :  43 - 0x2b
      12'hD92: dout <= 8'b00010101; // 3474 :  21 - 0x15
      12'hD93: dout <= 8'b00101010; // 3475 :  42 - 0x2a
      12'hD94: dout <= 8'b01010110; // 3476 :  86 - 0x56
      12'hD95: dout <= 8'b10101100; // 3477 : 172 - 0xac
      12'hD96: dout <= 8'b01010000; // 3478 :  80 - 0x50
      12'hD97: dout <= 8'b11100000; // 3479 : 224 - 0xe0
      12'hD98: dout <= 8'b11101010; // 3480 : 234 - 0xea -- plane 1
      12'hD99: dout <= 8'b11010100; // 3481 : 212 - 0xd4
      12'hD9A: dout <= 8'b11101010; // 3482 : 234 - 0xea
      12'hD9B: dout <= 8'b11010100; // 3483 : 212 - 0xd4
      12'hD9C: dout <= 8'b10101000; // 3484 : 168 - 0xa8
      12'hD9D: dout <= 8'b01010000; // 3485 :  80 - 0x50
      12'hD9E: dout <= 8'b10100000; // 3486 : 160 - 0xa0
      12'hD9F: dout <= 8'b00000000; // 3487 :   0 - 0x0
      12'hDA0: dout <= 8'b00000001; // 3488 :   1 - 0x1 -- Sprite 0xda
      12'hDA1: dout <= 8'b00001101; // 3489 :  13 - 0xd
      12'hDA2: dout <= 8'b00010011; // 3490 :  19 - 0x13
      12'hDA3: dout <= 8'b00001101; // 3491 :  13 - 0xd
      12'hDA4: dout <= 8'b00000001; // 3492 :   1 - 0x1
      12'hDA5: dout <= 8'b00000001; // 3493 :   1 - 0x1
      12'hDA6: dout <= 8'b00000001; // 3494 :   1 - 0x1
      12'hDA7: dout <= 8'b00000001; // 3495 :   1 - 0x1
      12'hDA8: dout <= 8'b00000000; // 3496 :   0 - 0x0 -- plane 1
      12'hDA9: dout <= 8'b00000000; // 3497 :   0 - 0x0
      12'hDAA: dout <= 8'b00001100; // 3498 :  12 - 0xc
      12'hDAB: dout <= 8'b00000000; // 3499 :   0 - 0x0
      12'hDAC: dout <= 8'b00000000; // 3500 :   0 - 0x0
      12'hDAD: dout <= 8'b00000000; // 3501 :   0 - 0x0
      12'hDAE: dout <= 8'b00000000; // 3502 :   0 - 0x0
      12'hDAF: dout <= 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout <= 8'b11000000; // 3504 : 192 - 0xc0 -- Sprite 0xdb
      12'hDB1: dout <= 8'b01000000; // 3505 :  64 - 0x40
      12'hDB2: dout <= 8'b01000000; // 3506 :  64 - 0x40
      12'hDB3: dout <= 8'b01011000; // 3507 :  88 - 0x58
      12'hDB4: dout <= 8'b01100100; // 3508 : 100 - 0x64
      12'hDB5: dout <= 8'b01011000; // 3509 :  88 - 0x58
      12'hDB6: dout <= 8'b01000000; // 3510 :  64 - 0x40
      12'hDB7: dout <= 8'b01000000; // 3511 :  64 - 0x40
      12'hDB8: dout <= 8'b00000000; // 3512 :   0 - 0x0 -- plane 1
      12'hDB9: dout <= 8'b10000000; // 3513 : 128 - 0x80
      12'hDBA: dout <= 8'b10000000; // 3514 : 128 - 0x80
      12'hDBB: dout <= 8'b10000000; // 3515 : 128 - 0x80
      12'hDBC: dout <= 8'b10011000; // 3516 : 152 - 0x98
      12'hDBD: dout <= 8'b10000000; // 3517 : 128 - 0x80
      12'hDBE: dout <= 8'b10000000; // 3518 : 128 - 0x80
      12'hDBF: dout <= 8'b10000000; // 3519 : 128 - 0x80
      12'hDC0: dout <= 8'b00000000; // 3520 :   0 - 0x0 -- Sprite 0xdc
      12'hDC1: dout <= 8'b00000000; // 3521 :   0 - 0x0
      12'hDC2: dout <= 8'b00000000; // 3522 :   0 - 0x0
      12'hDC3: dout <= 8'b00000110; // 3523 :   6 - 0x6
      12'hDC4: dout <= 8'b00000111; // 3524 :   7 - 0x7
      12'hDC5: dout <= 8'b00000111; // 3525 :   7 - 0x7
      12'hDC6: dout <= 8'b00000111; // 3526 :   7 - 0x7
      12'hDC7: dout <= 8'b00000011; // 3527 :   3 - 0x3
      12'hDC8: dout <= 8'b00000000; // 3528 :   0 - 0x0 -- plane 1
      12'hDC9: dout <= 8'b00000000; // 3529 :   0 - 0x0
      12'hDCA: dout <= 8'b00000000; // 3530 :   0 - 0x0
      12'hDCB: dout <= 8'b00000000; // 3531 :   0 - 0x0
      12'hDCC: dout <= 8'b00000010; // 3532 :   2 - 0x2
      12'hDCD: dout <= 8'b00000011; // 3533 :   3 - 0x3
      12'hDCE: dout <= 8'b00000011; // 3534 :   3 - 0x3
      12'hDCF: dout <= 8'b00000001; // 3535 :   1 - 0x1
      12'hDD0: dout <= 8'b00000000; // 3536 :   0 - 0x0 -- Sprite 0xdd
      12'hDD1: dout <= 8'b00000000; // 3537 :   0 - 0x0
      12'hDD2: dout <= 8'b00000000; // 3538 :   0 - 0x0
      12'hDD3: dout <= 8'b10110000; // 3539 : 176 - 0xb0
      12'hDD4: dout <= 8'b11110000; // 3540 : 240 - 0xf0
      12'hDD5: dout <= 8'b11110000; // 3541 : 240 - 0xf0
      12'hDD6: dout <= 8'b11110000; // 3542 : 240 - 0xf0
      12'hDD7: dout <= 8'b11100000; // 3543 : 224 - 0xe0
      12'hDD8: dout <= 8'b00000000; // 3544 :   0 - 0x0 -- plane 1
      12'hDD9: dout <= 8'b00000000; // 3545 :   0 - 0x0
      12'hDDA: dout <= 8'b00000000; // 3546 :   0 - 0x0
      12'hDDB: dout <= 8'b00000000; // 3547 :   0 - 0x0
      12'hDDC: dout <= 8'b10100000; // 3548 : 160 - 0xa0
      12'hDDD: dout <= 8'b11100000; // 3549 : 224 - 0xe0
      12'hDDE: dout <= 8'b11100000; // 3550 : 224 - 0xe0
      12'hDDF: dout <= 8'b11000000; // 3551 : 192 - 0xc0
      12'hDE0: dout <= 8'b11001111; // 3552 : 207 - 0xcf -- Sprite 0xde
      12'hDE1: dout <= 8'b10000000; // 3553 : 128 - 0x80
      12'hDE2: dout <= 8'b11001111; // 3554 : 207 - 0xcf
      12'hDE3: dout <= 8'b01001000; // 3555 :  72 - 0x48
      12'hDE4: dout <= 8'b01001000; // 3556 :  72 - 0x48
      12'hDE5: dout <= 8'b01001000; // 3557 :  72 - 0x48
      12'hDE6: dout <= 8'b01001000; // 3558 :  72 - 0x48
      12'hDE7: dout <= 8'b01001000; // 3559 :  72 - 0x48
      12'hDE8: dout <= 8'b00110000; // 3560 :  48 - 0x30 -- plane 1
      12'hDE9: dout <= 8'b01111111; // 3561 : 127 - 0x7f
      12'hDEA: dout <= 8'b00110000; // 3562 :  48 - 0x30
      12'hDEB: dout <= 8'b00110000; // 3563 :  48 - 0x30
      12'hDEC: dout <= 8'b00110000; // 3564 :  48 - 0x30
      12'hDED: dout <= 8'b00110000; // 3565 :  48 - 0x30
      12'hDEE: dout <= 8'b00110000; // 3566 :  48 - 0x30
      12'hDEF: dout <= 8'b00110000; // 3567 :  48 - 0x30
      12'hDF0: dout <= 8'b11110011; // 3568 : 243 - 0xf3 -- Sprite 0xdf
      12'hDF1: dout <= 8'b00000001; // 3569 :   1 - 0x1
      12'hDF2: dout <= 8'b11110011; // 3570 : 243 - 0xf3
      12'hDF3: dout <= 8'b00010010; // 3571 :  18 - 0x12
      12'hDF4: dout <= 8'b00010010; // 3572 :  18 - 0x12
      12'hDF5: dout <= 8'b00010010; // 3573 :  18 - 0x12
      12'hDF6: dout <= 8'b00010010; // 3574 :  18 - 0x12
      12'hDF7: dout <= 8'b00010010; // 3575 :  18 - 0x12
      12'hDF8: dout <= 8'b00001100; // 3576 :  12 - 0xc -- plane 1
      12'hDF9: dout <= 8'b11111110; // 3577 : 254 - 0xfe
      12'hDFA: dout <= 8'b00001100; // 3578 :  12 - 0xc
      12'hDFB: dout <= 8'b00001100; // 3579 :  12 - 0xc
      12'hDFC: dout <= 8'b00001100; // 3580 :  12 - 0xc
      12'hDFD: dout <= 8'b00001100; // 3581 :  12 - 0xc
      12'hDFE: dout <= 8'b00001100; // 3582 :  12 - 0xc
      12'hDFF: dout <= 8'b00001100; // 3583 :  12 - 0xc
      12'hE00: dout <= 8'b00000000; // 3584 :   0 - 0x0 -- Sprite 0xe0
      12'hE01: dout <= 8'b00000000; // 3585 :   0 - 0x0
      12'hE02: dout <= 8'b00000000; // 3586 :   0 - 0x0
      12'hE03: dout <= 8'b00000000; // 3587 :   0 - 0x0
      12'hE04: dout <= 8'b00000000; // 3588 :   0 - 0x0
      12'hE05: dout <= 8'b00000000; // 3589 :   0 - 0x0
      12'hE06: dout <= 8'b00000000; // 3590 :   0 - 0x0
      12'hE07: dout <= 8'b00000000; // 3591 :   0 - 0x0
      12'hE08: dout <= 8'b00000000; // 3592 :   0 - 0x0 -- plane 1
      12'hE09: dout <= 8'b00000000; // 3593 :   0 - 0x0
      12'hE0A: dout <= 8'b00000000; // 3594 :   0 - 0x0
      12'hE0B: dout <= 8'b00000000; // 3595 :   0 - 0x0
      12'hE0C: dout <= 8'b00000000; // 3596 :   0 - 0x0
      12'hE0D: dout <= 8'b00000000; // 3597 :   0 - 0x0
      12'hE0E: dout <= 8'b00000000; // 3598 :   0 - 0x0
      12'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout <= 8'b00000000; // 3600 :   0 - 0x0 -- Sprite 0xe1
      12'hE11: dout <= 8'b00000000; // 3601 :   0 - 0x0
      12'hE12: dout <= 8'b00000000; // 3602 :   0 - 0x0
      12'hE13: dout <= 8'b00000000; // 3603 :   0 - 0x0
      12'hE14: dout <= 8'b00000000; // 3604 :   0 - 0x0
      12'hE15: dout <= 8'b00000000; // 3605 :   0 - 0x0
      12'hE16: dout <= 8'b00000000; // 3606 :   0 - 0x0
      12'hE17: dout <= 8'b00000000; // 3607 :   0 - 0x0
      12'hE18: dout <= 8'b00000000; // 3608 :   0 - 0x0 -- plane 1
      12'hE19: dout <= 8'b00000000; // 3609 :   0 - 0x0
      12'hE1A: dout <= 8'b00000000; // 3610 :   0 - 0x0
      12'hE1B: dout <= 8'b00000000; // 3611 :   0 - 0x0
      12'hE1C: dout <= 8'b00000000; // 3612 :   0 - 0x0
      12'hE1D: dout <= 8'b00000000; // 3613 :   0 - 0x0
      12'hE1E: dout <= 8'b00000000; // 3614 :   0 - 0x0
      12'hE1F: dout <= 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout <= 8'b00000000; // 3616 :   0 - 0x0 -- Sprite 0xe2
      12'hE21: dout <= 8'b00000000; // 3617 :   0 - 0x0
      12'hE22: dout <= 8'b00000000; // 3618 :   0 - 0x0
      12'hE23: dout <= 8'b00000000; // 3619 :   0 - 0x0
      12'hE24: dout <= 8'b00000000; // 3620 :   0 - 0x0
      12'hE25: dout <= 8'b00000000; // 3621 :   0 - 0x0
      12'hE26: dout <= 8'b00000000; // 3622 :   0 - 0x0
      12'hE27: dout <= 8'b00000000; // 3623 :   0 - 0x0
      12'hE28: dout <= 8'b00000000; // 3624 :   0 - 0x0 -- plane 1
      12'hE29: dout <= 8'b00000000; // 3625 :   0 - 0x0
      12'hE2A: dout <= 8'b00000000; // 3626 :   0 - 0x0
      12'hE2B: dout <= 8'b00000000; // 3627 :   0 - 0x0
      12'hE2C: dout <= 8'b00000000; // 3628 :   0 - 0x0
      12'hE2D: dout <= 8'b00000000; // 3629 :   0 - 0x0
      12'hE2E: dout <= 8'b00000000; // 3630 :   0 - 0x0
      12'hE2F: dout <= 8'b00000000; // 3631 :   0 - 0x0
      12'hE30: dout <= 8'b00000000; // 3632 :   0 - 0x0 -- Sprite 0xe3
      12'hE31: dout <= 8'b00000000; // 3633 :   0 - 0x0
      12'hE32: dout <= 8'b00000000; // 3634 :   0 - 0x0
      12'hE33: dout <= 8'b00000000; // 3635 :   0 - 0x0
      12'hE34: dout <= 8'b00000000; // 3636 :   0 - 0x0
      12'hE35: dout <= 8'b00000000; // 3637 :   0 - 0x0
      12'hE36: dout <= 8'b00000000; // 3638 :   0 - 0x0
      12'hE37: dout <= 8'b00000000; // 3639 :   0 - 0x0
      12'hE38: dout <= 8'b00000000; // 3640 :   0 - 0x0 -- plane 1
      12'hE39: dout <= 8'b00000000; // 3641 :   0 - 0x0
      12'hE3A: dout <= 8'b00000000; // 3642 :   0 - 0x0
      12'hE3B: dout <= 8'b00000000; // 3643 :   0 - 0x0
      12'hE3C: dout <= 8'b00000000; // 3644 :   0 - 0x0
      12'hE3D: dout <= 8'b00000000; // 3645 :   0 - 0x0
      12'hE3E: dout <= 8'b00000000; // 3646 :   0 - 0x0
      12'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout <= 8'b00000000; // 3648 :   0 - 0x0 -- Sprite 0xe4
      12'hE41: dout <= 8'b00000000; // 3649 :   0 - 0x0
      12'hE42: dout <= 8'b00000000; // 3650 :   0 - 0x0
      12'hE43: dout <= 8'b00000000; // 3651 :   0 - 0x0
      12'hE44: dout <= 8'b00000000; // 3652 :   0 - 0x0
      12'hE45: dout <= 8'b00000000; // 3653 :   0 - 0x0
      12'hE46: dout <= 8'b00000000; // 3654 :   0 - 0x0
      12'hE47: dout <= 8'b00000000; // 3655 :   0 - 0x0
      12'hE48: dout <= 8'b00000000; // 3656 :   0 - 0x0 -- plane 1
      12'hE49: dout <= 8'b00000000; // 3657 :   0 - 0x0
      12'hE4A: dout <= 8'b00000000; // 3658 :   0 - 0x0
      12'hE4B: dout <= 8'b00000000; // 3659 :   0 - 0x0
      12'hE4C: dout <= 8'b00000000; // 3660 :   0 - 0x0
      12'hE4D: dout <= 8'b00000000; // 3661 :   0 - 0x0
      12'hE4E: dout <= 8'b00000000; // 3662 :   0 - 0x0
      12'hE4F: dout <= 8'b00000000; // 3663 :   0 - 0x0
      12'hE50: dout <= 8'b00000000; // 3664 :   0 - 0x0 -- Sprite 0xe5
      12'hE51: dout <= 8'b00000000; // 3665 :   0 - 0x0
      12'hE52: dout <= 8'b00000000; // 3666 :   0 - 0x0
      12'hE53: dout <= 8'b00000000; // 3667 :   0 - 0x0
      12'hE54: dout <= 8'b00000000; // 3668 :   0 - 0x0
      12'hE55: dout <= 8'b00000000; // 3669 :   0 - 0x0
      12'hE56: dout <= 8'b00000000; // 3670 :   0 - 0x0
      12'hE57: dout <= 8'b00000000; // 3671 :   0 - 0x0
      12'hE58: dout <= 8'b00000000; // 3672 :   0 - 0x0 -- plane 1
      12'hE59: dout <= 8'b00000000; // 3673 :   0 - 0x0
      12'hE5A: dout <= 8'b00000000; // 3674 :   0 - 0x0
      12'hE5B: dout <= 8'b00000000; // 3675 :   0 - 0x0
      12'hE5C: dout <= 8'b00000000; // 3676 :   0 - 0x0
      12'hE5D: dout <= 8'b00000000; // 3677 :   0 - 0x0
      12'hE5E: dout <= 8'b00000000; // 3678 :   0 - 0x0
      12'hE5F: dout <= 8'b00000000; // 3679 :   0 - 0x0
      12'hE60: dout <= 8'b00000000; // 3680 :   0 - 0x0 -- Sprite 0xe6
      12'hE61: dout <= 8'b00000000; // 3681 :   0 - 0x0
      12'hE62: dout <= 8'b00000000; // 3682 :   0 - 0x0
      12'hE63: dout <= 8'b00000000; // 3683 :   0 - 0x0
      12'hE64: dout <= 8'b00000000; // 3684 :   0 - 0x0
      12'hE65: dout <= 8'b00000000; // 3685 :   0 - 0x0
      12'hE66: dout <= 8'b00000000; // 3686 :   0 - 0x0
      12'hE67: dout <= 8'b00000000; // 3687 :   0 - 0x0
      12'hE68: dout <= 8'b00000000; // 3688 :   0 - 0x0 -- plane 1
      12'hE69: dout <= 8'b00000000; // 3689 :   0 - 0x0
      12'hE6A: dout <= 8'b00000000; // 3690 :   0 - 0x0
      12'hE6B: dout <= 8'b00000000; // 3691 :   0 - 0x0
      12'hE6C: dout <= 8'b00000000; // 3692 :   0 - 0x0
      12'hE6D: dout <= 8'b00000000; // 3693 :   0 - 0x0
      12'hE6E: dout <= 8'b00000000; // 3694 :   0 - 0x0
      12'hE6F: dout <= 8'b00000000; // 3695 :   0 - 0x0
      12'hE70: dout <= 8'b00000000; // 3696 :   0 - 0x0 -- Sprite 0xe7
      12'hE71: dout <= 8'b00000000; // 3697 :   0 - 0x0
      12'hE72: dout <= 8'b00000000; // 3698 :   0 - 0x0
      12'hE73: dout <= 8'b00000000; // 3699 :   0 - 0x0
      12'hE74: dout <= 8'b00000000; // 3700 :   0 - 0x0
      12'hE75: dout <= 8'b00000000; // 3701 :   0 - 0x0
      12'hE76: dout <= 8'b00000000; // 3702 :   0 - 0x0
      12'hE77: dout <= 8'b00000000; // 3703 :   0 - 0x0
      12'hE78: dout <= 8'b00000000; // 3704 :   0 - 0x0 -- plane 1
      12'hE79: dout <= 8'b00000000; // 3705 :   0 - 0x0
      12'hE7A: dout <= 8'b00000000; // 3706 :   0 - 0x0
      12'hE7B: dout <= 8'b00000000; // 3707 :   0 - 0x0
      12'hE7C: dout <= 8'b00000000; // 3708 :   0 - 0x0
      12'hE7D: dout <= 8'b00000000; // 3709 :   0 - 0x0
      12'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout <= 8'b00000000; // 3712 :   0 - 0x0 -- Sprite 0xe8
      12'hE81: dout <= 8'b00000000; // 3713 :   0 - 0x0
      12'hE82: dout <= 8'b00000000; // 3714 :   0 - 0x0
      12'hE83: dout <= 8'b00000000; // 3715 :   0 - 0x0
      12'hE84: dout <= 8'b00000000; // 3716 :   0 - 0x0
      12'hE85: dout <= 8'b00000000; // 3717 :   0 - 0x0
      12'hE86: dout <= 8'b00000000; // 3718 :   0 - 0x0
      12'hE87: dout <= 8'b00000000; // 3719 :   0 - 0x0
      12'hE88: dout <= 8'b00000000; // 3720 :   0 - 0x0 -- plane 1
      12'hE89: dout <= 8'b00000000; // 3721 :   0 - 0x0
      12'hE8A: dout <= 8'b00000000; // 3722 :   0 - 0x0
      12'hE8B: dout <= 8'b00000000; // 3723 :   0 - 0x0
      12'hE8C: dout <= 8'b00000000; // 3724 :   0 - 0x0
      12'hE8D: dout <= 8'b00000000; // 3725 :   0 - 0x0
      12'hE8E: dout <= 8'b00000000; // 3726 :   0 - 0x0
      12'hE8F: dout <= 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout <= 8'b00000000; // 3728 :   0 - 0x0 -- Sprite 0xe9
      12'hE91: dout <= 8'b00000000; // 3729 :   0 - 0x0
      12'hE92: dout <= 8'b00000000; // 3730 :   0 - 0x0
      12'hE93: dout <= 8'b00000000; // 3731 :   0 - 0x0
      12'hE94: dout <= 8'b00000000; // 3732 :   0 - 0x0
      12'hE95: dout <= 8'b00000000; // 3733 :   0 - 0x0
      12'hE96: dout <= 8'b00000000; // 3734 :   0 - 0x0
      12'hE97: dout <= 8'b00000000; // 3735 :   0 - 0x0
      12'hE98: dout <= 8'b00000000; // 3736 :   0 - 0x0 -- plane 1
      12'hE99: dout <= 8'b00000000; // 3737 :   0 - 0x0
      12'hE9A: dout <= 8'b00000000; // 3738 :   0 - 0x0
      12'hE9B: dout <= 8'b00000000; // 3739 :   0 - 0x0
      12'hE9C: dout <= 8'b00000000; // 3740 :   0 - 0x0
      12'hE9D: dout <= 8'b00000000; // 3741 :   0 - 0x0
      12'hE9E: dout <= 8'b00000000; // 3742 :   0 - 0x0
      12'hE9F: dout <= 8'b00000000; // 3743 :   0 - 0x0
      12'hEA0: dout <= 8'b00000000; // 3744 :   0 - 0x0 -- Sprite 0xea
      12'hEA1: dout <= 8'b00000000; // 3745 :   0 - 0x0
      12'hEA2: dout <= 8'b00000000; // 3746 :   0 - 0x0
      12'hEA3: dout <= 8'b00000000; // 3747 :   0 - 0x0
      12'hEA4: dout <= 8'b00000000; // 3748 :   0 - 0x0
      12'hEA5: dout <= 8'b00000000; // 3749 :   0 - 0x0
      12'hEA6: dout <= 8'b00000000; // 3750 :   0 - 0x0
      12'hEA7: dout <= 8'b00000000; // 3751 :   0 - 0x0
      12'hEA8: dout <= 8'b00000000; // 3752 :   0 - 0x0 -- plane 1
      12'hEA9: dout <= 8'b00000000; // 3753 :   0 - 0x0
      12'hEAA: dout <= 8'b00000000; // 3754 :   0 - 0x0
      12'hEAB: dout <= 8'b00000000; // 3755 :   0 - 0x0
      12'hEAC: dout <= 8'b00000000; // 3756 :   0 - 0x0
      12'hEAD: dout <= 8'b00000000; // 3757 :   0 - 0x0
      12'hEAE: dout <= 8'b00000000; // 3758 :   0 - 0x0
      12'hEAF: dout <= 8'b00000000; // 3759 :   0 - 0x0
      12'hEB0: dout <= 8'b00000000; // 3760 :   0 - 0x0 -- Sprite 0xeb
      12'hEB1: dout <= 8'b00000000; // 3761 :   0 - 0x0
      12'hEB2: dout <= 8'b00000000; // 3762 :   0 - 0x0
      12'hEB3: dout <= 8'b00000000; // 3763 :   0 - 0x0
      12'hEB4: dout <= 8'b00000000; // 3764 :   0 - 0x0
      12'hEB5: dout <= 8'b00000000; // 3765 :   0 - 0x0
      12'hEB6: dout <= 8'b00000000; // 3766 :   0 - 0x0
      12'hEB7: dout <= 8'b00000000; // 3767 :   0 - 0x0
      12'hEB8: dout <= 8'b00000000; // 3768 :   0 - 0x0 -- plane 1
      12'hEB9: dout <= 8'b00000000; // 3769 :   0 - 0x0
      12'hEBA: dout <= 8'b00000000; // 3770 :   0 - 0x0
      12'hEBB: dout <= 8'b00000000; // 3771 :   0 - 0x0
      12'hEBC: dout <= 8'b00000000; // 3772 :   0 - 0x0
      12'hEBD: dout <= 8'b00000000; // 3773 :   0 - 0x0
      12'hEBE: dout <= 8'b00000000; // 3774 :   0 - 0x0
      12'hEBF: dout <= 8'b00000000; // 3775 :   0 - 0x0
      12'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Sprite 0xec
      12'hEC1: dout <= 8'b00000000; // 3777 :   0 - 0x0
      12'hEC2: dout <= 8'b00000000; // 3778 :   0 - 0x0
      12'hEC3: dout <= 8'b00000000; // 3779 :   0 - 0x0
      12'hEC4: dout <= 8'b00000000; // 3780 :   0 - 0x0
      12'hEC5: dout <= 8'b00000000; // 3781 :   0 - 0x0
      12'hEC6: dout <= 8'b00000000; // 3782 :   0 - 0x0
      12'hEC7: dout <= 8'b00000000; // 3783 :   0 - 0x0
      12'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0 -- plane 1
      12'hEC9: dout <= 8'b00000000; // 3785 :   0 - 0x0
      12'hECA: dout <= 8'b00000000; // 3786 :   0 - 0x0
      12'hECB: dout <= 8'b00000000; // 3787 :   0 - 0x0
      12'hECC: dout <= 8'b00000000; // 3788 :   0 - 0x0
      12'hECD: dout <= 8'b00000000; // 3789 :   0 - 0x0
      12'hECE: dout <= 8'b00000000; // 3790 :   0 - 0x0
      12'hECF: dout <= 8'b00000000; // 3791 :   0 - 0x0
      12'hED0: dout <= 8'b00000000; // 3792 :   0 - 0x0 -- Sprite 0xed
      12'hED1: dout <= 8'b00000000; // 3793 :   0 - 0x0
      12'hED2: dout <= 8'b00000000; // 3794 :   0 - 0x0
      12'hED3: dout <= 8'b00000000; // 3795 :   0 - 0x0
      12'hED4: dout <= 8'b00000000; // 3796 :   0 - 0x0
      12'hED5: dout <= 8'b00000000; // 3797 :   0 - 0x0
      12'hED6: dout <= 8'b00000000; // 3798 :   0 - 0x0
      12'hED7: dout <= 8'b00000000; // 3799 :   0 - 0x0
      12'hED8: dout <= 8'b00000000; // 3800 :   0 - 0x0 -- plane 1
      12'hED9: dout <= 8'b00000000; // 3801 :   0 - 0x0
      12'hEDA: dout <= 8'b00000000; // 3802 :   0 - 0x0
      12'hEDB: dout <= 8'b00000000; // 3803 :   0 - 0x0
      12'hEDC: dout <= 8'b00000000; // 3804 :   0 - 0x0
      12'hEDD: dout <= 8'b00000000; // 3805 :   0 - 0x0
      12'hEDE: dout <= 8'b00000000; // 3806 :   0 - 0x0
      12'hEDF: dout <= 8'b00000000; // 3807 :   0 - 0x0
      12'hEE0: dout <= 8'b00000000; // 3808 :   0 - 0x0 -- Sprite 0xee
      12'hEE1: dout <= 8'b00000000; // 3809 :   0 - 0x0
      12'hEE2: dout <= 8'b00000000; // 3810 :   0 - 0x0
      12'hEE3: dout <= 8'b00000000; // 3811 :   0 - 0x0
      12'hEE4: dout <= 8'b00000000; // 3812 :   0 - 0x0
      12'hEE5: dout <= 8'b00000000; // 3813 :   0 - 0x0
      12'hEE6: dout <= 8'b00000000; // 3814 :   0 - 0x0
      12'hEE7: dout <= 8'b00000000; // 3815 :   0 - 0x0
      12'hEE8: dout <= 8'b00000000; // 3816 :   0 - 0x0 -- plane 1
      12'hEE9: dout <= 8'b00000000; // 3817 :   0 - 0x0
      12'hEEA: dout <= 8'b00000000; // 3818 :   0 - 0x0
      12'hEEB: dout <= 8'b00000000; // 3819 :   0 - 0x0
      12'hEEC: dout <= 8'b00000000; // 3820 :   0 - 0x0
      12'hEED: dout <= 8'b00000000; // 3821 :   0 - 0x0
      12'hEEE: dout <= 8'b00000000; // 3822 :   0 - 0x0
      12'hEEF: dout <= 8'b00000000; // 3823 :   0 - 0x0
      12'hEF0: dout <= 8'b00000000; // 3824 :   0 - 0x0 -- Sprite 0xef
      12'hEF1: dout <= 8'b00000000; // 3825 :   0 - 0x0
      12'hEF2: dout <= 8'b00000000; // 3826 :   0 - 0x0
      12'hEF3: dout <= 8'b00000000; // 3827 :   0 - 0x0
      12'hEF4: dout <= 8'b00000000; // 3828 :   0 - 0x0
      12'hEF5: dout <= 8'b00000000; // 3829 :   0 - 0x0
      12'hEF6: dout <= 8'b00000000; // 3830 :   0 - 0x0
      12'hEF7: dout <= 8'b00000000; // 3831 :   0 - 0x0
      12'hEF8: dout <= 8'b00000000; // 3832 :   0 - 0x0 -- plane 1
      12'hEF9: dout <= 8'b00000000; // 3833 :   0 - 0x0
      12'hEFA: dout <= 8'b00000000; // 3834 :   0 - 0x0
      12'hEFB: dout <= 8'b00000000; // 3835 :   0 - 0x0
      12'hEFC: dout <= 8'b00000000; // 3836 :   0 - 0x0
      12'hEFD: dout <= 8'b00000000; // 3837 :   0 - 0x0
      12'hEFE: dout <= 8'b00000000; // 3838 :   0 - 0x0
      12'hEFF: dout <= 8'b00000000; // 3839 :   0 - 0x0
      12'hF00: dout <= 8'b00000000; // 3840 :   0 - 0x0 -- Sprite 0xf0
      12'hF01: dout <= 8'b00000000; // 3841 :   0 - 0x0
      12'hF02: dout <= 8'b00000000; // 3842 :   0 - 0x0
      12'hF03: dout <= 8'b00000000; // 3843 :   0 - 0x0
      12'hF04: dout <= 8'b00000000; // 3844 :   0 - 0x0
      12'hF05: dout <= 8'b00000000; // 3845 :   0 - 0x0
      12'hF06: dout <= 8'b00000000; // 3846 :   0 - 0x0
      12'hF07: dout <= 8'b00000000; // 3847 :   0 - 0x0
      12'hF08: dout <= 8'b00000000; // 3848 :   0 - 0x0 -- plane 1
      12'hF09: dout <= 8'b00000000; // 3849 :   0 - 0x0
      12'hF0A: dout <= 8'b00000000; // 3850 :   0 - 0x0
      12'hF0B: dout <= 8'b00000000; // 3851 :   0 - 0x0
      12'hF0C: dout <= 8'b00000000; // 3852 :   0 - 0x0
      12'hF0D: dout <= 8'b00000000; // 3853 :   0 - 0x0
      12'hF0E: dout <= 8'b00000000; // 3854 :   0 - 0x0
      12'hF0F: dout <= 8'b00000000; // 3855 :   0 - 0x0
      12'hF10: dout <= 8'b00000000; // 3856 :   0 - 0x0 -- Sprite 0xf1
      12'hF11: dout <= 8'b00000000; // 3857 :   0 - 0x0
      12'hF12: dout <= 8'b00000000; // 3858 :   0 - 0x0
      12'hF13: dout <= 8'b00000000; // 3859 :   0 - 0x0
      12'hF14: dout <= 8'b00000000; // 3860 :   0 - 0x0
      12'hF15: dout <= 8'b00000000; // 3861 :   0 - 0x0
      12'hF16: dout <= 8'b00000000; // 3862 :   0 - 0x0
      12'hF17: dout <= 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout <= 8'b00000000; // 3864 :   0 - 0x0 -- plane 1
      12'hF19: dout <= 8'b00000000; // 3865 :   0 - 0x0
      12'hF1A: dout <= 8'b00000000; // 3866 :   0 - 0x0
      12'hF1B: dout <= 8'b00000000; // 3867 :   0 - 0x0
      12'hF1C: dout <= 8'b00000000; // 3868 :   0 - 0x0
      12'hF1D: dout <= 8'b00000000; // 3869 :   0 - 0x0
      12'hF1E: dout <= 8'b00000000; // 3870 :   0 - 0x0
      12'hF1F: dout <= 8'b00000000; // 3871 :   0 - 0x0
      12'hF20: dout <= 8'b00000000; // 3872 :   0 - 0x0 -- Sprite 0xf2
      12'hF21: dout <= 8'b00000000; // 3873 :   0 - 0x0
      12'hF22: dout <= 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout <= 8'b00000000; // 3875 :   0 - 0x0
      12'hF24: dout <= 8'b00000000; // 3876 :   0 - 0x0
      12'hF25: dout <= 8'b00000000; // 3877 :   0 - 0x0
      12'hF26: dout <= 8'b00000000; // 3878 :   0 - 0x0
      12'hF27: dout <= 8'b00000000; // 3879 :   0 - 0x0
      12'hF28: dout <= 8'b00000000; // 3880 :   0 - 0x0 -- plane 1
      12'hF29: dout <= 8'b00000000; // 3881 :   0 - 0x0
      12'hF2A: dout <= 8'b00000000; // 3882 :   0 - 0x0
      12'hF2B: dout <= 8'b00000000; // 3883 :   0 - 0x0
      12'hF2C: dout <= 8'b00000000; // 3884 :   0 - 0x0
      12'hF2D: dout <= 8'b00000000; // 3885 :   0 - 0x0
      12'hF2E: dout <= 8'b00000000; // 3886 :   0 - 0x0
      12'hF2F: dout <= 8'b00000000; // 3887 :   0 - 0x0
      12'hF30: dout <= 8'b00000000; // 3888 :   0 - 0x0 -- Sprite 0xf3
      12'hF31: dout <= 8'b00000000; // 3889 :   0 - 0x0
      12'hF32: dout <= 8'b00000000; // 3890 :   0 - 0x0
      12'hF33: dout <= 8'b00000000; // 3891 :   0 - 0x0
      12'hF34: dout <= 8'b00000000; // 3892 :   0 - 0x0
      12'hF35: dout <= 8'b00000000; // 3893 :   0 - 0x0
      12'hF36: dout <= 8'b00000000; // 3894 :   0 - 0x0
      12'hF37: dout <= 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout <= 8'b00000000; // 3896 :   0 - 0x0 -- plane 1
      12'hF39: dout <= 8'b00000000; // 3897 :   0 - 0x0
      12'hF3A: dout <= 8'b00000000; // 3898 :   0 - 0x0
      12'hF3B: dout <= 8'b00000000; // 3899 :   0 - 0x0
      12'hF3C: dout <= 8'b00000000; // 3900 :   0 - 0x0
      12'hF3D: dout <= 8'b00000000; // 3901 :   0 - 0x0
      12'hF3E: dout <= 8'b00000000; // 3902 :   0 - 0x0
      12'hF3F: dout <= 8'b00000000; // 3903 :   0 - 0x0
      12'hF40: dout <= 8'b00000000; // 3904 :   0 - 0x0 -- Sprite 0xf4
      12'hF41: dout <= 8'b00000000; // 3905 :   0 - 0x0
      12'hF42: dout <= 8'b00000000; // 3906 :   0 - 0x0
      12'hF43: dout <= 8'b00000000; // 3907 :   0 - 0x0
      12'hF44: dout <= 8'b00000000; // 3908 :   0 - 0x0
      12'hF45: dout <= 8'b00000000; // 3909 :   0 - 0x0
      12'hF46: dout <= 8'b00000000; // 3910 :   0 - 0x0
      12'hF47: dout <= 8'b00000000; // 3911 :   0 - 0x0
      12'hF48: dout <= 8'b00000000; // 3912 :   0 - 0x0 -- plane 1
      12'hF49: dout <= 8'b00000000; // 3913 :   0 - 0x0
      12'hF4A: dout <= 8'b00000000; // 3914 :   0 - 0x0
      12'hF4B: dout <= 8'b00000000; // 3915 :   0 - 0x0
      12'hF4C: dout <= 8'b00000000; // 3916 :   0 - 0x0
      12'hF4D: dout <= 8'b00000000; // 3917 :   0 - 0x0
      12'hF4E: dout <= 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout <= 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout <= 8'b00000000; // 3920 :   0 - 0x0 -- Sprite 0xf5
      12'hF51: dout <= 8'b00000000; // 3921 :   0 - 0x0
      12'hF52: dout <= 8'b00000000; // 3922 :   0 - 0x0
      12'hF53: dout <= 8'b00000000; // 3923 :   0 - 0x0
      12'hF54: dout <= 8'b00000000; // 3924 :   0 - 0x0
      12'hF55: dout <= 8'b00000000; // 3925 :   0 - 0x0
      12'hF56: dout <= 8'b00000000; // 3926 :   0 - 0x0
      12'hF57: dout <= 8'b00000000; // 3927 :   0 - 0x0
      12'hF58: dout <= 8'b00000000; // 3928 :   0 - 0x0 -- plane 1
      12'hF59: dout <= 8'b00000000; // 3929 :   0 - 0x0
      12'hF5A: dout <= 8'b00000000; // 3930 :   0 - 0x0
      12'hF5B: dout <= 8'b00000000; // 3931 :   0 - 0x0
      12'hF5C: dout <= 8'b00000000; // 3932 :   0 - 0x0
      12'hF5D: dout <= 8'b00000000; // 3933 :   0 - 0x0
      12'hF5E: dout <= 8'b00000000; // 3934 :   0 - 0x0
      12'hF5F: dout <= 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Sprite 0xf6
      12'hF61: dout <= 8'b00000000; // 3937 :   0 - 0x0
      12'hF62: dout <= 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout <= 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout <= 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout <= 8'b00000000; // 3941 :   0 - 0x0
      12'hF66: dout <= 8'b00000000; // 3942 :   0 - 0x0
      12'hF67: dout <= 8'b00000000; // 3943 :   0 - 0x0
      12'hF68: dout <= 8'b00000000; // 3944 :   0 - 0x0 -- plane 1
      12'hF69: dout <= 8'b00000000; // 3945 :   0 - 0x0
      12'hF6A: dout <= 8'b00000000; // 3946 :   0 - 0x0
      12'hF6B: dout <= 8'b00000000; // 3947 :   0 - 0x0
      12'hF6C: dout <= 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout <= 8'b00000000; // 3949 :   0 - 0x0
      12'hF6E: dout <= 8'b00000000; // 3950 :   0 - 0x0
      12'hF6F: dout <= 8'b00000000; // 3951 :   0 - 0x0
      12'hF70: dout <= 8'b00000000; // 3952 :   0 - 0x0 -- Sprite 0xf7
      12'hF71: dout <= 8'b00000000; // 3953 :   0 - 0x0
      12'hF72: dout <= 8'b00000000; // 3954 :   0 - 0x0
      12'hF73: dout <= 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout <= 8'b00000000; // 3956 :   0 - 0x0
      12'hF75: dout <= 8'b00000000; // 3957 :   0 - 0x0
      12'hF76: dout <= 8'b00000000; // 3958 :   0 - 0x0
      12'hF77: dout <= 8'b00000000; // 3959 :   0 - 0x0
      12'hF78: dout <= 8'b00000000; // 3960 :   0 - 0x0 -- plane 1
      12'hF79: dout <= 8'b00000000; // 3961 :   0 - 0x0
      12'hF7A: dout <= 8'b00000000; // 3962 :   0 - 0x0
      12'hF7B: dout <= 8'b00000000; // 3963 :   0 - 0x0
      12'hF7C: dout <= 8'b00000000; // 3964 :   0 - 0x0
      12'hF7D: dout <= 8'b00000000; // 3965 :   0 - 0x0
      12'hF7E: dout <= 8'b00000000; // 3966 :   0 - 0x0
      12'hF7F: dout <= 8'b00000000; // 3967 :   0 - 0x0
      12'hF80: dout <= 8'b00000000; // 3968 :   0 - 0x0 -- Sprite 0xf8
      12'hF81: dout <= 8'b00000000; // 3969 :   0 - 0x0
      12'hF82: dout <= 8'b00000000; // 3970 :   0 - 0x0
      12'hF83: dout <= 8'b00000000; // 3971 :   0 - 0x0
      12'hF84: dout <= 8'b00000000; // 3972 :   0 - 0x0
      12'hF85: dout <= 8'b00000000; // 3973 :   0 - 0x0
      12'hF86: dout <= 8'b00000000; // 3974 :   0 - 0x0
      12'hF87: dout <= 8'b00000000; // 3975 :   0 - 0x0
      12'hF88: dout <= 8'b00000000; // 3976 :   0 - 0x0 -- plane 1
      12'hF89: dout <= 8'b00000000; // 3977 :   0 - 0x0
      12'hF8A: dout <= 8'b00000000; // 3978 :   0 - 0x0
      12'hF8B: dout <= 8'b00000000; // 3979 :   0 - 0x0
      12'hF8C: dout <= 8'b00000000; // 3980 :   0 - 0x0
      12'hF8D: dout <= 8'b00000000; // 3981 :   0 - 0x0
      12'hF8E: dout <= 8'b00000000; // 3982 :   0 - 0x0
      12'hF8F: dout <= 8'b00000000; // 3983 :   0 - 0x0
      12'hF90: dout <= 8'b00000000; // 3984 :   0 - 0x0 -- Sprite 0xf9
      12'hF91: dout <= 8'b00000000; // 3985 :   0 - 0x0
      12'hF92: dout <= 8'b00000000; // 3986 :   0 - 0x0
      12'hF93: dout <= 8'b00000000; // 3987 :   0 - 0x0
      12'hF94: dout <= 8'b00000000; // 3988 :   0 - 0x0
      12'hF95: dout <= 8'b00000000; // 3989 :   0 - 0x0
      12'hF96: dout <= 8'b00000000; // 3990 :   0 - 0x0
      12'hF97: dout <= 8'b00000000; // 3991 :   0 - 0x0
      12'hF98: dout <= 8'b00000000; // 3992 :   0 - 0x0 -- plane 1
      12'hF99: dout <= 8'b00000000; // 3993 :   0 - 0x0
      12'hF9A: dout <= 8'b00000000; // 3994 :   0 - 0x0
      12'hF9B: dout <= 8'b00000000; // 3995 :   0 - 0x0
      12'hF9C: dout <= 8'b00000000; // 3996 :   0 - 0x0
      12'hF9D: dout <= 8'b00000000; // 3997 :   0 - 0x0
      12'hF9E: dout <= 8'b00000000; // 3998 :   0 - 0x0
      12'hF9F: dout <= 8'b00000000; // 3999 :   0 - 0x0
      12'hFA0: dout <= 8'b00000000; // 4000 :   0 - 0x0 -- Sprite 0xfa
      12'hFA1: dout <= 8'b00000000; // 4001 :   0 - 0x0
      12'hFA2: dout <= 8'b00000000; // 4002 :   0 - 0x0
      12'hFA3: dout <= 8'b00000000; // 4003 :   0 - 0x0
      12'hFA4: dout <= 8'b00000000; // 4004 :   0 - 0x0
      12'hFA5: dout <= 8'b00000000; // 4005 :   0 - 0x0
      12'hFA6: dout <= 8'b00000000; // 4006 :   0 - 0x0
      12'hFA7: dout <= 8'b00000000; // 4007 :   0 - 0x0
      12'hFA8: dout <= 8'b00000000; // 4008 :   0 - 0x0 -- plane 1
      12'hFA9: dout <= 8'b00000000; // 4009 :   0 - 0x0
      12'hFAA: dout <= 8'b00000000; // 4010 :   0 - 0x0
      12'hFAB: dout <= 8'b00000000; // 4011 :   0 - 0x0
      12'hFAC: dout <= 8'b00000000; // 4012 :   0 - 0x0
      12'hFAD: dout <= 8'b00000000; // 4013 :   0 - 0x0
      12'hFAE: dout <= 8'b00000000; // 4014 :   0 - 0x0
      12'hFAF: dout <= 8'b00000000; // 4015 :   0 - 0x0
      12'hFB0: dout <= 8'b00000000; // 4016 :   0 - 0x0 -- Sprite 0xfb
      12'hFB1: dout <= 8'b00000000; // 4017 :   0 - 0x0
      12'hFB2: dout <= 8'b00000000; // 4018 :   0 - 0x0
      12'hFB3: dout <= 8'b00000000; // 4019 :   0 - 0x0
      12'hFB4: dout <= 8'b00000000; // 4020 :   0 - 0x0
      12'hFB5: dout <= 8'b00000000; // 4021 :   0 - 0x0
      12'hFB6: dout <= 8'b00000000; // 4022 :   0 - 0x0
      12'hFB7: dout <= 8'b00000000; // 4023 :   0 - 0x0
      12'hFB8: dout <= 8'b00000000; // 4024 :   0 - 0x0 -- plane 1
      12'hFB9: dout <= 8'b00000000; // 4025 :   0 - 0x0
      12'hFBA: dout <= 8'b00000000; // 4026 :   0 - 0x0
      12'hFBB: dout <= 8'b00000000; // 4027 :   0 - 0x0
      12'hFBC: dout <= 8'b00000000; // 4028 :   0 - 0x0
      12'hFBD: dout <= 8'b00000000; // 4029 :   0 - 0x0
      12'hFBE: dout <= 8'b00000000; // 4030 :   0 - 0x0
      12'hFBF: dout <= 8'b00000000; // 4031 :   0 - 0x0
      12'hFC0: dout <= 8'b00000000; // 4032 :   0 - 0x0 -- Sprite 0xfc
      12'hFC1: dout <= 8'b00000000; // 4033 :   0 - 0x0
      12'hFC2: dout <= 8'b10001110; // 4034 : 142 - 0x8e
      12'hFC3: dout <= 8'b10001010; // 4035 : 138 - 0x8a
      12'hFC4: dout <= 8'b10001010; // 4036 : 138 - 0x8a
      12'hFC5: dout <= 8'b10001010; // 4037 : 138 - 0x8a
      12'hFC6: dout <= 8'b10001010; // 4038 : 138 - 0x8a
      12'hFC7: dout <= 8'b11101110; // 4039 : 238 - 0xee
      12'hFC8: dout <= 8'b00000000; // 4040 :   0 - 0x0 -- plane 1
      12'hFC9: dout <= 8'b00000000; // 4041 :   0 - 0x0
      12'hFCA: dout <= 8'b00000000; // 4042 :   0 - 0x0
      12'hFCB: dout <= 8'b00000000; // 4043 :   0 - 0x0
      12'hFCC: dout <= 8'b00000000; // 4044 :   0 - 0x0
      12'hFCD: dout <= 8'b00000000; // 4045 :   0 - 0x0
      12'hFCE: dout <= 8'b00000000; // 4046 :   0 - 0x0
      12'hFCF: dout <= 8'b00000000; // 4047 :   0 - 0x0
      12'hFD0: dout <= 8'b00000000; // 4048 :   0 - 0x0 -- Sprite 0xfd
      12'hFD1: dout <= 8'b00000000; // 4049 :   0 - 0x0
      12'hFD2: dout <= 8'b01001100; // 4050 :  76 - 0x4c
      12'hFD3: dout <= 8'b10101010; // 4051 : 170 - 0xaa
      12'hFD4: dout <= 8'b10101010; // 4052 : 170 - 0xaa
      12'hFD5: dout <= 8'b11101010; // 4053 : 234 - 0xea
      12'hFD6: dout <= 8'b10101010; // 4054 : 170 - 0xaa
      12'hFD7: dout <= 8'b10101100; // 4055 : 172 - 0xac
      12'hFD8: dout <= 8'b00000000; // 4056 :   0 - 0x0 -- plane 1
      12'hFD9: dout <= 8'b00000000; // 4057 :   0 - 0x0
      12'hFDA: dout <= 8'b00000000; // 4058 :   0 - 0x0
      12'hFDB: dout <= 8'b00000000; // 4059 :   0 - 0x0
      12'hFDC: dout <= 8'b00000000; // 4060 :   0 - 0x0
      12'hFDD: dout <= 8'b00000000; // 4061 :   0 - 0x0
      12'hFDE: dout <= 8'b00000000; // 4062 :   0 - 0x0
      12'hFDF: dout <= 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout <= 8'b00000000; // 4064 :   0 - 0x0 -- Sprite 0xfe
      12'hFE1: dout <= 8'b00000000; // 4065 :   0 - 0x0
      12'hFE2: dout <= 8'b11101100; // 4066 : 236 - 0xec
      12'hFE3: dout <= 8'b01001010; // 4067 :  74 - 0x4a
      12'hFE4: dout <= 8'b01001010; // 4068 :  74 - 0x4a
      12'hFE5: dout <= 8'b01001010; // 4069 :  74 - 0x4a
      12'hFE6: dout <= 8'b01001010; // 4070 :  74 - 0x4a
      12'hFE7: dout <= 8'b11101010; // 4071 : 234 - 0xea
      12'hFE8: dout <= 8'b00000000; // 4072 :   0 - 0x0 -- plane 1
      12'hFE9: dout <= 8'b00000000; // 4073 :   0 - 0x0
      12'hFEA: dout <= 8'b00000000; // 4074 :   0 - 0x0
      12'hFEB: dout <= 8'b00000000; // 4075 :   0 - 0x0
      12'hFEC: dout <= 8'b00000000; // 4076 :   0 - 0x0
      12'hFED: dout <= 8'b00000000; // 4077 :   0 - 0x0
      12'hFEE: dout <= 8'b00000000; // 4078 :   0 - 0x0
      12'hFEF: dout <= 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout <= 8'b00000000; // 4080 :   0 - 0x0 -- Sprite 0xff
      12'hFF1: dout <= 8'b00000000; // 4081 :   0 - 0x0
      12'hFF2: dout <= 8'b01100000; // 4082 :  96 - 0x60
      12'hFF3: dout <= 8'b10001000; // 4083 : 136 - 0x88
      12'hFF4: dout <= 8'b10100000; // 4084 : 160 - 0xa0
      12'hFF5: dout <= 8'b10100000; // 4085 : 160 - 0xa0
      12'hFF6: dout <= 8'b10101000; // 4086 : 168 - 0xa8
      12'hFF7: dout <= 8'b01000000; // 4087 :  64 - 0x40
      12'hFF8: dout <= 8'b00000000; // 4088 :   0 - 0x0 -- plane 1
      12'hFF9: dout <= 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout <= 8'b00000000; // 4090 :   0 - 0x0
      12'hFFB: dout <= 8'b00000000; // 4091 :   0 - 0x0
      12'hFFC: dout <= 8'b00000000; // 4092 :   0 - 0x0
      12'hFFD: dout <= 8'b00000000; // 4093 :   0 - 0x0
      12'hFFE: dout <= 8'b00000000; // 4094 :   0 - 0x0
      12'hFFF: dout <= 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
