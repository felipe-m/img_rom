//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables
//- Only the first Name Table: 1KiB


//-  Original memory dump file name: donkeykong_ntable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_NTABLE_DONKEYKONG
  (
     input     clk,   // clock
     input      [10-1:0] addr,  //1024 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      10'h0: dout <= 8'b00100100; //    0 :  36 - 0x24 -- line 0x0
      10'h1: dout <= 8'b00100100; //    1 :  36 - 0x24
      10'h2: dout <= 8'b00100100; //    2 :  36 - 0x24
      10'h3: dout <= 8'b00100100; //    3 :  36 - 0x24
      10'h4: dout <= 8'b00100100; //    4 :  36 - 0x24
      10'h5: dout <= 8'b00100100; //    5 :  36 - 0x24
      10'h6: dout <= 8'b00100100; //    6 :  36 - 0x24
      10'h7: dout <= 8'b00100100; //    7 :  36 - 0x24
      10'h8: dout <= 8'b00100100; //    8 :  36 - 0x24
      10'h9: dout <= 8'b00100100; //    9 :  36 - 0x24
      10'hA: dout <= 8'b00100100; //   10 :  36 - 0x24
      10'hB: dout <= 8'b00100100; //   11 :  36 - 0x24
      10'hC: dout <= 8'b00100100; //   12 :  36 - 0x24
      10'hD: dout <= 8'b00100100; //   13 :  36 - 0x24
      10'hE: dout <= 8'b00100100; //   14 :  36 - 0x24
      10'hF: dout <= 8'b00100100; //   15 :  36 - 0x24
      10'h10: dout <= 8'b00100100; //   16 :  36 - 0x24
      10'h11: dout <= 8'b00100100; //   17 :  36 - 0x24
      10'h12: dout <= 8'b00100100; //   18 :  36 - 0x24
      10'h13: dout <= 8'b00100100; //   19 :  36 - 0x24
      10'h14: dout <= 8'b00100100; //   20 :  36 - 0x24
      10'h15: dout <= 8'b00100100; //   21 :  36 - 0x24
      10'h16: dout <= 8'b00100100; //   22 :  36 - 0x24
      10'h17: dout <= 8'b00100100; //   23 :  36 - 0x24
      10'h18: dout <= 8'b00100100; //   24 :  36 - 0x24
      10'h19: dout <= 8'b00100100; //   25 :  36 - 0x24
      10'h1A: dout <= 8'b00100100; //   26 :  36 - 0x24
      10'h1B: dout <= 8'b00100100; //   27 :  36 - 0x24
      10'h1C: dout <= 8'b00100100; //   28 :  36 - 0x24
      10'h1D: dout <= 8'b00100100; //   29 :  36 - 0x24
      10'h1E: dout <= 8'b00100100; //   30 :  36 - 0x24
      10'h1F: dout <= 8'b00100100; //   31 :  36 - 0x24
      10'h20: dout <= 8'b00100100; //   32 :  36 - 0x24 -- line 0x1
      10'h21: dout <= 8'b00100100; //   33 :  36 - 0x24
      10'h22: dout <= 8'b00100100; //   34 :  36 - 0x24
      10'h23: dout <= 8'b00100100; //   35 :  36 - 0x24
      10'h24: dout <= 8'b00100100; //   36 :  36 - 0x24
      10'h25: dout <= 8'b00100100; //   37 :  36 - 0x24
      10'h26: dout <= 8'b00100100; //   38 :  36 - 0x24
      10'h27: dout <= 8'b00100100; //   39 :  36 - 0x24
      10'h28: dout <= 8'b00100100; //   40 :  36 - 0x24
      10'h29: dout <= 8'b00100100; //   41 :  36 - 0x24
      10'h2A: dout <= 8'b00111111; //   42 :  63 - 0x3f
      10'h2B: dout <= 8'b00100100; //   43 :  36 - 0x24
      10'h2C: dout <= 8'b00111111; //   44 :  63 - 0x3f
      10'h2D: dout <= 8'b00100100; //   45 :  36 - 0x24
      10'h2E: dout <= 8'b00100100; //   46 :  36 - 0x24
      10'h2F: dout <= 8'b00100100; //   47 :  36 - 0x24
      10'h30: dout <= 8'b00100100; //   48 :  36 - 0x24
      10'h31: dout <= 8'b00100100; //   49 :  36 - 0x24
      10'h32: dout <= 8'b00100100; //   50 :  36 - 0x24
      10'h33: dout <= 8'b00100100; //   51 :  36 - 0x24
      10'h34: dout <= 8'b00100100; //   52 :  36 - 0x24
      10'h35: dout <= 8'b00100100; //   53 :  36 - 0x24
      10'h36: dout <= 8'b00100100; //   54 :  36 - 0x24
      10'h37: dout <= 8'b00100100; //   55 :  36 - 0x24
      10'h38: dout <= 8'b00100100; //   56 :  36 - 0x24
      10'h39: dout <= 8'b00100100; //   57 :  36 - 0x24
      10'h3A: dout <= 8'b00100100; //   58 :  36 - 0x24
      10'h3B: dout <= 8'b00100100; //   59 :  36 - 0x24
      10'h3C: dout <= 8'b00100100; //   60 :  36 - 0x24
      10'h3D: dout <= 8'b00100100; //   61 :  36 - 0x24
      10'h3E: dout <= 8'b00100100; //   62 :  36 - 0x24
      10'h3F: dout <= 8'b00100100; //   63 :  36 - 0x24
      10'h40: dout <= 8'b00100100; //   64 :  36 - 0x24 -- line 0x2
      10'h41: dout <= 8'b00100100; //   65 :  36 - 0x24
      10'h42: dout <= 8'b00100100; //   66 :  36 - 0x24
      10'h43: dout <= 8'b00100100; //   67 :  36 - 0x24
      10'h44: dout <= 8'b00100100; //   68 :  36 - 0x24
      10'h45: dout <= 8'b00100100; //   69 :  36 - 0x24
      10'h46: dout <= 8'b00100100; //   70 :  36 - 0x24
      10'h47: dout <= 8'b00100100; //   71 :  36 - 0x24
      10'h48: dout <= 8'b00100100; //   72 :  36 - 0x24
      10'h49: dout <= 8'b00100100; //   73 :  36 - 0x24
      10'h4A: dout <= 8'b00111111; //   74 :  63 - 0x3f
      10'h4B: dout <= 8'b00100100; //   75 :  36 - 0x24
      10'h4C: dout <= 8'b00111111; //   76 :  63 - 0x3f
      10'h4D: dout <= 8'b00100100; //   77 :  36 - 0x24
      10'h4E: dout <= 8'b00100100; //   78 :  36 - 0x24
      10'h4F: dout <= 8'b00100100; //   79 :  36 - 0x24
      10'h50: dout <= 8'b00100100; //   80 :  36 - 0x24
      10'h51: dout <= 8'b00100100; //   81 :  36 - 0x24
      10'h52: dout <= 8'b00100100; //   82 :  36 - 0x24
      10'h53: dout <= 8'b00100100; //   83 :  36 - 0x24
      10'h54: dout <= 8'b00100100; //   84 :  36 - 0x24
      10'h55: dout <= 8'b00100100; //   85 :  36 - 0x24
      10'h56: dout <= 8'b00100100; //   86 :  36 - 0x24
      10'h57: dout <= 8'b00100100; //   87 :  36 - 0x24
      10'h58: dout <= 8'b00100100; //   88 :  36 - 0x24
      10'h59: dout <= 8'b00100100; //   89 :  36 - 0x24
      10'h5A: dout <= 8'b00100100; //   90 :  36 - 0x24
      10'h5B: dout <= 8'b00100100; //   91 :  36 - 0x24
      10'h5C: dout <= 8'b00100100; //   92 :  36 - 0x24
      10'h5D: dout <= 8'b00100100; //   93 :  36 - 0x24
      10'h5E: dout <= 8'b00100100; //   94 :  36 - 0x24
      10'h5F: dout <= 8'b00100100; //   95 :  36 - 0x24
      10'h60: dout <= 8'b00100100; //   96 :  36 - 0x24 -- line 0x3
      10'h61: dout <= 8'b00100100; //   97 :  36 - 0x24
      10'h62: dout <= 8'b00100100; //   98 :  36 - 0x24
      10'h63: dout <= 8'b11111111; //   99 : 255 - 0xff
      10'h64: dout <= 8'b00000000; //  100 :   0 - 0x0
      10'h65: dout <= 8'b00000000; //  101 :   0 - 0x0
      10'h66: dout <= 8'b00000010; //  102 :   2 - 0x2
      10'h67: dout <= 8'b00000010; //  103 :   2 - 0x2
      10'h68: dout <= 8'b00000000; //  104 :   0 - 0x0
      10'h69: dout <= 8'b00000000; //  105 :   0 - 0x0
      10'h6A: dout <= 8'b00111111; //  106 :  63 - 0x3f
      10'h6B: dout <= 8'b00100100; //  107 :  36 - 0x24
      10'h6C: dout <= 8'b00111111; //  108 :  63 - 0x3f
      10'h6D: dout <= 8'b11010000; //  109 : 208 - 0xd0
      10'h6E: dout <= 8'b11010001; //  110 : 209 - 0xd1
      10'h6F: dout <= 8'b11010010; //  111 : 210 - 0xd2
      10'h70: dout <= 8'b00000000; //  112 :   0 - 0x0
      10'h71: dout <= 8'b00000000; //  113 :   0 - 0x0
      10'h72: dout <= 8'b00000010; //  114 :   2 - 0x2
      10'h73: dout <= 8'b00000010; //  115 :   2 - 0x2
      10'h74: dout <= 8'b00000000; //  116 :   0 - 0x0
      10'h75: dout <= 8'b00000000; //  117 :   0 - 0x0
      10'h76: dout <= 8'b00100100; //  118 :  36 - 0x24
      10'h77: dout <= 8'b00100100; //  119 :  36 - 0x24
      10'h78: dout <= 8'b00100100; //  120 :  36 - 0x24
      10'h79: dout <= 8'b00100100; //  121 :  36 - 0x24
      10'h7A: dout <= 8'b00100100; //  122 :  36 - 0x24
      10'h7B: dout <= 8'b00100100; //  123 :  36 - 0x24
      10'h7C: dout <= 8'b00100100; //  124 :  36 - 0x24
      10'h7D: dout <= 8'b00100100; //  125 :  36 - 0x24
      10'h7E: dout <= 8'b00100100; //  126 :  36 - 0x24
      10'h7F: dout <= 8'b00100100; //  127 :  36 - 0x24
      10'h80: dout <= 8'b00100100; //  128 :  36 - 0x24 -- line 0x4
      10'h81: dout <= 8'b01010000; //  129 :  80 - 0x50
      10'h82: dout <= 8'b01010100; //  130 :  84 - 0x54
      10'h83: dout <= 8'b01011000; //  131 :  88 - 0x58
      10'h84: dout <= 8'b00100100; //  132 :  36 - 0x24
      10'h85: dout <= 8'b00100100; //  133 :  36 - 0x24
      10'h86: dout <= 8'b10001100; //  134 : 140 - 0x8c
      10'h87: dout <= 8'b10010000; //  135 : 144 - 0x90
      10'h88: dout <= 8'b10010100; //  136 : 148 - 0x94
      10'h89: dout <= 8'b10011000; //  137 : 152 - 0x98
      10'h8A: dout <= 8'b00111111; //  138 :  63 - 0x3f
      10'h8B: dout <= 8'b00100100; //  139 :  36 - 0x24
      10'h8C: dout <= 8'b00111111; //  140 :  63 - 0x3f
      10'h8D: dout <= 8'b00100100; //  141 :  36 - 0x24
      10'h8E: dout <= 8'b00100100; //  142 :  36 - 0x24
      10'h8F: dout <= 8'b00100100; //  143 :  36 - 0x24
      10'h90: dout <= 8'b00100100; //  144 :  36 - 0x24
      10'h91: dout <= 8'b00100100; //  145 :  36 - 0x24
      10'h92: dout <= 8'b00100100; //  146 :  36 - 0x24
      10'h93: dout <= 8'b00100100; //  147 :  36 - 0x24
      10'h94: dout <= 8'b00100101; //  148 :  37 - 0x25
      10'h95: dout <= 8'b00010110; //  149 :  22 - 0x16
      10'h96: dout <= 8'b00101010; //  150 :  42 - 0x2a
      10'h97: dout <= 8'b00100110; //  151 :  38 - 0x26
      10'h98: dout <= 8'b00100111; //  152 :  39 - 0x27
      10'h99: dout <= 8'b00101000; //  153 :  40 - 0x28
      10'h9A: dout <= 8'b00101001; //  154 :  41 - 0x29
      10'h9B: dout <= 8'b00101010; //  155 :  42 - 0x2a
      10'h9C: dout <= 8'b00010101; //  156 :  21 - 0x15
      10'h9D: dout <= 8'b00101101; //  157 :  45 - 0x2d
      10'h9E: dout <= 8'b00100100; //  158 :  36 - 0x24
      10'h9F: dout <= 8'b00100100; //  159 :  36 - 0x24
      10'hA0: dout <= 8'b00100100; //  160 :  36 - 0x24 -- line 0x5
      10'hA1: dout <= 8'b01010001; //  161 :  81 - 0x51
      10'hA2: dout <= 8'b01010101; //  162 :  85 - 0x55
      10'hA3: dout <= 8'b01011001; //  163 :  89 - 0x59
      10'hA4: dout <= 8'b00100100; //  164 :  36 - 0x24
      10'hA5: dout <= 8'b00100100; //  165 :  36 - 0x24
      10'hA6: dout <= 8'b10001101; //  166 : 141 - 0x8d
      10'hA7: dout <= 8'b10010001; //  167 : 145 - 0x91
      10'hA8: dout <= 8'b10010101; //  168 : 149 - 0x95
      10'hA9: dout <= 8'b10011001; //  169 : 153 - 0x99
      10'hAA: dout <= 8'b00111111; //  170 :  63 - 0x3f
      10'hAB: dout <= 8'b00100100; //  171 :  36 - 0x24
      10'hAC: dout <= 8'b00111111; //  172 :  63 - 0x3f
      10'hAD: dout <= 8'b00110000; //  173 :  48 - 0x30
      10'hAE: dout <= 8'b00110000; //  174 :  48 - 0x30
      10'hAF: dout <= 8'b00110000; //  175 :  48 - 0x30
      10'hB0: dout <= 8'b00110000; //  176 :  48 - 0x30
      10'hB1: dout <= 8'b00110000; //  177 :  48 - 0x30
      10'hB2: dout <= 8'b00110000; //  178 :  48 - 0x30
      10'hB3: dout <= 8'b00100100; //  179 :  36 - 0x24
      10'hB4: dout <= 8'b00101011; //  180 :  43 - 0x2b
      10'hB5: dout <= 8'b00000010; //  181 :   2 - 0x2
      10'hB6: dout <= 8'b00101100; //  182 :  44 - 0x2c
      10'hB7: dout <= 8'b00000011; //  183 :   3 - 0x3
      10'hB8: dout <= 8'b00000000; //  184 :   0 - 0x0
      10'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      10'hBA: dout <= 8'b00000000; //  186 :   0 - 0x0
      10'hBB: dout <= 8'b00101100; //  187 :  44 - 0x2c
      10'hBC: dout <= 8'b00000001; //  188 :   1 - 0x1
      10'hBD: dout <= 8'b00101111; //  189 :  47 - 0x2f
      10'hBE: dout <= 8'b00100100; //  190 :  36 - 0x24
      10'hBF: dout <= 8'b00100100; //  191 :  36 - 0x24
      10'hC0: dout <= 8'b00100100; //  192 :  36 - 0x24 -- line 0x6
      10'hC1: dout <= 8'b01010010; //  193 :  82 - 0x52
      10'hC2: dout <= 8'b01010110; //  194 :  86 - 0x56
      10'hC3: dout <= 8'b01011010; //  195 :  90 - 0x5a
      10'hC4: dout <= 8'b00100100; //  196 :  36 - 0x24
      10'hC5: dout <= 8'b10001010; //  197 : 138 - 0x8a
      10'hC6: dout <= 8'b10001110; //  198 : 142 - 0x8e
      10'hC7: dout <= 8'b10010010; //  199 : 146 - 0x92
      10'hC8: dout <= 8'b10010110; //  200 : 150 - 0x96
      10'hC9: dout <= 8'b10011010; //  201 : 154 - 0x9a
      10'hCA: dout <= 8'b00110000; //  202 :  48 - 0x30
      10'hCB: dout <= 8'b00110000; //  203 :  48 - 0x30
      10'hCC: dout <= 8'b00110000; //  204 :  48 - 0x30
      10'hCD: dout <= 8'b00100100; //  205 :  36 - 0x24
      10'hCE: dout <= 8'b00100100; //  206 :  36 - 0x24
      10'hCF: dout <= 8'b00100100; //  207 :  36 - 0x24
      10'hD0: dout <= 8'b00100100; //  208 :  36 - 0x24
      10'hD1: dout <= 8'b00100100; //  209 :  36 - 0x24
      10'hD2: dout <= 8'b00111111; //  210 :  63 - 0x3f
      10'hD3: dout <= 8'b00100100; //  211 :  36 - 0x24
      10'hD4: dout <= 8'b00100100; //  212 :  36 - 0x24
      10'hD5: dout <= 8'b00100100; //  213 :  36 - 0x24
      10'hD6: dout <= 8'b00100100; //  214 :  36 - 0x24
      10'hD7: dout <= 8'b00100100; //  215 :  36 - 0x24
      10'hD8: dout <= 8'b00100100; //  216 :  36 - 0x24
      10'hD9: dout <= 8'b00100100; //  217 :  36 - 0x24
      10'hDA: dout <= 8'b00100100; //  218 :  36 - 0x24
      10'hDB: dout <= 8'b00100100; //  219 :  36 - 0x24
      10'hDC: dout <= 8'b00100100; //  220 :  36 - 0x24
      10'hDD: dout <= 8'b00100100; //  221 :  36 - 0x24
      10'hDE: dout <= 8'b00100100; //  222 :  36 - 0x24
      10'hDF: dout <= 8'b00100100; //  223 :  36 - 0x24
      10'hE0: dout <= 8'b00100100; //  224 :  36 - 0x24 -- line 0x7
      10'hE1: dout <= 8'b01010011; //  225 :  83 - 0x53
      10'hE2: dout <= 8'b01010111; //  226 :  87 - 0x57
      10'hE3: dout <= 8'b01011011; //  227 :  91 - 0x5b
      10'hE4: dout <= 8'b10001001; //  228 : 137 - 0x89
      10'hE5: dout <= 8'b10001011; //  229 : 139 - 0x8b
      10'hE6: dout <= 8'b10001111; //  230 : 143 - 0x8f
      10'hE7: dout <= 8'b10010011; //  231 : 147 - 0x93
      10'hE8: dout <= 8'b10010111; //  232 : 151 - 0x97
      10'hE9: dout <= 8'b10011011; //  233 : 155 - 0x9b
      10'hEA: dout <= 8'b00111111; //  234 :  63 - 0x3f
      10'hEB: dout <= 8'b00100100; //  235 :  36 - 0x24
      10'hEC: dout <= 8'b00111111; //  236 :  63 - 0x3f
      10'hED: dout <= 8'b00100100; //  237 :  36 - 0x24
      10'hEE: dout <= 8'b00100100; //  238 :  36 - 0x24
      10'hEF: dout <= 8'b00100100; //  239 :  36 - 0x24
      10'hF0: dout <= 8'b00100100; //  240 :  36 - 0x24
      10'hF1: dout <= 8'b00100100; //  241 :  36 - 0x24
      10'hF2: dout <= 8'b00111111; //  242 :  63 - 0x3f
      10'hF3: dout <= 8'b00100100; //  243 :  36 - 0x24
      10'hF4: dout <= 8'b00100100; //  244 :  36 - 0x24
      10'hF5: dout <= 8'b00100100; //  245 :  36 - 0x24
      10'hF6: dout <= 8'b00100100; //  246 :  36 - 0x24
      10'hF7: dout <= 8'b00100100; //  247 :  36 - 0x24
      10'hF8: dout <= 8'b00100100; //  248 :  36 - 0x24
      10'hF9: dout <= 8'b00100100; //  249 :  36 - 0x24
      10'hFA: dout <= 8'b00100100; //  250 :  36 - 0x24
      10'hFB: dout <= 8'b00100100; //  251 :  36 - 0x24
      10'hFC: dout <= 8'b00100100; //  252 :  36 - 0x24
      10'hFD: dout <= 8'b00100100; //  253 :  36 - 0x24
      10'hFE: dout <= 8'b00100100; //  254 :  36 - 0x24
      10'hFF: dout <= 8'b00100100; //  255 :  36 - 0x24
      10'h100: dout <= 8'b00100100; //  256 :  36 - 0x24 -- line 0x8
      10'h101: dout <= 8'b00100100; //  257 :  36 - 0x24
      10'h102: dout <= 8'b00110000; //  258 :  48 - 0x30
      10'h103: dout <= 8'b00110000; //  259 :  48 - 0x30
      10'h104: dout <= 8'b00110000; //  260 :  48 - 0x30
      10'h105: dout <= 8'b00110000; //  261 :  48 - 0x30
      10'h106: dout <= 8'b00110000; //  262 :  48 - 0x30
      10'h107: dout <= 8'b00110000; //  263 :  48 - 0x30
      10'h108: dout <= 8'b00110000; //  264 :  48 - 0x30
      10'h109: dout <= 8'b00110000; //  265 :  48 - 0x30
      10'h10A: dout <= 8'b00110000; //  266 :  48 - 0x30
      10'h10B: dout <= 8'b00110000; //  267 :  48 - 0x30
      10'h10C: dout <= 8'b00110000; //  268 :  48 - 0x30
      10'h10D: dout <= 8'b00110000; //  269 :  48 - 0x30
      10'h10E: dout <= 8'b00110000; //  270 :  48 - 0x30
      10'h10F: dout <= 8'b00110000; //  271 :  48 - 0x30
      10'h110: dout <= 8'b00111110; //  272 :  62 - 0x3e
      10'h111: dout <= 8'b00111110; //  273 :  62 - 0x3e
      10'h112: dout <= 8'b01000101; //  274 :  69 - 0x45
      10'h113: dout <= 8'b00111101; //  275 :  61 - 0x3d
      10'h114: dout <= 8'b00111101; //  276 :  61 - 0x3d
      10'h115: dout <= 8'b00111101; //  277 :  61 - 0x3d
      10'h116: dout <= 8'b00111100; //  278 :  60 - 0x3c
      10'h117: dout <= 8'b00111100; //  279 :  60 - 0x3c
      10'h118: dout <= 8'b00111100; //  280 :  60 - 0x3c
      10'h119: dout <= 8'b00111011; //  281 :  59 - 0x3b
      10'h11A: dout <= 8'b00111011; //  282 :  59 - 0x3b
      10'h11B: dout <= 8'b00111011; //  283 :  59 - 0x3b
      10'h11C: dout <= 8'b00100100; //  284 :  36 - 0x24
      10'h11D: dout <= 8'b00100100; //  285 :  36 - 0x24
      10'h11E: dout <= 8'b00100100; //  286 :  36 - 0x24
      10'h11F: dout <= 8'b00100100; //  287 :  36 - 0x24
      10'h120: dout <= 8'b00100100; //  288 :  36 - 0x24 -- line 0x9
      10'h121: dout <= 8'b00100100; //  289 :  36 - 0x24
      10'h122: dout <= 8'b00100100; //  290 :  36 - 0x24
      10'h123: dout <= 8'b00100100; //  291 :  36 - 0x24
      10'h124: dout <= 8'b00100100; //  292 :  36 - 0x24
      10'h125: dout <= 8'b00100100; //  293 :  36 - 0x24
      10'h126: dout <= 8'b00100100; //  294 :  36 - 0x24
      10'h127: dout <= 8'b00100100; //  295 :  36 - 0x24
      10'h128: dout <= 8'b00100100; //  296 :  36 - 0x24
      10'h129: dout <= 8'b00100100; //  297 :  36 - 0x24
      10'h12A: dout <= 8'b00100100; //  298 :  36 - 0x24
      10'h12B: dout <= 8'b00100100; //  299 :  36 - 0x24
      10'h12C: dout <= 8'b00100100; //  300 :  36 - 0x24
      10'h12D: dout <= 8'b00111111; //  301 :  63 - 0x3f
      10'h12E: dout <= 8'b00100100; //  302 :  36 - 0x24
      10'h12F: dout <= 8'b00100100; //  303 :  36 - 0x24
      10'h130: dout <= 8'b00110111; //  304 :  55 - 0x37
      10'h131: dout <= 8'b00110111; //  305 :  55 - 0x37
      10'h132: dout <= 8'b00110111; //  306 :  55 - 0x37
      10'h133: dout <= 8'b00110110; //  307 :  54 - 0x36
      10'h134: dout <= 8'b00110110; //  308 :  54 - 0x36
      10'h135: dout <= 8'b00110110; //  309 :  54 - 0x36
      10'h136: dout <= 8'b00110101; //  310 :  53 - 0x35
      10'h137: dout <= 8'b00110101; //  311 :  53 - 0x35
      10'h138: dout <= 8'b00110101; //  312 :  53 - 0x35
      10'h139: dout <= 8'b01001001; //  313 :  73 - 0x49
      10'h13A: dout <= 8'b00110100; //  314 :  52 - 0x34
      10'h13B: dout <= 8'b00110100; //  315 :  52 - 0x34
      10'h13C: dout <= 8'b00100100; //  316 :  36 - 0x24
      10'h13D: dout <= 8'b00100100; //  317 :  36 - 0x24
      10'h13E: dout <= 8'b00100100; //  318 :  36 - 0x24
      10'h13F: dout <= 8'b00100100; //  319 :  36 - 0x24
      10'h140: dout <= 8'b00100100; //  320 :  36 - 0x24 -- line 0xa
      10'h141: dout <= 8'b00100100; //  321 :  36 - 0x24
      10'h142: dout <= 8'b00100100; //  322 :  36 - 0x24
      10'h143: dout <= 8'b00100100; //  323 :  36 - 0x24
      10'h144: dout <= 8'b00100100; //  324 :  36 - 0x24
      10'h145: dout <= 8'b00100100; //  325 :  36 - 0x24
      10'h146: dout <= 8'b00100100; //  326 :  36 - 0x24
      10'h147: dout <= 8'b00100100; //  327 :  36 - 0x24
      10'h148: dout <= 8'b00100100; //  328 :  36 - 0x24
      10'h149: dout <= 8'b00100100; //  329 :  36 - 0x24
      10'h14A: dout <= 8'b00100100; //  330 :  36 - 0x24
      10'h14B: dout <= 8'b00100100; //  331 :  36 - 0x24
      10'h14C: dout <= 8'b00100100; //  332 :  36 - 0x24
      10'h14D: dout <= 8'b00100100; //  333 :  36 - 0x24
      10'h14E: dout <= 8'b00100100; //  334 :  36 - 0x24
      10'h14F: dout <= 8'b00100100; //  335 :  36 - 0x24
      10'h150: dout <= 8'b00100100; //  336 :  36 - 0x24
      10'h151: dout <= 8'b00100100; //  337 :  36 - 0x24
      10'h152: dout <= 8'b00100100; //  338 :  36 - 0x24
      10'h153: dout <= 8'b00100100; //  339 :  36 - 0x24
      10'h154: dout <= 8'b00100100; //  340 :  36 - 0x24
      10'h155: dout <= 8'b00100100; //  341 :  36 - 0x24
      10'h156: dout <= 8'b00100100; //  342 :  36 - 0x24
      10'h157: dout <= 8'b00100100; //  343 :  36 - 0x24
      10'h158: dout <= 8'b00100100; //  344 :  36 - 0x24
      10'h159: dout <= 8'b00111111; //  345 :  63 - 0x3f
      10'h15A: dout <= 8'b00100100; //  346 :  36 - 0x24
      10'h15B: dout <= 8'b00100100; //  347 :  36 - 0x24
      10'h15C: dout <= 8'b00100100; //  348 :  36 - 0x24
      10'h15D: dout <= 8'b00100100; //  349 :  36 - 0x24
      10'h15E: dout <= 8'b00100100; //  350 :  36 - 0x24
      10'h15F: dout <= 8'b00100100; //  351 :  36 - 0x24
      10'h160: dout <= 8'b00100100; //  352 :  36 - 0x24 -- line 0xb
      10'h161: dout <= 8'b00100100; //  353 :  36 - 0x24
      10'h162: dout <= 8'b00100100; //  354 :  36 - 0x24
      10'h163: dout <= 8'b00100100; //  355 :  36 - 0x24
      10'h164: dout <= 8'b00100100; //  356 :  36 - 0x24
      10'h165: dout <= 8'b00100100; //  357 :  36 - 0x24
      10'h166: dout <= 8'b00100100; //  358 :  36 - 0x24
      10'h167: dout <= 8'b00100100; //  359 :  36 - 0x24
      10'h168: dout <= 8'b00100100; //  360 :  36 - 0x24
      10'h169: dout <= 8'b00100100; //  361 :  36 - 0x24
      10'h16A: dout <= 8'b00100100; //  362 :  36 - 0x24
      10'h16B: dout <= 8'b00100100; //  363 :  36 - 0x24
      10'h16C: dout <= 8'b00100100; //  364 :  36 - 0x24
      10'h16D: dout <= 8'b01000000; //  365 :  64 - 0x40
      10'h16E: dout <= 8'b00111000; //  366 :  56 - 0x38
      10'h16F: dout <= 8'b00111000; //  367 :  56 - 0x38
      10'h170: dout <= 8'b00111001; //  368 :  57 - 0x39
      10'h171: dout <= 8'b00111001; //  369 :  57 - 0x39
      10'h172: dout <= 8'b00111001; //  370 :  57 - 0x39
      10'h173: dout <= 8'b00111010; //  371 :  58 - 0x3a
      10'h174: dout <= 8'b00111010; //  372 :  58 - 0x3a
      10'h175: dout <= 8'b00111010; //  373 :  58 - 0x3a
      10'h176: dout <= 8'b00111011; //  374 :  59 - 0x3b
      10'h177: dout <= 8'b00111011; //  375 :  59 - 0x3b
      10'h178: dout <= 8'b00111011; //  376 :  59 - 0x3b
      10'h179: dout <= 8'b01000011; //  377 :  67 - 0x43
      10'h17A: dout <= 8'b00111100; //  378 :  60 - 0x3c
      10'h17B: dout <= 8'b00111100; //  379 :  60 - 0x3c
      10'h17C: dout <= 8'b00111101; //  380 :  61 - 0x3d
      10'h17D: dout <= 8'b00111101; //  381 :  61 - 0x3d
      10'h17E: dout <= 8'b00100100; //  382 :  36 - 0x24
      10'h17F: dout <= 8'b00100100; //  383 :  36 - 0x24
      10'h180: dout <= 8'b00100100; //  384 :  36 - 0x24 -- line 0xc
      10'h181: dout <= 8'b00100100; //  385 :  36 - 0x24
      10'h182: dout <= 8'b00100100; //  386 :  36 - 0x24
      10'h183: dout <= 8'b00100100; //  387 :  36 - 0x24
      10'h184: dout <= 8'b00111101; //  388 :  61 - 0x3d
      10'h185: dout <= 8'b00111101; //  389 :  61 - 0x3d
      10'h186: dout <= 8'b00111101; //  390 :  61 - 0x3d
      10'h187: dout <= 8'b00111110; //  391 :  62 - 0x3e
      10'h188: dout <= 8'b00111110; //  392 :  62 - 0x3e
      10'h189: dout <= 8'b00111110; //  393 :  62 - 0x3e
      10'h18A: dout <= 8'b00110000; //  394 :  48 - 0x30
      10'h18B: dout <= 8'b00110000; //  395 :  48 - 0x30
      10'h18C: dout <= 8'b00110000; //  396 :  48 - 0x30
      10'h18D: dout <= 8'b00110001; //  397 :  49 - 0x31
      10'h18E: dout <= 8'b00110001; //  398 :  49 - 0x31
      10'h18F: dout <= 8'b00110001; //  399 :  49 - 0x31
      10'h190: dout <= 8'b00110010; //  400 :  50 - 0x32
      10'h191: dout <= 8'b00110010; //  401 :  50 - 0x32
      10'h192: dout <= 8'b00110010; //  402 :  50 - 0x32
      10'h193: dout <= 8'b00110011; //  403 :  51 - 0x33
      10'h194: dout <= 8'b00110011; //  404 :  51 - 0x33
      10'h195: dout <= 8'b00110011; //  405 :  51 - 0x33
      10'h196: dout <= 8'b00110100; //  406 :  52 - 0x34
      10'h197: dout <= 8'b01001001; //  407 :  73 - 0x49
      10'h198: dout <= 8'b00110100; //  408 :  52 - 0x34
      10'h199: dout <= 8'b00110101; //  409 :  53 - 0x35
      10'h19A: dout <= 8'b00110101; //  410 :  53 - 0x35
      10'h19B: dout <= 8'b00110101; //  411 :  53 - 0x35
      10'h19C: dout <= 8'b00110110; //  412 :  54 - 0x36
      10'h19D: dout <= 8'b00110110; //  413 :  54 - 0x36
      10'h19E: dout <= 8'b00100100; //  414 :  36 - 0x24
      10'h19F: dout <= 8'b00100100; //  415 :  36 - 0x24
      10'h1A0: dout <= 8'b00100100; //  416 :  36 - 0x24 -- line 0xd
      10'h1A1: dout <= 8'b00100100; //  417 :  36 - 0x24
      10'h1A2: dout <= 8'b00100100; //  418 :  36 - 0x24
      10'h1A3: dout <= 8'b00100100; //  419 :  36 - 0x24
      10'h1A4: dout <= 8'b00110110; //  420 :  54 - 0x36
      10'h1A5: dout <= 8'b00110110; //  421 :  54 - 0x36
      10'h1A6: dout <= 8'b01001011; //  422 :  75 - 0x4b
      10'h1A7: dout <= 8'b00110111; //  423 :  55 - 0x37
      10'h1A8: dout <= 8'b00110111; //  424 :  55 - 0x37
      10'h1A9: dout <= 8'b00110111; //  425 :  55 - 0x37
      10'h1AA: dout <= 8'b00100100; //  426 :  36 - 0x24
      10'h1AB: dout <= 8'b00111111; //  427 :  63 - 0x3f
      10'h1AC: dout <= 8'b00100100; //  428 :  36 - 0x24
      10'h1AD: dout <= 8'b00100100; //  429 :  36 - 0x24
      10'h1AE: dout <= 8'b00100100; //  430 :  36 - 0x24
      10'h1AF: dout <= 8'b00100100; //  431 :  36 - 0x24
      10'h1B0: dout <= 8'b00100100; //  432 :  36 - 0x24
      10'h1B1: dout <= 8'b00100100; //  433 :  36 - 0x24
      10'h1B2: dout <= 8'b00100100; //  434 :  36 - 0x24
      10'h1B3: dout <= 8'b00100100; //  435 :  36 - 0x24
      10'h1B4: dout <= 8'b00100100; //  436 :  36 - 0x24
      10'h1B5: dout <= 8'b00100100; //  437 :  36 - 0x24
      10'h1B6: dout <= 8'b00100100; //  438 :  36 - 0x24
      10'h1B7: dout <= 8'b00100100; //  439 :  36 - 0x24
      10'h1B8: dout <= 8'b00100100; //  440 :  36 - 0x24
      10'h1B9: dout <= 8'b00100100; //  441 :  36 - 0x24
      10'h1BA: dout <= 8'b00100100; //  442 :  36 - 0x24
      10'h1BB: dout <= 8'b00100100; //  443 :  36 - 0x24
      10'h1BC: dout <= 8'b00100100; //  444 :  36 - 0x24
      10'h1BD: dout <= 8'b00100100; //  445 :  36 - 0x24
      10'h1BE: dout <= 8'b00100100; //  446 :  36 - 0x24
      10'h1BF: dout <= 8'b00100100; //  447 :  36 - 0x24
      10'h1C0: dout <= 8'b00100100; //  448 :  36 - 0x24 -- line 0xe
      10'h1C1: dout <= 8'b00100100; //  449 :  36 - 0x24
      10'h1C2: dout <= 8'b00100100; //  450 :  36 - 0x24
      10'h1C3: dout <= 8'b00100100; //  451 :  36 - 0x24
      10'h1C4: dout <= 8'b00100100; //  452 :  36 - 0x24
      10'h1C5: dout <= 8'b00100100; //  453 :  36 - 0x24
      10'h1C6: dout <= 8'b00111111; //  454 :  63 - 0x3f
      10'h1C7: dout <= 8'b00100100; //  455 :  36 - 0x24
      10'h1C8: dout <= 8'b00100100; //  456 :  36 - 0x24
      10'h1C9: dout <= 8'b00100100; //  457 :  36 - 0x24
      10'h1CA: dout <= 8'b00100100; //  458 :  36 - 0x24
      10'h1CB: dout <= 8'b00111111; //  459 :  63 - 0x3f
      10'h1CC: dout <= 8'b00100100; //  460 :  36 - 0x24
      10'h1CD: dout <= 8'b00100100; //  461 :  36 - 0x24
      10'h1CE: dout <= 8'b00100100; //  462 :  36 - 0x24
      10'h1CF: dout <= 8'b00100100; //  463 :  36 - 0x24
      10'h1D0: dout <= 8'b00100100; //  464 :  36 - 0x24
      10'h1D1: dout <= 8'b00100100; //  465 :  36 - 0x24
      10'h1D2: dout <= 8'b00100100; //  466 :  36 - 0x24
      10'h1D3: dout <= 8'b00100100; //  467 :  36 - 0x24
      10'h1D4: dout <= 8'b00100100; //  468 :  36 - 0x24
      10'h1D5: dout <= 8'b00100100; //  469 :  36 - 0x24
      10'h1D6: dout <= 8'b00100100; //  470 :  36 - 0x24
      10'h1D7: dout <= 8'b00100100; //  471 :  36 - 0x24
      10'h1D8: dout <= 8'b00100100; //  472 :  36 - 0x24
      10'h1D9: dout <= 8'b00100100; //  473 :  36 - 0x24
      10'h1DA: dout <= 8'b00100100; //  474 :  36 - 0x24
      10'h1DB: dout <= 8'b00100100; //  475 :  36 - 0x24
      10'h1DC: dout <= 8'b00100100; //  476 :  36 - 0x24
      10'h1DD: dout <= 8'b00100100; //  477 :  36 - 0x24
      10'h1DE: dout <= 8'b00100100; //  478 :  36 - 0x24
      10'h1DF: dout <= 8'b00100100; //  479 :  36 - 0x24
      10'h1E0: dout <= 8'b00100100; //  480 :  36 - 0x24 -- line 0xf
      10'h1E1: dout <= 8'b00100100; //  481 :  36 - 0x24
      10'h1E2: dout <= 8'b00110000; //  482 :  48 - 0x30
      10'h1E3: dout <= 8'b00110000; //  483 :  48 - 0x30
      10'h1E4: dout <= 8'b00111110; //  484 :  62 - 0x3e
      10'h1E5: dout <= 8'b00111110; //  485 :  62 - 0x3e
      10'h1E6: dout <= 8'b01000101; //  486 :  69 - 0x45
      10'h1E7: dout <= 8'b00111101; //  487 :  61 - 0x3d
      10'h1E8: dout <= 8'b00111101; //  488 :  61 - 0x3d
      10'h1E9: dout <= 8'b00111101; //  489 :  61 - 0x3d
      10'h1EA: dout <= 8'b00111100; //  490 :  60 - 0x3c
      10'h1EB: dout <= 8'b01000011; //  491 :  67 - 0x43
      10'h1EC: dout <= 8'b00111100; //  492 :  60 - 0x3c
      10'h1ED: dout <= 8'b00111011; //  493 :  59 - 0x3b
      10'h1EE: dout <= 8'b00111011; //  494 :  59 - 0x3b
      10'h1EF: dout <= 8'b00111011; //  495 :  59 - 0x3b
      10'h1F0: dout <= 8'b00111010; //  496 :  58 - 0x3a
      10'h1F1: dout <= 8'b00111010; //  497 :  58 - 0x3a
      10'h1F2: dout <= 8'b00111010; //  498 :  58 - 0x3a
      10'h1F3: dout <= 8'b00111001; //  499 :  57 - 0x39
      10'h1F4: dout <= 8'b00111001; //  500 :  57 - 0x39
      10'h1F5: dout <= 8'b00111001; //  501 :  57 - 0x39
      10'h1F6: dout <= 8'b00111000; //  502 :  56 - 0x38
      10'h1F7: dout <= 8'b01000000; //  503 :  64 - 0x40
      10'h1F8: dout <= 8'b00111000; //  504 :  56 - 0x38
      10'h1F9: dout <= 8'b00100100; //  505 :  36 - 0x24
      10'h1FA: dout <= 8'b00100100; //  506 :  36 - 0x24
      10'h1FB: dout <= 8'b00100100; //  507 :  36 - 0x24
      10'h1FC: dout <= 8'b00100100; //  508 :  36 - 0x24
      10'h1FD: dout <= 8'b00100100; //  509 :  36 - 0x24
      10'h1FE: dout <= 8'b00100100; //  510 :  36 - 0x24
      10'h1FF: dout <= 8'b00100100; //  511 :  36 - 0x24
      10'h200: dout <= 8'b00100100; //  512 :  36 - 0x24 -- line 0x10
      10'h201: dout <= 8'b00100100; //  513 :  36 - 0x24
      10'h202: dout <= 8'b00100100; //  514 :  36 - 0x24
      10'h203: dout <= 8'b00100100; //  515 :  36 - 0x24
      10'h204: dout <= 8'b00110111; //  516 :  55 - 0x37
      10'h205: dout <= 8'b00110111; //  517 :  55 - 0x37
      10'h206: dout <= 8'b00110111; //  518 :  55 - 0x37
      10'h207: dout <= 8'b00110110; //  519 :  54 - 0x36
      10'h208: dout <= 8'b00110110; //  520 :  54 - 0x36
      10'h209: dout <= 8'b00110110; //  521 :  54 - 0x36
      10'h20A: dout <= 8'b01001010; //  522 :  74 - 0x4a
      10'h20B: dout <= 8'b00110101; //  523 :  53 - 0x35
      10'h20C: dout <= 8'b00110101; //  524 :  53 - 0x35
      10'h20D: dout <= 8'b00110100; //  525 :  52 - 0x34
      10'h20E: dout <= 8'b00110100; //  526 :  52 - 0x34
      10'h20F: dout <= 8'b00110100; //  527 :  52 - 0x34
      10'h210: dout <= 8'b01001000; //  528 :  72 - 0x48
      10'h211: dout <= 8'b00110011; //  529 :  51 - 0x33
      10'h212: dout <= 8'b00110011; //  530 :  51 - 0x33
      10'h213: dout <= 8'b00110010; //  531 :  50 - 0x32
      10'h214: dout <= 8'b00110010; //  532 :  50 - 0x32
      10'h215: dout <= 8'b00110010; //  533 :  50 - 0x32
      10'h216: dout <= 8'b00110001; //  534 :  49 - 0x31
      10'h217: dout <= 8'b00110001; //  535 :  49 - 0x31
      10'h218: dout <= 8'b00110001; //  536 :  49 - 0x31
      10'h219: dout <= 8'b00110000; //  537 :  48 - 0x30
      10'h21A: dout <= 8'b00110000; //  538 :  48 - 0x30
      10'h21B: dout <= 8'b00110000; //  539 :  48 - 0x30
      10'h21C: dout <= 8'b00100100; //  540 :  36 - 0x24
      10'h21D: dout <= 8'b00100100; //  541 :  36 - 0x24
      10'h21E: dout <= 8'b00100100; //  542 :  36 - 0x24
      10'h21F: dout <= 8'b00100100; //  543 :  36 - 0x24
      10'h220: dout <= 8'b00100100; //  544 :  36 - 0x24 -- line 0x11
      10'h221: dout <= 8'b00100100; //  545 :  36 - 0x24
      10'h222: dout <= 8'b00100100; //  546 :  36 - 0x24
      10'h223: dout <= 8'b00100100; //  547 :  36 - 0x24
      10'h224: dout <= 8'b00100100; //  548 :  36 - 0x24
      10'h225: dout <= 8'b00100100; //  549 :  36 - 0x24
      10'h226: dout <= 8'b00100100; //  550 :  36 - 0x24
      10'h227: dout <= 8'b00100100; //  551 :  36 - 0x24
      10'h228: dout <= 8'b00100100; //  552 :  36 - 0x24
      10'h229: dout <= 8'b00100100; //  553 :  36 - 0x24
      10'h22A: dout <= 8'b00100100; //  554 :  36 - 0x24
      10'h22B: dout <= 8'b00100100; //  555 :  36 - 0x24
      10'h22C: dout <= 8'b00100100; //  556 :  36 - 0x24
      10'h22D: dout <= 8'b00100100; //  557 :  36 - 0x24
      10'h22E: dout <= 8'b00100100; //  558 :  36 - 0x24
      10'h22F: dout <= 8'b00100100; //  559 :  36 - 0x24
      10'h230: dout <= 8'b00111111; //  560 :  63 - 0x3f
      10'h231: dout <= 8'b00100100; //  561 :  36 - 0x24
      10'h232: dout <= 8'b00100100; //  562 :  36 - 0x24
      10'h233: dout <= 8'b00100100; //  563 :  36 - 0x24
      10'h234: dout <= 8'b00100100; //  564 :  36 - 0x24
      10'h235: dout <= 8'b00100100; //  565 :  36 - 0x24
      10'h236: dout <= 8'b00100100; //  566 :  36 - 0x24
      10'h237: dout <= 8'b00100100; //  567 :  36 - 0x24
      10'h238: dout <= 8'b00100100; //  568 :  36 - 0x24
      10'h239: dout <= 8'b00111111; //  569 :  63 - 0x3f
      10'h23A: dout <= 8'b00100100; //  570 :  36 - 0x24
      10'h23B: dout <= 8'b00100100; //  571 :  36 - 0x24
      10'h23C: dout <= 8'b00100100; //  572 :  36 - 0x24
      10'h23D: dout <= 8'b00100100; //  573 :  36 - 0x24
      10'h23E: dout <= 8'b00100100; //  574 :  36 - 0x24
      10'h23F: dout <= 8'b00100100; //  575 :  36 - 0x24
      10'h240: dout <= 8'b00100100; //  576 :  36 - 0x24 -- line 0x12
      10'h241: dout <= 8'b00100100; //  577 :  36 - 0x24
      10'h242: dout <= 8'b00100100; //  578 :  36 - 0x24
      10'h243: dout <= 8'b00100100; //  579 :  36 - 0x24
      10'h244: dout <= 8'b00100100; //  580 :  36 - 0x24
      10'h245: dout <= 8'b00100100; //  581 :  36 - 0x24
      10'h246: dout <= 8'b00100100; //  582 :  36 - 0x24
      10'h247: dout <= 8'b00100100; //  583 :  36 - 0x24
      10'h248: dout <= 8'b00100100; //  584 :  36 - 0x24
      10'h249: dout <= 8'b00100100; //  585 :  36 - 0x24
      10'h24A: dout <= 8'b00111111; //  586 :  63 - 0x3f
      10'h24B: dout <= 8'b00100100; //  587 :  36 - 0x24
      10'h24C: dout <= 8'b00100100; //  588 :  36 - 0x24
      10'h24D: dout <= 8'b00100100; //  589 :  36 - 0x24
      10'h24E: dout <= 8'b00100100; //  590 :  36 - 0x24
      10'h24F: dout <= 8'b00100100; //  591 :  36 - 0x24
      10'h250: dout <= 8'b00111111; //  592 :  63 - 0x3f
      10'h251: dout <= 8'b00100100; //  593 :  36 - 0x24
      10'h252: dout <= 8'b00100100; //  594 :  36 - 0x24
      10'h253: dout <= 8'b00100100; //  595 :  36 - 0x24
      10'h254: dout <= 8'b00100100; //  596 :  36 - 0x24
      10'h255: dout <= 8'b00100100; //  597 :  36 - 0x24
      10'h256: dout <= 8'b00100100; //  598 :  36 - 0x24
      10'h257: dout <= 8'b00100100; //  599 :  36 - 0x24
      10'h258: dout <= 8'b00100100; //  600 :  36 - 0x24
      10'h259: dout <= 8'b01000000; //  601 :  64 - 0x40
      10'h25A: dout <= 8'b00111000; //  602 :  56 - 0x38
      10'h25B: dout <= 8'b00111000; //  603 :  56 - 0x38
      10'h25C: dout <= 8'b00111001; //  604 :  57 - 0x39
      10'h25D: dout <= 8'b00111001; //  605 :  57 - 0x39
      10'h25E: dout <= 8'b00100100; //  606 :  36 - 0x24
      10'h25F: dout <= 8'b00100100; //  607 :  36 - 0x24
      10'h260: dout <= 8'b00100100; //  608 :  36 - 0x24 -- line 0x13
      10'h261: dout <= 8'b00100100; //  609 :  36 - 0x24
      10'h262: dout <= 8'b00100100; //  610 :  36 - 0x24
      10'h263: dout <= 8'b00100100; //  611 :  36 - 0x24
      10'h264: dout <= 8'b00111001; //  612 :  57 - 0x39
      10'h265: dout <= 8'b00111001; //  613 :  57 - 0x39
      10'h266: dout <= 8'b00111001; //  614 :  57 - 0x39
      10'h267: dout <= 8'b00111010; //  615 :  58 - 0x3a
      10'h268: dout <= 8'b00111010; //  616 :  58 - 0x3a
      10'h269: dout <= 8'b00111010; //  617 :  58 - 0x3a
      10'h26A: dout <= 8'b01000010; //  618 :  66 - 0x42
      10'h26B: dout <= 8'b00111011; //  619 :  59 - 0x3b
      10'h26C: dout <= 8'b00111011; //  620 :  59 - 0x3b
      10'h26D: dout <= 8'b00111100; //  621 :  60 - 0x3c
      10'h26E: dout <= 8'b00111100; //  622 :  60 - 0x3c
      10'h26F: dout <= 8'b00111100; //  623 :  60 - 0x3c
      10'h270: dout <= 8'b01000100; //  624 :  68 - 0x44
      10'h271: dout <= 8'b00111101; //  625 :  61 - 0x3d
      10'h272: dout <= 8'b00111101; //  626 :  61 - 0x3d
      10'h273: dout <= 8'b00111110; //  627 :  62 - 0x3e
      10'h274: dout <= 8'b00111110; //  628 :  62 - 0x3e
      10'h275: dout <= 8'b00111110; //  629 :  62 - 0x3e
      10'h276: dout <= 8'b00110000; //  630 :  48 - 0x30
      10'h277: dout <= 8'b00110000; //  631 :  48 - 0x30
      10'h278: dout <= 8'b00110000; //  632 :  48 - 0x30
      10'h279: dout <= 8'b00110001; //  633 :  49 - 0x31
      10'h27A: dout <= 8'b00110001; //  634 :  49 - 0x31
      10'h27B: dout <= 8'b00110001; //  635 :  49 - 0x31
      10'h27C: dout <= 8'b00110010; //  636 :  50 - 0x32
      10'h27D: dout <= 8'b00110010; //  637 :  50 - 0x32
      10'h27E: dout <= 8'b00100100; //  638 :  36 - 0x24
      10'h27F: dout <= 8'b00100100; //  639 :  36 - 0x24
      10'h280: dout <= 8'b00100100; //  640 :  36 - 0x24 -- line 0x14
      10'h281: dout <= 8'b00100100; //  641 :  36 - 0x24
      10'h282: dout <= 8'b00100100; //  642 :  36 - 0x24
      10'h283: dout <= 8'b00100100; //  643 :  36 - 0x24
      10'h284: dout <= 8'b00110010; //  644 :  50 - 0x32
      10'h285: dout <= 8'b00110010; //  645 :  50 - 0x32
      10'h286: dout <= 8'b01000111; //  646 :  71 - 0x47
      10'h287: dout <= 8'b00110011; //  647 :  51 - 0x33
      10'h288: dout <= 8'b00110011; //  648 :  51 - 0x33
      10'h289: dout <= 8'b00110011; //  649 :  51 - 0x33
      10'h28A: dout <= 8'b00110100; //  650 :  52 - 0x34
      10'h28B: dout <= 8'b00110100; //  651 :  52 - 0x34
      10'h28C: dout <= 8'b00110100; //  652 :  52 - 0x34
      10'h28D: dout <= 8'b00110101; //  653 :  53 - 0x35
      10'h28E: dout <= 8'b01001010; //  654 :  74 - 0x4a
      10'h28F: dout <= 8'b00110101; //  655 :  53 - 0x35
      10'h290: dout <= 8'b00110110; //  656 :  54 - 0x36
      10'h291: dout <= 8'b00110110; //  657 :  54 - 0x36
      10'h292: dout <= 8'b00110110; //  658 :  54 - 0x36
      10'h293: dout <= 8'b00110111; //  659 :  55 - 0x37
      10'h294: dout <= 8'b00110111; //  660 :  55 - 0x37
      10'h295: dout <= 8'b00110111; //  661 :  55 - 0x37
      10'h296: dout <= 8'b00100100; //  662 :  36 - 0x24
      10'h297: dout <= 8'b00100100; //  663 :  36 - 0x24
      10'h298: dout <= 8'b00100100; //  664 :  36 - 0x24
      10'h299: dout <= 8'b00100100; //  665 :  36 - 0x24
      10'h29A: dout <= 8'b00100100; //  666 :  36 - 0x24
      10'h29B: dout <= 8'b00100100; //  667 :  36 - 0x24
      10'h29C: dout <= 8'b00100100; //  668 :  36 - 0x24
      10'h29D: dout <= 8'b00100100; //  669 :  36 - 0x24
      10'h29E: dout <= 8'b00100100; //  670 :  36 - 0x24
      10'h29F: dout <= 8'b00100100; //  671 :  36 - 0x24
      10'h2A0: dout <= 8'b00100100; //  672 :  36 - 0x24 -- line 0x15
      10'h2A1: dout <= 8'b00100100; //  673 :  36 - 0x24
      10'h2A2: dout <= 8'b00100100; //  674 :  36 - 0x24
      10'h2A3: dout <= 8'b00100100; //  675 :  36 - 0x24
      10'h2A4: dout <= 8'b00100100; //  676 :  36 - 0x24
      10'h2A5: dout <= 8'b00100100; //  677 :  36 - 0x24
      10'h2A6: dout <= 8'b00111111; //  678 :  63 - 0x3f
      10'h2A7: dout <= 8'b00100100; //  679 :  36 - 0x24
      10'h2A8: dout <= 8'b00100100; //  680 :  36 - 0x24
      10'h2A9: dout <= 8'b00100100; //  681 :  36 - 0x24
      10'h2AA: dout <= 8'b00100100; //  682 :  36 - 0x24
      10'h2AB: dout <= 8'b00100100; //  683 :  36 - 0x24
      10'h2AC: dout <= 8'b00100100; //  684 :  36 - 0x24
      10'h2AD: dout <= 8'b00100100; //  685 :  36 - 0x24
      10'h2AE: dout <= 8'b00111111; //  686 :  63 - 0x3f
      10'h2AF: dout <= 8'b00100100; //  687 :  36 - 0x24
      10'h2B0: dout <= 8'b00100100; //  688 :  36 - 0x24
      10'h2B1: dout <= 8'b00100100; //  689 :  36 - 0x24
      10'h2B2: dout <= 8'b00100100; //  690 :  36 - 0x24
      10'h2B3: dout <= 8'b00100100; //  691 :  36 - 0x24
      10'h2B4: dout <= 8'b00100100; //  692 :  36 - 0x24
      10'h2B5: dout <= 8'b00100100; //  693 :  36 - 0x24
      10'h2B6: dout <= 8'b00100100; //  694 :  36 - 0x24
      10'h2B7: dout <= 8'b00100100; //  695 :  36 - 0x24
      10'h2B8: dout <= 8'b00100100; //  696 :  36 - 0x24
      10'h2B9: dout <= 8'b00100100; //  697 :  36 - 0x24
      10'h2BA: dout <= 8'b00100100; //  698 :  36 - 0x24
      10'h2BB: dout <= 8'b00100100; //  699 :  36 - 0x24
      10'h2BC: dout <= 8'b00100100; //  700 :  36 - 0x24
      10'h2BD: dout <= 8'b00100100; //  701 :  36 - 0x24
      10'h2BE: dout <= 8'b00100100; //  702 :  36 - 0x24
      10'h2BF: dout <= 8'b00100100; //  703 :  36 - 0x24
      10'h2C0: dout <= 8'b00100100; //  704 :  36 - 0x24 -- line 0x16
      10'h2C1: dout <= 8'b00100100; //  705 :  36 - 0x24
      10'h2C2: dout <= 8'b00111011; //  706 :  59 - 0x3b
      10'h2C3: dout <= 8'b00111011; //  707 :  59 - 0x3b
      10'h2C4: dout <= 8'b00111010; //  708 :  58 - 0x3a
      10'h2C5: dout <= 8'b00111010; //  709 :  58 - 0x3a
      10'h2C6: dout <= 8'b01000001; //  710 :  65 - 0x41
      10'h2C7: dout <= 8'b00111001; //  711 :  57 - 0x39
      10'h2C8: dout <= 8'b00111001; //  712 :  57 - 0x39
      10'h2C9: dout <= 8'b00111001; //  713 :  57 - 0x39
      10'h2CA: dout <= 8'b00111000; //  714 :  56 - 0x38
      10'h2CB: dout <= 8'b00111000; //  715 :  56 - 0x38
      10'h2CC: dout <= 8'b00111000; //  716 :  56 - 0x38
      10'h2CD: dout <= 8'b00100100; //  717 :  36 - 0x24
      10'h2CE: dout <= 8'b00111111; //  718 :  63 - 0x3f
      10'h2CF: dout <= 8'b00100100; //  719 :  36 - 0x24
      10'h2D0: dout <= 8'b00100100; //  720 :  36 - 0x24
      10'h2D1: dout <= 8'b00100100; //  721 :  36 - 0x24
      10'h2D2: dout <= 8'b00100100; //  722 :  36 - 0x24
      10'h2D3: dout <= 8'b00100100; //  723 :  36 - 0x24
      10'h2D4: dout <= 8'b00100100; //  724 :  36 - 0x24
      10'h2D5: dout <= 8'b00100100; //  725 :  36 - 0x24
      10'h2D6: dout <= 8'b00100100; //  726 :  36 - 0x24
      10'h2D7: dout <= 8'b00100100; //  727 :  36 - 0x24
      10'h2D8: dout <= 8'b00100100; //  728 :  36 - 0x24
      10'h2D9: dout <= 8'b00100100; //  729 :  36 - 0x24
      10'h2DA: dout <= 8'b00100100; //  730 :  36 - 0x24
      10'h2DB: dout <= 8'b00100100; //  731 :  36 - 0x24
      10'h2DC: dout <= 8'b00100100; //  732 :  36 - 0x24
      10'h2DD: dout <= 8'b00100100; //  733 :  36 - 0x24
      10'h2DE: dout <= 8'b00100100; //  734 :  36 - 0x24
      10'h2DF: dout <= 8'b00100100; //  735 :  36 - 0x24
      10'h2E0: dout <= 8'b00100100; //  736 :  36 - 0x24 -- line 0x17
      10'h2E1: dout <= 8'b00100100; //  737 :  36 - 0x24
      10'h2E2: dout <= 8'b00110100; //  738 :  52 - 0x34
      10'h2E3: dout <= 8'b00110100; //  739 :  52 - 0x34
      10'h2E4: dout <= 8'b00110011; //  740 :  51 - 0x33
      10'h2E5: dout <= 8'b00110011; //  741 :  51 - 0x33
      10'h2E6: dout <= 8'b00110011; //  742 :  51 - 0x33
      10'h2E7: dout <= 8'b00110010; //  743 :  50 - 0x32
      10'h2E8: dout <= 8'b00110010; //  744 :  50 - 0x32
      10'h2E9: dout <= 8'b00110010; //  745 :  50 - 0x32
      10'h2EA: dout <= 8'b00110001; //  746 :  49 - 0x31
      10'h2EB: dout <= 8'b00110001; //  747 :  49 - 0x31
      10'h2EC: dout <= 8'b01000110; //  748 :  70 - 0x46
      10'h2ED: dout <= 8'b00110000; //  749 :  48 - 0x30
      10'h2EE: dout <= 8'b00110000; //  750 :  48 - 0x30
      10'h2EF: dout <= 8'b00110000; //  751 :  48 - 0x30
      10'h2F0: dout <= 8'b00111110; //  752 :  62 - 0x3e
      10'h2F1: dout <= 8'b00111110; //  753 :  62 - 0x3e
      10'h2F2: dout <= 8'b00111110; //  754 :  62 - 0x3e
      10'h2F3: dout <= 8'b00111101; //  755 :  61 - 0x3d
      10'h2F4: dout <= 8'b00111101; //  756 :  61 - 0x3d
      10'h2F5: dout <= 8'b00111101; //  757 :  61 - 0x3d
      10'h2F6: dout <= 8'b00111100; //  758 :  60 - 0x3c
      10'h2F7: dout <= 8'b00111100; //  759 :  60 - 0x3c
      10'h2F8: dout <= 8'b00111100; //  760 :  60 - 0x3c
      10'h2F9: dout <= 8'b00111011; //  761 :  59 - 0x3b
      10'h2FA: dout <= 8'b00111011; //  762 :  59 - 0x3b
      10'h2FB: dout <= 8'b00111011; //  763 :  59 - 0x3b
      10'h2FC: dout <= 8'b00100100; //  764 :  36 - 0x24
      10'h2FD: dout <= 8'b00100100; //  765 :  36 - 0x24
      10'h2FE: dout <= 8'b00100100; //  766 :  36 - 0x24
      10'h2FF: dout <= 8'b00100100; //  767 :  36 - 0x24
      10'h300: dout <= 8'b00100100; //  768 :  36 - 0x24 -- line 0x18
      10'h301: dout <= 8'b00100100; //  769 :  36 - 0x24
      10'h302: dout <= 8'b00100100; //  770 :  36 - 0x24
      10'h303: dout <= 8'b00100100; //  771 :  36 - 0x24
      10'h304: dout <= 8'b00100100; //  772 :  36 - 0x24
      10'h305: dout <= 8'b00100100; //  773 :  36 - 0x24
      10'h306: dout <= 8'b00100100; //  774 :  36 - 0x24
      10'h307: dout <= 8'b00100100; //  775 :  36 - 0x24
      10'h308: dout <= 8'b00100100; //  776 :  36 - 0x24
      10'h309: dout <= 8'b00100100; //  777 :  36 - 0x24
      10'h30A: dout <= 8'b00100100; //  778 :  36 - 0x24
      10'h30B: dout <= 8'b00100100; //  779 :  36 - 0x24
      10'h30C: dout <= 8'b00111111; //  780 :  63 - 0x3f
      10'h30D: dout <= 8'b00100100; //  781 :  36 - 0x24
      10'h30E: dout <= 8'b00100100; //  782 :  36 - 0x24
      10'h30F: dout <= 8'b00100100; //  783 :  36 - 0x24
      10'h310: dout <= 8'b00110111; //  784 :  55 - 0x37
      10'h311: dout <= 8'b00110111; //  785 :  55 - 0x37
      10'h312: dout <= 8'b00110111; //  786 :  55 - 0x37
      10'h313: dout <= 8'b00110110; //  787 :  54 - 0x36
      10'h314: dout <= 8'b00110110; //  788 :  54 - 0x36
      10'h315: dout <= 8'b00110110; //  789 :  54 - 0x36
      10'h316: dout <= 8'b00110101; //  790 :  53 - 0x35
      10'h317: dout <= 8'b00110101; //  791 :  53 - 0x35
      10'h318: dout <= 8'b00110101; //  792 :  53 - 0x35
      10'h319: dout <= 8'b01001001; //  793 :  73 - 0x49
      10'h31A: dout <= 8'b00110100; //  794 :  52 - 0x34
      10'h31B: dout <= 8'b00110100; //  795 :  52 - 0x34
      10'h31C: dout <= 8'b00100100; //  796 :  36 - 0x24
      10'h31D: dout <= 8'b00100100; //  797 :  36 - 0x24
      10'h31E: dout <= 8'b00100100; //  798 :  36 - 0x24
      10'h31F: dout <= 8'b00100100; //  799 :  36 - 0x24
      10'h320: dout <= 8'b00100100; //  800 :  36 - 0x24 -- line 0x19
      10'h321: dout <= 8'b00100100; //  801 :  36 - 0x24
      10'h322: dout <= 8'b00100100; //  802 :  36 - 0x24
      10'h323: dout <= 8'b00100100; //  803 :  36 - 0x24
      10'h324: dout <= 8'b01001100; //  804 :  76 - 0x4c
      10'h325: dout <= 8'b01001110; //  805 :  78 - 0x4e
      10'h326: dout <= 8'b00100100; //  806 :  36 - 0x24
      10'h327: dout <= 8'b00100100; //  807 :  36 - 0x24
      10'h328: dout <= 8'b00100100; //  808 :  36 - 0x24
      10'h329: dout <= 8'b00100100; //  809 :  36 - 0x24
      10'h32A: dout <= 8'b00100100; //  810 :  36 - 0x24
      10'h32B: dout <= 8'b00100100; //  811 :  36 - 0x24
      10'h32C: dout <= 8'b00100100; //  812 :  36 - 0x24
      10'h32D: dout <= 8'b00100100; //  813 :  36 - 0x24
      10'h32E: dout <= 8'b00100100; //  814 :  36 - 0x24
      10'h32F: dout <= 8'b00100100; //  815 :  36 - 0x24
      10'h330: dout <= 8'b00100100; //  816 :  36 - 0x24
      10'h331: dout <= 8'b00100100; //  817 :  36 - 0x24
      10'h332: dout <= 8'b00100100; //  818 :  36 - 0x24
      10'h333: dout <= 8'b00100100; //  819 :  36 - 0x24
      10'h334: dout <= 8'b00100100; //  820 :  36 - 0x24
      10'h335: dout <= 8'b00100100; //  821 :  36 - 0x24
      10'h336: dout <= 8'b00100100; //  822 :  36 - 0x24
      10'h337: dout <= 8'b00100100; //  823 :  36 - 0x24
      10'h338: dout <= 8'b00100100; //  824 :  36 - 0x24
      10'h339: dout <= 8'b00111111; //  825 :  63 - 0x3f
      10'h33A: dout <= 8'b00100100; //  826 :  36 - 0x24
      10'h33B: dout <= 8'b00100100; //  827 :  36 - 0x24
      10'h33C: dout <= 8'b00100100; //  828 :  36 - 0x24
      10'h33D: dout <= 8'b00100100; //  829 :  36 - 0x24
      10'h33E: dout <= 8'b00100100; //  830 :  36 - 0x24
      10'h33F: dout <= 8'b00100100; //  831 :  36 - 0x24
      10'h340: dout <= 8'b00100100; //  832 :  36 - 0x24 -- line 0x1a
      10'h341: dout <= 8'b00100100; //  833 :  36 - 0x24
      10'h342: dout <= 8'b00100100; //  834 :  36 - 0x24
      10'h343: dout <= 8'b00100100; //  835 :  36 - 0x24
      10'h344: dout <= 8'b01001101; //  836 :  77 - 0x4d
      10'h345: dout <= 8'b01001111; //  837 :  79 - 0x4f
      10'h346: dout <= 8'b00100100; //  838 :  36 - 0x24
      10'h347: dout <= 8'b00100100; //  839 :  36 - 0x24
      10'h348: dout <= 8'b00100100; //  840 :  36 - 0x24
      10'h349: dout <= 8'b00100100; //  841 :  36 - 0x24
      10'h34A: dout <= 8'b00100100; //  842 :  36 - 0x24
      10'h34B: dout <= 8'b00100100; //  843 :  36 - 0x24
      10'h34C: dout <= 8'b00111111; //  844 :  63 - 0x3f
      10'h34D: dout <= 8'b00100100; //  845 :  36 - 0x24
      10'h34E: dout <= 8'b00100100; //  846 :  36 - 0x24
      10'h34F: dout <= 8'b00100100; //  847 :  36 - 0x24
      10'h350: dout <= 8'b00111000; //  848 :  56 - 0x38
      10'h351: dout <= 8'b00111000; //  849 :  56 - 0x38
      10'h352: dout <= 8'b00111000; //  850 :  56 - 0x38
      10'h353: dout <= 8'b00111001; //  851 :  57 - 0x39
      10'h354: dout <= 8'b00111001; //  852 :  57 - 0x39
      10'h355: dout <= 8'b00111001; //  853 :  57 - 0x39
      10'h356: dout <= 8'b00111010; //  854 :  58 - 0x3a
      10'h357: dout <= 8'b00111010; //  855 :  58 - 0x3a
      10'h358: dout <= 8'b00111010; //  856 :  58 - 0x3a
      10'h359: dout <= 8'b01000010; //  857 :  66 - 0x42
      10'h35A: dout <= 8'b00111011; //  858 :  59 - 0x3b
      10'h35B: dout <= 8'b00111011; //  859 :  59 - 0x3b
      10'h35C: dout <= 8'b00111100; //  860 :  60 - 0x3c
      10'h35D: dout <= 8'b00111100; //  861 :  60 - 0x3c
      10'h35E: dout <= 8'b00111100; //  862 :  60 - 0x3c
      10'h35F: dout <= 8'b00100100; //  863 :  36 - 0x24
      10'h360: dout <= 8'b00100100; //  864 :  36 - 0x24 -- line 0x1b
      10'h361: dout <= 8'b00110000; //  865 :  48 - 0x30
      10'h362: dout <= 8'b00110000; //  866 :  48 - 0x30
      10'h363: dout <= 8'b00110000; //  867 :  48 - 0x30
      10'h364: dout <= 8'b00110000; //  868 :  48 - 0x30
      10'h365: dout <= 8'b00110000; //  869 :  48 - 0x30
      10'h366: dout <= 8'b00110000; //  870 :  48 - 0x30
      10'h367: dout <= 8'b00110000; //  871 :  48 - 0x30
      10'h368: dout <= 8'b00110000; //  872 :  48 - 0x30
      10'h369: dout <= 8'b00110000; //  873 :  48 - 0x30
      10'h36A: dout <= 8'b00110000; //  874 :  48 - 0x30
      10'h36B: dout <= 8'b00110000; //  875 :  48 - 0x30
      10'h36C: dout <= 8'b00110000; //  876 :  48 - 0x30
      10'h36D: dout <= 8'b00110000; //  877 :  48 - 0x30
      10'h36E: dout <= 8'b00110000; //  878 :  48 - 0x30
      10'h36F: dout <= 8'b00110000; //  879 :  48 - 0x30
      10'h370: dout <= 8'b00110001; //  880 :  49 - 0x31
      10'h371: dout <= 8'b00110001; //  881 :  49 - 0x31
      10'h372: dout <= 8'b00110001; //  882 :  49 - 0x31
      10'h373: dout <= 8'b00110010; //  883 :  50 - 0x32
      10'h374: dout <= 8'b00110010; //  884 :  50 - 0x32
      10'h375: dout <= 8'b00110010; //  885 :  50 - 0x32
      10'h376: dout <= 8'b00110011; //  886 :  51 - 0x33
      10'h377: dout <= 8'b00110011; //  887 :  51 - 0x33
      10'h378: dout <= 8'b00110011; //  888 :  51 - 0x33
      10'h379: dout <= 8'b00110100; //  889 :  52 - 0x34
      10'h37A: dout <= 8'b00110100; //  890 :  52 - 0x34
      10'h37B: dout <= 8'b00110100; //  891 :  52 - 0x34
      10'h37C: dout <= 8'b00110101; //  892 :  53 - 0x35
      10'h37D: dout <= 8'b00110101; //  893 :  53 - 0x35
      10'h37E: dout <= 8'b00110101; //  894 :  53 - 0x35
      10'h37F: dout <= 8'b00100100; //  895 :  36 - 0x24
      10'h380: dout <= 8'b00100100; //  896 :  36 - 0x24 -- line 0x1c
      10'h381: dout <= 8'b00100100; //  897 :  36 - 0x24
      10'h382: dout <= 8'b00100100; //  898 :  36 - 0x24
      10'h383: dout <= 8'b00100100; //  899 :  36 - 0x24
      10'h384: dout <= 8'b00100100; //  900 :  36 - 0x24
      10'h385: dout <= 8'b00100100; //  901 :  36 - 0x24
      10'h386: dout <= 8'b00100100; //  902 :  36 - 0x24
      10'h387: dout <= 8'b00100100; //  903 :  36 - 0x24
      10'h388: dout <= 8'b00100100; //  904 :  36 - 0x24
      10'h389: dout <= 8'b00100100; //  905 :  36 - 0x24
      10'h38A: dout <= 8'b00100100; //  906 :  36 - 0x24
      10'h38B: dout <= 8'b00100100; //  907 :  36 - 0x24
      10'h38C: dout <= 8'b00100100; //  908 :  36 - 0x24
      10'h38D: dout <= 8'b00100100; //  909 :  36 - 0x24
      10'h38E: dout <= 8'b00100100; //  910 :  36 - 0x24
      10'h38F: dout <= 8'b00100100; //  911 :  36 - 0x24
      10'h390: dout <= 8'b00100100; //  912 :  36 - 0x24
      10'h391: dout <= 8'b00100100; //  913 :  36 - 0x24
      10'h392: dout <= 8'b00100100; //  914 :  36 - 0x24
      10'h393: dout <= 8'b00100100; //  915 :  36 - 0x24
      10'h394: dout <= 8'b00100100; //  916 :  36 - 0x24
      10'h395: dout <= 8'b00100100; //  917 :  36 - 0x24
      10'h396: dout <= 8'b00100100; //  918 :  36 - 0x24
      10'h397: dout <= 8'b00100100; //  919 :  36 - 0x24
      10'h398: dout <= 8'b00100100; //  920 :  36 - 0x24
      10'h399: dout <= 8'b00100100; //  921 :  36 - 0x24
      10'h39A: dout <= 8'b00100100; //  922 :  36 - 0x24
      10'h39B: dout <= 8'b00100100; //  923 :  36 - 0x24
      10'h39C: dout <= 8'b00100100; //  924 :  36 - 0x24
      10'h39D: dout <= 8'b00100100; //  925 :  36 - 0x24
      10'h39E: dout <= 8'b00100100; //  926 :  36 - 0x24
      10'h39F: dout <= 8'b00100100; //  927 :  36 - 0x24
      10'h3A0: dout <= 8'b00100100; //  928 :  36 - 0x24 -- line 0x1d
      10'h3A1: dout <= 8'b00100100; //  929 :  36 - 0x24
      10'h3A2: dout <= 8'b00100100; //  930 :  36 - 0x24
      10'h3A3: dout <= 8'b00100100; //  931 :  36 - 0x24
      10'h3A4: dout <= 8'b00100100; //  932 :  36 - 0x24
      10'h3A5: dout <= 8'b00100100; //  933 :  36 - 0x24
      10'h3A6: dout <= 8'b00100100; //  934 :  36 - 0x24
      10'h3A7: dout <= 8'b00100100; //  935 :  36 - 0x24
      10'h3A8: dout <= 8'b00100100; //  936 :  36 - 0x24
      10'h3A9: dout <= 8'b00100100; //  937 :  36 - 0x24
      10'h3AA: dout <= 8'b00100100; //  938 :  36 - 0x24
      10'h3AB: dout <= 8'b00100100; //  939 :  36 - 0x24
      10'h3AC: dout <= 8'b00100100; //  940 :  36 - 0x24
      10'h3AD: dout <= 8'b00100100; //  941 :  36 - 0x24
      10'h3AE: dout <= 8'b00100100; //  942 :  36 - 0x24
      10'h3AF: dout <= 8'b00100100; //  943 :  36 - 0x24
      10'h3B0: dout <= 8'b00100100; //  944 :  36 - 0x24
      10'h3B1: dout <= 8'b00100100; //  945 :  36 - 0x24
      10'h3B2: dout <= 8'b00100100; //  946 :  36 - 0x24
      10'h3B3: dout <= 8'b00100100; //  947 :  36 - 0x24
      10'h3B4: dout <= 8'b00100100; //  948 :  36 - 0x24
      10'h3B5: dout <= 8'b00100100; //  949 :  36 - 0x24
      10'h3B6: dout <= 8'b00100100; //  950 :  36 - 0x24
      10'h3B7: dout <= 8'b00100100; //  951 :  36 - 0x24
      10'h3B8: dout <= 8'b00100100; //  952 :  36 - 0x24
      10'h3B9: dout <= 8'b00100100; //  953 :  36 - 0x24
      10'h3BA: dout <= 8'b00100100; //  954 :  36 - 0x24
      10'h3BB: dout <= 8'b00100100; //  955 :  36 - 0x24
      10'h3BC: dout <= 8'b00100100; //  956 :  36 - 0x24
      10'h3BD: dout <= 8'b00100100; //  957 :  36 - 0x24
      10'h3BE: dout <= 8'b00100100; //  958 :  36 - 0x24
      10'h3BF: dout <= 8'b00100100; //  959 :  36 - 0x24
        //-- Attribute Table 0----
      10'h3C0: dout <= 8'b11111111; //  960 : 255 - 0xff
      10'h3C1: dout <= 8'b11111111; //  961 : 255 - 0xff
      10'h3C2: dout <= 8'b11111111; //  962 : 255 - 0xff
      10'h3C3: dout <= 8'b11111111; //  963 : 255 - 0xff
      10'h3C4: dout <= 8'b11111111; //  964 : 255 - 0xff
      10'h3C5: dout <= 8'b11111111; //  965 : 255 - 0xff
      10'h3C6: dout <= 8'b11111111; //  966 : 255 - 0xff
      10'h3C7: dout <= 8'b11111111; //  967 : 255 - 0xff
      10'h3C8: dout <= 8'b01010101; //  968 :  85 - 0x55
      10'h3C9: dout <= 8'b10101010; //  969 : 170 - 0xaa
      10'h3CA: dout <= 8'b00100010; //  970 :  34 - 0x22
      10'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      10'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      10'h3CD: dout <= 8'b00001111; //  973 :  15 - 0xf
      10'h3CE: dout <= 8'b00001111; //  974 :  15 - 0xf
      10'h3CF: dout <= 8'b00001111; //  975 :  15 - 0xf
      10'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0
      10'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      10'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      10'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      10'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      10'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      10'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      10'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      10'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0
      10'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      10'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      10'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      10'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      10'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      10'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      10'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      10'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0
      10'h3E1: dout <= 8'b00000000; //  993 :   0 - 0x0
      10'h3E2: dout <= 8'b00000000; //  994 :   0 - 0x0
      10'h3E3: dout <= 8'b00000000; //  995 :   0 - 0x0
      10'h3E4: dout <= 8'b00000000; //  996 :   0 - 0x0
      10'h3E5: dout <= 8'b00000000; //  997 :   0 - 0x0
      10'h3E6: dout <= 8'b00000000; //  998 :   0 - 0x0
      10'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      10'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0
      10'h3E9: dout <= 8'b00000000; // 1001 :   0 - 0x0
      10'h3EA: dout <= 8'b00000000; // 1002 :   0 - 0x0
      10'h3EB: dout <= 8'b00000000; // 1003 :   0 - 0x0
      10'h3EC: dout <= 8'b00000000; // 1004 :   0 - 0x0
      10'h3ED: dout <= 8'b00000000; // 1005 :   0 - 0x0
      10'h3EE: dout <= 8'b00000000; // 1006 :   0 - 0x0
      10'h3EF: dout <= 8'b00000000; // 1007 :   0 - 0x0
      10'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0
      10'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      10'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      10'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      10'h3F4: dout <= 8'b00000000; // 1012 :   0 - 0x0
      10'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      10'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      10'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      10'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0
      10'h3F9: dout <= 8'b00000000; // 1017 :   0 - 0x0
      10'h3FA: dout <= 8'b00000000; // 1018 :   0 - 0x0
      10'h3FB: dout <= 8'b00000000; // 1019 :   0 - 0x0
      10'h3FC: dout <= 8'b00000000; // 1020 :   0 - 0x0
      10'h3FD: dout <= 8'b00000000; // 1021 :   0 - 0x0
      10'h3FE: dout <= 8'b00000000; // 1022 :   0 - 0x0
      10'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
    endcase
  end

endmodule
