---   Background Pattern table COLOR PLANE 1
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: smario_traspas_patron.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_MARIO_TRASPAS_BG_PLN1 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_MARIO_TRASPAS_BG_PLN1;

architecture BEHAVIORAL of ROM_PTABLE_MARIO_TRASPAS_BG_PLN1 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table COLOR PLANE 1
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Background 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Background 0x1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Background 0x2
    "00000000", --   17 - 0x11  :    0 - 0x0
    "00000000", --   18 - 0x12  :    0 - 0x0
    "00000000", --   19 - 0x13  :    0 - 0x0
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00000000", --   21 - 0x15  :    0 - 0x0
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- Background 0x3
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Background 0x4
    "00000000", --   33 - 0x21  :    0 - 0x0
    "00000000", --   34 - 0x22  :    0 - 0x0
    "00000000", --   35 - 0x23  :    0 - 0x0
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- Background 0x5
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Background 0x6
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00000000", --   51 - 0x33  :    0 - 0x0
    "00000000", --   52 - 0x34  :    0 - 0x0
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000000", --   54 - 0x36  :    0 - 0x0
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0 -- Background 0x7
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Background 0x8
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0 -- Background 0x9
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Background 0xa
    "00000000", --   81 - 0x51  :    0 - 0x0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00000000", --   88 - 0x58  :    0 - 0x0 -- Background 0xb
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Background 0xc
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0 -- Background 0xd
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Background 0xe
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0 -- Background 0xf
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Background 0x10
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0 -- Background 0x11
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Background 0x12
    "00000000", --  145 - 0x91  :    0 - 0x0
    "00000000", --  146 - 0x92  :    0 - 0x0
    "00000000", --  147 - 0x93  :    0 - 0x0
    "00000000", --  148 - 0x94  :    0 - 0x0
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- Background 0x13
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Background 0x14
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "00000000", --  164 - 0xa4  :    0 - 0x0
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0 -- Background 0x15
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Background 0x16
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0 -- Background 0x17
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Background 0x18
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "00000000", --  194 - 0xc2  :    0 - 0x0
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00000000", --  196 - 0xc4  :    0 - 0x0
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- Background 0x19
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Background 0x1a
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00000000", --  211 - 0xd3  :    0 - 0x0
    "00000000", --  212 - 0xd4  :    0 - 0x0
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Background 0x1b
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Background 0x1c
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00000000", --  228 - 0xe4  :    0 - 0x0
    "00000000", --  229 - 0xe5  :    0 - 0x0
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- Background 0x1d
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Background 0x1e
    "00000000", --  241 - 0xf1  :    0 - 0x0
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "00000000", --  243 - 0xf3  :    0 - 0x0
    "00000000", --  244 - 0xf4  :    0 - 0x0
    "00000000", --  245 - 0xf5  :    0 - 0x0
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- Background 0x1f
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Background 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Background 0x21
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00000000", --  272 - 0x110  :    0 - 0x0 -- Background 0x22
    "00000000", --  273 - 0x111  :    0 - 0x0
    "00000000", --  274 - 0x112  :    0 - 0x0
    "00000000", --  275 - 0x113  :    0 - 0x0
    "00000000", --  276 - 0x114  :    0 - 0x0
    "00000000", --  277 - 0x115  :    0 - 0x0
    "00000000", --  278 - 0x116  :    0 - 0x0
    "00000000", --  279 - 0x117  :    0 - 0x0
    "00000000", --  280 - 0x118  :    0 - 0x0 -- Background 0x23
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00000000", --  283 - 0x11b  :    0 - 0x0
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Background 0x24
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0 -- Background 0x25
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000000", --  298 - 0x12a  :    0 - 0x0
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "11111111", --  304 - 0x130  :  255 - 0xff -- Background 0x26
    "11111111", --  305 - 0x131  :  255 - 0xff
    "11111111", --  306 - 0x132  :  255 - 0xff
    "11111111", --  307 - 0x133  :  255 - 0xff
    "11111111", --  308 - 0x134  :  255 - 0xff
    "11111111", --  309 - 0x135  :  255 - 0xff
    "11111111", --  310 - 0x136  :  255 - 0xff
    "11111111", --  311 - 0x137  :  255 - 0xff
    "11111111", --  312 - 0x138  :  255 - 0xff -- Background 0x27
    "11111111", --  313 - 0x139  :  255 - 0xff
    "11111111", --  314 - 0x13a  :  255 - 0xff
    "11111111", --  315 - 0x13b  :  255 - 0xff
    "11111111", --  316 - 0x13c  :  255 - 0xff
    "11111111", --  317 - 0x13d  :  255 - 0xff
    "11111111", --  318 - 0x13e  :  255 - 0xff
    "11111111", --  319 - 0x13f  :  255 - 0xff
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Background 0x28
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "00000000", --  324 - 0x144  :    0 - 0x0
    "00000000", --  325 - 0x145  :    0 - 0x0
    "00000000", --  326 - 0x146  :    0 - 0x0
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00000000", --  328 - 0x148  :    0 - 0x0 -- Background 0x29
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000000", --  330 - 0x14a  :    0 - 0x0
    "00000000", --  331 - 0x14b  :    0 - 0x0
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "01111111", --  336 - 0x150  :  127 - 0x7f -- Background 0x2a
    "01111111", --  337 - 0x151  :  127 - 0x7f
    "01111111", --  338 - 0x152  :  127 - 0x7f
    "01111111", --  339 - 0x153  :  127 - 0x7f
    "01111111", --  340 - 0x154  :  127 - 0x7f
    "01111111", --  341 - 0x155  :  127 - 0x7f
    "01111111", --  342 - 0x156  :  127 - 0x7f
    "01111111", --  343 - 0x157  :  127 - 0x7f
    "00000000", --  344 - 0x158  :    0 - 0x0 -- Background 0x2b
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "11111111", --  352 - 0x160  :  255 - 0xff -- Background 0x2c
    "10000000", --  353 - 0x161  :  128 - 0x80
    "10000000", --  354 - 0x162  :  128 - 0x80
    "10000000", --  355 - 0x163  :  128 - 0x80
    "10000000", --  356 - 0x164  :  128 - 0x80
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00011100", --  358 - 0x166  :   28 - 0x1c
    "00111110", --  359 - 0x167  :   62 - 0x3e
    "01111111", --  360 - 0x168  :  127 - 0x7f -- Background 0x2d
    "01111111", --  361 - 0x169  :  127 - 0x7f
    "01111111", --  362 - 0x16a  :  127 - 0x7f
    "00111110", --  363 - 0x16b  :   62 - 0x3e
    "00011100", --  364 - 0x16c  :   28 - 0x1c
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "11111111", --  367 - 0x16f  :  255 - 0xff
    "00001000", --  368 - 0x170  :    8 - 0x8 -- Background 0x2e
    "00000100", --  369 - 0x171  :    4 - 0x4
    "00000100", --  370 - 0x172  :    4 - 0x4
    "00000100", --  371 - 0x173  :    4 - 0x4
    "00000100", --  372 - 0x174  :    4 - 0x4
    "00000100", --  373 - 0x175  :    4 - 0x4
    "00001000", --  374 - 0x176  :    8 - 0x8
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000011", --  376 - 0x178  :    3 - 0x3 -- Background 0x2f
    "00000101", --  377 - 0x179  :    5 - 0x5
    "00001011", --  378 - 0x17a  :   11 - 0xb
    "00001011", --  379 - 0x17b  :   11 - 0xb
    "00001111", --  380 - 0x17c  :   15 - 0xf
    "00001111", --  381 - 0x17d  :   15 - 0xf
    "00000111", --  382 - 0x17e  :    7 - 0x7
    "00000011", --  383 - 0x17f  :    3 - 0x3
    "00000001", --  384 - 0x180  :    1 - 0x1 -- Background 0x30
    "00000011", --  385 - 0x181  :    3 - 0x3
    "00000111", --  386 - 0x182  :    7 - 0x7
    "00001111", --  387 - 0x183  :   15 - 0xf
    "00011111", --  388 - 0x184  :   31 - 0x1f
    "00111111", --  389 - 0x185  :   63 - 0x3f
    "01111111", --  390 - 0x186  :  127 - 0x7f
    "11111111", --  391 - 0x187  :  255 - 0xff
    "00000000", --  392 - 0x188  :    0 - 0x0 -- Background 0x31
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000111", --  397 - 0x18d  :    7 - 0x7
    "00111111", --  398 - 0x18e  :   63 - 0x3f
    "11111111", --  399 - 0x18f  :  255 - 0xff
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Background 0x32
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000000", --  403 - 0x193  :    0 - 0x0
    "00000000", --  404 - 0x194  :    0 - 0x0
    "11100000", --  405 - 0x195  :  224 - 0xe0
    "11111100", --  406 - 0x196  :  252 - 0xfc
    "11111111", --  407 - 0x197  :  255 - 0xff
    "10000000", --  408 - 0x198  :  128 - 0x80 -- Background 0x33
    "11000000", --  409 - 0x199  :  192 - 0xc0
    "11100000", --  410 - 0x19a  :  224 - 0xe0
    "11110000", --  411 - 0x19b  :  240 - 0xf0
    "11111000", --  412 - 0x19c  :  248 - 0xf8
    "11111100", --  413 - 0x19d  :  252 - 0xfc
    "11111110", --  414 - 0x19e  :  254 - 0xfe
    "11111111", --  415 - 0x19f  :  255 - 0xff
    "11111111", --  416 - 0x1a0  :  255 - 0xff -- Background 0x34
    "11111111", --  417 - 0x1a1  :  255 - 0xff
    "11111111", --  418 - 0x1a2  :  255 - 0xff
    "11111111", --  419 - 0x1a3  :  255 - 0xff
    "11111111", --  420 - 0x1a4  :  255 - 0xff
    "11111111", --  421 - 0x1a5  :  255 - 0xff
    "11111111", --  422 - 0x1a6  :  255 - 0xff
    "11111111", --  423 - 0x1a7  :  255 - 0xff
    "00000111", --  424 - 0x1a8  :    7 - 0x7 -- Background 0x35
    "00001000", --  425 - 0x1a9  :    8 - 0x8
    "00010000", --  426 - 0x1aa  :   16 - 0x10
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "01100000", --  428 - 0x1ac  :   96 - 0x60
    "10000000", --  429 - 0x1ad  :  128 - 0x80
    "10000000", --  430 - 0x1ae  :  128 - 0x80
    "01000000", --  431 - 0x1af  :   64 - 0x40
    "00000011", --  432 - 0x1b0  :    3 - 0x3 -- Background 0x36
    "00000100", --  433 - 0x1b1  :    4 - 0x4
    "00011000", --  434 - 0x1b2  :   24 - 0x18
    "00100000", --  435 - 0x1b3  :   32 - 0x20
    "00100000", --  436 - 0x1b4  :   32 - 0x20
    "00100000", --  437 - 0x1b5  :   32 - 0x20
    "01000110", --  438 - 0x1b6  :   70 - 0x46
    "10001000", --  439 - 0x1b7  :  136 - 0x88
    "11000000", --  440 - 0x1b8  :  192 - 0xc0 -- Background 0x37
    "00100000", --  441 - 0x1b9  :   32 - 0x20
    "00010000", --  442 - 0x1ba  :   16 - 0x10
    "00010100", --  443 - 0x1bb  :   20 - 0x14
    "00001010", --  444 - 0x1bc  :   10 - 0xa
    "01000001", --  445 - 0x1bd  :   65 - 0x41
    "00100001", --  446 - 0x1be  :   33 - 0x21
    "00000001", --  447 - 0x1bf  :    1 - 0x1
    "10010000", --  448 - 0x1c0  :  144 - 0x90 -- Background 0x38
    "10101000", --  449 - 0x1c1  :  168 - 0xa8
    "01001000", --  450 - 0x1c2  :   72 - 0x48
    "00001010", --  451 - 0x1c3  :   10 - 0xa
    "00000101", --  452 - 0x1c4  :    5 - 0x5
    "00000001", --  453 - 0x1c5  :    1 - 0x1
    "00000001", --  454 - 0x1c6  :    1 - 0x1
    "00000010", --  455 - 0x1c7  :    2 - 0x2
    "00100100", --  456 - 0x1c8  :   36 - 0x24 -- Background 0x39
    "00010010", --  457 - 0x1c9  :   18 - 0x12
    "00001001", --  458 - 0x1ca  :    9 - 0x9
    "00001000", --  459 - 0x1cb  :    8 - 0x8
    "00000111", --  460 - 0x1cc  :    7 - 0x7
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Background 0x3a
    "01000000", --  465 - 0x1d1  :   64 - 0x40
    "11100011", --  466 - 0x1d2  :  227 - 0xe3
    "00111111", --  467 - 0x1d3  :   63 - 0x3f
    "00001100", --  468 - 0x1d4  :   12 - 0xc
    "10000001", --  469 - 0x1d5  :  129 - 0x81
    "01100010", --  470 - 0x1d6  :   98 - 0x62
    "00011100", --  471 - 0x1d7  :   28 - 0x1c
    "01000000", --  472 - 0x1d8  :   64 - 0x40 -- Background 0x3b
    "10000000", --  473 - 0x1d9  :  128 - 0x80
    "11000010", --  474 - 0x1da  :  194 - 0xc2
    "01111100", --  475 - 0x1db  :  124 - 0x7c
    "00111000", --  476 - 0x1dc  :   56 - 0x38
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "11000011", --  478 - 0x1de  :  195 - 0xc3
    "00111100", --  479 - 0x1df  :   60 - 0x3c
    "00000100", --  480 - 0x1e0  :    4 - 0x4 -- Background 0x3c
    "00000010", --  481 - 0x1e1  :    2 - 0x2
    "00000001", --  482 - 0x1e2  :    1 - 0x1
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000110", --  484 - 0x1e4  :    6 - 0x6
    "10011000", --  485 - 0x1e5  :  152 - 0x98
    "01100000", --  486 - 0x1e6  :   96 - 0x60
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "11000000", --  488 - 0x1e8  :  192 - 0xc0 -- Background 0x3d
    "11100000", --  489 - 0x1e9  :  224 - 0xe0
    "11110000", --  490 - 0x1ea  :  240 - 0xf0
    "11110000", --  491 - 0x1eb  :  240 - 0xf0
    "11110000", --  492 - 0x1ec  :  240 - 0xf0
    "11110000", --  493 - 0x1ed  :  240 - 0xf0
    "11100000", --  494 - 0x1ee  :  224 - 0xe0
    "11000000", --  495 - 0x1ef  :  192 - 0xc0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Background 0x3e
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00000000", --  500 - 0x1f4  :    0 - 0x0
    "00000000", --  501 - 0x1f5  :    0 - 0x0
    "00011100", --  502 - 0x1f6  :   28 - 0x1c
    "00111110", --  503 - 0x1f7  :   62 - 0x3e
    "01111111", --  504 - 0x1f8  :  127 - 0x7f -- Background 0x3f
    "01111111", --  505 - 0x1f9  :  127 - 0x7f
    "01111111", --  506 - 0x1fa  :  127 - 0x7f
    "00111110", --  507 - 0x1fb  :   62 - 0x3e
    "00011100", --  508 - 0x1fc  :   28 - 0x1c
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "11111111", --  512 - 0x200  :  255 - 0xff -- Background 0x40
    "11111111", --  513 - 0x201  :  255 - 0xff
    "11111111", --  514 - 0x202  :  255 - 0xff
    "11111111", --  515 - 0x203  :  255 - 0xff
    "11111111", --  516 - 0x204  :  255 - 0xff
    "11111111", --  517 - 0x205  :  255 - 0xff
    "11111111", --  518 - 0x206  :  255 - 0xff
    "11111111", --  519 - 0x207  :  255 - 0xff
    "00000000", --  520 - 0x208  :    0 - 0x0 -- Background 0x41
    "00001000", --  521 - 0x209  :    8 - 0x8
    "00011000", --  522 - 0x20a  :   24 - 0x18
    "00111000", --  523 - 0x20b  :   56 - 0x38
    "11111100", --  524 - 0x20c  :  252 - 0xfc
    "10111111", --  525 - 0x20d  :  191 - 0xbf
    "01011110", --  526 - 0x20e  :   94 - 0x5e
    "11011001", --  527 - 0x20f  :  217 - 0xd9
    "10000001", --  528 - 0x210  :  129 - 0x81 -- Background 0x42
    "10000001", --  529 - 0x211  :  129 - 0x81
    "10000001", --  530 - 0x212  :  129 - 0x81
    "10000001", --  531 - 0x213  :  129 - 0x81
    "10000001", --  532 - 0x214  :  129 - 0x81
    "10000001", --  533 - 0x215  :  129 - 0x81
    "10000001", --  534 - 0x216  :  129 - 0x81
    "10000001", --  535 - 0x217  :  129 - 0x81
    "00000001", --  536 - 0x218  :    1 - 0x1 -- Background 0x43
    "00000001", --  537 - 0x219  :    1 - 0x1
    "00000001", --  538 - 0x21a  :    1 - 0x1
    "00000001", --  539 - 0x21b  :    1 - 0x1
    "00000001", --  540 - 0x21c  :    1 - 0x1
    "00000001", --  541 - 0x21d  :    1 - 0x1
    "00000001", --  542 - 0x21e  :    1 - 0x1
    "00000001", --  543 - 0x21f  :    1 - 0x1
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Background 0x44
    "01111111", --  545 - 0x221  :  127 - 0x7f
    "01111111", --  546 - 0x222  :  127 - 0x7f
    "01100111", --  547 - 0x223  :  103 - 0x67
    "01100111", --  548 - 0x224  :  103 - 0x67
    "01111111", --  549 - 0x225  :  127 - 0x7f
    "01111111", --  550 - 0x226  :  127 - 0x7f
    "01111111", --  551 - 0x227  :  127 - 0x7f
    "00000000", --  552 - 0x228  :    0 - 0x0 -- Background 0x45
    "11111111", --  553 - 0x229  :  255 - 0xff
    "11111111", --  554 - 0x22a  :  255 - 0xff
    "11111111", --  555 - 0x22b  :  255 - 0xff
    "11111111", --  556 - 0x22c  :  255 - 0xff
    "11111111", --  557 - 0x22d  :  255 - 0xff
    "11111111", --  558 - 0x22e  :  255 - 0xff
    "11111111", --  559 - 0x22f  :  255 - 0xff
    "01111111", --  560 - 0x230  :  127 - 0x7f -- Background 0x46
    "01111111", --  561 - 0x231  :  127 - 0x7f
    "01111111", --  562 - 0x232  :  127 - 0x7f
    "01111111", --  563 - 0x233  :  127 - 0x7f
    "01111111", --  564 - 0x234  :  127 - 0x7f
    "01111111", --  565 - 0x235  :  127 - 0x7f
    "01111111", --  566 - 0x236  :  127 - 0x7f
    "01111111", --  567 - 0x237  :  127 - 0x7f
    "11111111", --  568 - 0x238  :  255 - 0xff -- Background 0x47
    "11111111", --  569 - 0x239  :  255 - 0xff
    "11111111", --  570 - 0x23a  :  255 - 0xff
    "11111111", --  571 - 0x23b  :  255 - 0xff
    "11111111", --  572 - 0x23c  :  255 - 0xff
    "11111111", --  573 - 0x23d  :  255 - 0xff
    "11111111", --  574 - 0x23e  :  255 - 0xff
    "11111111", --  575 - 0x23f  :  255 - 0xff
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Background 0x48
    "11111111", --  577 - 0x241  :  255 - 0xff
    "11111111", --  578 - 0x242  :  255 - 0xff
    "11111111", --  579 - 0x243  :  255 - 0xff
    "11111111", --  580 - 0x244  :  255 - 0xff
    "11111111", --  581 - 0x245  :  255 - 0xff
    "11111111", --  582 - 0x246  :  255 - 0xff
    "11111111", --  583 - 0x247  :  255 - 0xff
    "00000000", --  584 - 0x248  :    0 - 0x0 -- Background 0x49
    "11111111", --  585 - 0x249  :  255 - 0xff
    "11111111", --  586 - 0x24a  :  255 - 0xff
    "11100111", --  587 - 0x24b  :  231 - 0xe7
    "11100111", --  588 - 0x24c  :  231 - 0xe7
    "11111111", --  589 - 0x24d  :  255 - 0xff
    "11111111", --  590 - 0x24e  :  255 - 0xff
    "11111111", --  591 - 0x24f  :  255 - 0xff
    "11111111", --  592 - 0x250  :  255 - 0xff -- Background 0x4a
    "11111111", --  593 - 0x251  :  255 - 0xff
    "11111111", --  594 - 0x252  :  255 - 0xff
    "11111111", --  595 - 0x253  :  255 - 0xff
    "11111111", --  596 - 0x254  :  255 - 0xff
    "11111111", --  597 - 0x255  :  255 - 0xff
    "11111111", --  598 - 0x256  :  255 - 0xff
    "11111111", --  599 - 0x257  :  255 - 0xff
    "00111111", --  600 - 0x258  :   63 - 0x3f -- Background 0x4b
    "01100000", --  601 - 0x259  :   96 - 0x60
    "01000000", --  602 - 0x25a  :   64 - 0x40
    "11000000", --  603 - 0x25b  :  192 - 0xc0
    "10000000", --  604 - 0x25c  :  128 - 0x80
    "10000000", --  605 - 0x25d  :  128 - 0x80
    "10000000", --  606 - 0x25e  :  128 - 0x80
    "10000000", --  607 - 0x25f  :  128 - 0x80
    "10000000", --  608 - 0x260  :  128 - 0x80 -- Background 0x4c
    "10000000", --  609 - 0x261  :  128 - 0x80
    "10000000", --  610 - 0x262  :  128 - 0x80
    "10000000", --  611 - 0x263  :  128 - 0x80
    "10000000", --  612 - 0x264  :  128 - 0x80
    "10000001", --  613 - 0x265  :  129 - 0x81
    "01000010", --  614 - 0x266  :   66 - 0x42
    "00111100", --  615 - 0x267  :   60 - 0x3c
    "11111111", --  616 - 0x268  :  255 - 0xff -- Background 0x4d
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Background 0x4e
    "00000000", --  625 - 0x271  :    0 - 0x0
    "00000000", --  626 - 0x272  :    0 - 0x0
    "00000000", --  627 - 0x273  :    0 - 0x0
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000001", --  629 - 0x275  :    1 - 0x1
    "10000010", --  630 - 0x276  :  130 - 0x82
    "01111100", --  631 - 0x277  :  124 - 0x7c
    "00000000", --  632 - 0x278  :    0 - 0x0 -- Background 0x4f
    "00000000", --  633 - 0x279  :    0 - 0x0
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "00000000", --  635 - 0x27b  :    0 - 0x0
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000001", --  637 - 0x27d  :    1 - 0x1
    "10000011", --  638 - 0x27e  :  131 - 0x83
    "11111111", --  639 - 0x27f  :  255 - 0xff
    "11111000", --  640 - 0x280  :  248 - 0xf8 -- Background 0x50
    "00000100", --  641 - 0x281  :    4 - 0x4
    "00000010", --  642 - 0x282  :    2 - 0x2
    "00000010", --  643 - 0x283  :    2 - 0x2
    "00000001", --  644 - 0x284  :    1 - 0x1
    "00000001", --  645 - 0x285  :    1 - 0x1
    "00000001", --  646 - 0x286  :    1 - 0x1
    "00000001", --  647 - 0x287  :    1 - 0x1
    "00000001", --  648 - 0x288  :    1 - 0x1 -- Background 0x51
    "00000001", --  649 - 0x289  :    1 - 0x1
    "00000001", --  650 - 0x28a  :    1 - 0x1
    "00000001", --  651 - 0x28b  :    1 - 0x1
    "00000001", --  652 - 0x28c  :    1 - 0x1
    "10000001", --  653 - 0x28d  :  129 - 0x81
    "01000010", --  654 - 0x28e  :   66 - 0x42
    "00111100", --  655 - 0x28f  :   60 - 0x3c
    "11111111", --  656 - 0x290  :  255 - 0xff -- Background 0x52
    "11111111", --  657 - 0x291  :  255 - 0xff
    "11111111", --  658 - 0x292  :  255 - 0xff
    "11111111", --  659 - 0x293  :  255 - 0xff
    "11111111", --  660 - 0x294  :  255 - 0xff
    "11111111", --  661 - 0x295  :  255 - 0xff
    "11111111", --  662 - 0x296  :  255 - 0xff
    "11111111", --  663 - 0x297  :  255 - 0xff
    "01111111", --  664 - 0x298  :  127 - 0x7f -- Background 0x53
    "10000000", --  665 - 0x299  :  128 - 0x80
    "10100000", --  666 - 0x29a  :  160 - 0xa0
    "10000111", --  667 - 0x29b  :  135 - 0x87
    "10001111", --  668 - 0x29c  :  143 - 0x8f
    "10001110", --  669 - 0x29d  :  142 - 0x8e
    "10001110", --  670 - 0x29e  :  142 - 0x8e
    "10000110", --  671 - 0x29f  :  134 - 0x86
    "11111110", --  672 - 0x2a0  :  254 - 0xfe -- Background 0x54
    "00000001", --  673 - 0x2a1  :    1 - 0x1
    "00000101", --  674 - 0x2a2  :    5 - 0x5
    "11000001", --  675 - 0x2a3  :  193 - 0xc1
    "11100001", --  676 - 0x2a4  :  225 - 0xe1
    "01110001", --  677 - 0x2a5  :  113 - 0x71
    "01110001", --  678 - 0x2a6  :  113 - 0x71
    "11110001", --  679 - 0x2a7  :  241 - 0xf1
    "10000001", --  680 - 0x2a8  :  129 - 0x81 -- Background 0x55
    "10000001", --  681 - 0x2a9  :  129 - 0x81
    "10000000", --  682 - 0x2aa  :  128 - 0x80
    "10000001", --  683 - 0x2ab  :  129 - 0x81
    "10000001", --  684 - 0x2ac  :  129 - 0x81
    "10100000", --  685 - 0x2ad  :  160 - 0xa0
    "10000000", --  686 - 0x2ae  :  128 - 0x80
    "11111111", --  687 - 0x2af  :  255 - 0xff
    "11110001", --  688 - 0x2b0  :  241 - 0xf1 -- Background 0x56
    "11000001", --  689 - 0x2b1  :  193 - 0xc1
    "11000001", --  690 - 0x2b2  :  193 - 0xc1
    "10000001", --  691 - 0x2b3  :  129 - 0x81
    "11000001", --  692 - 0x2b4  :  193 - 0xc1
    "11000101", --  693 - 0x2b5  :  197 - 0xc5
    "00000001", --  694 - 0x2b6  :    1 - 0x1
    "11111111", --  695 - 0x2b7  :  255 - 0xff
    "01111111", --  696 - 0x2b8  :  127 - 0x7f -- Background 0x57
    "11111111", --  697 - 0x2b9  :  255 - 0xff
    "11111111", --  698 - 0x2ba  :  255 - 0xff
    "11111111", --  699 - 0x2bb  :  255 - 0xff
    "11111111", --  700 - 0x2bc  :  255 - 0xff
    "11111111", --  701 - 0x2bd  :  255 - 0xff
    "11111111", --  702 - 0x2be  :  255 - 0xff
    "11111111", --  703 - 0x2bf  :  255 - 0xff
    "11111110", --  704 - 0x2c0  :  254 - 0xfe -- Background 0x58
    "11111111", --  705 - 0x2c1  :  255 - 0xff
    "11111111", --  706 - 0x2c2  :  255 - 0xff
    "11111111", --  707 - 0x2c3  :  255 - 0xff
    "11111111", --  708 - 0x2c4  :  255 - 0xff
    "11111111", --  709 - 0x2c5  :  255 - 0xff
    "11111111", --  710 - 0x2c6  :  255 - 0xff
    "11111111", --  711 - 0x2c7  :  255 - 0xff
    "11111111", --  712 - 0x2c8  :  255 - 0xff -- Background 0x59
    "11111111", --  713 - 0x2c9  :  255 - 0xff
    "11111111", --  714 - 0x2ca  :  255 - 0xff
    "11111111", --  715 - 0x2cb  :  255 - 0xff
    "11111111", --  716 - 0x2cc  :  255 - 0xff
    "11111111", --  717 - 0x2cd  :  255 - 0xff
    "11111111", --  718 - 0x2ce  :  255 - 0xff
    "01111111", --  719 - 0x2cf  :  127 - 0x7f
    "11111111", --  720 - 0x2d0  :  255 - 0xff -- Background 0x5a
    "11111111", --  721 - 0x2d1  :  255 - 0xff
    "11111111", --  722 - 0x2d2  :  255 - 0xff
    "11111111", --  723 - 0x2d3  :  255 - 0xff
    "11111111", --  724 - 0x2d4  :  255 - 0xff
    "11111111", --  725 - 0x2d5  :  255 - 0xff
    "11111111", --  726 - 0x2d6  :  255 - 0xff
    "11111110", --  727 - 0x2d7  :  254 - 0xfe
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Background 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00111000", --  734 - 0x2de  :   56 - 0x38
    "01111100", --  735 - 0x2df  :  124 - 0x7c
    "11111110", --  736 - 0x2e0  :  254 - 0xfe -- Background 0x5c
    "11111110", --  737 - 0x2e1  :  254 - 0xfe
    "11111110", --  738 - 0x2e2  :  254 - 0xfe
    "01111100", --  739 - 0x2e3  :  124 - 0x7c
    "00111000", --  740 - 0x2e4  :   56 - 0x38
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00100000", --  744 - 0x2e8  :   32 - 0x20 -- Background 0x5d
    "11100111", --  745 - 0x2e9  :  231 - 0xe7
    "11100111", --  746 - 0x2ea  :  231 - 0xe7
    "11100111", --  747 - 0x2eb  :  231 - 0xe7
    "11100111", --  748 - 0x2ec  :  231 - 0xe7
    "11100111", --  749 - 0x2ed  :  231 - 0xe7
    "11101111", --  750 - 0x2ee  :  239 - 0xef
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000010", --  752 - 0x2f0  :    2 - 0x2 -- Background 0x5e
    "01111110", --  753 - 0x2f1  :  126 - 0x7e
    "01111110", --  754 - 0x2f2  :  126 - 0x7e
    "01111110", --  755 - 0x2f3  :  126 - 0x7e
    "01111110", --  756 - 0x2f4  :  126 - 0x7e
    "01111110", --  757 - 0x2f5  :  126 - 0x7e
    "11111110", --  758 - 0x2f6  :  254 - 0xfe
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "01111111", --  760 - 0x2f8  :  127 - 0x7f -- Background 0x5f
    "01111111", --  761 - 0x2f9  :  127 - 0x7f
    "01111111", --  762 - 0x2fa  :  127 - 0x7f
    "01100111", --  763 - 0x2fb  :  103 - 0x67
    "01100111", --  764 - 0x2fc  :  103 - 0x67
    "01111111", --  765 - 0x2fd  :  127 - 0x7f
    "01111111", --  766 - 0x2fe  :  127 - 0x7f
    "01111111", --  767 - 0x2ff  :  127 - 0x7f
    "11111111", --  768 - 0x300  :  255 - 0xff -- Background 0x60
    "10000000", --  769 - 0x301  :  128 - 0x80
    "11111100", --  770 - 0x302  :  252 - 0xfc
    "10001100", --  771 - 0x303  :  140 - 0x8c
    "10001100", --  772 - 0x304  :  140 - 0x8c
    "10001100", --  773 - 0x305  :  140 - 0x8c
    "10001100", --  774 - 0x306  :  140 - 0x8c
    "10001100", --  775 - 0x307  :  140 - 0x8c
    "11111111", --  776 - 0x308  :  255 - 0xff -- Background 0x61
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00001111", --  778 - 0x30a  :   15 - 0xf
    "00001001", --  779 - 0x30b  :    9 - 0x9
    "00001001", --  780 - 0x30c  :    9 - 0x9
    "00001001", --  781 - 0x30d  :    9 - 0x9
    "00001001", --  782 - 0x30e  :    9 - 0x9
    "00001001", --  783 - 0x30f  :    9 - 0x9
    "11111111", --  784 - 0x310  :  255 - 0xff -- Background 0x62
    "00000000", --  785 - 0x311  :    0 - 0x0
    "11111111", --  786 - 0x312  :  255 - 0xff
    "11111111", --  787 - 0x313  :  255 - 0xff
    "11111111", --  788 - 0x314  :  255 - 0xff
    "11111111", --  789 - 0x315  :  255 - 0xff
    "11111111", --  790 - 0x316  :  255 - 0xff
    "11111111", --  791 - 0x317  :  255 - 0xff
    "11111111", --  792 - 0x318  :  255 - 0xff -- Background 0x63
    "00000001", --  793 - 0x319  :    1 - 0x1
    "11111111", --  794 - 0x31a  :  255 - 0xff
    "10101001", --  795 - 0x31b  :  169 - 0xa9
    "11010001", --  796 - 0x31c  :  209 - 0xd1
    "10101001", --  797 - 0x31d  :  169 - 0xa9
    "11010001", --  798 - 0x31e  :  209 - 0xd1
    "10101001", --  799 - 0x31f  :  169 - 0xa9
    "10001100", --  800 - 0x320  :  140 - 0x8c -- Background 0x64
    "10001100", --  801 - 0x321  :  140 - 0x8c
    "10001100", --  802 - 0x322  :  140 - 0x8c
    "10001100", --  803 - 0x323  :  140 - 0x8c
    "10001100", --  804 - 0x324  :  140 - 0x8c
    "10001100", --  805 - 0x325  :  140 - 0x8c
    "11111111", --  806 - 0x326  :  255 - 0xff
    "00111111", --  807 - 0x327  :   63 - 0x3f
    "00001001", --  808 - 0x328  :    9 - 0x9 -- Background 0x65
    "00001001", --  809 - 0x329  :    9 - 0x9
    "00001001", --  810 - 0x32a  :    9 - 0x9
    "00001001", --  811 - 0x32b  :    9 - 0x9
    "00001001", --  812 - 0x32c  :    9 - 0x9
    "00001001", --  813 - 0x32d  :    9 - 0x9
    "11111111", --  814 - 0x32e  :  255 - 0xff
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "11111111", --  816 - 0x330  :  255 - 0xff -- Background 0x66
    "11111111", --  817 - 0x331  :  255 - 0xff
    "11111111", --  818 - 0x332  :  255 - 0xff
    "11111111", --  819 - 0x333  :  255 - 0xff
    "11111111", --  820 - 0x334  :  255 - 0xff
    "11111111", --  821 - 0x335  :  255 - 0xff
    "11111111", --  822 - 0x336  :  255 - 0xff
    "11111111", --  823 - 0x337  :  255 - 0xff
    "11010001", --  824 - 0x338  :  209 - 0xd1 -- Background 0x67
    "10101001", --  825 - 0x339  :  169 - 0xa9
    "11010001", --  826 - 0x33a  :  209 - 0xd1
    "10101001", --  827 - 0x33b  :  169 - 0xa9
    "11010001", --  828 - 0x33c  :  209 - 0xd1
    "10101001", --  829 - 0x33d  :  169 - 0xa9
    "11111111", --  830 - 0x33e  :  255 - 0xff
    "11111100", --  831 - 0x33f  :  252 - 0xfc
    "00100011", --  832 - 0x340  :   35 - 0x23 -- Background 0x68
    "00100011", --  833 - 0x341  :   35 - 0x23
    "00100011", --  834 - 0x342  :   35 - 0x23
    "00100011", --  835 - 0x343  :   35 - 0x23
    "00100011", --  836 - 0x344  :   35 - 0x23
    "00100011", --  837 - 0x345  :   35 - 0x23
    "00100011", --  838 - 0x346  :   35 - 0x23
    "00100011", --  839 - 0x347  :   35 - 0x23
    "00000100", --  840 - 0x348  :    4 - 0x4 -- Background 0x69
    "00000100", --  841 - 0x349  :    4 - 0x4
    "00000100", --  842 - 0x34a  :    4 - 0x4
    "00000100", --  843 - 0x34b  :    4 - 0x4
    "00000100", --  844 - 0x34c  :    4 - 0x4
    "00000100", --  845 - 0x34d  :    4 - 0x4
    "00000100", --  846 - 0x34e  :    4 - 0x4
    "00000100", --  847 - 0x34f  :    4 - 0x4
    "01000100", --  848 - 0x350  :   68 - 0x44 -- Background 0x6a
    "10100100", --  849 - 0x351  :  164 - 0xa4
    "01000100", --  850 - 0x352  :   68 - 0x44
    "10100100", --  851 - 0x353  :  164 - 0xa4
    "01000100", --  852 - 0x354  :   68 - 0x44
    "10100100", --  853 - 0x355  :  164 - 0xa4
    "01000100", --  854 - 0x356  :   68 - 0x44
    "10100100", --  855 - 0x357  :  164 - 0xa4
    "00011111", --  856 - 0x358  :   31 - 0x1f -- Background 0x6b
    "00111111", --  857 - 0x359  :   63 - 0x3f
    "01111111", --  858 - 0x35a  :  127 - 0x7f
    "01111111", --  859 - 0x35b  :  127 - 0x7f
    "11111111", --  860 - 0x35c  :  255 - 0xff
    "11111111", --  861 - 0x35d  :  255 - 0xff
    "11111111", --  862 - 0x35e  :  255 - 0xff
    "11111110", --  863 - 0x35f  :  254 - 0xfe
    "11111111", --  864 - 0x360  :  255 - 0xff -- Background 0x6c
    "01111111", --  865 - 0x361  :  127 - 0x7f
    "01111111", --  866 - 0x362  :  127 - 0x7f
    "00111111", --  867 - 0x363  :   63 - 0x3f
    "00000000", --  868 - 0x364  :    0 - 0x0
    "00000000", --  869 - 0x365  :    0 - 0x0
    "00000001", --  870 - 0x366  :    1 - 0x1
    "00000001", --  871 - 0x367  :    1 - 0x1
    "11111111", --  872 - 0x368  :  255 - 0xff -- Background 0x6d
    "10000000", --  873 - 0x369  :  128 - 0x80
    "10000000", --  874 - 0x36a  :  128 - 0x80
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "11111000", --  877 - 0x36d  :  248 - 0xf8
    "11111100", --  878 - 0x36e  :  252 - 0xfc
    "11111100", --  879 - 0x36f  :  252 - 0xfc
    "11111111", --  880 - 0x370  :  255 - 0xff -- Background 0x6e
    "11111111", --  881 - 0x371  :  255 - 0xff
    "11111111", --  882 - 0x372  :  255 - 0xff
    "11111111", --  883 - 0x373  :  255 - 0xff
    "11111111", --  884 - 0x374  :  255 - 0xff
    "01111110", --  885 - 0x375  :  126 - 0x7e
    "00111100", --  886 - 0x376  :   60 - 0x3c
    "00000000", --  887 - 0x377  :    0 - 0x0
    "11111000", --  888 - 0x378  :  248 - 0xf8 -- Background 0x6f
    "00000100", --  889 - 0x379  :    4 - 0x4
    "00000010", --  890 - 0x37a  :    2 - 0x2
    "00000010", --  891 - 0x37b  :    2 - 0x2
    "00011101", --  892 - 0x37c  :   29 - 0x1d
    "00111111", --  893 - 0x37d  :   63 - 0x3f
    "01111111", --  894 - 0x37e  :  127 - 0x7f
    "01111111", --  895 - 0x37f  :  127 - 0x7f
    "11111100", --  896 - 0x380  :  252 - 0xfc -- Background 0x70
    "10000000", --  897 - 0x381  :  128 - 0x80
    "10000000", --  898 - 0x382  :  128 - 0x80
    "10000000", --  899 - 0x383  :  128 - 0x80
    "10000000", --  900 - 0x384  :  128 - 0x80
    "10000000", --  901 - 0x385  :  128 - 0x80
    "01100000", --  902 - 0x386  :   96 - 0x60
    "00011111", --  903 - 0x387  :   31 - 0x1f
    "00000011", --  904 - 0x388  :    3 - 0x3 -- Background 0x71
    "00000011", --  905 - 0x389  :    3 - 0x3
    "00000011", --  906 - 0x38a  :    3 - 0x3
    "00000011", --  907 - 0x38b  :    3 - 0x3
    "00000001", --  908 - 0x38c  :    1 - 0x1
    "00000001", --  909 - 0x38d  :    1 - 0x1
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "11111111", --  911 - 0x38f  :  255 - 0xff
    "11111110", --  912 - 0x390  :  254 - 0xfe -- Background 0x72
    "11111110", --  913 - 0x391  :  254 - 0xfe
    "11111110", --  914 - 0x392  :  254 - 0xfe
    "11111110", --  915 - 0x393  :  254 - 0xfe
    "11111100", --  916 - 0x394  :  252 - 0xfc
    "11111100", --  917 - 0x395  :  252 - 0xfc
    "11111000", --  918 - 0x396  :  248 - 0xf8
    "11111111", --  919 - 0x397  :  255 - 0xff
    "00000000", --  920 - 0x398  :    0 - 0x0 -- Background 0x73
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "11111111", --  927 - 0x39f  :  255 - 0xff
    "01111111", --  928 - 0x3a0  :  127 - 0x7f -- Background 0x74
    "00111111", --  929 - 0x3a1  :   63 - 0x3f
    "00011101", --  930 - 0x3a2  :   29 - 0x1d
    "00000001", --  931 - 0x3a3  :    1 - 0x1
    "00000001", --  932 - 0x3a4  :    1 - 0x1
    "00000001", --  933 - 0x3a5  :    1 - 0x1
    "00000011", --  934 - 0x3a6  :    3 - 0x3
    "11111110", --  935 - 0x3a7  :  254 - 0xfe
    "10000000", --  936 - 0x3a8  :  128 - 0x80 -- Background 0x75
    "10000000", --  937 - 0x3a9  :  128 - 0x80
    "10000000", --  938 - 0x3aa  :  128 - 0x80
    "10000000", --  939 - 0x3ab  :  128 - 0x80
    "10000000", --  940 - 0x3ac  :  128 - 0x80
    "10000100", --  941 - 0x3ad  :  132 - 0x84
    "11001010", --  942 - 0x3ae  :  202 - 0xca
    "10110001", --  943 - 0x3af  :  177 - 0xb1
    "00000001", --  944 - 0x3b0  :    1 - 0x1 -- Background 0x76
    "00000001", --  945 - 0x3b1  :    1 - 0x1
    "00000001", --  946 - 0x3b2  :    1 - 0x1
    "00000001", --  947 - 0x3b3  :    1 - 0x1
    "00000001", --  948 - 0x3b4  :    1 - 0x1
    "00100001", --  949 - 0x3b5  :   33 - 0x21
    "01010011", --  950 - 0x3b6  :   83 - 0x53
    "10001101", --  951 - 0x3b7  :  141 - 0x8d
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- Background 0x77
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "01110111", --  956 - 0x3bc  :  119 - 0x77
    "11111111", --  957 - 0x3bd  :  255 - 0xff
    "11111111", --  958 - 0x3be  :  255 - 0xff
    "11111111", --  959 - 0x3bf  :  255 - 0xff
    "11111111", --  960 - 0x3c0  :  255 - 0xff -- Background 0x78
    "11111111", --  961 - 0x3c1  :  255 - 0xff
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "11111111", --  963 - 0x3c3  :  255 - 0xff
    "11111111", --  964 - 0x3c4  :  255 - 0xff
    "11111111", --  965 - 0x3c5  :  255 - 0xff
    "11111111", --  966 - 0x3c6  :  255 - 0xff
    "11111111", --  967 - 0x3c7  :  255 - 0xff
    "11111111", --  968 - 0x3c8  :  255 - 0xff -- Background 0x79
    "11111111", --  969 - 0x3c9  :  255 - 0xff
    "11111111", --  970 - 0x3ca  :  255 - 0xff
    "01110111", --  971 - 0x3cb  :  119 - 0x77
    "01110111", --  972 - 0x3cc  :  119 - 0x77
    "01110111", --  973 - 0x3cd  :  119 - 0x77
    "01110111", --  974 - 0x3ce  :  119 - 0x77
    "01110111", --  975 - 0x3cf  :  119 - 0x77
    "11111111", --  976 - 0x3d0  :  255 - 0xff -- Background 0x7a
    "11111111", --  977 - 0x3d1  :  255 - 0xff
    "11111111", --  978 - 0x3d2  :  255 - 0xff
    "11100111", --  979 - 0x3d3  :  231 - 0xe7
    "11100111", --  980 - 0x3d4  :  231 - 0xe7
    "11111111", --  981 - 0x3d5  :  255 - 0xff
    "11111111", --  982 - 0x3d6  :  255 - 0xff
    "11111110", --  983 - 0x3d7  :  254 - 0xfe
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Background 0x7b
    "00100001", --  985 - 0x3d9  :   33 - 0x21
    "00100001", --  986 - 0x3da  :   33 - 0x21
    "01000001", --  987 - 0x3db  :   65 - 0x41
    "01000001", --  988 - 0x3dc  :   65 - 0x41
    "01000001", --  989 - 0x3dd  :   65 - 0x41
    "01000001", --  990 - 0x3de  :   65 - 0x41
    "01000001", --  991 - 0x3df  :   65 - 0x41
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Background 0x7c
    "10000000", --  993 - 0x3e1  :  128 - 0x80
    "10000000", --  994 - 0x3e2  :  128 - 0x80
    "10000000", --  995 - 0x3e3  :  128 - 0x80
    "10000000", --  996 - 0x3e4  :  128 - 0x80
    "10000000", --  997 - 0x3e5  :  128 - 0x80
    "10000000", --  998 - 0x3e6  :  128 - 0x80
    "10000000", --  999 - 0x3e7  :  128 - 0x80
    "00100001", -- 1000 - 0x3e8  :   33 - 0x21 -- Background 0x7d
    "00100001", -- 1001 - 0x3e9  :   33 - 0x21
    "00000001", -- 1002 - 0x3ea  :    1 - 0x1
    "00000001", -- 1003 - 0x3eb  :    1 - 0x1
    "00000001", -- 1004 - 0x3ec  :    1 - 0x1
    "00000001", -- 1005 - 0x3ed  :    1 - 0x1
    "00000001", -- 1006 - 0x3ee  :    1 - 0x1
    "00000001", -- 1007 - 0x3ef  :    1 - 0x1
    "10000000", -- 1008 - 0x3f0  :  128 - 0x80 -- Background 0x7e
    "10000000", -- 1009 - 0x3f1  :  128 - 0x80
    "10000000", -- 1010 - 0x3f2  :  128 - 0x80
    "10000000", -- 1011 - 0x3f3  :  128 - 0x80
    "10000000", -- 1012 - 0x3f4  :  128 - 0x80
    "10000000", -- 1013 - 0x3f5  :  128 - 0x80
    "10000000", -- 1014 - 0x3f6  :  128 - 0x80
    "10000000", -- 1015 - 0x3f7  :  128 - 0x80
    "00000001", -- 1016 - 0x3f8  :    1 - 0x1 -- Background 0x7f
    "00000001", -- 1017 - 0x3f9  :    1 - 0x1
    "00000110", -- 1018 - 0x3fa  :    6 - 0x6
    "00001000", -- 1019 - 0x3fb  :    8 - 0x8
    "00011000", -- 1020 - 0x3fc  :   24 - 0x18
    "00100000", -- 1021 - 0x3fd  :   32 - 0x20
    "00100000", -- 1022 - 0x3fe  :   32 - 0x20
    "11000000", -- 1023 - 0x3ff  :  192 - 0xc0
    "00000100", -- 1024 - 0x400  :    4 - 0x4 -- Background 0x80
    "00000100", -- 1025 - 0x401  :    4 - 0x4
    "11000100", -- 1026 - 0x402  :  196 - 0xc4
    "11110100", -- 1027 - 0x403  :  244 - 0xf4
    "11110100", -- 1028 - 0x404  :  244 - 0xf4
    "00000100", -- 1029 - 0x405  :    4 - 0x4
    "00000100", -- 1030 - 0x406  :    4 - 0x4
    "00000101", -- 1031 - 0x407  :    5 - 0x5
    "01110000", -- 1032 - 0x408  :  112 - 0x70 -- Background 0x81
    "11110000", -- 1033 - 0x409  :  240 - 0xf0
    "11110000", -- 1034 - 0x40a  :  240 - 0xf0
    "11111111", -- 1035 - 0x40b  :  255 - 0xff
    "11111111", -- 1036 - 0x40c  :  255 - 0xff
    "11110000", -- 1037 - 0x40d  :  240 - 0xf0
    "11110000", -- 1038 - 0x40e  :  240 - 0xf0
    "01110000", -- 1039 - 0x40f  :  112 - 0x70
    "11000000", -- 1040 - 0x410  :  192 - 0xc0 -- Background 0x82
    "10000111", -- 1041 - 0x411  :  135 - 0x87
    "00011000", -- 1042 - 0x412  :   24 - 0x18
    "10110000", -- 1043 - 0x413  :  176 - 0xb0
    "11100111", -- 1044 - 0x414  :  231 - 0xe7
    "11100111", -- 1045 - 0x415  :  231 - 0xe7
    "11101111", -- 1046 - 0x416  :  239 - 0xef
    "11101111", -- 1047 - 0x417  :  239 - 0xef
    "01101111", -- 1048 - 0x418  :  111 - 0x6f -- Background 0x83
    "01000011", -- 1049 - 0x419  :   67 - 0x43
    "01011101", -- 1050 - 0x41a  :   93 - 0x5d
    "00111111", -- 1051 - 0x41b  :   63 - 0x3f
    "00111111", -- 1052 - 0x41c  :   63 - 0x3f
    "01111111", -- 1053 - 0x41d  :  127 - 0x7f
    "01111111", -- 1054 - 0x41e  :  127 - 0x7f
    "11111111", -- 1055 - 0x41f  :  255 - 0xff
    "00000011", -- 1056 - 0x420  :    3 - 0x3 -- Background 0x84
    "11111111", -- 1057 - 0x421  :  255 - 0xff
    "11110001", -- 1058 - 0x422  :  241 - 0xf1
    "01101110", -- 1059 - 0x423  :  110 - 0x6e
    "11001111", -- 1060 - 0x424  :  207 - 0xcf
    "11011111", -- 1061 - 0x425  :  223 - 0xdf
    "11111111", -- 1062 - 0x426  :  255 - 0xff
    "11111111", -- 1063 - 0x427  :  255 - 0xff
    "11111101", -- 1064 - 0x428  :  253 - 0xfd -- Background 0x85
    "11111011", -- 1065 - 0x429  :  251 - 0xfb
    "11111011", -- 1066 - 0x42a  :  251 - 0xfb
    "11110111", -- 1067 - 0x42b  :  247 - 0xf7
    "11110111", -- 1068 - 0x42c  :  247 - 0xf7
    "00001111", -- 1069 - 0x42d  :   15 - 0xf
    "01111111", -- 1070 - 0x42e  :  127 - 0x7f
    "11111111", -- 1071 - 0x42f  :  255 - 0xff
    "11111111", -- 1072 - 0x430  :  255 - 0xff -- Background 0x86
    "10000000", -- 1073 - 0x431  :  128 - 0x80
    "10000000", -- 1074 - 0x432  :  128 - 0x80
    "10000000", -- 1075 - 0x433  :  128 - 0x80
    "10000000", -- 1076 - 0x434  :  128 - 0x80
    "11111111", -- 1077 - 0x435  :  255 - 0xff
    "11111111", -- 1078 - 0x436  :  255 - 0xff
    "10000000", -- 1079 - 0x437  :  128 - 0x80
    "11111110", -- 1080 - 0x438  :  254 - 0xfe -- Background 0x87
    "00000011", -- 1081 - 0x439  :    3 - 0x3
    "00000011", -- 1082 - 0x43a  :    3 - 0x3
    "00000011", -- 1083 - 0x43b  :    3 - 0x3
    "00000011", -- 1084 - 0x43c  :    3 - 0x3
    "11111111", -- 1085 - 0x43d  :  255 - 0xff
    "11111111", -- 1086 - 0x43e  :  255 - 0xff
    "00000011", -- 1087 - 0x43f  :    3 - 0x3
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Background 0x88
    "11111111", -- 1089 - 0x441  :  255 - 0xff
    "00000000", -- 1090 - 0x442  :    0 - 0x0
    "00000000", -- 1091 - 0x443  :    0 - 0x0
    "00000000", -- 1092 - 0x444  :    0 - 0x0
    "00000000", -- 1093 - 0x445  :    0 - 0x0
    "11111111", -- 1094 - 0x446  :  255 - 0xff
    "11111111", -- 1095 - 0x447  :  255 - 0xff
    "00100011", -- 1096 - 0x448  :   35 - 0x23 -- Background 0x89
    "11110011", -- 1097 - 0x449  :  243 - 0xf3
    "00001011", -- 1098 - 0x44a  :   11 - 0xb
    "00001011", -- 1099 - 0x44b  :   11 - 0xb
    "00001011", -- 1100 - 0x44c  :   11 - 0xb
    "00000111", -- 1101 - 0x44d  :    7 - 0x7
    "11111111", -- 1102 - 0x44e  :  255 - 0xff
    "11111111", -- 1103 - 0x44f  :  255 - 0xff
    "10000000", -- 1104 - 0x450  :  128 - 0x80 -- Background 0x8a
    "10000000", -- 1105 - 0x451  :  128 - 0x80
    "10000000", -- 1106 - 0x452  :  128 - 0x80
    "10000000", -- 1107 - 0x453  :  128 - 0x80
    "11111111", -- 1108 - 0x454  :  255 - 0xff
    "10000000", -- 1109 - 0x455  :  128 - 0x80
    "10000000", -- 1110 - 0x456  :  128 - 0x80
    "10000000", -- 1111 - 0x457  :  128 - 0x80
    "00000011", -- 1112 - 0x458  :    3 - 0x3 -- Background 0x8b
    "00000011", -- 1113 - 0x459  :    3 - 0x3
    "00000011", -- 1114 - 0x45a  :    3 - 0x3
    "00000011", -- 1115 - 0x45b  :    3 - 0x3
    "11111111", -- 1116 - 0x45c  :  255 - 0xff
    "00000011", -- 1117 - 0x45d  :    3 - 0x3
    "00000011", -- 1118 - 0x45e  :    3 - 0x3
    "00000011", -- 1119 - 0x45f  :    3 - 0x3
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Background 0x8c
    "00000000", -- 1121 - 0x461  :    0 - 0x0
    "00000000", -- 1122 - 0x462  :    0 - 0x0
    "00000000", -- 1123 - 0x463  :    0 - 0x0
    "00000000", -- 1124 - 0x464  :    0 - 0x0
    "11111111", -- 1125 - 0x465  :  255 - 0xff
    "00000000", -- 1126 - 0x466  :    0 - 0x0
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000111", -- 1128 - 0x468  :    7 - 0x7 -- Background 0x8d
    "00000111", -- 1129 - 0x469  :    7 - 0x7
    "00000011", -- 1130 - 0x46a  :    3 - 0x3
    "00000011", -- 1131 - 0x46b  :    3 - 0x3
    "00000011", -- 1132 - 0x46c  :    3 - 0x3
    "11111111", -- 1133 - 0x46d  :  255 - 0xff
    "00000011", -- 1134 - 0x46e  :    3 - 0x3
    "00000011", -- 1135 - 0x46f  :    3 - 0x3
    "10000000", -- 1136 - 0x470  :  128 - 0x80 -- Background 0x8e
    "11111111", -- 1137 - 0x471  :  255 - 0xff
    "11111111", -- 1138 - 0x472  :  255 - 0xff
    "11111111", -- 1139 - 0x473  :  255 - 0xff
    "11111111", -- 1140 - 0x474  :  255 - 0xff
    "11111111", -- 1141 - 0x475  :  255 - 0xff
    "11111111", -- 1142 - 0x476  :  255 - 0xff
    "11111111", -- 1143 - 0x477  :  255 - 0xff
    "00000011", -- 1144 - 0x478  :    3 - 0x3 -- Background 0x8f
    "11111111", -- 1145 - 0x479  :  255 - 0xff
    "11111111", -- 1146 - 0x47a  :  255 - 0xff
    "11111111", -- 1147 - 0x47b  :  255 - 0xff
    "11111111", -- 1148 - 0x47c  :  255 - 0xff
    "11111111", -- 1149 - 0x47d  :  255 - 0xff
    "11111111", -- 1150 - 0x47e  :  255 - 0xff
    "11111111", -- 1151 - 0x47f  :  255 - 0xff
    "11111111", -- 1152 - 0x480  :  255 - 0xff -- Background 0x90
    "11111111", -- 1153 - 0x481  :  255 - 0xff
    "11111111", -- 1154 - 0x482  :  255 - 0xff
    "11111111", -- 1155 - 0x483  :  255 - 0xff
    "11111111", -- 1156 - 0x484  :  255 - 0xff
    "11111111", -- 1157 - 0x485  :  255 - 0xff
    "11111111", -- 1158 - 0x486  :  255 - 0xff
    "11111111", -- 1159 - 0x487  :  255 - 0xff
    "11111111", -- 1160 - 0x488  :  255 - 0xff -- Background 0x91
    "11111111", -- 1161 - 0x489  :  255 - 0xff
    "11010101", -- 1162 - 0x48a  :  213 - 0xd5
    "10101010", -- 1163 - 0x48b  :  170 - 0xaa
    "11010101", -- 1164 - 0x48c  :  213 - 0xd5
    "10000000", -- 1165 - 0x48d  :  128 - 0x80
    "10000000", -- 1166 - 0x48e  :  128 - 0x80
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "11111111", -- 1168 - 0x490  :  255 - 0xff -- Background 0x92
    "11111111", -- 1169 - 0x491  :  255 - 0xff
    "01010111", -- 1170 - 0x492  :   87 - 0x57
    "10101011", -- 1171 - 0x493  :  171 - 0xab
    "01010111", -- 1172 - 0x494  :   87 - 0x57
    "00000011", -- 1173 - 0x495  :    3 - 0x3
    "00000011", -- 1174 - 0x496  :    3 - 0x3
    "11111110", -- 1175 - 0x497  :  254 - 0xfe
    "11111111", -- 1176 - 0x498  :  255 - 0xff -- Background 0x93
    "10101010", -- 1177 - 0x499  :  170 - 0xaa
    "01010101", -- 1178 - 0x49a  :   85 - 0x55
    "10101010", -- 1179 - 0x49b  :  170 - 0xaa
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "11111111", -- 1182 - 0x49e  :  255 - 0xff
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "11111111", -- 1184 - 0x4a0  :  255 - 0xff -- Background 0x94
    "10101111", -- 1185 - 0x4a1  :  175 - 0xaf
    "01010111", -- 1186 - 0x4a2  :   87 - 0x57
    "10101011", -- 1187 - 0x4a3  :  171 - 0xab
    "00001011", -- 1188 - 0x4a4  :   11 - 0xb
    "00001011", -- 1189 - 0x4a5  :   11 - 0xb
    "11110011", -- 1190 - 0x4a6  :  243 - 0xf3
    "00100011", -- 1191 - 0x4a7  :   35 - 0x23
    "11111111", -- 1192 - 0x4a8  :  255 - 0xff -- Background 0x95
    "11111111", -- 1193 - 0x4a9  :  255 - 0xff
    "11111111", -- 1194 - 0x4aa  :  255 - 0xff
    "11111111", -- 1195 - 0x4ab  :  255 - 0xff
    "11111111", -- 1196 - 0x4ac  :  255 - 0xff
    "11111111", -- 1197 - 0x4ad  :  255 - 0xff
    "11111111", -- 1198 - 0x4ae  :  255 - 0xff
    "11111111", -- 1199 - 0x4af  :  255 - 0xff
    "11111111", -- 1200 - 0x4b0  :  255 - 0xff -- Background 0x96
    "11111111", -- 1201 - 0x4b1  :  255 - 0xff
    "11111111", -- 1202 - 0x4b2  :  255 - 0xff
    "11111111", -- 1203 - 0x4b3  :  255 - 0xff
    "11111111", -- 1204 - 0x4b4  :  255 - 0xff
    "11111111", -- 1205 - 0x4b5  :  255 - 0xff
    "11111111", -- 1206 - 0x4b6  :  255 - 0xff
    "11111111", -- 1207 - 0x4b7  :  255 - 0xff
    "11111111", -- 1208 - 0x4b8  :  255 - 0xff -- Background 0x97
    "11111111", -- 1209 - 0x4b9  :  255 - 0xff
    "11111111", -- 1210 - 0x4ba  :  255 - 0xff
    "11111111", -- 1211 - 0x4bb  :  255 - 0xff
    "11111111", -- 1212 - 0x4bc  :  255 - 0xff
    "11111111", -- 1213 - 0x4bd  :  255 - 0xff
    "11111111", -- 1214 - 0x4be  :  255 - 0xff
    "11111111", -- 1215 - 0x4bf  :  255 - 0xff
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Background 0x98
    "11111111", -- 1217 - 0x4c1  :  255 - 0xff
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111111", -- 1219 - 0x4c3  :  255 - 0xff
    "11111111", -- 1220 - 0x4c4  :  255 - 0xff
    "11111111", -- 1221 - 0x4c5  :  255 - 0xff
    "11111111", -- 1222 - 0x4c6  :  255 - 0xff
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0 -- Background 0x99
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "00000000", -- 1228 - 0x4cc  :    0 - 0x0
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Background 0x9a
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00000000", -- 1235 - 0x4d3  :    0 - 0x0
    "00000000", -- 1236 - 0x4d4  :    0 - 0x0
    "00000000", -- 1237 - 0x4d5  :    0 - 0x0
    "00000000", -- 1238 - 0x4d6  :    0 - 0x0
    "00000000", -- 1239 - 0x4d7  :    0 - 0x0
    "11111111", -- 1240 - 0x4d8  :  255 - 0xff -- Background 0x9b
    "11111111", -- 1241 - 0x4d9  :  255 - 0xff
    "11111111", -- 1242 - 0x4da  :  255 - 0xff
    "11111111", -- 1243 - 0x4db  :  255 - 0xff
    "11111111", -- 1244 - 0x4dc  :  255 - 0xff
    "11111111", -- 1245 - 0x4dd  :  255 - 0xff
    "11111111", -- 1246 - 0x4de  :  255 - 0xff
    "11111111", -- 1247 - 0x4df  :  255 - 0xff
    "11111111", -- 1248 - 0x4e0  :  255 - 0xff -- Background 0x9c
    "11111111", -- 1249 - 0x4e1  :  255 - 0xff
    "11111111", -- 1250 - 0x4e2  :  255 - 0xff
    "11111111", -- 1251 - 0x4e3  :  255 - 0xff
    "11111111", -- 1252 - 0x4e4  :  255 - 0xff
    "11111111", -- 1253 - 0x4e5  :  255 - 0xff
    "11111111", -- 1254 - 0x4e6  :  255 - 0xff
    "11111111", -- 1255 - 0x4e7  :  255 - 0xff
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0 -- Background 0x9d
    "11100000", -- 1257 - 0x4e9  :  224 - 0xe0
    "11100000", -- 1258 - 0x4ea  :  224 - 0xe0
    "11100000", -- 1259 - 0x4eb  :  224 - 0xe0
    "11100000", -- 1260 - 0x4ec  :  224 - 0xe0
    "11100000", -- 1261 - 0x4ed  :  224 - 0xe0
    "11100000", -- 1262 - 0x4ee  :  224 - 0xe0
    "11100000", -- 1263 - 0x4ef  :  224 - 0xe0
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0 -- Background 0x9e
    "00001111", -- 1265 - 0x4f1  :   15 - 0xf
    "00001111", -- 1266 - 0x4f2  :   15 - 0xf
    "00001111", -- 1267 - 0x4f3  :   15 - 0xf
    "00001111", -- 1268 - 0x4f4  :   15 - 0xf
    "00001111", -- 1269 - 0x4f5  :   15 - 0xf
    "00001111", -- 1270 - 0x4f6  :   15 - 0xf
    "00001111", -- 1271 - 0x4f7  :   15 - 0xf
    "01001000", -- 1272 - 0x4f8  :   72 - 0x48 -- Background 0x9f
    "01001000", -- 1273 - 0x4f9  :   72 - 0x48
    "01101100", -- 1274 - 0x4fa  :  108 - 0x6c
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "11111110", -- 1278 - 0x4fe  :  254 - 0xfe
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000101", -- 1280 - 0x500  :    5 - 0x5 -- Background 0xa0
    "00000101", -- 1281 - 0x501  :    5 - 0x5
    "11000101", -- 1282 - 0x502  :  197 - 0xc5
    "11110101", -- 1283 - 0x503  :  245 - 0xf5
    "11110100", -- 1284 - 0x504  :  244 - 0xf4
    "00000100", -- 1285 - 0x505  :    4 - 0x4
    "00000100", -- 1286 - 0x506  :    4 - 0x4
    "00000100", -- 1287 - 0x507  :    4 - 0x4
    "01110000", -- 1288 - 0x508  :  112 - 0x70 -- Background 0xa1
    "01110000", -- 1289 - 0x509  :  112 - 0x70
    "01110000", -- 1290 - 0x50a  :  112 - 0x70
    "01111111", -- 1291 - 0x50b  :  127 - 0x7f
    "01111111", -- 1292 - 0x50c  :  127 - 0x7f
    "01110000", -- 1293 - 0x50d  :  112 - 0x70
    "01110000", -- 1294 - 0x50e  :  112 - 0x70
    "01110000", -- 1295 - 0x50f  :  112 - 0x70
    "00000000", -- 1296 - 0x510  :    0 - 0x0 -- Background 0xa2
    "00000000", -- 1297 - 0x511  :    0 - 0x0
    "00000000", -- 1298 - 0x512  :    0 - 0x0
    "00000000", -- 1299 - 0x513  :    0 - 0x0
    "00000000", -- 1300 - 0x514  :    0 - 0x0
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "00000000", -- 1302 - 0x516  :    0 - 0x0
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "00000000", -- 1304 - 0x518  :    0 - 0x0 -- Background 0xa3
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "00000000", -- 1306 - 0x51a  :    0 - 0x0
    "00000000", -- 1307 - 0x51b  :    0 - 0x0
    "00000000", -- 1308 - 0x51c  :    0 - 0x0
    "00000000", -- 1309 - 0x51d  :    0 - 0x0
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "11111111", -- 1312 - 0x520  :  255 - 0xff -- Background 0xa4
    "11111111", -- 1313 - 0x521  :  255 - 0xff
    "11111111", -- 1314 - 0x522  :  255 - 0xff
    "11111111", -- 1315 - 0x523  :  255 - 0xff
    "11111111", -- 1316 - 0x524  :  255 - 0xff
    "11111110", -- 1317 - 0x525  :  254 - 0xfe
    "10111110", -- 1318 - 0x526  :  190 - 0xbe
    "11001110", -- 1319 - 0x527  :  206 - 0xce
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- Background 0xa5
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "00000011", -- 1324 - 0x52c  :    3 - 0x3
    "00000100", -- 1325 - 0x52d  :    4 - 0x4
    "00000100", -- 1326 - 0x52e  :    4 - 0x4
    "00000100", -- 1327 - 0x52f  :    4 - 0x4
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Background 0xa6
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "01100000", -- 1330 - 0x532  :   96 - 0x60
    "00110000", -- 1331 - 0x533  :   48 - 0x30
    "00110000", -- 1332 - 0x534  :   48 - 0x30
    "10011000", -- 1333 - 0x535  :  152 - 0x98
    "10011000", -- 1334 - 0x536  :  152 - 0x98
    "10011000", -- 1335 - 0x537  :  152 - 0x98
    "00000100", -- 1336 - 0x538  :    4 - 0x4 -- Background 0xa7
    "00000100", -- 1337 - 0x539  :    4 - 0x4
    "00000100", -- 1338 - 0x53a  :    4 - 0x4
    "00000100", -- 1339 - 0x53b  :    4 - 0x4
    "00000100", -- 1340 - 0x53c  :    4 - 0x4
    "00000011", -- 1341 - 0x53d  :    3 - 0x3
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "10011000", -- 1344 - 0x540  :  152 - 0x98 -- Background 0xa8
    "10011000", -- 1345 - 0x541  :  152 - 0x98
    "10011000", -- 1346 - 0x542  :  152 - 0x98
    "10011000", -- 1347 - 0x543  :  152 - 0x98
    "10011000", -- 1348 - 0x544  :  152 - 0x98
    "00110000", -- 1349 - 0x545  :   48 - 0x30
    "00110000", -- 1350 - 0x546  :   48 - 0x30
    "01100000", -- 1351 - 0x547  :   96 - 0x60
    "00001111", -- 1352 - 0x548  :   15 - 0xf -- Background 0xa9
    "11101111", -- 1353 - 0x549  :  239 - 0xef
    "11101111", -- 1354 - 0x54a  :  239 - 0xef
    "11101111", -- 1355 - 0x54b  :  239 - 0xef
    "11101111", -- 1356 - 0x54c  :  239 - 0xef
    "11101111", -- 1357 - 0x54d  :  239 - 0xef
    "11101111", -- 1358 - 0x54e  :  239 - 0xef
    "11100000", -- 1359 - 0x54f  :  224 - 0xe0
    "11100000", -- 1360 - 0x550  :  224 - 0xe0 -- Background 0xaa
    "11101111", -- 1361 - 0x551  :  239 - 0xef
    "11101111", -- 1362 - 0x552  :  239 - 0xef
    "11101111", -- 1363 - 0x553  :  239 - 0xef
    "11101111", -- 1364 - 0x554  :  239 - 0xef
    "11101111", -- 1365 - 0x555  :  239 - 0xef
    "11101111", -- 1366 - 0x556  :  239 - 0xef
    "00001111", -- 1367 - 0x557  :   15 - 0xf
    "10000000", -- 1368 - 0x558  :  128 - 0x80 -- Background 0xab
    "01000000", -- 1369 - 0x559  :   64 - 0x40
    "00100000", -- 1370 - 0x55a  :   32 - 0x20
    "00010000", -- 1371 - 0x55b  :   16 - 0x10
    "00001111", -- 1372 - 0x55c  :   15 - 0xf
    "00001111", -- 1373 - 0x55d  :   15 - 0xf
    "00001111", -- 1374 - 0x55e  :   15 - 0xf
    "00001111", -- 1375 - 0x55f  :   15 - 0xf
    "00001111", -- 1376 - 0x560  :   15 - 0xf -- Background 0xac
    "00001111", -- 1377 - 0x561  :   15 - 0xf
    "00001111", -- 1378 - 0x562  :   15 - 0xf
    "00001111", -- 1379 - 0x563  :   15 - 0xf
    "00011111", -- 1380 - 0x564  :   31 - 0x1f
    "00111111", -- 1381 - 0x565  :   63 - 0x3f
    "01111111", -- 1382 - 0x566  :  127 - 0x7f
    "11111111", -- 1383 - 0x567  :  255 - 0xff
    "00000001", -- 1384 - 0x568  :    1 - 0x1 -- Background 0xad
    "00000011", -- 1385 - 0x569  :    3 - 0x3
    "00000111", -- 1386 - 0x56a  :    7 - 0x7
    "00001111", -- 1387 - 0x56b  :   15 - 0xf
    "11111111", -- 1388 - 0x56c  :  255 - 0xff
    "11111111", -- 1389 - 0x56d  :  255 - 0xff
    "11111111", -- 1390 - 0x56e  :  255 - 0xff
    "11111111", -- 1391 - 0x56f  :  255 - 0xff
    "11111111", -- 1392 - 0x570  :  255 - 0xff -- Background 0xae
    "11111111", -- 1393 - 0x571  :  255 - 0xff
    "11111111", -- 1394 - 0x572  :  255 - 0xff
    "11111111", -- 1395 - 0x573  :  255 - 0xff
    "11111111", -- 1396 - 0x574  :  255 - 0xff
    "11111111", -- 1397 - 0x575  :  255 - 0xff
    "11111111", -- 1398 - 0x576  :  255 - 0xff
    "11111111", -- 1399 - 0x577  :  255 - 0xff
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Background 0xaf
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "00011111", -- 1408 - 0x580  :   31 - 0x1f -- Background 0xb0
    "00100000", -- 1409 - 0x581  :   32 - 0x20
    "01000000", -- 1410 - 0x582  :   64 - 0x40
    "01000000", -- 1411 - 0x583  :   64 - 0x40
    "01000000", -- 1412 - 0x584  :   64 - 0x40
    "10000000", -- 1413 - 0x585  :  128 - 0x80
    "10000010", -- 1414 - 0x586  :  130 - 0x82
    "10000010", -- 1415 - 0x587  :  130 - 0x82
    "10000010", -- 1416 - 0x588  :  130 - 0x82 -- Background 0xb1
    "10000000", -- 1417 - 0x589  :  128 - 0x80
    "10100000", -- 1418 - 0x58a  :  160 - 0xa0
    "01000100", -- 1419 - 0x58b  :   68 - 0x44
    "01000011", -- 1420 - 0x58c  :   67 - 0x43
    "01000000", -- 1421 - 0x58d  :   64 - 0x40
    "00100001", -- 1422 - 0x58e  :   33 - 0x21
    "00011110", -- 1423 - 0x58f  :   30 - 0x1e
    "11111000", -- 1424 - 0x590  :  248 - 0xf8 -- Background 0xb2
    "00000100", -- 1425 - 0x591  :    4 - 0x4
    "00000010", -- 1426 - 0x592  :    2 - 0x2
    "00000010", -- 1427 - 0x593  :    2 - 0x2
    "00000010", -- 1428 - 0x594  :    2 - 0x2
    "00000001", -- 1429 - 0x595  :    1 - 0x1
    "01000001", -- 1430 - 0x596  :   65 - 0x41
    "01000001", -- 1431 - 0x597  :   65 - 0x41
    "01000001", -- 1432 - 0x598  :   65 - 0x41 -- Background 0xb3
    "00000001", -- 1433 - 0x599  :    1 - 0x1
    "00000101", -- 1434 - 0x59a  :    5 - 0x5
    "00100010", -- 1435 - 0x59b  :   34 - 0x22
    "11000010", -- 1436 - 0x59c  :  194 - 0xc2
    "00000010", -- 1437 - 0x59d  :    2 - 0x2
    "10000100", -- 1438 - 0x59e  :  132 - 0x84
    "01111000", -- 1439 - 0x59f  :  120 - 0x78
    "10000000", -- 1440 - 0x5a0  :  128 - 0x80 -- Background 0xb4
    "01111111", -- 1441 - 0x5a1  :  127 - 0x7f
    "01111111", -- 1442 - 0x5a2  :  127 - 0x7f
    "01111111", -- 1443 - 0x5a3  :  127 - 0x7f
    "01111111", -- 1444 - 0x5a4  :  127 - 0x7f
    "01111111", -- 1445 - 0x5a5  :  127 - 0x7f
    "01111111", -- 1446 - 0x5a6  :  127 - 0x7f
    "01111111", -- 1447 - 0x5a7  :  127 - 0x7f
    "01100001", -- 1448 - 0x5a8  :   97 - 0x61 -- Background 0xb5
    "11011111", -- 1449 - 0x5a9  :  223 - 0xdf
    "11011111", -- 1450 - 0x5aa  :  223 - 0xdf
    "11011111", -- 1451 - 0x5ab  :  223 - 0xdf
    "11011111", -- 1452 - 0x5ac  :  223 - 0xdf
    "11111111", -- 1453 - 0x5ad  :  255 - 0xff
    "11000001", -- 1454 - 0x5ae  :  193 - 0xc1
    "11011111", -- 1455 - 0x5af  :  223 - 0xdf
    "01111111", -- 1456 - 0x5b0  :  127 - 0x7f -- Background 0xb6
    "01111111", -- 1457 - 0x5b1  :  127 - 0x7f
    "11111111", -- 1458 - 0x5b2  :  255 - 0xff
    "00111111", -- 1459 - 0x5b3  :   63 - 0x3f
    "01001111", -- 1460 - 0x5b4  :   79 - 0x4f
    "01110001", -- 1461 - 0x5b5  :  113 - 0x71
    "01111111", -- 1462 - 0x5b6  :  127 - 0x7f
    "11111111", -- 1463 - 0x5b7  :  255 - 0xff
    "11011111", -- 1464 - 0x5b8  :  223 - 0xdf -- Background 0xb7
    "11011111", -- 1465 - 0x5b9  :  223 - 0xdf
    "10111111", -- 1466 - 0x5ba  :  191 - 0xbf
    "10111111", -- 1467 - 0x5bb  :  191 - 0xbf
    "01111111", -- 1468 - 0x5bc  :  127 - 0x7f
    "01111111", -- 1469 - 0x5bd  :  127 - 0x7f
    "01111111", -- 1470 - 0x5be  :  127 - 0x7f
    "01111111", -- 1471 - 0x5bf  :  127 - 0x7f
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Background 0xb8
    "00000000", -- 1473 - 0x5c1  :    0 - 0x0
    "00000011", -- 1474 - 0x5c2  :    3 - 0x3
    "00001100", -- 1475 - 0x5c3  :   12 - 0xc
    "00010000", -- 1476 - 0x5c4  :   16 - 0x10
    "00100000", -- 1477 - 0x5c5  :   32 - 0x20
    "01000000", -- 1478 - 0x5c6  :   64 - 0x40
    "01000000", -- 1479 - 0x5c7  :   64 - 0x40
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0 -- Background 0xb9
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "11000000", -- 1482 - 0x5ca  :  192 - 0xc0
    "00110000", -- 1483 - 0x5cb  :   48 - 0x30
    "00001000", -- 1484 - 0x5cc  :    8 - 0x8
    "00000100", -- 1485 - 0x5cd  :    4 - 0x4
    "00000010", -- 1486 - 0x5ce  :    2 - 0x2
    "00000010", -- 1487 - 0x5cf  :    2 - 0x2
    "10000000", -- 1488 - 0x5d0  :  128 - 0x80 -- Background 0xba
    "10000000", -- 1489 - 0x5d1  :  128 - 0x80
    "10000000", -- 1490 - 0x5d2  :  128 - 0x80
    "10000000", -- 1491 - 0x5d3  :  128 - 0x80
    "10000000", -- 1492 - 0x5d4  :  128 - 0x80
    "10000000", -- 1493 - 0x5d5  :  128 - 0x80
    "10000000", -- 1494 - 0x5d6  :  128 - 0x80
    "10000000", -- 1495 - 0x5d7  :  128 - 0x80
    "00000001", -- 1496 - 0x5d8  :    1 - 0x1 -- Background 0xbb
    "00000001", -- 1497 - 0x5d9  :    1 - 0x1
    "00000001", -- 1498 - 0x5da  :    1 - 0x1
    "00000001", -- 1499 - 0x5db  :    1 - 0x1
    "00000001", -- 1500 - 0x5dc  :    1 - 0x1
    "00000001", -- 1501 - 0x5dd  :    1 - 0x1
    "00000001", -- 1502 - 0x5de  :    1 - 0x1
    "00000001", -- 1503 - 0x5df  :    1 - 0x1
    "01000000", -- 1504 - 0x5e0  :   64 - 0x40 -- Background 0xbc
    "01000000", -- 1505 - 0x5e1  :   64 - 0x40
    "01000000", -- 1506 - 0x5e2  :   64 - 0x40
    "00100000", -- 1507 - 0x5e3  :   32 - 0x20
    "00110000", -- 1508 - 0x5e4  :   48 - 0x30
    "00011100", -- 1509 - 0x5e5  :   28 - 0x1c
    "00001111", -- 1510 - 0x5e6  :   15 - 0xf
    "00000111", -- 1511 - 0x5e7  :    7 - 0x7
    "00000010", -- 1512 - 0x5e8  :    2 - 0x2 -- Background 0xbd
    "00000010", -- 1513 - 0x5e9  :    2 - 0x2
    "00000010", -- 1514 - 0x5ea  :    2 - 0x2
    "00000100", -- 1515 - 0x5eb  :    4 - 0x4
    "00001100", -- 1516 - 0x5ec  :   12 - 0xc
    "00111000", -- 1517 - 0x5ed  :   56 - 0x38
    "11110000", -- 1518 - 0x5ee  :  240 - 0xf0
    "11110000", -- 1519 - 0x5ef  :  240 - 0xf0
    "00001000", -- 1520 - 0x5f0  :    8 - 0x8 -- Background 0xbe
    "00001000", -- 1521 - 0x5f1  :    8 - 0x8
    "00001000", -- 1522 - 0x5f2  :    8 - 0x8
    "00001000", -- 1523 - 0x5f3  :    8 - 0x8
    "00001000", -- 1524 - 0x5f4  :    8 - 0x8
    "00001100", -- 1525 - 0x5f5  :   12 - 0xc
    "00000101", -- 1526 - 0x5f6  :    5 - 0x5
    "00001010", -- 1527 - 0x5f7  :   10 - 0xa
    "00010000", -- 1528 - 0x5f8  :   16 - 0x10 -- Background 0xbf
    "01010000", -- 1529 - 0x5f9  :   80 - 0x50
    "01010000", -- 1530 - 0x5fa  :   80 - 0x50
    "01010000", -- 1531 - 0x5fb  :   80 - 0x50
    "01010000", -- 1532 - 0x5fc  :   80 - 0x50
    "00110000", -- 1533 - 0x5fd  :   48 - 0x30
    "10100000", -- 1534 - 0x5fe  :  160 - 0xa0
    "01010000", -- 1535 - 0x5ff  :   80 - 0x50
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Background 0xc0
    "01000001", -- 1537 - 0x601  :   65 - 0x41
    "00100010", -- 1538 - 0x602  :   34 - 0x22
    "00100010", -- 1539 - 0x603  :   34 - 0x22
    "00011100", -- 1540 - 0x604  :   28 - 0x1c
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000000", -- 1542 - 0x606  :    0 - 0x0
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "11100011", -- 1544 - 0x608  :  227 - 0xe3 -- Background 0xc1
    "00010100", -- 1545 - 0x609  :   20 - 0x14
    "00111110", -- 1546 - 0x60a  :   62 - 0x3e
    "00111110", -- 1547 - 0x60b  :   62 - 0x3e
    "00111110", -- 1548 - 0x60c  :   62 - 0x3e
    "00111110", -- 1549 - 0x60d  :   62 - 0x3e
    "00010100", -- 1550 - 0x60e  :   20 - 0x14
    "11100011", -- 1551 - 0x60f  :  227 - 0xe3
    "11111111", -- 1552 - 0x610  :  255 - 0xff -- Background 0xc2
    "11111111", -- 1553 - 0x611  :  255 - 0xff
    "11111000", -- 1554 - 0x612  :  248 - 0xf8
    "11110000", -- 1555 - 0x613  :  240 - 0xf0
    "11110000", -- 1556 - 0x614  :  240 - 0xf0
    "11100000", -- 1557 - 0x615  :  224 - 0xe0
    "11100000", -- 1558 - 0x616  :  224 - 0xe0
    "11100000", -- 1559 - 0x617  :  224 - 0xe0
    "11111111", -- 1560 - 0x618  :  255 - 0xff -- Background 0xc3
    "11111111", -- 1561 - 0x619  :  255 - 0xff
    "01111111", -- 1562 - 0x61a  :  127 - 0x7f
    "00111111", -- 1563 - 0x61b  :   63 - 0x3f
    "00111111", -- 1564 - 0x61c  :   63 - 0x3f
    "10011111", -- 1565 - 0x61d  :  159 - 0x9f
    "10011111", -- 1566 - 0x61e  :  159 - 0x9f
    "10011111", -- 1567 - 0x61f  :  159 - 0x9f
    "11100000", -- 1568 - 0x620  :  224 - 0xe0 -- Background 0xc4
    "11100000", -- 1569 - 0x621  :  224 - 0xe0
    "11100000", -- 1570 - 0x622  :  224 - 0xe0
    "11100000", -- 1571 - 0x623  :  224 - 0xe0
    "11100000", -- 1572 - 0x624  :  224 - 0xe0
    "11110011", -- 1573 - 0x625  :  243 - 0xf3
    "11110000", -- 1574 - 0x626  :  240 - 0xf0
    "11111000", -- 1575 - 0x627  :  248 - 0xf8
    "10011111", -- 1576 - 0x628  :  159 - 0x9f -- Background 0xc5
    "10011111", -- 1577 - 0x629  :  159 - 0x9f
    "10011111", -- 1578 - 0x62a  :  159 - 0x9f
    "10011111", -- 1579 - 0x62b  :  159 - 0x9f
    "10011111", -- 1580 - 0x62c  :  159 - 0x9f
    "00111111", -- 1581 - 0x62d  :   63 - 0x3f
    "00111111", -- 1582 - 0x62e  :   63 - 0x3f
    "01111111", -- 1583 - 0x62f  :  127 - 0x7f
    "00000000", -- 1584 - 0x630  :    0 - 0x0 -- Background 0xc6
    "01110000", -- 1585 - 0x631  :  112 - 0x70
    "00011111", -- 1586 - 0x632  :   31 - 0x1f
    "00010000", -- 1587 - 0x633  :   16 - 0x10
    "01110000", -- 1588 - 0x634  :  112 - 0x70
    "01111111", -- 1589 - 0x635  :  127 - 0x7f
    "01111111", -- 1590 - 0x636  :  127 - 0x7f
    "01111111", -- 1591 - 0x637  :  127 - 0x7f
    "00000000", -- 1592 - 0x638  :    0 - 0x0 -- Background 0xc7
    "00000011", -- 1593 - 0x639  :    3 - 0x3
    "11111000", -- 1594 - 0x63a  :  248 - 0xf8
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "00000011", -- 1596 - 0x63c  :    3 - 0x3
    "11111011", -- 1597 - 0x63d  :  251 - 0xfb
    "11111011", -- 1598 - 0x63e  :  251 - 0xfb
    "11111011", -- 1599 - 0x63f  :  251 - 0xfb
    "01111100", -- 1600 - 0x640  :  124 - 0x7c -- Background 0xc8
    "01111011", -- 1601 - 0x641  :  123 - 0x7b
    "01110110", -- 1602 - 0x642  :  118 - 0x76
    "01110101", -- 1603 - 0x643  :  117 - 0x75
    "01110101", -- 1604 - 0x644  :  117 - 0x75
    "01110111", -- 1605 - 0x645  :  119 - 0x77
    "00010111", -- 1606 - 0x646  :   23 - 0x17
    "01100111", -- 1607 - 0x647  :  103 - 0x67
    "00111011", -- 1608 - 0x648  :   59 - 0x3b -- Background 0xc9
    "11111011", -- 1609 - 0x649  :  251 - 0xfb
    "01111011", -- 1610 - 0x64a  :  123 - 0x7b
    "11111011", -- 1611 - 0x64b  :  251 - 0xfb
    "11111011", -- 1612 - 0x64c  :  251 - 0xfb
    "11110011", -- 1613 - 0x64d  :  243 - 0xf3
    "11111000", -- 1614 - 0x64e  :  248 - 0xf8
    "11110011", -- 1615 - 0x64f  :  243 - 0xf3
    "00001111", -- 1616 - 0x650  :   15 - 0xf -- Background 0xca
    "00001111", -- 1617 - 0x651  :   15 - 0xf
    "00011111", -- 1618 - 0x652  :   31 - 0x1f
    "00011111", -- 1619 - 0x653  :   31 - 0x1f
    "00111111", -- 1620 - 0x654  :   63 - 0x3f
    "00111100", -- 1621 - 0x655  :   60 - 0x3c
    "01111000", -- 1622 - 0x656  :  120 - 0x78
    "01111010", -- 1623 - 0x657  :  122 - 0x7a
    "11111000", -- 1624 - 0x658  :  248 - 0xf8 -- Background 0xcb
    "11111000", -- 1625 - 0x659  :  248 - 0xf8
    "11111100", -- 1626 - 0x65a  :  252 - 0xfc
    "11111100", -- 1627 - 0x65b  :  252 - 0xfc
    "11111110", -- 1628 - 0x65c  :  254 - 0xfe
    "00111110", -- 1629 - 0x65d  :   62 - 0x3e
    "00011110", -- 1630 - 0x65e  :   30 - 0x1e
    "01011111", -- 1631 - 0x65f  :   95 - 0x5f
    "01110110", -- 1632 - 0x660  :  118 - 0x76 -- Background 0xcc
    "01110110", -- 1633 - 0x661  :  118 - 0x76
    "01110110", -- 1634 - 0x662  :  118 - 0x76
    "01110000", -- 1635 - 0x663  :  112 - 0x70
    "01111101", -- 1636 - 0x664  :  125 - 0x7d
    "01111100", -- 1637 - 0x665  :  124 - 0x7c
    "01111111", -- 1638 - 0x666  :  127 - 0x7f
    "01111111", -- 1639 - 0x667  :  127 - 0x7f
    "01101111", -- 1640 - 0x668  :  111 - 0x6f -- Background 0xcd
    "01101111", -- 1641 - 0x669  :  111 - 0x6f
    "01101111", -- 1642 - 0x66a  :  111 - 0x6f
    "00001111", -- 1643 - 0x66b  :   15 - 0xf
    "10111111", -- 1644 - 0x66c  :  191 - 0xbf
    "00111111", -- 1645 - 0x66d  :   63 - 0x3f
    "11111111", -- 1646 - 0x66e  :  255 - 0xff
    "11111111", -- 1647 - 0x66f  :  255 - 0xff
    "00111100", -- 1648 - 0x670  :   60 - 0x3c -- Background 0xce
    "01111110", -- 1649 - 0x671  :  126 - 0x7e
    "01111110", -- 1650 - 0x672  :  126 - 0x7e
    "11111111", -- 1651 - 0x673  :  255 - 0xff
    "11111111", -- 1652 - 0x674  :  255 - 0xff
    "11111111", -- 1653 - 0x675  :  255 - 0xff
    "01000010", -- 1654 - 0x676  :   66 - 0x42
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "11110000", -- 1664 - 0x680  :  240 - 0xf0 -- Background 0xd0
    "11100000", -- 1665 - 0x681  :  224 - 0xe0
    "11100000", -- 1666 - 0x682  :  224 - 0xe0
    "11000000", -- 1667 - 0x683  :  192 - 0xc0
    "11000000", -- 1668 - 0x684  :  192 - 0xc0
    "10000000", -- 1669 - 0x685  :  128 - 0x80
    "10000000", -- 1670 - 0x686  :  128 - 0x80
    "10000000", -- 1671 - 0x687  :  128 - 0x80
    "00001111", -- 1672 - 0x688  :   15 - 0xf -- Background 0xd1
    "00000111", -- 1673 - 0x689  :    7 - 0x7
    "00000111", -- 1674 - 0x68a  :    7 - 0x7
    "00000011", -- 1675 - 0x68b  :    3 - 0x3
    "00000011", -- 1676 - 0x68c  :    3 - 0x3
    "00000001", -- 1677 - 0x68d  :    1 - 0x1
    "00000001", -- 1678 - 0x68e  :    1 - 0x1
    "00000001", -- 1679 - 0x68f  :    1 - 0x1
    "10000000", -- 1680 - 0x690  :  128 - 0x80 -- Background 0xd2
    "10000000", -- 1681 - 0x691  :  128 - 0x80
    "11000000", -- 1682 - 0x692  :  192 - 0xc0
    "11000000", -- 1683 - 0x693  :  192 - 0xc0
    "11100000", -- 1684 - 0x694  :  224 - 0xe0
    "11111000", -- 1685 - 0x695  :  248 - 0xf8
    "11111110", -- 1686 - 0x696  :  254 - 0xfe
    "11111111", -- 1687 - 0x697  :  255 - 0xff
    "11111111", -- 1688 - 0x698  :  255 - 0xff -- Background 0xd3
    "01111111", -- 1689 - 0x699  :  127 - 0x7f
    "00011111", -- 1690 - 0x69a  :   31 - 0x1f
    "00000111", -- 1691 - 0x69b  :    7 - 0x7
    "00000011", -- 1692 - 0x69c  :    3 - 0x3
    "00000011", -- 1693 - 0x69d  :    3 - 0x3
    "00000001", -- 1694 - 0x69e  :    1 - 0x1
    "10000001", -- 1695 - 0x69f  :  129 - 0x81
    "10000000", -- 1696 - 0x6a0  :  128 - 0x80 -- Background 0xd4
    "10000000", -- 1697 - 0x6a1  :  128 - 0x80
    "10000000", -- 1698 - 0x6a2  :  128 - 0x80
    "11000000", -- 1699 - 0x6a3  :  192 - 0xc0
    "11000000", -- 1700 - 0x6a4  :  192 - 0xc0
    "11100000", -- 1701 - 0x6a5  :  224 - 0xe0
    "11100000", -- 1702 - 0x6a6  :  224 - 0xe0
    "11110000", -- 1703 - 0x6a7  :  240 - 0xf0
    "00000001", -- 1704 - 0x6a8  :    1 - 0x1 -- Background 0xd5
    "00000001", -- 1705 - 0x6a9  :    1 - 0x1
    "00000001", -- 1706 - 0x6aa  :    1 - 0x1
    "00000011", -- 1707 - 0x6ab  :    3 - 0x3
    "00000011", -- 1708 - 0x6ac  :    3 - 0x3
    "00000111", -- 1709 - 0x6ad  :    7 - 0x7
    "00000111", -- 1710 - 0x6ae  :    7 - 0x7
    "00001111", -- 1711 - 0x6af  :   15 - 0xf
    "11111111", -- 1712 - 0x6b0  :  255 - 0xff -- Background 0xd6
    "11111111", -- 1713 - 0x6b1  :  255 - 0xff
    "11111111", -- 1714 - 0x6b2  :  255 - 0xff
    "11111111", -- 1715 - 0x6b3  :  255 - 0xff
    "11111111", -- 1716 - 0x6b4  :  255 - 0xff
    "11111111", -- 1717 - 0x6b5  :  255 - 0xff
    "11111111", -- 1718 - 0x6b6  :  255 - 0xff
    "11111111", -- 1719 - 0x6b7  :  255 - 0xff
    "11111111", -- 1720 - 0x6b8  :  255 - 0xff -- Background 0xd7
    "11111111", -- 1721 - 0x6b9  :  255 - 0xff
    "11111111", -- 1722 - 0x6ba  :  255 - 0xff
    "11111111", -- 1723 - 0x6bb  :  255 - 0xff
    "11111111", -- 1724 - 0x6bc  :  255 - 0xff
    "11111111", -- 1725 - 0x6bd  :  255 - 0xff
    "11111111", -- 1726 - 0x6be  :  255 - 0xff
    "11111111", -- 1727 - 0x6bf  :  255 - 0xff
    "10000001", -- 1728 - 0x6c0  :  129 - 0x81 -- Background 0xd8
    "10000001", -- 1729 - 0x6c1  :  129 - 0x81
    "10000001", -- 1730 - 0x6c2  :  129 - 0x81
    "10000001", -- 1731 - 0x6c3  :  129 - 0x81
    "10000001", -- 1732 - 0x6c4  :  129 - 0x81
    "10000001", -- 1733 - 0x6c5  :  129 - 0x81
    "10000001", -- 1734 - 0x6c6  :  129 - 0x81
    "10000001", -- 1735 - 0x6c7  :  129 - 0x81
    "00000001", -- 1736 - 0x6c8  :    1 - 0x1 -- Background 0xd9
    "00000001", -- 1737 - 0x6c9  :    1 - 0x1
    "00000001", -- 1738 - 0x6ca  :    1 - 0x1
    "00000011", -- 1739 - 0x6cb  :    3 - 0x3
    "00000011", -- 1740 - 0x6cc  :    3 - 0x3
    "00000111", -- 1741 - 0x6cd  :    7 - 0x7
    "00000111", -- 1742 - 0x6ce  :    7 - 0x7
    "00001111", -- 1743 - 0x6cf  :   15 - 0xf
    "00000001", -- 1744 - 0x6d0  :    1 - 0x1 -- Background 0xda
    "00000001", -- 1745 - 0x6d1  :    1 - 0x1
    "00000001", -- 1746 - 0x6d2  :    1 - 0x1
    "00000001", -- 1747 - 0x6d3  :    1 - 0x1
    "00000001", -- 1748 - 0x6d4  :    1 - 0x1
    "00000001", -- 1749 - 0x6d5  :    1 - 0x1
    "00000001", -- 1750 - 0x6d6  :    1 - 0x1
    "00000001", -- 1751 - 0x6d7  :    1 - 0x1
    "10000001", -- 1752 - 0x6d8  :  129 - 0x81 -- Background 0xdb
    "10000001", -- 1753 - 0x6d9  :  129 - 0x81
    "10000001", -- 1754 - 0x6da  :  129 - 0x81
    "10000001", -- 1755 - 0x6db  :  129 - 0x81
    "10000001", -- 1756 - 0x6dc  :  129 - 0x81
    "10000001", -- 1757 - 0x6dd  :  129 - 0x81
    "10000001", -- 1758 - 0x6de  :  129 - 0x81
    "10000001", -- 1759 - 0x6df  :  129 - 0x81
    "11111111", -- 1760 - 0x6e0  :  255 - 0xff -- Background 0xdc
    "00000011", -- 1761 - 0x6e1  :    3 - 0x3
    "00000011", -- 1762 - 0x6e2  :    3 - 0x3
    "00000011", -- 1763 - 0x6e3  :    3 - 0x3
    "00000011", -- 1764 - 0x6e4  :    3 - 0x3
    "00000011", -- 1765 - 0x6e5  :    3 - 0x3
    "00000011", -- 1766 - 0x6e6  :    3 - 0x3
    "11111111", -- 1767 - 0x6e7  :  255 - 0xff
    "11111111", -- 1768 - 0x6e8  :  255 - 0xff -- Background 0xdd
    "11111111", -- 1769 - 0x6e9  :  255 - 0xff
    "11111111", -- 1770 - 0x6ea  :  255 - 0xff
    "11111111", -- 1771 - 0x6eb  :  255 - 0xff
    "11111111", -- 1772 - 0x6ec  :  255 - 0xff
    "11111111", -- 1773 - 0x6ed  :  255 - 0xff
    "11111111", -- 1774 - 0x6ee  :  255 - 0xff
    "11111111", -- 1775 - 0x6ef  :  255 - 0xff
    "10000000", -- 1776 - 0x6f0  :  128 - 0x80 -- Background 0xde
    "10000000", -- 1777 - 0x6f1  :  128 - 0x80
    "10000000", -- 1778 - 0x6f2  :  128 - 0x80
    "10000000", -- 1779 - 0x6f3  :  128 - 0x80
    "10000000", -- 1780 - 0x6f4  :  128 - 0x80
    "10000000", -- 1781 - 0x6f5  :  128 - 0x80
    "10000000", -- 1782 - 0x6f6  :  128 - 0x80
    "10000000", -- 1783 - 0x6f7  :  128 - 0x80
    "00000001", -- 1784 - 0x6f8  :    1 - 0x1 -- Background 0xdf
    "00000001", -- 1785 - 0x6f9  :    1 - 0x1
    "00000001", -- 1786 - 0x6fa  :    1 - 0x1
    "00000011", -- 1787 - 0x6fb  :    3 - 0x3
    "00000111", -- 1788 - 0x6fc  :    7 - 0x7
    "00000011", -- 1789 - 0x6fd  :    3 - 0x3
    "00000001", -- 1790 - 0x6fe  :    1 - 0x1
    "00000001", -- 1791 - 0x6ff  :    1 - 0x1
    "10000001", -- 1792 - 0x700  :  129 - 0x81 -- Background 0xe0
    "10000001", -- 1793 - 0x701  :  129 - 0x81
    "10000001", -- 1794 - 0x702  :  129 - 0x81
    "10000001", -- 1795 - 0x703  :  129 - 0x81
    "10000001", -- 1796 - 0x704  :  129 - 0x81
    "10000001", -- 1797 - 0x705  :  129 - 0x81
    "10000001", -- 1798 - 0x706  :  129 - 0x81
    "10000001", -- 1799 - 0x707  :  129 - 0x81
    "11111111", -- 1800 - 0x708  :  255 - 0xff -- Background 0xe1
    "11111111", -- 1801 - 0x709  :  255 - 0xff
    "11111111", -- 1802 - 0x70a  :  255 - 0xff
    "11111111", -- 1803 - 0x70b  :  255 - 0xff
    "11111111", -- 1804 - 0x70c  :  255 - 0xff
    "11111111", -- 1805 - 0x70d  :  255 - 0xff
    "11111111", -- 1806 - 0x70e  :  255 - 0xff
    "11111111", -- 1807 - 0x70f  :  255 - 0xff
    "11111111", -- 1808 - 0x710  :  255 - 0xff -- Background 0xe2
    "11111111", -- 1809 - 0x711  :  255 - 0xff
    "11111111", -- 1810 - 0x712  :  255 - 0xff
    "11111111", -- 1811 - 0x713  :  255 - 0xff
    "11111111", -- 1812 - 0x714  :  255 - 0xff
    "11111111", -- 1813 - 0x715  :  255 - 0xff
    "11111111", -- 1814 - 0x716  :  255 - 0xff
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "10000001", -- 1816 - 0x718  :  129 - 0x81 -- Background 0xe3
    "10000001", -- 1817 - 0x719  :  129 - 0x81
    "10000001", -- 1818 - 0x71a  :  129 - 0x81
    "10000001", -- 1819 - 0x71b  :  129 - 0x81
    "10000001", -- 1820 - 0x71c  :  129 - 0x81
    "10000001", -- 1821 - 0x71d  :  129 - 0x81
    "10000001", -- 1822 - 0x71e  :  129 - 0x81
    "10000001", -- 1823 - 0x71f  :  129 - 0x81
    "10000000", -- 1824 - 0x720  :  128 - 0x80 -- Background 0xe4
    "10000000", -- 1825 - 0x721  :  128 - 0x80
    "11000000", -- 1826 - 0x722  :  192 - 0xc0
    "11000000", -- 1827 - 0x723  :  192 - 0xc0
    "11100000", -- 1828 - 0x724  :  224 - 0xe0
    "11111000", -- 1829 - 0x725  :  248 - 0xf8
    "11111110", -- 1830 - 0x726  :  254 - 0xfe
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "11111111", -- 1832 - 0x728  :  255 - 0xff -- Background 0xe5
    "01111111", -- 1833 - 0x729  :  127 - 0x7f
    "00011111", -- 1834 - 0x72a  :   31 - 0x1f
    "00000111", -- 1835 - 0x72b  :    7 - 0x7
    "00000011", -- 1836 - 0x72c  :    3 - 0x3
    "00000011", -- 1837 - 0x72d  :    3 - 0x3
    "00000001", -- 1838 - 0x72e  :    1 - 0x1
    "10000001", -- 1839 - 0x72f  :  129 - 0x81
    "10000001", -- 1840 - 0x730  :  129 - 0x81 -- Background 0xe6
    "10000001", -- 1841 - 0x731  :  129 - 0x81
    "10000001", -- 1842 - 0x732  :  129 - 0x81
    "10000001", -- 1843 - 0x733  :  129 - 0x81
    "10000001", -- 1844 - 0x734  :  129 - 0x81
    "10000001", -- 1845 - 0x735  :  129 - 0x81
    "10000001", -- 1846 - 0x736  :  129 - 0x81
    "10000001", -- 1847 - 0x737  :  129 - 0x81
    "10000001", -- 1848 - 0x738  :  129 - 0x81 -- Background 0xe7
    "10000001", -- 1849 - 0x739  :  129 - 0x81
    "10000001", -- 1850 - 0x73a  :  129 - 0x81
    "10000001", -- 1851 - 0x73b  :  129 - 0x81
    "10000001", -- 1852 - 0x73c  :  129 - 0x81
    "10000001", -- 1853 - 0x73d  :  129 - 0x81
    "10000001", -- 1854 - 0x73e  :  129 - 0x81
    "10000001", -- 1855 - 0x73f  :  129 - 0x81
    "01111110", -- 1856 - 0x740  :  126 - 0x7e -- Background 0xe8
    "00111100", -- 1857 - 0x741  :   60 - 0x3c
    "00111100", -- 1858 - 0x742  :   60 - 0x3c
    "00011000", -- 1859 - 0x743  :   24 - 0x18
    "00011000", -- 1860 - 0x744  :   24 - 0x18
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "11110010", -- 1864 - 0x748  :  242 - 0xf2 -- Background 0xe9
    "11111110", -- 1865 - 0x749  :  254 - 0xfe
    "11111110", -- 1866 - 0x74a  :  254 - 0xfe
    "11111111", -- 1867 - 0x74b  :  255 - 0xff
    "11111111", -- 1868 - 0x74c  :  255 - 0xff
    "11101111", -- 1869 - 0x74d  :  239 - 0xef
    "11110111", -- 1870 - 0x74e  :  247 - 0xf7
    "11111000", -- 1871 - 0x74f  :  248 - 0xf8
    "10111111", -- 1872 - 0x750  :  191 - 0xbf -- Background 0xea
    "10111110", -- 1873 - 0x751  :  190 - 0xbe
    "10111101", -- 1874 - 0x752  :  189 - 0xbd
    "01111011", -- 1875 - 0x753  :  123 - 0x7b
    "01111011", -- 1876 - 0x754  :  123 - 0x7b
    "00000111", -- 1877 - 0x755  :    7 - 0x7
    "11110011", -- 1878 - 0x756  :  243 - 0xf3
    "11111101", -- 1879 - 0x757  :  253 - 0xfd
    "11111111", -- 1880 - 0x758  :  255 - 0xff -- Background 0xeb
    "11111111", -- 1881 - 0x759  :  255 - 0xff
    "11111111", -- 1882 - 0x75a  :  255 - 0xff
    "01100111", -- 1883 - 0x75b  :  103 - 0x67
    "01011001", -- 1884 - 0x75c  :   89 - 0x59
    "10011110", -- 1885 - 0x75d  :  158 - 0x9e
    "10111111", -- 1886 - 0x75e  :  191 - 0xbf
    "10111111", -- 1887 - 0x75f  :  191 - 0xbf
    "00100000", -- 1888 - 0x760  :   32 - 0x20 -- Background 0xec
    "11100110", -- 1889 - 0x761  :  230 - 0xe6
    "01010100", -- 1890 - 0x762  :   84 - 0x54
    "00100110", -- 1891 - 0x763  :   38 - 0x26
    "00100001", -- 1892 - 0x764  :   33 - 0x21
    "00000110", -- 1893 - 0x765  :    6 - 0x6
    "01010100", -- 1894 - 0x766  :   84 - 0x54
    "00100110", -- 1895 - 0x767  :   38 - 0x26
    "00100000", -- 1896 - 0x768  :   32 - 0x20 -- Background 0xed
    "10011010", -- 1897 - 0x769  :  154 - 0x9a
    "00000001", -- 1898 - 0x76a  :    1 - 0x1
    "01001001", -- 1899 - 0x76b  :   73 - 0x49
    "00100000", -- 1900 - 0x76c  :   32 - 0x20
    "10100101", -- 1901 - 0x76d  :  165 - 0xa5
    "11001001", -- 1902 - 0x76e  :  201 - 0xc9
    "01000110", -- 1903 - 0x76f  :   70 - 0x46
    "11010001", -- 1904 - 0x770  :  209 - 0xd1 -- Background 0xee
    "11011000", -- 1905 - 0x771  :  216 - 0xd8
    "11011000", -- 1906 - 0x772  :  216 - 0xd8
    "11011110", -- 1907 - 0x773  :  222 - 0xde
    "11010001", -- 1908 - 0x774  :  209 - 0xd1
    "11010000", -- 1909 - 0x775  :  208 - 0xd0
    "11011010", -- 1910 - 0x776  :  218 - 0xda
    "11011110", -- 1911 - 0x777  :  222 - 0xde
    "11011011", -- 1912 - 0x778  :  219 - 0xdb -- Background 0xef
    "11011001", -- 1913 - 0x779  :  217 - 0xd9
    "11011011", -- 1914 - 0x77a  :  219 - 0xdb
    "11011100", -- 1915 - 0x77b  :  220 - 0xdc
    "11011011", -- 1916 - 0x77c  :  219 - 0xdb
    "11011111", -- 1917 - 0x77d  :  223 - 0xdf
    "00100000", -- 1918 - 0x77e  :   32 - 0x20
    "11100110", -- 1919 - 0x77f  :  230 - 0xe6
    "11011010", -- 1920 - 0x780  :  218 - 0xda -- Background 0xf0
    "11011011", -- 1921 - 0x781  :  219 - 0xdb
    "11100000", -- 1922 - 0x782  :  224 - 0xe0
    "00100001", -- 1923 - 0x783  :   33 - 0x21
    "00000110", -- 1924 - 0x784  :    6 - 0x6
    "00001010", -- 1925 - 0x785  :   10 - 0xa
    "11010110", -- 1926 - 0x786  :  214 - 0xd6
    "11010111", -- 1927 - 0x787  :  215 - 0xd7
    "00100001", -- 1928 - 0x788  :   33 - 0x21 -- Background 0xf1
    "00100110", -- 1929 - 0x789  :   38 - 0x26
    "00010100", -- 1930 - 0x78a  :   20 - 0x14
    "11010000", -- 1931 - 0x78b  :  208 - 0xd0
    "11101000", -- 1932 - 0x78c  :  232 - 0xe8
    "11010001", -- 1933 - 0x78d  :  209 - 0xd1
    "11010000", -- 1934 - 0x78e  :  208 - 0xd0
    "11010001", -- 1935 - 0x78f  :  209 - 0xd1
    "11011110", -- 1936 - 0x790  :  222 - 0xde -- Background 0xf2
    "11010001", -- 1937 - 0x791  :  209 - 0xd1
    "11010000", -- 1938 - 0x792  :  208 - 0xd0
    "11010001", -- 1939 - 0x793  :  209 - 0xd1
    "11010000", -- 1940 - 0x794  :  208 - 0xd0
    "11010001", -- 1941 - 0x795  :  209 - 0xd1
    "00100110", -- 1942 - 0x796  :   38 - 0x26
    "00100001", -- 1943 - 0x797  :   33 - 0x21
    "01000010", -- 1944 - 0x798  :   66 - 0x42 -- Background 0xf3
    "11011011", -- 1945 - 0x799  :  219 - 0xdb
    "11011011", -- 1946 - 0x79a  :  219 - 0xdb
    "01000010", -- 1947 - 0x79b  :   66 - 0x42
    "00100110", -- 1948 - 0x79c  :   38 - 0x26
    "11011011", -- 1949 - 0x79d  :  219 - 0xdb
    "01000010", -- 1950 - 0x79e  :   66 - 0x42
    "11011011", -- 1951 - 0x79f  :  219 - 0xdb
    "01000110", -- 1952 - 0x7a0  :   70 - 0x46 -- Background 0xf4
    "11011011", -- 1953 - 0x7a1  :  219 - 0xdb
    "00100001", -- 1954 - 0x7a2  :   33 - 0x21
    "01101100", -- 1955 - 0x7a3  :  108 - 0x6c
    "00001110", -- 1956 - 0x7a4  :   14 - 0xe
    "11011111", -- 1957 - 0x7a5  :  223 - 0xdf
    "11011011", -- 1958 - 0x7a6  :  219 - 0xdb
    "11011011", -- 1959 - 0x7a7  :  219 - 0xdb
    "11100100", -- 1960 - 0x7a8  :  228 - 0xe4 -- Background 0xf5
    "11100101", -- 1961 - 0x7a9  :  229 - 0xe5
    "00100110", -- 1962 - 0x7aa  :   38 - 0x26
    "00100001", -- 1963 - 0x7ab  :   33 - 0x21
    "10000110", -- 1964 - 0x7ac  :  134 - 0x86
    "00010100", -- 1965 - 0x7ad  :   20 - 0x14
    "11011011", -- 1966 - 0x7ae  :  219 - 0xdb
    "11011011", -- 1967 - 0x7af  :  219 - 0xdb
    "00100110", -- 1968 - 0x7b0  :   38 - 0x26 -- Background 0xf6
    "11011011", -- 1969 - 0x7b1  :  219 - 0xdb
    "11100011", -- 1970 - 0x7b2  :  227 - 0xe3
    "11011011", -- 1971 - 0x7b3  :  219 - 0xdb
    "11100000", -- 1972 - 0x7b4  :  224 - 0xe0
    "11011011", -- 1973 - 0x7b5  :  219 - 0xdb
    "11011011", -- 1974 - 0x7b6  :  219 - 0xdb
    "11100110", -- 1975 - 0x7b7  :  230 - 0xe6
    "11011011", -- 1976 - 0x7b8  :  219 - 0xdb -- Background 0xf7
    "01000010", -- 1977 - 0x7b9  :   66 - 0x42
    "11011011", -- 1978 - 0x7ba  :  219 - 0xdb
    "11011011", -- 1979 - 0x7bb  :  219 - 0xdb
    "11011011", -- 1980 - 0x7bc  :  219 - 0xdb
    "11010100", -- 1981 - 0x7bd  :  212 - 0xd4
    "11011001", -- 1982 - 0x7be  :  217 - 0xd9
    "00100110", -- 1983 - 0x7bf  :   38 - 0x26
    "11100111", -- 1984 - 0x7c0  :  231 - 0xe7 -- Background 0xf8
    "00100001", -- 1985 - 0x7c1  :   33 - 0x21
    "11000101", -- 1986 - 0x7c2  :  197 - 0xc5
    "00010110", -- 1987 - 0x7c3  :   22 - 0x16
    "01011111", -- 1988 - 0x7c4  :   95 - 0x5f
    "10010101", -- 1989 - 0x7c5  :  149 - 0x95
    "10010101", -- 1990 - 0x7c6  :  149 - 0x95
    "10010101", -- 1991 - 0x7c7  :  149 - 0x95
    "10010101", -- 1992 - 0x7c8  :  149 - 0x95 -- Background 0xf9
    "10010110", -- 1993 - 0x7c9  :  150 - 0x96
    "10010101", -- 1994 - 0x7ca  :  149 - 0x95
    "10010101", -- 1995 - 0x7cb  :  149 - 0x95
    "10010111", -- 1996 - 0x7cc  :  151 - 0x97
    "10011000", -- 1997 - 0x7cd  :  152 - 0x98
    "10010111", -- 1998 - 0x7ce  :  151 - 0x97
    "10011000", -- 1999 - 0x7cf  :  152 - 0x98
    "00001000", -- 2000 - 0x7d0  :    8 - 0x8 -- Background 0xfa
    "00000101", -- 2001 - 0x7d1  :    5 - 0x5
    "00100100", -- 2002 - 0x7d2  :   36 - 0x24
    "00010111", -- 2003 - 0x7d3  :   23 - 0x17
    "00010010", -- 2004 - 0x7d4  :   18 - 0x12
    "00010111", -- 2005 - 0x7d5  :   23 - 0x17
    "00011101", -- 2006 - 0x7d6  :   29 - 0x1d
    "00001110", -- 2007 - 0x7d7  :   14 - 0xe
    "00011001", -- 2008 - 0x7d8  :   25 - 0x19 -- Background 0xfb
    "00010101", -- 2009 - 0x7d9  :   21 - 0x15
    "00001010", -- 2010 - 0x7da  :   10 - 0xa
    "00100010", -- 2011 - 0x7db  :   34 - 0x22
    "00001110", -- 2012 - 0x7dc  :   14 - 0xe
    "00011011", -- 2013 - 0x7dd  :   27 - 0x1b
    "00100100", -- 2014 - 0x7de  :   36 - 0x24
    "00010000", -- 2015 - 0x7df  :   16 - 0x10
    "00011001", -- 2016 - 0x7e0  :   25 - 0x19 -- Background 0xfc
    "00010101", -- 2017 - 0x7e1  :   21 - 0x15
    "00001010", -- 2018 - 0x7e2  :   10 - 0xa
    "00100010", -- 2019 - 0x7e3  :   34 - 0x22
    "00001110", -- 2020 - 0x7e4  :   14 - 0xe
    "00011011", -- 2021 - 0x7e5  :   27 - 0x1b
    "00100100", -- 2022 - 0x7e6  :   36 - 0x24
    "00010000", -- 2023 - 0x7e7  :   16 - 0x10
    "00011001", -- 2024 - 0x7e8  :   25 - 0x19 -- Background 0xfd
    "00101000", -- 2025 - 0x7e9  :   40 - 0x28
    "00100010", -- 2026 - 0x7ea  :   34 - 0x22
    "11110110", -- 2027 - 0x7eb  :  246 - 0xf6
    "00000001", -- 2028 - 0x7ec  :    1 - 0x1
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00100011", -- 2030 - 0x7ee  :   35 - 0x23
    "11001001", -- 2031 - 0x7ef  :  201 - 0xc9
    "10101010", -- 2032 - 0x7f0  :  170 - 0xaa -- Background 0xfe
    "00100011", -- 2033 - 0x7f1  :   35 - 0x23
    "11101010", -- 2034 - 0x7f2  :  234 - 0xea
    "00000100", -- 2035 - 0x7f3  :    4 - 0x4
    "10011001", -- 2036 - 0x7f4  :  153 - 0x99
    "10101010", -- 2037 - 0x7f5  :  170 - 0xaa
    "10101010", -- 2038 - 0x7f6  :  170 - 0xaa
    "10101010", -- 2039 - 0x7f7  :  170 - 0xaa
    "11111111", -- 2040 - 0x7f8  :  255 - 0xff -- Background 0xff
    "11111111", -- 2041 - 0x7f9  :  255 - 0xff
    "11111111", -- 2042 - 0x7fa  :  255 - 0xff
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111111", -- 2044 - 0x7fc  :  255 - 0xff
    "11111111", -- 2045 - 0x7fd  :  255 - 0xff
    "11111111", -- 2046 - 0x7fe  :  255 - 0xff
    "11111111"  -- 2047 - 0x7ff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
