//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: pacman_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_PACMAN
  (
     input     clk,   // clock
     input      [13-1:0] addr,  //8192 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Pattern Table 0---------
      13'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      13'h1: dout <= 8'b00000011; //    1 :   3 - 0x3
      13'h2: dout <= 8'b00001111; //    2 :  15 - 0xf
      13'h3: dout <= 8'b00011111; //    3 :  31 - 0x1f
      13'h4: dout <= 8'b00111111; //    4 :  63 - 0x3f
      13'h5: dout <= 8'b00111111; //    5 :  63 - 0x3f
      13'h6: dout <= 8'b01111111; //    6 : 127 - 0x7f
      13'h7: dout <= 8'b01111111; //    7 : 127 - 0x7f
      13'h8: dout <= 8'b00000000; //    8 :   0 - 0x0
      13'h9: dout <= 8'b00000000; //    9 :   0 - 0x0
      13'hA: dout <= 8'b00000000; //   10 :   0 - 0x0
      13'hB: dout <= 8'b00000000; //   11 :   0 - 0x0
      13'hC: dout <= 8'b00000000; //   12 :   0 - 0x0
      13'hD: dout <= 8'b00000000; //   13 :   0 - 0x0
      13'hE: dout <= 8'b00000000; //   14 :   0 - 0x0
      13'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      13'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x1
      13'h11: dout <= 8'b11000000; //   17 : 192 - 0xc0
      13'h12: dout <= 8'b11110000; //   18 : 240 - 0xf0
      13'h13: dout <= 8'b11111000; //   19 : 248 - 0xf8
      13'h14: dout <= 8'b11111000; //   20 : 248 - 0xf8
      13'h15: dout <= 8'b11111100; //   21 : 252 - 0xfc
      13'h16: dout <= 8'b11111100; //   22 : 252 - 0xfc
      13'h17: dout <= 8'b11111100; //   23 : 252 - 0xfc
      13'h18: dout <= 8'b00000000; //   24 :   0 - 0x0
      13'h19: dout <= 8'b00000000; //   25 :   0 - 0x0
      13'h1A: dout <= 8'b00000000; //   26 :   0 - 0x0
      13'h1B: dout <= 8'b00000000; //   27 :   0 - 0x0
      13'h1C: dout <= 8'b00000000; //   28 :   0 - 0x0
      13'h1D: dout <= 8'b00000000; //   29 :   0 - 0x0
      13'h1E: dout <= 8'b00000000; //   30 :   0 - 0x0
      13'h1F: dout <= 8'b00000000; //   31 :   0 - 0x0
      13'h20: dout <= 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x2
      13'h21: dout <= 8'b00000111; //   33 :   7 - 0x7
      13'h22: dout <= 8'b00011111; //   34 :  31 - 0x1f
      13'h23: dout <= 8'b00111111; //   35 :  63 - 0x3f
      13'h24: dout <= 8'b00111111; //   36 :  63 - 0x3f
      13'h25: dout <= 8'b00001111; //   37 :  15 - 0xf
      13'h26: dout <= 8'b00000011; //   38 :   3 - 0x3
      13'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      13'h28: dout <= 8'b00000000; //   40 :   0 - 0x0
      13'h29: dout <= 8'b00000000; //   41 :   0 - 0x0
      13'h2A: dout <= 8'b00000000; //   42 :   0 - 0x0
      13'h2B: dout <= 8'b00000000; //   43 :   0 - 0x0
      13'h2C: dout <= 8'b00000000; //   44 :   0 - 0x0
      13'h2D: dout <= 8'b00000000; //   45 :   0 - 0x0
      13'h2E: dout <= 8'b00000000; //   46 :   0 - 0x0
      13'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      13'h30: dout <= 8'b00000000; //   48 :   0 - 0x0 -- Sprite 0x3
      13'h31: dout <= 8'b00000000; //   49 :   0 - 0x0
      13'h32: dout <= 8'b00000111; //   50 :   7 - 0x7
      13'h33: dout <= 8'b00011111; //   51 :  31 - 0x1f
      13'h34: dout <= 8'b00111111; //   52 :  63 - 0x3f
      13'h35: dout <= 8'b00111111; //   53 :  63 - 0x3f
      13'h36: dout <= 8'b01111111; //   54 : 127 - 0x7f
      13'h37: dout <= 8'b01111111; //   55 : 127 - 0x7f
      13'h38: dout <= 8'b00000000; //   56 :   0 - 0x0
      13'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      13'h3A: dout <= 8'b00000000; //   58 :   0 - 0x0
      13'h3B: dout <= 8'b00000000; //   59 :   0 - 0x0
      13'h3C: dout <= 8'b00000000; //   60 :   0 - 0x0
      13'h3D: dout <= 8'b00000000; //   61 :   0 - 0x0
      13'h3E: dout <= 8'b00000000; //   62 :   0 - 0x0
      13'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      13'h40: dout <= 8'b01111110; //   64 : 126 - 0x7e -- Sprite 0x4
      13'h41: dout <= 8'b01111110; //   65 : 126 - 0x7e
      13'h42: dout <= 8'b01111100; //   66 : 124 - 0x7c
      13'h43: dout <= 8'b00111100; //   67 :  60 - 0x3c
      13'h44: dout <= 8'b00111000; //   68 :  56 - 0x38
      13'h45: dout <= 8'b00011000; //   69 :  24 - 0x18
      13'h46: dout <= 8'b00000000; //   70 :   0 - 0x0
      13'h47: dout <= 8'b00000000; //   71 :   0 - 0x0
      13'h48: dout <= 8'b00000000; //   72 :   0 - 0x0
      13'h49: dout <= 8'b00000000; //   73 :   0 - 0x0
      13'h4A: dout <= 8'b00000000; //   74 :   0 - 0x0
      13'h4B: dout <= 8'b00000000; //   75 :   0 - 0x0
      13'h4C: dout <= 8'b00000000; //   76 :   0 - 0x0
      13'h4D: dout <= 8'b00000000; //   77 :   0 - 0x0
      13'h4E: dout <= 8'b00000000; //   78 :   0 - 0x0
      13'h4F: dout <= 8'b00000000; //   79 :   0 - 0x0
      13'h50: dout <= 8'b00000000; //   80 :   0 - 0x0 -- Sprite 0x5
      13'h51: dout <= 8'b11000000; //   81 : 192 - 0xc0
      13'h52: dout <= 8'b11110000; //   82 : 240 - 0xf0
      13'h53: dout <= 8'b11111000; //   83 : 248 - 0xf8
      13'h54: dout <= 8'b11111000; //   84 : 248 - 0xf8
      13'h55: dout <= 8'b11111100; //   85 : 252 - 0xfc
      13'h56: dout <= 8'b01111100; //   86 : 124 - 0x7c
      13'h57: dout <= 8'b00111100; //   87 :  60 - 0x3c
      13'h58: dout <= 8'b00000000; //   88 :   0 - 0x0
      13'h59: dout <= 8'b00000000; //   89 :   0 - 0x0
      13'h5A: dout <= 8'b00000000; //   90 :   0 - 0x0
      13'h5B: dout <= 8'b00000000; //   91 :   0 - 0x0
      13'h5C: dout <= 8'b00000000; //   92 :   0 - 0x0
      13'h5D: dout <= 8'b00000000; //   93 :   0 - 0x0
      13'h5E: dout <= 8'b00000000; //   94 :   0 - 0x0
      13'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      13'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0x6
      13'h61: dout <= 8'b00000111; //   97 :   7 - 0x7
      13'h62: dout <= 8'b00000111; //   98 :   7 - 0x7
      13'h63: dout <= 8'b00000011; //   99 :   3 - 0x3
      13'h64: dout <= 8'b00000001; //  100 :   1 - 0x1
      13'h65: dout <= 8'b00000000; //  101 :   0 - 0x0
      13'h66: dout <= 8'b00000000; //  102 :   0 - 0x0
      13'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      13'h68: dout <= 8'b00000000; //  104 :   0 - 0x0
      13'h69: dout <= 8'b00000000; //  105 :   0 - 0x0
      13'h6A: dout <= 8'b00000000; //  106 :   0 - 0x0
      13'h6B: dout <= 8'b00000000; //  107 :   0 - 0x0
      13'h6C: dout <= 8'b00000000; //  108 :   0 - 0x0
      13'h6D: dout <= 8'b00000000; //  109 :   0 - 0x0
      13'h6E: dout <= 8'b00000000; //  110 :   0 - 0x0
      13'h6F: dout <= 8'b00000000; //  111 :   0 - 0x0
      13'h70: dout <= 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0x7
      13'h71: dout <= 8'b00000000; //  113 :   0 - 0x0
      13'h72: dout <= 8'b00000111; //  114 :   7 - 0x7
      13'h73: dout <= 8'b00011111; //  115 :  31 - 0x1f
      13'h74: dout <= 8'b00111111; //  116 :  63 - 0x3f
      13'h75: dout <= 8'b00111111; //  117 :  63 - 0x3f
      13'h76: dout <= 8'b01111110; //  118 : 126 - 0x7e
      13'h77: dout <= 8'b01111100; //  119 : 124 - 0x7c
      13'h78: dout <= 8'b00000000; //  120 :   0 - 0x0
      13'h79: dout <= 8'b00000000; //  121 :   0 - 0x0
      13'h7A: dout <= 8'b00000000; //  122 :   0 - 0x0
      13'h7B: dout <= 8'b00000000; //  123 :   0 - 0x0
      13'h7C: dout <= 8'b00000000; //  124 :   0 - 0x0
      13'h7D: dout <= 8'b00000000; //  125 :   0 - 0x0
      13'h7E: dout <= 8'b00000000; //  126 :   0 - 0x0
      13'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      13'h80: dout <= 8'b01111000; //  128 : 120 - 0x78 -- Sprite 0x8
      13'h81: dout <= 8'b01110000; //  129 : 112 - 0x70
      13'h82: dout <= 8'b01100000; //  130 :  96 - 0x60
      13'h83: dout <= 8'b00000000; //  131 :   0 - 0x0
      13'h84: dout <= 8'b00000000; //  132 :   0 - 0x0
      13'h85: dout <= 8'b00000000; //  133 :   0 - 0x0
      13'h86: dout <= 8'b00000000; //  134 :   0 - 0x0
      13'h87: dout <= 8'b00000000; //  135 :   0 - 0x0
      13'h88: dout <= 8'b00000000; //  136 :   0 - 0x0
      13'h89: dout <= 8'b00000000; //  137 :   0 - 0x0
      13'h8A: dout <= 8'b00000000; //  138 :   0 - 0x0
      13'h8B: dout <= 8'b00000000; //  139 :   0 - 0x0
      13'h8C: dout <= 8'b00000000; //  140 :   0 - 0x0
      13'h8D: dout <= 8'b00000000; //  141 :   0 - 0x0
      13'h8E: dout <= 8'b00000000; //  142 :   0 - 0x0
      13'h8F: dout <= 8'b00000000; //  143 :   0 - 0x0
      13'h90: dout <= 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x9
      13'h91: dout <= 8'b00000000; //  145 :   0 - 0x0
      13'h92: dout <= 8'b00000000; //  146 :   0 - 0x0
      13'h93: dout <= 8'b00000000; //  147 :   0 - 0x0
      13'h94: dout <= 8'b00000000; //  148 :   0 - 0x0
      13'h95: dout <= 8'b01000000; //  149 :  64 - 0x40
      13'h96: dout <= 8'b11110000; //  150 : 240 - 0xf0
      13'h97: dout <= 8'b11111000; //  151 : 248 - 0xf8
      13'h98: dout <= 8'b00000000; //  152 :   0 - 0x0
      13'h99: dout <= 8'b00000000; //  153 :   0 - 0x0
      13'h9A: dout <= 8'b00000000; //  154 :   0 - 0x0
      13'h9B: dout <= 8'b00000000; //  155 :   0 - 0x0
      13'h9C: dout <= 8'b00000000; //  156 :   0 - 0x0
      13'h9D: dout <= 8'b00000000; //  157 :   0 - 0x0
      13'h9E: dout <= 8'b00000000; //  158 :   0 - 0x0
      13'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      13'hA0: dout <= 8'b11111110; //  160 : 254 - 0xfe -- Sprite 0xa
      13'hA1: dout <= 8'b01111111; //  161 : 127 - 0x7f
      13'hA2: dout <= 8'b01111111; //  162 : 127 - 0x7f
      13'hA3: dout <= 8'b00111111; //  163 :  63 - 0x3f
      13'hA4: dout <= 8'b00001110; //  164 :  14 - 0xe
      13'hA5: dout <= 8'b00000000; //  165 :   0 - 0x0
      13'hA6: dout <= 8'b00000000; //  166 :   0 - 0x0
      13'hA7: dout <= 8'b00000000; //  167 :   0 - 0x0
      13'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0
      13'hA9: dout <= 8'b00000000; //  169 :   0 - 0x0
      13'hAA: dout <= 8'b00000000; //  170 :   0 - 0x0
      13'hAB: dout <= 8'b00000000; //  171 :   0 - 0x0
      13'hAC: dout <= 8'b00000000; //  172 :   0 - 0x0
      13'hAD: dout <= 8'b00000000; //  173 :   0 - 0x0
      13'hAE: dout <= 8'b00000000; //  174 :   0 - 0x0
      13'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      13'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0xb
      13'hB1: dout <= 8'b00000000; //  177 :   0 - 0x0
      13'hB2: dout <= 8'b00000000; //  178 :   0 - 0x0
      13'hB3: dout <= 8'b00000000; //  179 :   0 - 0x0
      13'hB4: dout <= 8'b00000000; //  180 :   0 - 0x0
      13'hB5: dout <= 8'b00000000; //  181 :   0 - 0x0
      13'hB6: dout <= 8'b00000000; //  182 :   0 - 0x0
      13'hB7: dout <= 8'b11100000; //  183 : 224 - 0xe0
      13'hB8: dout <= 8'b00000000; //  184 :   0 - 0x0
      13'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      13'hBA: dout <= 8'b00000000; //  186 :   0 - 0x0
      13'hBB: dout <= 8'b00000000; //  187 :   0 - 0x0
      13'hBC: dout <= 8'b00000000; //  188 :   0 - 0x0
      13'hBD: dout <= 8'b00000000; //  189 :   0 - 0x0
      13'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      13'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      13'hC0: dout <= 8'b11111100; //  192 : 252 - 0xfc -- Sprite 0xc
      13'hC1: dout <= 8'b11111111; //  193 : 255 - 0xff
      13'hC2: dout <= 8'b01111111; //  194 : 127 - 0x7f
      13'hC3: dout <= 8'b00111111; //  195 :  63 - 0x3f
      13'hC4: dout <= 8'b00001110; //  196 :  14 - 0xe
      13'hC5: dout <= 8'b00000000; //  197 :   0 - 0x0
      13'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      13'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      13'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0
      13'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      13'hCA: dout <= 8'b00000000; //  202 :   0 - 0x0
      13'hCB: dout <= 8'b00000000; //  203 :   0 - 0x0
      13'hCC: dout <= 8'b00000000; //  204 :   0 - 0x0
      13'hCD: dout <= 8'b00000000; //  205 :   0 - 0x0
      13'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      13'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      13'hD0: dout <= 8'b11110000; //  208 : 240 - 0xf0 -- Sprite 0xd
      13'hD1: dout <= 8'b11111111; //  209 : 255 - 0xff
      13'hD2: dout <= 8'b11111111; //  210 : 255 - 0xff
      13'hD3: dout <= 8'b01111111; //  211 : 127 - 0x7f
      13'hD4: dout <= 8'b00011110; //  212 :  30 - 0x1e
      13'hD5: dout <= 8'b00000000; //  213 :   0 - 0x0
      13'hD6: dout <= 8'b00000000; //  214 :   0 - 0x0
      13'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      13'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0
      13'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      13'hDA: dout <= 8'b00000000; //  218 :   0 - 0x0
      13'hDB: dout <= 8'b00000000; //  219 :   0 - 0x0
      13'hDC: dout <= 8'b00000000; //  220 :   0 - 0x0
      13'hDD: dout <= 8'b00000000; //  221 :   0 - 0x0
      13'hDE: dout <= 8'b00000000; //  222 :   0 - 0x0
      13'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      13'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0xe
      13'hE1: dout <= 8'b00001111; //  225 :  15 - 0xf
      13'hE2: dout <= 8'b11111111; //  226 : 255 - 0xff
      13'hE3: dout <= 8'b11111111; //  227 : 255 - 0xff
      13'hE4: dout <= 8'b01111111; //  228 : 127 - 0x7f
      13'hE5: dout <= 8'b00011110; //  229 :  30 - 0x1e
      13'hE6: dout <= 8'b00000000; //  230 :   0 - 0x0
      13'hE7: dout <= 8'b00000000; //  231 :   0 - 0x0
      13'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0
      13'hE9: dout <= 8'b00000000; //  233 :   0 - 0x0
      13'hEA: dout <= 8'b00000000; //  234 :   0 - 0x0
      13'hEB: dout <= 8'b00000000; //  235 :   0 - 0x0
      13'hEC: dout <= 8'b00000000; //  236 :   0 - 0x0
      13'hED: dout <= 8'b00000000; //  237 :   0 - 0x0
      13'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      13'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      13'hF0: dout <= 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0xf
      13'hF1: dout <= 8'b00000011; //  241 :   3 - 0x3
      13'hF2: dout <= 8'b00001111; //  242 :  15 - 0xf
      13'hF3: dout <= 8'b01111111; //  243 : 127 - 0x7f
      13'hF4: dout <= 8'b11111111; //  244 : 255 - 0xff
      13'hF5: dout <= 8'b01111110; //  245 : 126 - 0x7e
      13'hF6: dout <= 8'b00011100; //  246 :  28 - 0x1c
      13'hF7: dout <= 8'b00000000; //  247 :   0 - 0x0
      13'hF8: dout <= 8'b00000000; //  248 :   0 - 0x0
      13'hF9: dout <= 8'b00000000; //  249 :   0 - 0x0
      13'hFA: dout <= 8'b00000000; //  250 :   0 - 0x0
      13'hFB: dout <= 8'b00000000; //  251 :   0 - 0x0
      13'hFC: dout <= 8'b00000000; //  252 :   0 - 0x0
      13'hFD: dout <= 8'b00000000; //  253 :   0 - 0x0
      13'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      13'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      13'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x10
      13'h101: dout <= 8'b00000001; //  257 :   1 - 0x1
      13'h102: dout <= 8'b00000011; //  258 :   3 - 0x3
      13'h103: dout <= 8'b00001111; //  259 :  15 - 0xf
      13'h104: dout <= 8'b00011111; //  260 :  31 - 0x1f
      13'h105: dout <= 8'b01111111; //  261 : 127 - 0x7f
      13'h106: dout <= 8'b01111110; //  262 : 126 - 0x7e
      13'h107: dout <= 8'b00111100; //  263 :  60 - 0x3c
      13'h108: dout <= 8'b00000000; //  264 :   0 - 0x0
      13'h109: dout <= 8'b00000000; //  265 :   0 - 0x0
      13'h10A: dout <= 8'b00000000; //  266 :   0 - 0x0
      13'h10B: dout <= 8'b00000000; //  267 :   0 - 0x0
      13'h10C: dout <= 8'b00000000; //  268 :   0 - 0x0
      13'h10D: dout <= 8'b00000000; //  269 :   0 - 0x0
      13'h10E: dout <= 8'b00000000; //  270 :   0 - 0x0
      13'h10F: dout <= 8'b00000000; //  271 :   0 - 0x0
      13'h110: dout <= 8'b00000000; //  272 :   0 - 0x0 -- Sprite 0x11
      13'h111: dout <= 8'b00000001; //  273 :   1 - 0x1
      13'h112: dout <= 8'b00000011; //  274 :   3 - 0x3
      13'h113: dout <= 8'b00000111; //  275 :   7 - 0x7
      13'h114: dout <= 8'b00000111; //  276 :   7 - 0x7
      13'h115: dout <= 8'b00001111; //  277 :  15 - 0xf
      13'h116: dout <= 8'b00011111; //  278 :  31 - 0x1f
      13'h117: dout <= 8'b00001110; //  279 :  14 - 0xe
      13'h118: dout <= 8'b00000000; //  280 :   0 - 0x0
      13'h119: dout <= 8'b00000000; //  281 :   0 - 0x0
      13'h11A: dout <= 8'b00000000; //  282 :   0 - 0x0
      13'h11B: dout <= 8'b00000000; //  283 :   0 - 0x0
      13'h11C: dout <= 8'b00000000; //  284 :   0 - 0x0
      13'h11D: dout <= 8'b00000000; //  285 :   0 - 0x0
      13'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      13'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      13'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x12
      13'h121: dout <= 8'b00000000; //  289 :   0 - 0x0
      13'h122: dout <= 8'b00000001; //  290 :   1 - 0x1
      13'h123: dout <= 8'b00000011; //  291 :   3 - 0x3
      13'h124: dout <= 8'b00000011; //  292 :   3 - 0x3
      13'h125: dout <= 8'b00000011; //  293 :   3 - 0x3
      13'h126: dout <= 8'b00000111; //  294 :   7 - 0x7
      13'h127: dout <= 8'b00000010; //  295 :   2 - 0x2
      13'h128: dout <= 8'b00000000; //  296 :   0 - 0x0
      13'h129: dout <= 8'b00000000; //  297 :   0 - 0x0
      13'h12A: dout <= 8'b00000000; //  298 :   0 - 0x0
      13'h12B: dout <= 8'b00000000; //  299 :   0 - 0x0
      13'h12C: dout <= 8'b00000000; //  300 :   0 - 0x0
      13'h12D: dout <= 8'b00000000; //  301 :   0 - 0x0
      13'h12E: dout <= 8'b00000000; //  302 :   0 - 0x0
      13'h12F: dout <= 8'b00000000; //  303 :   0 - 0x0
      13'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x13
      13'h131: dout <= 8'b00000000; //  305 :   0 - 0x0
      13'h132: dout <= 8'b00000001; //  306 :   1 - 0x1
      13'h133: dout <= 8'b00000001; //  307 :   1 - 0x1
      13'h134: dout <= 8'b00000001; //  308 :   1 - 0x1
      13'h135: dout <= 8'b00000001; //  309 :   1 - 0x1
      13'h136: dout <= 8'b00000001; //  310 :   1 - 0x1
      13'h137: dout <= 8'b00000001; //  311 :   1 - 0x1
      13'h138: dout <= 8'b00000000; //  312 :   0 - 0x0
      13'h139: dout <= 8'b00000000; //  313 :   0 - 0x0
      13'h13A: dout <= 8'b00000000; //  314 :   0 - 0x0
      13'h13B: dout <= 8'b00000000; //  315 :   0 - 0x0
      13'h13C: dout <= 8'b00000000; //  316 :   0 - 0x0
      13'h13D: dout <= 8'b00000000; //  317 :   0 - 0x0
      13'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      13'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      13'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x14
      13'h141: dout <= 8'b00000000; //  321 :   0 - 0x0
      13'h142: dout <= 8'b00000000; //  322 :   0 - 0x0
      13'h143: dout <= 8'b00000000; //  323 :   0 - 0x0
      13'h144: dout <= 8'b00000000; //  324 :   0 - 0x0
      13'h145: dout <= 8'b00000000; //  325 :   0 - 0x0
      13'h146: dout <= 8'b00000100; //  326 :   4 - 0x4
      13'h147: dout <= 8'b00000010; //  327 :   2 - 0x2
      13'h148: dout <= 8'b00000000; //  328 :   0 - 0x0
      13'h149: dout <= 8'b00000000; //  329 :   0 - 0x0
      13'h14A: dout <= 8'b00000000; //  330 :   0 - 0x0
      13'h14B: dout <= 8'b00000000; //  331 :   0 - 0x0
      13'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      13'h14D: dout <= 8'b00000000; //  333 :   0 - 0x0
      13'h14E: dout <= 8'b00000000; //  334 :   0 - 0x0
      13'h14F: dout <= 8'b00000000; //  335 :   0 - 0x0
      13'h150: dout <= 8'b00000000; //  336 :   0 - 0x0 -- Sprite 0x15
      13'h151: dout <= 8'b00000000; //  337 :   0 - 0x0
      13'h152: dout <= 8'b00000000; //  338 :   0 - 0x0
      13'h153: dout <= 8'b00000000; //  339 :   0 - 0x0
      13'h154: dout <= 8'b00000000; //  340 :   0 - 0x0
      13'h155: dout <= 8'b00000000; //  341 :   0 - 0x0
      13'h156: dout <= 8'b00100000; //  342 :  32 - 0x20
      13'h157: dout <= 8'b01001000; //  343 :  72 - 0x48
      13'h158: dout <= 8'b00000000; //  344 :   0 - 0x0
      13'h159: dout <= 8'b00000000; //  345 :   0 - 0x0
      13'h15A: dout <= 8'b00000000; //  346 :   0 - 0x0
      13'h15B: dout <= 8'b00000000; //  347 :   0 - 0x0
      13'h15C: dout <= 8'b00000000; //  348 :   0 - 0x0
      13'h15D: dout <= 8'b00000000; //  349 :   0 - 0x0
      13'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      13'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      13'h160: dout <= 8'b00010000; //  352 :  16 - 0x10 -- Sprite 0x16
      13'h161: dout <= 8'b00001000; //  353 :   8 - 0x8
      13'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      13'h163: dout <= 8'b00110000; //  355 :  48 - 0x30
      13'h164: dout <= 8'b00000000; //  356 :   0 - 0x0
      13'h165: dout <= 8'b00001000; //  357 :   8 - 0x8
      13'h166: dout <= 8'b00010010; //  358 :  18 - 0x12
      13'h167: dout <= 8'b00000100; //  359 :   4 - 0x4
      13'h168: dout <= 8'b00000000; //  360 :   0 - 0x0
      13'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      13'h16A: dout <= 8'b00000000; //  362 :   0 - 0x0
      13'h16B: dout <= 8'b00000000; //  363 :   0 - 0x0
      13'h16C: dout <= 8'b00000000; //  364 :   0 - 0x0
      13'h16D: dout <= 8'b00000000; //  365 :   0 - 0x0
      13'h16E: dout <= 8'b00000000; //  366 :   0 - 0x0
      13'h16F: dout <= 8'b00000000; //  367 :   0 - 0x0
      13'h170: dout <= 8'b00010000; //  368 :  16 - 0x10 -- Sprite 0x17
      13'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      13'h172: dout <= 8'b00001100; //  370 :  12 - 0xc
      13'h173: dout <= 8'b00000000; //  371 :   0 - 0x0
      13'h174: dout <= 8'b00010000; //  372 :  16 - 0x10
      13'h175: dout <= 8'b00001000; //  373 :   8 - 0x8
      13'h176: dout <= 8'b01000000; //  374 :  64 - 0x40
      13'h177: dout <= 8'b00100000; //  375 :  32 - 0x20
      13'h178: dout <= 8'b00000000; //  376 :   0 - 0x0
      13'h179: dout <= 8'b00000000; //  377 :   0 - 0x0
      13'h17A: dout <= 8'b00000000; //  378 :   0 - 0x0
      13'h17B: dout <= 8'b00000000; //  379 :   0 - 0x0
      13'h17C: dout <= 8'b00000000; //  380 :   0 - 0x0
      13'h17D: dout <= 8'b00000000; //  381 :   0 - 0x0
      13'h17E: dout <= 8'b00000000; //  382 :   0 - 0x0
      13'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      13'h180: dout <= 8'b00000000; //  384 :   0 - 0x0 -- Sprite 0x18
      13'h181: dout <= 8'b00000000; //  385 :   0 - 0x0
      13'h182: dout <= 8'b00000011; //  386 :   3 - 0x3
      13'h183: dout <= 8'b00000011; //  387 :   3 - 0x3
      13'h184: dout <= 8'b00000001; //  388 :   1 - 0x1
      13'h185: dout <= 8'b00100001; //  389 :  33 - 0x21
      13'h186: dout <= 8'b00100001; //  390 :  33 - 0x21
      13'h187: dout <= 8'b01110011; //  391 : 115 - 0x73
      13'h188: dout <= 8'b00000000; //  392 :   0 - 0x0
      13'h189: dout <= 8'b00000000; //  393 :   0 - 0x0
      13'h18A: dout <= 8'b00000011; //  394 :   3 - 0x3
      13'h18B: dout <= 8'b00000011; //  395 :   3 - 0x3
      13'h18C: dout <= 8'b00010011; //  396 :  19 - 0x13
      13'h18D: dout <= 8'b00111111; //  397 :  63 - 0x3f
      13'h18E: dout <= 8'b00111111; //  398 :  63 - 0x3f
      13'h18F: dout <= 8'b01111111; //  399 : 127 - 0x7f
      13'h190: dout <= 8'b01111111; //  400 : 127 - 0x7f -- Sprite 0x19
      13'h191: dout <= 8'b01111111; //  401 : 127 - 0x7f
      13'h192: dout <= 8'b01111111; //  402 : 127 - 0x7f
      13'h193: dout <= 8'b01111111; //  403 : 127 - 0x7f
      13'h194: dout <= 8'b01101110; //  404 : 110 - 0x6e
      13'h195: dout <= 8'b01000110; //  405 :  70 - 0x46
      13'h196: dout <= 8'b00000000; //  406 :   0 - 0x0
      13'h197: dout <= 8'b00000000; //  407 :   0 - 0x0
      13'h198: dout <= 8'b01111111; //  408 : 127 - 0x7f
      13'h199: dout <= 8'b01111111; //  409 : 127 - 0x7f
      13'h19A: dout <= 8'b01111111; //  410 : 127 - 0x7f
      13'h19B: dout <= 8'b01111111; //  411 : 127 - 0x7f
      13'h19C: dout <= 8'b01101110; //  412 : 110 - 0x6e
      13'h19D: dout <= 8'b01000110; //  413 :  70 - 0x46
      13'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      13'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      13'h1A0: dout <= 8'b01111111; //  416 : 127 - 0x7f -- Sprite 0x1a
      13'h1A1: dout <= 8'b01111111; //  417 : 127 - 0x7f
      13'h1A2: dout <= 8'b01111111; //  418 : 127 - 0x7f
      13'h1A3: dout <= 8'b01111111; //  419 : 127 - 0x7f
      13'h1A4: dout <= 8'b01111011; //  420 : 123 - 0x7b
      13'h1A5: dout <= 8'b00110001; //  421 :  49 - 0x31
      13'h1A6: dout <= 8'b00000000; //  422 :   0 - 0x0
      13'h1A7: dout <= 8'b00000000; //  423 :   0 - 0x0
      13'h1A8: dout <= 8'b01111111; //  424 : 127 - 0x7f
      13'h1A9: dout <= 8'b01111111; //  425 : 127 - 0x7f
      13'h1AA: dout <= 8'b01111111; //  426 : 127 - 0x7f
      13'h1AB: dout <= 8'b01111111; //  427 : 127 - 0x7f
      13'h1AC: dout <= 8'b01111011; //  428 : 123 - 0x7b
      13'h1AD: dout <= 8'b00110001; //  429 :  49 - 0x31
      13'h1AE: dout <= 8'b00000000; //  430 :   0 - 0x0
      13'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      13'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x1b
      13'h1B1: dout <= 8'b00000011; //  433 :   3 - 0x3
      13'h1B2: dout <= 8'b00001111; //  434 :  15 - 0xf
      13'h1B3: dout <= 8'b00011111; //  435 :  31 - 0x1f
      13'h1B4: dout <= 8'b00100111; //  436 :  39 - 0x27
      13'h1B5: dout <= 8'b00000011; //  437 :   3 - 0x3
      13'h1B6: dout <= 8'b00000011; //  438 :   3 - 0x3
      13'h1B7: dout <= 8'b01000011; //  439 :  67 - 0x43
      13'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0
      13'h1B9: dout <= 8'b00000011; //  441 :   3 - 0x3
      13'h1BA: dout <= 8'b00001111; //  442 :  15 - 0xf
      13'h1BB: dout <= 8'b00011111; //  443 :  31 - 0x1f
      13'h1BC: dout <= 8'b00111111; //  444 :  63 - 0x3f
      13'h1BD: dout <= 8'b00111111; //  445 :  63 - 0x3f
      13'h1BE: dout <= 8'b00001111; //  446 :  15 - 0xf
      13'h1BF: dout <= 8'b01001111; //  447 :  79 - 0x4f
      13'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x1c
      13'h1C1: dout <= 8'b11000000; //  449 : 192 - 0xc0
      13'h1C2: dout <= 8'b11110000; //  450 : 240 - 0xf0
      13'h1C3: dout <= 8'b11111000; //  451 : 248 - 0xf8
      13'h1C4: dout <= 8'b10011100; //  452 : 156 - 0x9c
      13'h1C5: dout <= 8'b00001100; //  453 :  12 - 0xc
      13'h1C6: dout <= 8'b00001100; //  454 :  12 - 0xc
      13'h1C7: dout <= 8'b00001110; //  455 :  14 - 0xe
      13'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0
      13'h1C9: dout <= 8'b11000000; //  457 : 192 - 0xc0
      13'h1CA: dout <= 8'b11110000; //  458 : 240 - 0xf0
      13'h1CB: dout <= 8'b11111000; //  459 : 248 - 0xf8
      13'h1CC: dout <= 8'b11111100; //  460 : 252 - 0xfc
      13'h1CD: dout <= 8'b11111100; //  461 : 252 - 0xfc
      13'h1CE: dout <= 8'b00111100; //  462 :  60 - 0x3c
      13'h1CF: dout <= 8'b00111110; //  463 :  62 - 0x3e
      13'h1D0: dout <= 8'b01100111; //  464 : 103 - 0x67 -- Sprite 0x1d
      13'h1D1: dout <= 8'b01111111; //  465 : 127 - 0x7f
      13'h1D2: dout <= 8'b01111111; //  466 : 127 - 0x7f
      13'h1D3: dout <= 8'b01111111; //  467 : 127 - 0x7f
      13'h1D4: dout <= 8'b01101110; //  468 : 110 - 0x6e
      13'h1D5: dout <= 8'b01000110; //  469 :  70 - 0x46
      13'h1D6: dout <= 8'b00000000; //  470 :   0 - 0x0
      13'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      13'h1D8: dout <= 8'b01111111; //  472 : 127 - 0x7f
      13'h1D9: dout <= 8'b01111111; //  473 : 127 - 0x7f
      13'h1DA: dout <= 8'b01111111; //  474 : 127 - 0x7f
      13'h1DB: dout <= 8'b01111111; //  475 : 127 - 0x7f
      13'h1DC: dout <= 8'b01101110; //  476 : 110 - 0x6e
      13'h1DD: dout <= 8'b01000110; //  477 :  70 - 0x46
      13'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      13'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      13'h1E0: dout <= 8'b01100111; //  480 : 103 - 0x67 -- Sprite 0x1e
      13'h1E1: dout <= 8'b01111111; //  481 : 127 - 0x7f
      13'h1E2: dout <= 8'b01111111; //  482 : 127 - 0x7f
      13'h1E3: dout <= 8'b01111111; //  483 : 127 - 0x7f
      13'h1E4: dout <= 8'b01111011; //  484 : 123 - 0x7b
      13'h1E5: dout <= 8'b00110001; //  485 :  49 - 0x31
      13'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      13'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      13'h1E8: dout <= 8'b01111111; //  488 : 127 - 0x7f
      13'h1E9: dout <= 8'b01111111; //  489 : 127 - 0x7f
      13'h1EA: dout <= 8'b01111111; //  490 : 127 - 0x7f
      13'h1EB: dout <= 8'b01111111; //  491 : 127 - 0x7f
      13'h1EC: dout <= 8'b01111011; //  492 : 123 - 0x7b
      13'h1ED: dout <= 8'b00110001; //  493 :  49 - 0x31
      13'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      13'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      13'h1F0: dout <= 8'b10011110; //  496 : 158 - 0x9e -- Sprite 0x1f
      13'h1F1: dout <= 8'b11111110; //  497 : 254 - 0xfe
      13'h1F2: dout <= 8'b11111110; //  498 : 254 - 0xfe
      13'h1F3: dout <= 8'b11111110; //  499 : 254 - 0xfe
      13'h1F4: dout <= 8'b01110110; //  500 : 118 - 0x76
      13'h1F5: dout <= 8'b01100010; //  501 :  98 - 0x62
      13'h1F6: dout <= 8'b00000000; //  502 :   0 - 0x0
      13'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      13'h1F8: dout <= 8'b11111110; //  504 : 254 - 0xfe
      13'h1F9: dout <= 8'b11111110; //  505 : 254 - 0xfe
      13'h1FA: dout <= 8'b11111110; //  506 : 254 - 0xfe
      13'h1FB: dout <= 8'b11111110; //  507 : 254 - 0xfe
      13'h1FC: dout <= 8'b01110110; //  508 : 118 - 0x76
      13'h1FD: dout <= 8'b01100010; //  509 :  98 - 0x62
      13'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      13'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      13'h200: dout <= 8'b10011110; //  512 : 158 - 0x9e -- Sprite 0x20
      13'h201: dout <= 8'b11111110; //  513 : 254 - 0xfe
      13'h202: dout <= 8'b11111110; //  514 : 254 - 0xfe
      13'h203: dout <= 8'b11111110; //  515 : 254 - 0xfe
      13'h204: dout <= 8'b11011110; //  516 : 222 - 0xde
      13'h205: dout <= 8'b10001100; //  517 : 140 - 0x8c
      13'h206: dout <= 8'b00000000; //  518 :   0 - 0x0
      13'h207: dout <= 8'b00000000; //  519 :   0 - 0x0
      13'h208: dout <= 8'b11111110; //  520 : 254 - 0xfe
      13'h209: dout <= 8'b11111110; //  521 : 254 - 0xfe
      13'h20A: dout <= 8'b11111110; //  522 : 254 - 0xfe
      13'h20B: dout <= 8'b11111110; //  523 : 254 - 0xfe
      13'h20C: dout <= 8'b11011110; //  524 : 222 - 0xde
      13'h20D: dout <= 8'b10001100; //  525 : 140 - 0x8c
      13'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      13'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      13'h210: dout <= 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x21
      13'h211: dout <= 8'b00000011; //  529 :   3 - 0x3
      13'h212: dout <= 8'b00001111; //  530 :  15 - 0xf
      13'h213: dout <= 8'b00011111; //  531 :  31 - 0x1f
      13'h214: dout <= 8'b00111111; //  532 :  63 - 0x3f
      13'h215: dout <= 8'b00110011; //  533 :  51 - 0x33
      13'h216: dout <= 8'b00100001; //  534 :  33 - 0x21
      13'h217: dout <= 8'b01100001; //  535 :  97 - 0x61
      13'h218: dout <= 8'b00000000; //  536 :   0 - 0x0
      13'h219: dout <= 8'b00000011; //  537 :   3 - 0x3
      13'h21A: dout <= 8'b00001111; //  538 :  15 - 0xf
      13'h21B: dout <= 8'b00011111; //  539 :  31 - 0x1f
      13'h21C: dout <= 8'b00111111; //  540 :  63 - 0x3f
      13'h21D: dout <= 8'b00111111; //  541 :  63 - 0x3f
      13'h21E: dout <= 8'b00111111; //  542 :  63 - 0x3f
      13'h21F: dout <= 8'b01111111; //  543 : 127 - 0x7f
      13'h220: dout <= 8'b01100001; //  544 :  97 - 0x61 -- Sprite 0x22
      13'h221: dout <= 8'b01110011; //  545 : 115 - 0x73
      13'h222: dout <= 8'b01111111; //  546 : 127 - 0x7f
      13'h223: dout <= 8'b01111111; //  547 : 127 - 0x7f
      13'h224: dout <= 8'b01101110; //  548 : 110 - 0x6e
      13'h225: dout <= 8'b01000110; //  549 :  70 - 0x46
      13'h226: dout <= 8'b00000000; //  550 :   0 - 0x0
      13'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      13'h228: dout <= 8'b01110011; //  552 : 115 - 0x73
      13'h229: dout <= 8'b01110011; //  553 : 115 - 0x73
      13'h22A: dout <= 8'b01111111; //  554 : 127 - 0x7f
      13'h22B: dout <= 8'b01111111; //  555 : 127 - 0x7f
      13'h22C: dout <= 8'b01101110; //  556 : 110 - 0x6e
      13'h22D: dout <= 8'b01000110; //  557 :  70 - 0x46
      13'h22E: dout <= 8'b00000000; //  558 :   0 - 0x0
      13'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      13'h230: dout <= 8'b01100001; //  560 :  97 - 0x61 -- Sprite 0x23
      13'h231: dout <= 8'b01110011; //  561 : 115 - 0x73
      13'h232: dout <= 8'b01111111; //  562 : 127 - 0x7f
      13'h233: dout <= 8'b01111111; //  563 : 127 - 0x7f
      13'h234: dout <= 8'b01110111; //  564 : 119 - 0x77
      13'h235: dout <= 8'b00100011; //  565 :  35 - 0x23
      13'h236: dout <= 8'b00000000; //  566 :   0 - 0x0
      13'h237: dout <= 8'b00000000; //  567 :   0 - 0x0
      13'h238: dout <= 8'b01110011; //  568 : 115 - 0x73
      13'h239: dout <= 8'b01110011; //  569 : 115 - 0x73
      13'h23A: dout <= 8'b01111111; //  570 : 127 - 0x7f
      13'h23B: dout <= 8'b01111111; //  571 : 127 - 0x7f
      13'h23C: dout <= 8'b01110111; //  572 : 119 - 0x77
      13'h23D: dout <= 8'b00100011; //  573 :  35 - 0x23
      13'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      13'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      13'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x24
      13'h241: dout <= 8'b00000011; //  577 :   3 - 0x3
      13'h242: dout <= 8'b00001111; //  578 :  15 - 0xf
      13'h243: dout <= 8'b00011111; //  579 :  31 - 0x1f
      13'h244: dout <= 8'b00111111; //  580 :  63 - 0x3f
      13'h245: dout <= 8'b00111111; //  581 :  63 - 0x3f
      13'h246: dout <= 8'b00111111; //  582 :  63 - 0x3f
      13'h247: dout <= 8'b01111111; //  583 : 127 - 0x7f
      13'h248: dout <= 8'b00000000; //  584 :   0 - 0x0
      13'h249: dout <= 8'b00000000; //  585 :   0 - 0x0
      13'h24A: dout <= 8'b00000000; //  586 :   0 - 0x0
      13'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      13'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      13'h24D: dout <= 8'b00000110; //  589 :   6 - 0x6
      13'h24E: dout <= 8'b00000110; //  590 :   6 - 0x6
      13'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      13'h250: dout <= 8'b01111111; //  592 : 127 - 0x7f -- Sprite 0x25
      13'h251: dout <= 8'b01111111; //  593 : 127 - 0x7f
      13'h252: dout <= 8'b01111111; //  594 : 127 - 0x7f
      13'h253: dout <= 8'b01111111; //  595 : 127 - 0x7f
      13'h254: dout <= 8'b01101110; //  596 : 110 - 0x6e
      13'h255: dout <= 8'b01000110; //  597 :  70 - 0x46
      13'h256: dout <= 8'b00000000; //  598 :   0 - 0x0
      13'h257: dout <= 8'b00000000; //  599 :   0 - 0x0
      13'h258: dout <= 8'b00000000; //  600 :   0 - 0x0
      13'h259: dout <= 8'b00011001; //  601 :  25 - 0x19
      13'h25A: dout <= 8'b00100110; //  602 :  38 - 0x26
      13'h25B: dout <= 8'b00000000; //  603 :   0 - 0x0
      13'h25C: dout <= 8'b00000000; //  604 :   0 - 0x0
      13'h25D: dout <= 8'b00000000; //  605 :   0 - 0x0
      13'h25E: dout <= 8'b00000000; //  606 :   0 - 0x0
      13'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      13'h260: dout <= 8'b01111111; //  608 : 127 - 0x7f -- Sprite 0x26
      13'h261: dout <= 8'b01111111; //  609 : 127 - 0x7f
      13'h262: dout <= 8'b01111111; //  610 : 127 - 0x7f
      13'h263: dout <= 8'b01111111; //  611 : 127 - 0x7f
      13'h264: dout <= 8'b01111011; //  612 : 123 - 0x7b
      13'h265: dout <= 8'b00110001; //  613 :  49 - 0x31
      13'h266: dout <= 8'b00000000; //  614 :   0 - 0x0
      13'h267: dout <= 8'b00000000; //  615 :   0 - 0x0
      13'h268: dout <= 8'b00000000; //  616 :   0 - 0x0
      13'h269: dout <= 8'b00011001; //  617 :  25 - 0x19
      13'h26A: dout <= 8'b00100110; //  618 :  38 - 0x26
      13'h26B: dout <= 8'b00000000; //  619 :   0 - 0x0
      13'h26C: dout <= 8'b00000000; //  620 :   0 - 0x0
      13'h26D: dout <= 8'b00000000; //  621 :   0 - 0x0
      13'h26E: dout <= 8'b00000000; //  622 :   0 - 0x0
      13'h26F: dout <= 8'b00000000; //  623 :   0 - 0x0
      13'h270: dout <= 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x27
      13'h271: dout <= 8'b00000000; //  625 :   0 - 0x0
      13'h272: dout <= 8'b00000000; //  626 :   0 - 0x0
      13'h273: dout <= 8'b00000000; //  627 :   0 - 0x0
      13'h274: dout <= 8'b00000000; //  628 :   0 - 0x0
      13'h275: dout <= 8'b00000000; //  629 :   0 - 0x0
      13'h276: dout <= 8'b00000000; //  630 :   0 - 0x0
      13'h277: dout <= 8'b00000000; //  631 :   0 - 0x0
      13'h278: dout <= 8'b00000000; //  632 :   0 - 0x0
      13'h279: dout <= 8'b00001100; //  633 :  12 - 0xc
      13'h27A: dout <= 8'b00010010; //  634 :  18 - 0x12
      13'h27B: dout <= 8'b00010010; //  635 :  18 - 0x12
      13'h27C: dout <= 8'b00011110; //  636 :  30 - 0x1e
      13'h27D: dout <= 8'b00001100; //  637 :  12 - 0xc
      13'h27E: dout <= 8'b00000000; //  638 :   0 - 0x0
      13'h27F: dout <= 8'b00000000; //  639 :   0 - 0x0
      13'h280: dout <= 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x28
      13'h281: dout <= 8'b00000000; //  641 :   0 - 0x0
      13'h282: dout <= 8'b00000000; //  642 :   0 - 0x0
      13'h283: dout <= 8'b00000000; //  643 :   0 - 0x0
      13'h284: dout <= 8'b00000000; //  644 :   0 - 0x0
      13'h285: dout <= 8'b00000000; //  645 :   0 - 0x0
      13'h286: dout <= 8'b00000000; //  646 :   0 - 0x0
      13'h287: dout <= 8'b00000000; //  647 :   0 - 0x0
      13'h288: dout <= 8'b00000000; //  648 :   0 - 0x0
      13'h289: dout <= 8'b00000000; //  649 :   0 - 0x0
      13'h28A: dout <= 8'b00000000; //  650 :   0 - 0x0
      13'h28B: dout <= 8'b00000000; //  651 :   0 - 0x0
      13'h28C: dout <= 8'b00000000; //  652 :   0 - 0x0
      13'h28D: dout <= 8'b00111000; //  653 :  56 - 0x38
      13'h28E: dout <= 8'b01001101; //  654 :  77 - 0x4d
      13'h28F: dout <= 8'b01001101; //  655 :  77 - 0x4d
      13'h290: dout <= 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x29
      13'h291: dout <= 8'b00000000; //  657 :   0 - 0x0
      13'h292: dout <= 8'b00000000; //  658 :   0 - 0x0
      13'h293: dout <= 8'b00000000; //  659 :   0 - 0x0
      13'h294: dout <= 8'b00000000; //  660 :   0 - 0x0
      13'h295: dout <= 8'b00000000; //  661 :   0 - 0x0
      13'h296: dout <= 8'b00000000; //  662 :   0 - 0x0
      13'h297: dout <= 8'b00000000; //  663 :   0 - 0x0
      13'h298: dout <= 8'b00000000; //  664 :   0 - 0x0
      13'h299: dout <= 8'b00000000; //  665 :   0 - 0x0
      13'h29A: dout <= 8'b00000000; //  666 :   0 - 0x0
      13'h29B: dout <= 8'b00000000; //  667 :   0 - 0x0
      13'h29C: dout <= 8'b00000000; //  668 :   0 - 0x0
      13'h29D: dout <= 8'b11100000; //  669 : 224 - 0xe0
      13'h29E: dout <= 8'b00110000; //  670 :  48 - 0x30
      13'h29F: dout <= 8'b00110000; //  671 :  48 - 0x30
      13'h2A0: dout <= 8'b00000000; //  672 :   0 - 0x0 -- Sprite 0x2a
      13'h2A1: dout <= 8'b00000000; //  673 :   0 - 0x0
      13'h2A2: dout <= 8'b00000000; //  674 :   0 - 0x0
      13'h2A3: dout <= 8'b00000000; //  675 :   0 - 0x0
      13'h2A4: dout <= 8'b00000000; //  676 :   0 - 0x0
      13'h2A5: dout <= 8'b00000000; //  677 :   0 - 0x0
      13'h2A6: dout <= 8'b00000000; //  678 :   0 - 0x0
      13'h2A7: dout <= 8'b00000000; //  679 :   0 - 0x0
      13'h2A8: dout <= 8'b00111000; //  680 :  56 - 0x38
      13'h2A9: dout <= 8'b00000000; //  681 :   0 - 0x0
      13'h2AA: dout <= 8'b00000000; //  682 :   0 - 0x0
      13'h2AB: dout <= 8'b00000000; //  683 :   0 - 0x0
      13'h2AC: dout <= 8'b00000000; //  684 :   0 - 0x0
      13'h2AD: dout <= 8'b00000000; //  685 :   0 - 0x0
      13'h2AE: dout <= 8'b00000000; //  686 :   0 - 0x0
      13'h2AF: dout <= 8'b00000000; //  687 :   0 - 0x0
      13'h2B0: dout <= 8'b00000000; //  688 :   0 - 0x0 -- Sprite 0x2b
      13'h2B1: dout <= 8'b00000000; //  689 :   0 - 0x0
      13'h2B2: dout <= 8'b00000000; //  690 :   0 - 0x0
      13'h2B3: dout <= 8'b00000000; //  691 :   0 - 0x0
      13'h2B4: dout <= 8'b00000000; //  692 :   0 - 0x0
      13'h2B5: dout <= 8'b00000000; //  693 :   0 - 0x0
      13'h2B6: dout <= 8'b00000000; //  694 :   0 - 0x0
      13'h2B7: dout <= 8'b00000000; //  695 :   0 - 0x0
      13'h2B8: dout <= 8'b11100000; //  696 : 224 - 0xe0
      13'h2B9: dout <= 8'b00000000; //  697 :   0 - 0x0
      13'h2BA: dout <= 8'b00000000; //  698 :   0 - 0x0
      13'h2BB: dout <= 8'b00000000; //  699 :   0 - 0x0
      13'h2BC: dout <= 8'b00000000; //  700 :   0 - 0x0
      13'h2BD: dout <= 8'b00000000; //  701 :   0 - 0x0
      13'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      13'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      13'h2C0: dout <= 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x2c
      13'h2C1: dout <= 8'b00000000; //  705 :   0 - 0x0
      13'h2C2: dout <= 8'b00000000; //  706 :   0 - 0x0
      13'h2C3: dout <= 8'b00000000; //  707 :   0 - 0x0
      13'h2C4: dout <= 8'b00000000; //  708 :   0 - 0x0
      13'h2C5: dout <= 8'b00000000; //  709 :   0 - 0x0
      13'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      13'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      13'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0
      13'h2C9: dout <= 8'b00000000; //  713 :   0 - 0x0
      13'h2CA: dout <= 8'b00000000; //  714 :   0 - 0x0
      13'h2CB: dout <= 8'b00000000; //  715 :   0 - 0x0
      13'h2CC: dout <= 8'b00000000; //  716 :   0 - 0x0
      13'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      13'h2CE: dout <= 8'b00001100; //  718 :  12 - 0xc
      13'h2CF: dout <= 8'b00011110; //  719 :  30 - 0x1e
      13'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x2d
      13'h2D1: dout <= 8'b00000000; //  721 :   0 - 0x0
      13'h2D2: dout <= 8'b00000000; //  722 :   0 - 0x0
      13'h2D3: dout <= 8'b00000000; //  723 :   0 - 0x0
      13'h2D4: dout <= 8'b00000000; //  724 :   0 - 0x0
      13'h2D5: dout <= 8'b00000000; //  725 :   0 - 0x0
      13'h2D6: dout <= 8'b00000000; //  726 :   0 - 0x0
      13'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      13'h2D8: dout <= 8'b00010010; //  728 :  18 - 0x12
      13'h2D9: dout <= 8'b00010010; //  729 :  18 - 0x12
      13'h2DA: dout <= 8'b00001100; //  730 :  12 - 0xc
      13'h2DB: dout <= 8'b00000000; //  731 :   0 - 0x0
      13'h2DC: dout <= 8'b00000000; //  732 :   0 - 0x0
      13'h2DD: dout <= 8'b00000000; //  733 :   0 - 0x0
      13'h2DE: dout <= 8'b00000000; //  734 :   0 - 0x0
      13'h2DF: dout <= 8'b00000000; //  735 :   0 - 0x0
      13'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x2e
      13'h2E1: dout <= 8'b00000000; //  737 :   0 - 0x0
      13'h2E2: dout <= 8'b00000000; //  738 :   0 - 0x0
      13'h2E3: dout <= 8'b00000000; //  739 :   0 - 0x0
      13'h2E4: dout <= 8'b00000000; //  740 :   0 - 0x0
      13'h2E5: dout <= 8'b00000000; //  741 :   0 - 0x0
      13'h2E6: dout <= 8'b00000000; //  742 :   0 - 0x0
      13'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      13'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0
      13'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      13'h2EA: dout <= 8'b00000000; //  746 :   0 - 0x0
      13'h2EB: dout <= 8'b00010001; //  747 :  17 - 0x11
      13'h2EC: dout <= 8'b00110010; //  748 :  50 - 0x32
      13'h2ED: dout <= 8'b00010010; //  749 :  18 - 0x12
      13'h2EE: dout <= 8'b00010010; //  750 :  18 - 0x12
      13'h2EF: dout <= 8'b00010010; //  751 :  18 - 0x12
      13'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x2f
      13'h2F1: dout <= 8'b00000000; //  753 :   0 - 0x0
      13'h2F2: dout <= 8'b00000000; //  754 :   0 - 0x0
      13'h2F3: dout <= 8'b00000000; //  755 :   0 - 0x0
      13'h2F4: dout <= 8'b00000000; //  756 :   0 - 0x0
      13'h2F5: dout <= 8'b00000000; //  757 :   0 - 0x0
      13'h2F6: dout <= 8'b00000000; //  758 :   0 - 0x0
      13'h2F7: dout <= 8'b00000000; //  759 :   0 - 0x0
      13'h2F8: dout <= 8'b00000000; //  760 :   0 - 0x0
      13'h2F9: dout <= 8'b00000000; //  761 :   0 - 0x0
      13'h2FA: dout <= 8'b00000000; //  762 :   0 - 0x0
      13'h2FB: dout <= 8'b10001100; //  763 : 140 - 0x8c
      13'h2FC: dout <= 8'b01010010; //  764 :  82 - 0x52
      13'h2FD: dout <= 8'b01010010; //  765 :  82 - 0x52
      13'h2FE: dout <= 8'b01010010; //  766 :  82 - 0x52
      13'h2FF: dout <= 8'b01010010; //  767 :  82 - 0x52
      13'h300: dout <= 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x30
      13'h301: dout <= 8'b00000000; //  769 :   0 - 0x0
      13'h302: dout <= 8'b00000000; //  770 :   0 - 0x0
      13'h303: dout <= 8'b00000000; //  771 :   0 - 0x0
      13'h304: dout <= 8'b00000000; //  772 :   0 - 0x0
      13'h305: dout <= 8'b00000000; //  773 :   0 - 0x0
      13'h306: dout <= 8'b00000000; //  774 :   0 - 0x0
      13'h307: dout <= 8'b00000000; //  775 :   0 - 0x0
      13'h308: dout <= 8'b00010010; //  776 :  18 - 0x12
      13'h309: dout <= 8'b00111001; //  777 :  57 - 0x39
      13'h30A: dout <= 8'b00000000; //  778 :   0 - 0x0
      13'h30B: dout <= 8'b00000000; //  779 :   0 - 0x0
      13'h30C: dout <= 8'b00000000; //  780 :   0 - 0x0
      13'h30D: dout <= 8'b00000000; //  781 :   0 - 0x0
      13'h30E: dout <= 8'b00000000; //  782 :   0 - 0x0
      13'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      13'h310: dout <= 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x31
      13'h311: dout <= 8'b00000000; //  785 :   0 - 0x0
      13'h312: dout <= 8'b00000000; //  786 :   0 - 0x0
      13'h313: dout <= 8'b00000000; //  787 :   0 - 0x0
      13'h314: dout <= 8'b00000000; //  788 :   0 - 0x0
      13'h315: dout <= 8'b00000000; //  789 :   0 - 0x0
      13'h316: dout <= 8'b00000000; //  790 :   0 - 0x0
      13'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      13'h318: dout <= 8'b01010010; //  792 :  82 - 0x52
      13'h319: dout <= 8'b10001100; //  793 : 140 - 0x8c
      13'h31A: dout <= 8'b00000000; //  794 :   0 - 0x0
      13'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      13'h31C: dout <= 8'b00000000; //  796 :   0 - 0x0
      13'h31D: dout <= 8'b00000000; //  797 :   0 - 0x0
      13'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      13'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      13'h320: dout <= 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x32
      13'h321: dout <= 8'b00000000; //  801 :   0 - 0x0
      13'h322: dout <= 8'b00000000; //  802 :   0 - 0x0
      13'h323: dout <= 8'b00000000; //  803 :   0 - 0x0
      13'h324: dout <= 8'b00000000; //  804 :   0 - 0x0
      13'h325: dout <= 8'b00000000; //  805 :   0 - 0x0
      13'h326: dout <= 8'b00000000; //  806 :   0 - 0x0
      13'h327: dout <= 8'b00000000; //  807 :   0 - 0x0
      13'h328: dout <= 8'b00000000; //  808 :   0 - 0x0
      13'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      13'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      13'h32B: dout <= 8'b01110001; //  811 : 113 - 0x71
      13'h32C: dout <= 8'b10001010; //  812 : 138 - 0x8a
      13'h32D: dout <= 8'b00001010; //  813 :  10 - 0xa
      13'h32E: dout <= 8'b00010010; //  814 :  18 - 0x12
      13'h32F: dout <= 8'b00100010; //  815 :  34 - 0x22
      13'h330: dout <= 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x33
      13'h331: dout <= 8'b00000000; //  817 :   0 - 0x0
      13'h332: dout <= 8'b00000000; //  818 :   0 - 0x0
      13'h333: dout <= 8'b00000000; //  819 :   0 - 0x0
      13'h334: dout <= 8'b00000000; //  820 :   0 - 0x0
      13'h335: dout <= 8'b00000000; //  821 :   0 - 0x0
      13'h336: dout <= 8'b00000000; //  822 :   0 - 0x0
      13'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      13'h338: dout <= 8'b01000010; //  824 :  66 - 0x42
      13'h339: dout <= 8'b11111001; //  825 : 249 - 0xf9
      13'h33A: dout <= 8'b00000000; //  826 :   0 - 0x0
      13'h33B: dout <= 8'b00000000; //  827 :   0 - 0x0
      13'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      13'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      13'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      13'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      13'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x34
      13'h341: dout <= 8'b00000000; //  833 :   0 - 0x0
      13'h342: dout <= 8'b00000000; //  834 :   0 - 0x0
      13'h343: dout <= 8'b00000000; //  835 :   0 - 0x0
      13'h344: dout <= 8'b00000000; //  836 :   0 - 0x0
      13'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      13'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      13'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      13'h348: dout <= 8'b00000000; //  840 :   0 - 0x0
      13'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      13'h34A: dout <= 8'b00000000; //  842 :   0 - 0x0
      13'h34B: dout <= 8'b00110001; //  843 :  49 - 0x31
      13'h34C: dout <= 8'b01001010; //  844 :  74 - 0x4a
      13'h34D: dout <= 8'b00001010; //  845 :  10 - 0xa
      13'h34E: dout <= 8'b00110010; //  846 :  50 - 0x32
      13'h34F: dout <= 8'b00001010; //  847 :  10 - 0xa
      13'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x35
      13'h351: dout <= 8'b00000000; //  849 :   0 - 0x0
      13'h352: dout <= 8'b00000000; //  850 :   0 - 0x0
      13'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      13'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      13'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      13'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      13'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      13'h358: dout <= 8'b01001010; //  856 :  74 - 0x4a
      13'h359: dout <= 8'b00110001; //  857 :  49 - 0x31
      13'h35A: dout <= 8'b00000000; //  858 :   0 - 0x0
      13'h35B: dout <= 8'b00000000; //  859 :   0 - 0x0
      13'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      13'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      13'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      13'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      13'h360: dout <= 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x36
      13'h361: dout <= 8'b00000000; //  865 :   0 - 0x0
      13'h362: dout <= 8'b00000000; //  866 :   0 - 0x0
      13'h363: dout <= 8'b00000000; //  867 :   0 - 0x0
      13'h364: dout <= 8'b00000000; //  868 :   0 - 0x0
      13'h365: dout <= 8'b00000000; //  869 :   0 - 0x0
      13'h366: dout <= 8'b00000000; //  870 :   0 - 0x0
      13'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      13'h368: dout <= 8'b00000000; //  872 :   0 - 0x0
      13'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      13'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      13'h36B: dout <= 8'b00010001; //  875 :  17 - 0x11
      13'h36C: dout <= 8'b00110010; //  876 :  50 - 0x32
      13'h36D: dout <= 8'b01010010; //  877 :  82 - 0x52
      13'h36E: dout <= 8'b10010010; //  878 : 146 - 0x92
      13'h36F: dout <= 8'b11111010; //  879 : 250 - 0xfa
      13'h370: dout <= 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x37
      13'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      13'h372: dout <= 8'b00000000; //  882 :   0 - 0x0
      13'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      13'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      13'h375: dout <= 8'b00000000; //  885 :   0 - 0x0
      13'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      13'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      13'h378: dout <= 8'b00010010; //  888 :  18 - 0x12
      13'h379: dout <= 8'b00010001; //  889 :  17 - 0x11
      13'h37A: dout <= 8'b00000000; //  890 :   0 - 0x0
      13'h37B: dout <= 8'b00000000; //  891 :   0 - 0x0
      13'h37C: dout <= 8'b00000000; //  892 :   0 - 0x0
      13'h37D: dout <= 8'b00000000; //  893 :   0 - 0x0
      13'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      13'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      13'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x38
      13'h381: dout <= 8'b00000000; //  897 :   0 - 0x0
      13'h382: dout <= 8'b00000000; //  898 :   0 - 0x0
      13'h383: dout <= 8'b00000000; //  899 :   0 - 0x0
      13'h384: dout <= 8'b00000000; //  900 :   0 - 0x0
      13'h385: dout <= 8'b00000000; //  901 :   0 - 0x0
      13'h386: dout <= 8'b00000000; //  902 :   0 - 0x0
      13'h387: dout <= 8'b00000000; //  903 :   0 - 0x0
      13'h388: dout <= 8'b00000000; //  904 :   0 - 0x0
      13'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      13'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      13'h38B: dout <= 8'b01110001; //  907 : 113 - 0x71
      13'h38C: dout <= 8'b01000010; //  908 :  66 - 0x42
      13'h38D: dout <= 8'b01000010; //  909 :  66 - 0x42
      13'h38E: dout <= 8'b01110010; //  910 : 114 - 0x72
      13'h38F: dout <= 8'b00001010; //  911 :  10 - 0xa
      13'h390: dout <= 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x39
      13'h391: dout <= 8'b00000000; //  913 :   0 - 0x0
      13'h392: dout <= 8'b00000000; //  914 :   0 - 0x0
      13'h393: dout <= 8'b00000000; //  915 :   0 - 0x0
      13'h394: dout <= 8'b00000000; //  916 :   0 - 0x0
      13'h395: dout <= 8'b00000000; //  917 :   0 - 0x0
      13'h396: dout <= 8'b00000000; //  918 :   0 - 0x0
      13'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      13'h398: dout <= 8'b00001010; //  920 :  10 - 0xa
      13'h399: dout <= 8'b01110001; //  921 : 113 - 0x71
      13'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      13'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      13'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      13'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      13'h39E: dout <= 8'b00000000; //  926 :   0 - 0x0
      13'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      13'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x3a
      13'h3A1: dout <= 8'b00000000; //  929 :   0 - 0x0
      13'h3A2: dout <= 8'b00000000; //  930 :   0 - 0x0
      13'h3A3: dout <= 8'b00000000; //  931 :   0 - 0x0
      13'h3A4: dout <= 8'b00000000; //  932 :   0 - 0x0
      13'h3A5: dout <= 8'b00000000; //  933 :   0 - 0x0
      13'h3A6: dout <= 8'b00000000; //  934 :   0 - 0x0
      13'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      13'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0
      13'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      13'h3AA: dout <= 8'b00000000; //  938 :   0 - 0x0
      13'h3AB: dout <= 8'b01110001; //  939 : 113 - 0x71
      13'h3AC: dout <= 8'b00001010; //  940 :  10 - 0xa
      13'h3AD: dout <= 8'b00010010; //  941 :  18 - 0x12
      13'h3AE: dout <= 8'b00010010; //  942 :  18 - 0x12
      13'h3AF: dout <= 8'b00100010; //  943 :  34 - 0x22
      13'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x3b
      13'h3B1: dout <= 8'b00000000; //  945 :   0 - 0x0
      13'h3B2: dout <= 8'b00000000; //  946 :   0 - 0x0
      13'h3B3: dout <= 8'b00000000; //  947 :   0 - 0x0
      13'h3B4: dout <= 8'b00000000; //  948 :   0 - 0x0
      13'h3B5: dout <= 8'b00000000; //  949 :   0 - 0x0
      13'h3B6: dout <= 8'b00000000; //  950 :   0 - 0x0
      13'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      13'h3B8: dout <= 8'b00100010; //  952 :  34 - 0x22
      13'h3B9: dout <= 8'b00100001; //  953 :  33 - 0x21
      13'h3BA: dout <= 8'b00000000; //  954 :   0 - 0x0
      13'h3BB: dout <= 8'b00000000; //  955 :   0 - 0x0
      13'h3BC: dout <= 8'b00000000; //  956 :   0 - 0x0
      13'h3BD: dout <= 8'b00000000; //  957 :   0 - 0x0
      13'h3BE: dout <= 8'b00000000; //  958 :   0 - 0x0
      13'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      13'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x3c
      13'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      13'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      13'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      13'h3C4: dout <= 8'b00000000; //  964 :   0 - 0x0
      13'h3C5: dout <= 8'b00000000; //  965 :   0 - 0x0
      13'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      13'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      13'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0
      13'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      13'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      13'h3CB: dout <= 8'b01110001; //  971 : 113 - 0x71
      13'h3CC: dout <= 8'b10001010; //  972 : 138 - 0x8a
      13'h3CD: dout <= 8'b10001010; //  973 : 138 - 0x8a
      13'h3CE: dout <= 8'b01110010; //  974 : 114 - 0x72
      13'h3CF: dout <= 8'b10001010; //  975 : 138 - 0x8a
      13'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x3d
      13'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      13'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      13'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      13'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      13'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      13'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      13'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      13'h3D8: dout <= 8'b10001010; //  984 : 138 - 0x8a
      13'h3D9: dout <= 8'b01110001; //  985 : 113 - 0x71
      13'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      13'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      13'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      13'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      13'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      13'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      13'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x3e
      13'h3E1: dout <= 8'b00000000; //  993 :   0 - 0x0
      13'h3E2: dout <= 8'b00000000; //  994 :   0 - 0x0
      13'h3E3: dout <= 8'b00000000; //  995 :   0 - 0x0
      13'h3E4: dout <= 8'b00000000; //  996 :   0 - 0x0
      13'h3E5: dout <= 8'b00000000; //  997 :   0 - 0x0
      13'h3E6: dout <= 8'b00000000; //  998 :   0 - 0x0
      13'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      13'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0
      13'h3E9: dout <= 8'b00000000; // 1001 :   0 - 0x0
      13'h3EA: dout <= 8'b00000000; // 1002 :   0 - 0x0
      13'h3EB: dout <= 8'b10011000; // 1003 : 152 - 0x98
      13'h3EC: dout <= 8'b10100101; // 1004 : 165 - 0xa5
      13'h3ED: dout <= 8'b10100101; // 1005 : 165 - 0xa5
      13'h3EE: dout <= 8'b10100101; // 1006 : 165 - 0xa5
      13'h3EF: dout <= 8'b10100101; // 1007 : 165 - 0xa5
      13'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x3f
      13'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      13'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      13'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      13'h3F4: dout <= 8'b00000000; // 1012 :   0 - 0x0
      13'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      13'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      13'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      13'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0
      13'h3F9: dout <= 8'b00000000; // 1017 :   0 - 0x0
      13'h3FA: dout <= 8'b00000000; // 1018 :   0 - 0x0
      13'h3FB: dout <= 8'b11000110; // 1019 : 198 - 0xc6
      13'h3FC: dout <= 8'b00101001; // 1020 :  41 - 0x29
      13'h3FD: dout <= 8'b00101001; // 1021 :  41 - 0x29
      13'h3FE: dout <= 8'b00101001; // 1022 :  41 - 0x29
      13'h3FF: dout <= 8'b00101001; // 1023 :  41 - 0x29
      13'h400: dout <= 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x40
      13'h401: dout <= 8'b00000000; // 1025 :   0 - 0x0
      13'h402: dout <= 8'b00000000; // 1026 :   0 - 0x0
      13'h403: dout <= 8'b00000000; // 1027 :   0 - 0x0
      13'h404: dout <= 8'b00000000; // 1028 :   0 - 0x0
      13'h405: dout <= 8'b00000000; // 1029 :   0 - 0x0
      13'h406: dout <= 8'b00000000; // 1030 :   0 - 0x0
      13'h407: dout <= 8'b00000000; // 1031 :   0 - 0x0
      13'h408: dout <= 8'b10100101; // 1032 : 165 - 0xa5
      13'h409: dout <= 8'b10011000; // 1033 : 152 - 0x98
      13'h40A: dout <= 8'b00000000; // 1034 :   0 - 0x0
      13'h40B: dout <= 8'b00000000; // 1035 :   0 - 0x0
      13'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      13'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      13'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      13'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      13'h410: dout <= 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x41
      13'h411: dout <= 8'b00000000; // 1041 :   0 - 0x0
      13'h412: dout <= 8'b00000000; // 1042 :   0 - 0x0
      13'h413: dout <= 8'b00000000; // 1043 :   0 - 0x0
      13'h414: dout <= 8'b00000000; // 1044 :   0 - 0x0
      13'h415: dout <= 8'b00000000; // 1045 :   0 - 0x0
      13'h416: dout <= 8'b00000000; // 1046 :   0 - 0x0
      13'h417: dout <= 8'b00000000; // 1047 :   0 - 0x0
      13'h418: dout <= 8'b00101001; // 1048 :  41 - 0x29
      13'h419: dout <= 8'b11000110; // 1049 : 198 - 0xc6
      13'h41A: dout <= 8'b00000000; // 1050 :   0 - 0x0
      13'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      13'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      13'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      13'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      13'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      13'h420: dout <= 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x42
      13'h421: dout <= 8'b00000000; // 1057 :   0 - 0x0
      13'h422: dout <= 8'b00000000; // 1058 :   0 - 0x0
      13'h423: dout <= 8'b00000000; // 1059 :   0 - 0x0
      13'h424: dout <= 8'b00000000; // 1060 :   0 - 0x0
      13'h425: dout <= 8'b00000000; // 1061 :   0 - 0x0
      13'h426: dout <= 8'b00000000; // 1062 :   0 - 0x0
      13'h427: dout <= 8'b00000000; // 1063 :   0 - 0x0
      13'h428: dout <= 8'b00000000; // 1064 :   0 - 0x0
      13'h429: dout <= 8'b00000000; // 1065 :   0 - 0x0
      13'h42A: dout <= 8'b00000000; // 1066 :   0 - 0x0
      13'h42B: dout <= 8'b10011100; // 1067 : 156 - 0x9c
      13'h42C: dout <= 8'b10100001; // 1068 : 161 - 0xa1
      13'h42D: dout <= 8'b10100001; // 1069 : 161 - 0xa1
      13'h42E: dout <= 8'b10111101; // 1070 : 189 - 0xbd
      13'h42F: dout <= 8'b10100101; // 1071 : 165 - 0xa5
      13'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x43
      13'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      13'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      13'h433: dout <= 8'b00000000; // 1075 :   0 - 0x0
      13'h434: dout <= 8'b00000000; // 1076 :   0 - 0x0
      13'h435: dout <= 8'b00000000; // 1077 :   0 - 0x0
      13'h436: dout <= 8'b00000000; // 1078 :   0 - 0x0
      13'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      13'h438: dout <= 8'b10100101; // 1080 : 165 - 0xa5
      13'h439: dout <= 8'b10011000; // 1081 : 152 - 0x98
      13'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      13'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      13'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      13'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      13'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      13'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      13'h440: dout <= 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x44
      13'h441: dout <= 8'b00000000; // 1089 :   0 - 0x0
      13'h442: dout <= 8'b00000000; // 1090 :   0 - 0x0
      13'h443: dout <= 8'b00000000; // 1091 :   0 - 0x0
      13'h444: dout <= 8'b00000000; // 1092 :   0 - 0x0
      13'h445: dout <= 8'b00000000; // 1093 :   0 - 0x0
      13'h446: dout <= 8'b00000000; // 1094 :   0 - 0x0
      13'h447: dout <= 8'b00000000; // 1095 :   0 - 0x0
      13'h448: dout <= 8'b00000000; // 1096 :   0 - 0x0
      13'h449: dout <= 8'b00000000; // 1097 :   0 - 0x0
      13'h44A: dout <= 8'b00000000; // 1098 :   0 - 0x0
      13'h44B: dout <= 8'b01100010; // 1099 :  98 - 0x62
      13'h44C: dout <= 8'b10010101; // 1100 : 149 - 0x95
      13'h44D: dout <= 8'b00010101; // 1101 :  21 - 0x15
      13'h44E: dout <= 8'b00100101; // 1102 :  37 - 0x25
      13'h44F: dout <= 8'b01000101; // 1103 :  69 - 0x45
      13'h450: dout <= 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x45
      13'h451: dout <= 8'b00000000; // 1105 :   0 - 0x0
      13'h452: dout <= 8'b00000000; // 1106 :   0 - 0x0
      13'h453: dout <= 8'b00000000; // 1107 :   0 - 0x0
      13'h454: dout <= 8'b00000000; // 1108 :   0 - 0x0
      13'h455: dout <= 8'b00000000; // 1109 :   0 - 0x0
      13'h456: dout <= 8'b00000000; // 1110 :   0 - 0x0
      13'h457: dout <= 8'b00000000; // 1111 :   0 - 0x0
      13'h458: dout <= 8'b00000000; // 1112 :   0 - 0x0
      13'h459: dout <= 8'b00000000; // 1113 :   0 - 0x0
      13'h45A: dout <= 8'b00000000; // 1114 :   0 - 0x0
      13'h45B: dout <= 8'b00100010; // 1115 :  34 - 0x22
      13'h45C: dout <= 8'b01010101; // 1116 :  85 - 0x55
      13'h45D: dout <= 8'b01010101; // 1117 :  85 - 0x55
      13'h45E: dout <= 8'b01010101; // 1118 :  85 - 0x55
      13'h45F: dout <= 8'b01010101; // 1119 :  85 - 0x55
      13'h460: dout <= 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x46
      13'h461: dout <= 8'b00000000; // 1121 :   0 - 0x0
      13'h462: dout <= 8'b00000000; // 1122 :   0 - 0x0
      13'h463: dout <= 8'b00000000; // 1123 :   0 - 0x0
      13'h464: dout <= 8'b00000000; // 1124 :   0 - 0x0
      13'h465: dout <= 8'b00000000; // 1125 :   0 - 0x0
      13'h466: dout <= 8'b00000000; // 1126 :   0 - 0x0
      13'h467: dout <= 8'b00000000; // 1127 :   0 - 0x0
      13'h468: dout <= 8'b10000101; // 1128 : 133 - 0x85
      13'h469: dout <= 8'b11110010; // 1129 : 242 - 0xf2
      13'h46A: dout <= 8'b00000000; // 1130 :   0 - 0x0
      13'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      13'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      13'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      13'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      13'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      13'h470: dout <= 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x47
      13'h471: dout <= 8'b00000000; // 1137 :   0 - 0x0
      13'h472: dout <= 8'b00000000; // 1138 :   0 - 0x0
      13'h473: dout <= 8'b00000000; // 1139 :   0 - 0x0
      13'h474: dout <= 8'b00000000; // 1140 :   0 - 0x0
      13'h475: dout <= 8'b00000000; // 1141 :   0 - 0x0
      13'h476: dout <= 8'b00000000; // 1142 :   0 - 0x0
      13'h477: dout <= 8'b00000000; // 1143 :   0 - 0x0
      13'h478: dout <= 8'b01010101; // 1144 :  85 - 0x55
      13'h479: dout <= 8'b00100010; // 1145 :  34 - 0x22
      13'h47A: dout <= 8'b00000000; // 1146 :   0 - 0x0
      13'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      13'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      13'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      13'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      13'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      13'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x48
      13'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      13'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      13'h483: dout <= 8'b00000000; // 1155 :   0 - 0x0
      13'h484: dout <= 8'b00000000; // 1156 :   0 - 0x0
      13'h485: dout <= 8'b00000000; // 1157 :   0 - 0x0
      13'h486: dout <= 8'b00000000; // 1158 :   0 - 0x0
      13'h487: dout <= 8'b00000000; // 1159 :   0 - 0x0
      13'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0
      13'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      13'h48A: dout <= 8'b00000000; // 1162 :   0 - 0x0
      13'h48B: dout <= 8'b01100010; // 1163 :  98 - 0x62
      13'h48C: dout <= 8'b10010101; // 1164 : 149 - 0x95
      13'h48D: dout <= 8'b00010101; // 1165 :  21 - 0x15
      13'h48E: dout <= 8'b01100101; // 1166 : 101 - 0x65
      13'h48F: dout <= 8'b00010101; // 1167 :  21 - 0x15
      13'h490: dout <= 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x49
      13'h491: dout <= 8'b00000000; // 1169 :   0 - 0x0
      13'h492: dout <= 8'b00000000; // 1170 :   0 - 0x0
      13'h493: dout <= 8'b00000000; // 1171 :   0 - 0x0
      13'h494: dout <= 8'b00000000; // 1172 :   0 - 0x0
      13'h495: dout <= 8'b00000000; // 1173 :   0 - 0x0
      13'h496: dout <= 8'b00000000; // 1174 :   0 - 0x0
      13'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      13'h498: dout <= 8'b10010101; // 1176 : 149 - 0x95
      13'h499: dout <= 8'b01100010; // 1177 :  98 - 0x62
      13'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      13'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      13'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      13'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      13'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      13'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      13'h4A0: dout <= 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x4a
      13'h4A1: dout <= 8'b00000000; // 1185 :   0 - 0x0
      13'h4A2: dout <= 8'b00000000; // 1186 :   0 - 0x0
      13'h4A3: dout <= 8'b00000000; // 1187 :   0 - 0x0
      13'h4A4: dout <= 8'b00000000; // 1188 :   0 - 0x0
      13'h4A5: dout <= 8'b00000000; // 1189 :   0 - 0x0
      13'h4A6: dout <= 8'b00000000; // 1190 :   0 - 0x0
      13'h4A7: dout <= 8'b00000000; // 1191 :   0 - 0x0
      13'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0
      13'h4A9: dout <= 8'b00000000; // 1193 :   0 - 0x0
      13'h4AA: dout <= 8'b00000000; // 1194 :   0 - 0x0
      13'h4AB: dout <= 8'b11100010; // 1195 : 226 - 0xe2
      13'h4AC: dout <= 8'b10000101; // 1196 : 133 - 0x85
      13'h4AD: dout <= 8'b10000101; // 1197 : 133 - 0x85
      13'h4AE: dout <= 8'b11100101; // 1198 : 229 - 0xe5
      13'h4AF: dout <= 8'b00010101; // 1199 :  21 - 0x15
      13'h4B0: dout <= 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x4b
      13'h4B1: dout <= 8'b00000000; // 1201 :   0 - 0x0
      13'h4B2: dout <= 8'b00000000; // 1202 :   0 - 0x0
      13'h4B3: dout <= 8'b00000000; // 1203 :   0 - 0x0
      13'h4B4: dout <= 8'b00000000; // 1204 :   0 - 0x0
      13'h4B5: dout <= 8'b00000000; // 1205 :   0 - 0x0
      13'h4B6: dout <= 8'b00000000; // 1206 :   0 - 0x0
      13'h4B7: dout <= 8'b00000000; // 1207 :   0 - 0x0
      13'h4B8: dout <= 8'b00010101; // 1208 :  21 - 0x15
      13'h4B9: dout <= 8'b11100010; // 1209 : 226 - 0xe2
      13'h4BA: dout <= 8'b00000000; // 1210 :   0 - 0x0
      13'h4BB: dout <= 8'b00000000; // 1211 :   0 - 0x0
      13'h4BC: dout <= 8'b00000000; // 1212 :   0 - 0x0
      13'h4BD: dout <= 8'b00000000; // 1213 :   0 - 0x0
      13'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      13'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      13'h4C0: dout <= 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x4c
      13'h4C1: dout <= 8'b00000000; // 1217 :   0 - 0x0
      13'h4C2: dout <= 8'b00000000; // 1218 :   0 - 0x0
      13'h4C3: dout <= 8'b00000000; // 1219 :   0 - 0x0
      13'h4C4: dout <= 8'b00000000; // 1220 :   0 - 0x0
      13'h4C5: dout <= 8'b00000000; // 1221 :   0 - 0x0
      13'h4C6: dout <= 8'b00000000; // 1222 :   0 - 0x0
      13'h4C7: dout <= 8'b00000000; // 1223 :   0 - 0x0
      13'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0
      13'h4C9: dout <= 8'b00000000; // 1225 :   0 - 0x0
      13'h4CA: dout <= 8'b00000000; // 1226 :   0 - 0x0
      13'h4CB: dout <= 8'b00000000; // 1227 :   0 - 0x0
      13'h4CC: dout <= 8'b00000000; // 1228 :   0 - 0x0
      13'h4CD: dout <= 8'b00000000; // 1229 :   0 - 0x0
      13'h4CE: dout <= 8'b00000000; // 1230 :   0 - 0x0
      13'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      13'h4D0: dout <= 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x4d
      13'h4D1: dout <= 8'b00000000; // 1233 :   0 - 0x0
      13'h4D2: dout <= 8'b00000000; // 1234 :   0 - 0x0
      13'h4D3: dout <= 8'b00000001; // 1235 :   1 - 0x1
      13'h4D4: dout <= 8'b00000011; // 1236 :   3 - 0x3
      13'h4D5: dout <= 8'b00000111; // 1237 :   7 - 0x7
      13'h4D6: dout <= 8'b00001111; // 1238 :  15 - 0xf
      13'h4D7: dout <= 8'b00011111; // 1239 :  31 - 0x1f
      13'h4D8: dout <= 8'b00000000; // 1240 :   0 - 0x0
      13'h4D9: dout <= 8'b00000000; // 1241 :   0 - 0x0
      13'h4DA: dout <= 8'b00000000; // 1242 :   0 - 0x0
      13'h4DB: dout <= 8'b00000000; // 1243 :   0 - 0x0
      13'h4DC: dout <= 8'b00000000; // 1244 :   0 - 0x0
      13'h4DD: dout <= 8'b00000000; // 1245 :   0 - 0x0
      13'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      13'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      13'h4E0: dout <= 8'b00000000; // 1248 :   0 - 0x0 -- Sprite 0x4e
      13'h4E1: dout <= 8'b00001111; // 1249 :  15 - 0xf
      13'h4E2: dout <= 8'b01111111; // 1250 : 127 - 0x7f
      13'h4E3: dout <= 8'b11111111; // 1251 : 255 - 0xff
      13'h4E4: dout <= 8'b11111111; // 1252 : 255 - 0xff
      13'h4E5: dout <= 8'b11111111; // 1253 : 255 - 0xff
      13'h4E6: dout <= 8'b11111111; // 1254 : 255 - 0xff
      13'h4E7: dout <= 8'b11111111; // 1255 : 255 - 0xff
      13'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0
      13'h4E9: dout <= 8'b00000000; // 1257 :   0 - 0x0
      13'h4EA: dout <= 8'b00000000; // 1258 :   0 - 0x0
      13'h4EB: dout <= 8'b00000000; // 1259 :   0 - 0x0
      13'h4EC: dout <= 8'b00000000; // 1260 :   0 - 0x0
      13'h4ED: dout <= 8'b00000000; // 1261 :   0 - 0x0
      13'h4EE: dout <= 8'b00000000; // 1262 :   0 - 0x0
      13'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      13'h4F0: dout <= 8'b00011111; // 1264 :  31 - 0x1f -- Sprite 0x4f
      13'h4F1: dout <= 8'b00111111; // 1265 :  63 - 0x3f
      13'h4F2: dout <= 8'b00111111; // 1266 :  63 - 0x3f
      13'h4F3: dout <= 8'b00111111; // 1267 :  63 - 0x3f
      13'h4F4: dout <= 8'b01111111; // 1268 : 127 - 0x7f
      13'h4F5: dout <= 8'b01111111; // 1269 : 127 - 0x7f
      13'h4F6: dout <= 8'b01111111; // 1270 : 127 - 0x7f
      13'h4F7: dout <= 8'b01111111; // 1271 : 127 - 0x7f
      13'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0
      13'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      13'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      13'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      13'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      13'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      13'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      13'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      13'h500: dout <= 8'b11111111; // 1280 : 255 - 0xff -- Sprite 0x50
      13'h501: dout <= 8'b11111111; // 1281 : 255 - 0xff
      13'h502: dout <= 8'b11111111; // 1282 : 255 - 0xff
      13'h503: dout <= 8'b11111111; // 1283 : 255 - 0xff
      13'h504: dout <= 8'b11111111; // 1284 : 255 - 0xff
      13'h505: dout <= 8'b11111111; // 1285 : 255 - 0xff
      13'h506: dout <= 8'b11111111; // 1286 : 255 - 0xff
      13'h507: dout <= 8'b11111111; // 1287 : 255 - 0xff
      13'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0
      13'h509: dout <= 8'b00000000; // 1289 :   0 - 0x0
      13'h50A: dout <= 8'b00000000; // 1290 :   0 - 0x0
      13'h50B: dout <= 8'b00000000; // 1291 :   0 - 0x0
      13'h50C: dout <= 8'b00000000; // 1292 :   0 - 0x0
      13'h50D: dout <= 8'b00000000; // 1293 :   0 - 0x0
      13'h50E: dout <= 8'b00000000; // 1294 :   0 - 0x0
      13'h50F: dout <= 8'b00000000; // 1295 :   0 - 0x0
      13'h510: dout <= 8'b11111111; // 1296 : 255 - 0xff -- Sprite 0x51
      13'h511: dout <= 8'b11111111; // 1297 : 255 - 0xff
      13'h512: dout <= 8'b11111111; // 1298 : 255 - 0xff
      13'h513: dout <= 8'b11111111; // 1299 : 255 - 0xff
      13'h514: dout <= 8'b11111111; // 1300 : 255 - 0xff
      13'h515: dout <= 8'b11111111; // 1301 : 255 - 0xff
      13'h516: dout <= 8'b11111111; // 1302 : 255 - 0xff
      13'h517: dout <= 8'b11111110; // 1303 : 254 - 0xfe
      13'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0
      13'h519: dout <= 8'b00000000; // 1305 :   0 - 0x0
      13'h51A: dout <= 8'b00000000; // 1306 :   0 - 0x0
      13'h51B: dout <= 8'b00000000; // 1307 :   0 - 0x0
      13'h51C: dout <= 8'b00000000; // 1308 :   0 - 0x0
      13'h51D: dout <= 8'b00000000; // 1309 :   0 - 0x0
      13'h51E: dout <= 8'b00000000; // 1310 :   0 - 0x0
      13'h51F: dout <= 8'b00000000; // 1311 :   0 - 0x0
      13'h520: dout <= 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0x52
      13'h521: dout <= 8'b00000000; // 1313 :   0 - 0x0
      13'h522: dout <= 8'b00000000; // 1314 :   0 - 0x0
      13'h523: dout <= 8'b10000000; // 1315 : 128 - 0x80
      13'h524: dout <= 8'b11000000; // 1316 : 192 - 0xc0
      13'h525: dout <= 8'b11100000; // 1317 : 224 - 0xe0
      13'h526: dout <= 8'b11110000; // 1318 : 240 - 0xf0
      13'h527: dout <= 8'b11110000; // 1319 : 240 - 0xf0
      13'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0
      13'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      13'h52A: dout <= 8'b00000000; // 1322 :   0 - 0x0
      13'h52B: dout <= 8'b00000000; // 1323 :   0 - 0x0
      13'h52C: dout <= 8'b00000000; // 1324 :   0 - 0x0
      13'h52D: dout <= 8'b00000000; // 1325 :   0 - 0x0
      13'h52E: dout <= 8'b00000000; // 1326 :   0 - 0x0
      13'h52F: dout <= 8'b00000000; // 1327 :   0 - 0x0
      13'h530: dout <= 8'b11111111; // 1328 : 255 - 0xff -- Sprite 0x53
      13'h531: dout <= 8'b11111111; // 1329 : 255 - 0xff
      13'h532: dout <= 8'b11111110; // 1330 : 254 - 0xfe
      13'h533: dout <= 8'b11111100; // 1331 : 252 - 0xfc
      13'h534: dout <= 8'b11110000; // 1332 : 240 - 0xf0
      13'h535: dout <= 8'b11100000; // 1333 : 224 - 0xe0
      13'h536: dout <= 8'b10000000; // 1334 : 128 - 0x80
      13'h537: dout <= 8'b00000000; // 1335 :   0 - 0x0
      13'h538: dout <= 8'b00000000; // 1336 :   0 - 0x0
      13'h539: dout <= 8'b00000000; // 1337 :   0 - 0x0
      13'h53A: dout <= 8'b00000000; // 1338 :   0 - 0x0
      13'h53B: dout <= 8'b00000000; // 1339 :   0 - 0x0
      13'h53C: dout <= 8'b00000000; // 1340 :   0 - 0x0
      13'h53D: dout <= 8'b00000000; // 1341 :   0 - 0x0
      13'h53E: dout <= 8'b00000000; // 1342 :   0 - 0x0
      13'h53F: dout <= 8'b00000000; // 1343 :   0 - 0x0
      13'h540: dout <= 8'b11000000; // 1344 : 192 - 0xc0 -- Sprite 0x54
      13'h541: dout <= 8'b10000000; // 1345 : 128 - 0x80
      13'h542: dout <= 8'b00000000; // 1346 :   0 - 0x0
      13'h543: dout <= 8'b00000000; // 1347 :   0 - 0x0
      13'h544: dout <= 8'b00000000; // 1348 :   0 - 0x0
      13'h545: dout <= 8'b00000000; // 1349 :   0 - 0x0
      13'h546: dout <= 8'b00000000; // 1350 :   0 - 0x0
      13'h547: dout <= 8'b00000000; // 1351 :   0 - 0x0
      13'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0
      13'h549: dout <= 8'b00000000; // 1353 :   0 - 0x0
      13'h54A: dout <= 8'b00000000; // 1354 :   0 - 0x0
      13'h54B: dout <= 8'b00000000; // 1355 :   0 - 0x0
      13'h54C: dout <= 8'b00000000; // 1356 :   0 - 0x0
      13'h54D: dout <= 8'b00000000; // 1357 :   0 - 0x0
      13'h54E: dout <= 8'b00000000; // 1358 :   0 - 0x0
      13'h54F: dout <= 8'b00000000; // 1359 :   0 - 0x0
      13'h550: dout <= 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0x55
      13'h551: dout <= 8'b11110000; // 1361 : 240 - 0xf0
      13'h552: dout <= 8'b11111110; // 1362 : 254 - 0xfe
      13'h553: dout <= 8'b11111110; // 1363 : 254 - 0xfe
      13'h554: dout <= 8'b11111110; // 1364 : 254 - 0xfe
      13'h555: dout <= 8'b11111100; // 1365 : 252 - 0xfc
      13'h556: dout <= 8'b11111000; // 1366 : 248 - 0xf8
      13'h557: dout <= 8'b11111000; // 1367 : 248 - 0xf8
      13'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0
      13'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      13'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      13'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      13'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      13'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      13'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      13'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      13'h560: dout <= 8'b11110000; // 1376 : 240 - 0xf0 -- Sprite 0x56
      13'h561: dout <= 8'b11100000; // 1377 : 224 - 0xe0
      13'h562: dout <= 8'b11100000; // 1378 : 224 - 0xe0
      13'h563: dout <= 8'b11000000; // 1379 : 192 - 0xc0
      13'h564: dout <= 8'b10000000; // 1380 : 128 - 0x80
      13'h565: dout <= 8'b10000000; // 1381 : 128 - 0x80
      13'h566: dout <= 8'b00000000; // 1382 :   0 - 0x0
      13'h567: dout <= 8'b00000000; // 1383 :   0 - 0x0
      13'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0
      13'h569: dout <= 8'b00000000; // 1385 :   0 - 0x0
      13'h56A: dout <= 8'b00000000; // 1386 :   0 - 0x0
      13'h56B: dout <= 8'b00000000; // 1387 :   0 - 0x0
      13'h56C: dout <= 8'b00000000; // 1388 :   0 - 0x0
      13'h56D: dout <= 8'b00000000; // 1389 :   0 - 0x0
      13'h56E: dout <= 8'b00000000; // 1390 :   0 - 0x0
      13'h56F: dout <= 8'b00000000; // 1391 :   0 - 0x0
      13'h570: dout <= 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0x57
      13'h571: dout <= 8'b00000000; // 1393 :   0 - 0x0
      13'h572: dout <= 8'b00000000; // 1394 :   0 - 0x0
      13'h573: dout <= 8'b00000000; // 1395 :   0 - 0x0
      13'h574: dout <= 8'b00000000; // 1396 :   0 - 0x0
      13'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      13'h576: dout <= 8'b00000000; // 1398 :   0 - 0x0
      13'h577: dout <= 8'b00000100; // 1399 :   4 - 0x4
      13'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0
      13'h579: dout <= 8'b00000000; // 1401 :   0 - 0x0
      13'h57A: dout <= 8'b00000000; // 1402 :   0 - 0x0
      13'h57B: dout <= 8'b00000000; // 1403 :   0 - 0x0
      13'h57C: dout <= 8'b00000000; // 1404 :   0 - 0x0
      13'h57D: dout <= 8'b00000000; // 1405 :   0 - 0x0
      13'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      13'h57F: dout <= 8'b00000100; // 1407 :   4 - 0x4
      13'h580: dout <= 8'b00000110; // 1408 :   6 - 0x6 -- Sprite 0x58
      13'h581: dout <= 8'b00000110; // 1409 :   6 - 0x6
      13'h582: dout <= 8'b00000111; // 1410 :   7 - 0x7
      13'h583: dout <= 8'b00000111; // 1411 :   7 - 0x7
      13'h584: dout <= 8'b00000111; // 1412 :   7 - 0x7
      13'h585: dout <= 8'b00000111; // 1413 :   7 - 0x7
      13'h586: dout <= 8'b00000000; // 1414 :   0 - 0x0
      13'h587: dout <= 8'b00000000; // 1415 :   0 - 0x0
      13'h588: dout <= 8'b00000110; // 1416 :   6 - 0x6
      13'h589: dout <= 8'b00000110; // 1417 :   6 - 0x6
      13'h58A: dout <= 8'b00000111; // 1418 :   7 - 0x7
      13'h58B: dout <= 8'b00000111; // 1419 :   7 - 0x7
      13'h58C: dout <= 8'b00000111; // 1420 :   7 - 0x7
      13'h58D: dout <= 8'b00000111; // 1421 :   7 - 0x7
      13'h58E: dout <= 8'b00000000; // 1422 :   0 - 0x0
      13'h58F: dout <= 8'b00000000; // 1423 :   0 - 0x0
      13'h590: dout <= 8'b00000000; // 1424 :   0 - 0x0 -- Sprite 0x59
      13'h591: dout <= 8'b00000000; // 1425 :   0 - 0x0
      13'h592: dout <= 8'b00000000; // 1426 :   0 - 0x0
      13'h593: dout <= 8'b00000000; // 1427 :   0 - 0x0
      13'h594: dout <= 8'b00000000; // 1428 :   0 - 0x0
      13'h595: dout <= 8'b00000000; // 1429 :   0 - 0x0
      13'h596: dout <= 8'b00000000; // 1430 :   0 - 0x0
      13'h597: dout <= 8'b00010000; // 1431 :  16 - 0x10
      13'h598: dout <= 8'b00000000; // 1432 :   0 - 0x0
      13'h599: dout <= 8'b00000000; // 1433 :   0 - 0x0
      13'h59A: dout <= 8'b00000000; // 1434 :   0 - 0x0
      13'h59B: dout <= 8'b00000000; // 1435 :   0 - 0x0
      13'h59C: dout <= 8'b00000000; // 1436 :   0 - 0x0
      13'h59D: dout <= 8'b00000000; // 1437 :   0 - 0x0
      13'h59E: dout <= 8'b00000000; // 1438 :   0 - 0x0
      13'h59F: dout <= 8'b00010000; // 1439 :  16 - 0x10
      13'h5A0: dout <= 8'b00011100; // 1440 :  28 - 0x1c -- Sprite 0x5a
      13'h5A1: dout <= 8'b00011110; // 1441 :  30 - 0x1e
      13'h5A2: dout <= 8'b00011111; // 1442 :  31 - 0x1f
      13'h5A3: dout <= 8'b00011111; // 1443 :  31 - 0x1f
      13'h5A4: dout <= 8'b00011111; // 1444 :  31 - 0x1f
      13'h5A5: dout <= 8'b00011111; // 1445 :  31 - 0x1f
      13'h5A6: dout <= 8'b00000000; // 1446 :   0 - 0x0
      13'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      13'h5A8: dout <= 8'b00011100; // 1448 :  28 - 0x1c
      13'h5A9: dout <= 8'b00011110; // 1449 :  30 - 0x1e
      13'h5AA: dout <= 8'b00011111; // 1450 :  31 - 0x1f
      13'h5AB: dout <= 8'b00011111; // 1451 :  31 - 0x1f
      13'h5AC: dout <= 8'b00011111; // 1452 :  31 - 0x1f
      13'h5AD: dout <= 8'b00011111; // 1453 :  31 - 0x1f
      13'h5AE: dout <= 8'b00000000; // 1454 :   0 - 0x0
      13'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      13'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0x5b
      13'h5B1: dout <= 8'b00000000; // 1457 :   0 - 0x0
      13'h5B2: dout <= 8'b00000000; // 1458 :   0 - 0x0
      13'h5B3: dout <= 8'b00000000; // 1459 :   0 - 0x0
      13'h5B4: dout <= 8'b00000000; // 1460 :   0 - 0x0
      13'h5B5: dout <= 8'b00000000; // 1461 :   0 - 0x0
      13'h5B6: dout <= 8'b00000000; // 1462 :   0 - 0x0
      13'h5B7: dout <= 8'b11000000; // 1463 : 192 - 0xc0
      13'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0
      13'h5B9: dout <= 8'b00000000; // 1465 :   0 - 0x0
      13'h5BA: dout <= 8'b00000000; // 1466 :   0 - 0x0
      13'h5BB: dout <= 8'b00000000; // 1467 :   0 - 0x0
      13'h5BC: dout <= 8'b00000000; // 1468 :   0 - 0x0
      13'h5BD: dout <= 8'b00000000; // 1469 :   0 - 0x0
      13'h5BE: dout <= 8'b00000000; // 1470 :   0 - 0x0
      13'h5BF: dout <= 8'b11000000; // 1471 : 192 - 0xc0
      13'h5C0: dout <= 8'b11110000; // 1472 : 240 - 0xf0 -- Sprite 0x5c
      13'h5C1: dout <= 8'b11111100; // 1473 : 252 - 0xfc
      13'h5C2: dout <= 8'b11111111; // 1474 : 255 - 0xff
      13'h5C3: dout <= 8'b11111111; // 1475 : 255 - 0xff
      13'h5C4: dout <= 8'b11111111; // 1476 : 255 - 0xff
      13'h5C5: dout <= 8'b11111111; // 1477 : 255 - 0xff
      13'h5C6: dout <= 8'b00000000; // 1478 :   0 - 0x0
      13'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      13'h5C8: dout <= 8'b11110000; // 1480 : 240 - 0xf0
      13'h5C9: dout <= 8'b11111100; // 1481 : 252 - 0xfc
      13'h5CA: dout <= 8'b11111111; // 1482 : 255 - 0xff
      13'h5CB: dout <= 8'b11111111; // 1483 : 255 - 0xff
      13'h5CC: dout <= 8'b11111111; // 1484 : 255 - 0xff
      13'h5CD: dout <= 8'b11111111; // 1485 : 255 - 0xff
      13'h5CE: dout <= 8'b00000000; // 1486 :   0 - 0x0
      13'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      13'h5D0: dout <= 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0x5d
      13'h5D1: dout <= 8'b00000000; // 1489 :   0 - 0x0
      13'h5D2: dout <= 8'b00000001; // 1490 :   1 - 0x1
      13'h5D3: dout <= 8'b00000011; // 1491 :   3 - 0x3
      13'h5D4: dout <= 8'b00001111; // 1492 :  15 - 0xf
      13'h5D5: dout <= 8'b00001111; // 1493 :  15 - 0xf
      13'h5D6: dout <= 8'b00000000; // 1494 :   0 - 0x0
      13'h5D7: dout <= 8'b00000000; // 1495 :   0 - 0x0
      13'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0
      13'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      13'h5DA: dout <= 8'b00000001; // 1498 :   1 - 0x1
      13'h5DB: dout <= 8'b00000011; // 1499 :   3 - 0x3
      13'h5DC: dout <= 8'b00001111; // 1500 :  15 - 0xf
      13'h5DD: dout <= 8'b00001111; // 1501 :  15 - 0xf
      13'h5DE: dout <= 8'b00000000; // 1502 :   0 - 0x0
      13'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      13'h5E0: dout <= 8'b11111100; // 1504 : 252 - 0xfc -- Sprite 0x5e
      13'h5E1: dout <= 8'b11111100; // 1505 : 252 - 0xfc
      13'h5E2: dout <= 8'b11111100; // 1506 : 252 - 0xfc
      13'h5E3: dout <= 8'b11111100; // 1507 : 252 - 0xfc
      13'h5E4: dout <= 8'b11111000; // 1508 : 248 - 0xf8
      13'h5E5: dout <= 8'b11111100; // 1509 : 252 - 0xfc
      13'h5E6: dout <= 8'b00111100; // 1510 :  60 - 0x3c
      13'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      13'h5E8: dout <= 8'b11111000; // 1512 : 248 - 0xf8
      13'h5E9: dout <= 8'b11110000; // 1513 : 240 - 0xf0
      13'h5EA: dout <= 8'b11100000; // 1514 : 224 - 0xe0
      13'h5EB: dout <= 8'b11110000; // 1515 : 240 - 0xf0
      13'h5EC: dout <= 8'b11100000; // 1516 : 224 - 0xe0
      13'h5ED: dout <= 8'b11000000; // 1517 : 192 - 0xc0
      13'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      13'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      13'h5F0: dout <= 8'b00000100; // 1520 :   4 - 0x4 -- Sprite 0x5f
      13'h5F1: dout <= 8'b00001100; // 1521 :  12 - 0xc
      13'h5F2: dout <= 8'b00011100; // 1522 :  28 - 0x1c
      13'h5F3: dout <= 8'b00001100; // 1523 :  12 - 0xc
      13'h5F4: dout <= 8'b00011000; // 1524 :  24 - 0x18
      13'h5F5: dout <= 8'b00111100; // 1525 :  60 - 0x3c
      13'h5F6: dout <= 8'b00111100; // 1526 :  60 - 0x3c
      13'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      13'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0
      13'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      13'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      13'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      13'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      13'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      13'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      13'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      13'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0x60
      13'h601: dout <= 8'b00000011; // 1537 :   3 - 0x3
      13'h602: dout <= 8'b00001111; // 1538 :  15 - 0xf
      13'h603: dout <= 8'b00010011; // 1539 :  19 - 0x13
      13'h604: dout <= 8'b00100001; // 1540 :  33 - 0x21
      13'h605: dout <= 8'b00100001; // 1541 :  33 - 0x21
      13'h606: dout <= 8'b00100001; // 1542 :  33 - 0x21
      13'h607: dout <= 8'b01110011; // 1543 : 115 - 0x73
      13'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0
      13'h609: dout <= 8'b00000011; // 1545 :   3 - 0x3
      13'h60A: dout <= 8'b00001111; // 1546 :  15 - 0xf
      13'h60B: dout <= 8'b00011111; // 1547 :  31 - 0x1f
      13'h60C: dout <= 8'b00111111; // 1548 :  63 - 0x3f
      13'h60D: dout <= 8'b00111111; // 1549 :  63 - 0x3f
      13'h60E: dout <= 8'b00111001; // 1550 :  57 - 0x39
      13'h60F: dout <= 8'b01111011; // 1551 : 123 - 0x7b
      13'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0x61
      13'h611: dout <= 8'b11000000; // 1553 : 192 - 0xc0
      13'h612: dout <= 8'b11110000; // 1554 : 240 - 0xf0
      13'h613: dout <= 8'b11001000; // 1555 : 200 - 0xc8
      13'h614: dout <= 8'b10000100; // 1556 : 132 - 0x84
      13'h615: dout <= 8'b10000100; // 1557 : 132 - 0x84
      13'h616: dout <= 8'b10000100; // 1558 : 132 - 0x84
      13'h617: dout <= 8'b11001110; // 1559 : 206 - 0xce
      13'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0
      13'h619: dout <= 8'b11000000; // 1561 : 192 - 0xc0
      13'h61A: dout <= 8'b11110000; // 1562 : 240 - 0xf0
      13'h61B: dout <= 8'b11111000; // 1563 : 248 - 0xf8
      13'h61C: dout <= 8'b11111100; // 1564 : 252 - 0xfc
      13'h61D: dout <= 8'b11111100; // 1565 : 252 - 0xfc
      13'h61E: dout <= 8'b11100100; // 1566 : 228 - 0xe4
      13'h61F: dout <= 8'b11101110; // 1567 : 238 - 0xee
      13'h620: dout <= 8'b10010100; // 1568 : 148 - 0x94 -- Sprite 0x62
      13'h621: dout <= 8'b11101010; // 1569 : 234 - 0xea
      13'h622: dout <= 8'b11011110; // 1570 : 222 - 0xde
      13'h623: dout <= 8'b11101110; // 1571 : 238 - 0xee
      13'h624: dout <= 8'b11011110; // 1572 : 222 - 0xde
      13'h625: dout <= 8'b01100110; // 1573 : 102 - 0x66
      13'h626: dout <= 8'b01000010; // 1574 :  66 - 0x42
      13'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      13'h628: dout <= 8'b11111110; // 1576 : 254 - 0xfe
      13'h629: dout <= 8'b11111110; // 1577 : 254 - 0xfe
      13'h62A: dout <= 8'b11111110; // 1578 : 254 - 0xfe
      13'h62B: dout <= 8'b11111110; // 1579 : 254 - 0xfe
      13'h62C: dout <= 8'b11111110; // 1580 : 254 - 0xfe
      13'h62D: dout <= 8'b01100110; // 1581 : 102 - 0x66
      13'h62E: dout <= 8'b01000010; // 1582 :  66 - 0x42
      13'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      13'h630: dout <= 8'b10010100; // 1584 : 148 - 0x94 -- Sprite 0x63
      13'h631: dout <= 8'b11101010; // 1585 : 234 - 0xea
      13'h632: dout <= 8'b11011110; // 1586 : 222 - 0xde
      13'h633: dout <= 8'b11101110; // 1587 : 238 - 0xee
      13'h634: dout <= 8'b11011110; // 1588 : 222 - 0xde
      13'h635: dout <= 8'b11001110; // 1589 : 206 - 0xce
      13'h636: dout <= 8'b10001100; // 1590 : 140 - 0x8c
      13'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      13'h638: dout <= 8'b11111110; // 1592 : 254 - 0xfe
      13'h639: dout <= 8'b11111110; // 1593 : 254 - 0xfe
      13'h63A: dout <= 8'b11111110; // 1594 : 254 - 0xfe
      13'h63B: dout <= 8'b11111110; // 1595 : 254 - 0xfe
      13'h63C: dout <= 8'b11111110; // 1596 : 254 - 0xfe
      13'h63D: dout <= 8'b11011110; // 1597 : 222 - 0xde
      13'h63E: dout <= 8'b10001100; // 1598 : 140 - 0x8c
      13'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      13'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0x64
      13'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      13'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      13'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      13'h644: dout <= 8'b00000000; // 1604 :   0 - 0x0
      13'h645: dout <= 8'b00000000; // 1605 :   0 - 0x0
      13'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      13'h647: dout <= 8'b00000001; // 1607 :   1 - 0x1
      13'h648: dout <= 8'b00000000; // 1608 :   0 - 0x0
      13'h649: dout <= 8'b00000000; // 1609 :   0 - 0x0
      13'h64A: dout <= 8'b00000000; // 1610 :   0 - 0x0
      13'h64B: dout <= 8'b00000000; // 1611 :   0 - 0x0
      13'h64C: dout <= 8'b00000000; // 1612 :   0 - 0x0
      13'h64D: dout <= 8'b00000000; // 1613 :   0 - 0x0
      13'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      13'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      13'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0x65
      13'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      13'h652: dout <= 8'b00000000; // 1618 :   0 - 0x0
      13'h653: dout <= 8'b00000000; // 1619 :   0 - 0x0
      13'h654: dout <= 8'b00000000; // 1620 :   0 - 0x0
      13'h655: dout <= 8'b00110110; // 1621 :  54 - 0x36
      13'h656: dout <= 8'b00110110; // 1622 :  54 - 0x36
      13'h657: dout <= 8'b10010000; // 1623 : 144 - 0x90
      13'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0
      13'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      13'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      13'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      13'h65C: dout <= 8'b01101100; // 1628 : 108 - 0x6c
      13'h65D: dout <= 8'b11111110; // 1629 : 254 - 0xfe
      13'h65E: dout <= 8'b11111110; // 1630 : 254 - 0xfe
      13'h65F: dout <= 8'b11111100; // 1631 : 252 - 0xfc
      13'h660: dout <= 8'b00000001; // 1632 :   1 - 0x1 -- Sprite 0x66
      13'h661: dout <= 8'b00000011; // 1633 :   3 - 0x3
      13'h662: dout <= 8'b00000111; // 1634 :   7 - 0x7
      13'h663: dout <= 8'b00000111; // 1635 :   7 - 0x7
      13'h664: dout <= 8'b00011111; // 1636 :  31 - 0x1f
      13'h665: dout <= 8'b00011111; // 1637 :  31 - 0x1f
      13'h666: dout <= 8'b00011100; // 1638 :  28 - 0x1c
      13'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      13'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0
      13'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      13'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      13'h66B: dout <= 8'b00000000; // 1643 :   0 - 0x0
      13'h66C: dout <= 8'b00000000; // 1644 :   0 - 0x0
      13'h66D: dout <= 8'b00000000; // 1645 :   0 - 0x0
      13'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      13'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      13'h670: dout <= 8'b11111000; // 1648 : 248 - 0xf8 -- Sprite 0x67
      13'h671: dout <= 8'b11111000; // 1649 : 248 - 0xf8
      13'h672: dout <= 8'b11111000; // 1650 : 248 - 0xf8
      13'h673: dout <= 8'b11111000; // 1651 : 248 - 0xf8
      13'h674: dout <= 8'b11111110; // 1652 : 254 - 0xfe
      13'h675: dout <= 8'b11111110; // 1653 : 254 - 0xfe
      13'h676: dout <= 8'b00001110; // 1654 :  14 - 0xe
      13'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      13'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0
      13'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      13'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      13'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      13'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      13'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      13'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      13'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      13'h680: dout <= 8'b00000111; // 1664 :   7 - 0x7 -- Sprite 0x68
      13'h681: dout <= 8'b00001111; // 1665 :  15 - 0xf
      13'h682: dout <= 8'b00011111; // 1666 :  31 - 0x1f
      13'h683: dout <= 8'b00011111; // 1667 :  31 - 0x1f
      13'h684: dout <= 8'b00111111; // 1668 :  63 - 0x3f
      13'h685: dout <= 8'b00111111; // 1669 :  63 - 0x3f
      13'h686: dout <= 8'b00111000; // 1670 :  56 - 0x38
      13'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      13'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0
      13'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      13'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      13'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      13'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      13'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      13'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      13'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      13'h690: dout <= 8'b11111000; // 1680 : 248 - 0xf8 -- Sprite 0x69
      13'h691: dout <= 8'b11110000; // 1681 : 240 - 0xf0
      13'h692: dout <= 8'b11110000; // 1682 : 240 - 0xf0
      13'h693: dout <= 8'b11100000; // 1683 : 224 - 0xe0
      13'h694: dout <= 8'b11111000; // 1684 : 248 - 0xf8
      13'h695: dout <= 8'b11111000; // 1685 : 248 - 0xf8
      13'h696: dout <= 8'b00111000; // 1686 :  56 - 0x38
      13'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      13'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0
      13'h699: dout <= 8'b00000000; // 1689 :   0 - 0x0
      13'h69A: dout <= 8'b00000000; // 1690 :   0 - 0x0
      13'h69B: dout <= 8'b00000000; // 1691 :   0 - 0x0
      13'h69C: dout <= 8'b00000000; // 1692 :   0 - 0x0
      13'h69D: dout <= 8'b00000000; // 1693 :   0 - 0x0
      13'h69E: dout <= 8'b00000000; // 1694 :   0 - 0x0
      13'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      13'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0x6a
      13'h6A1: dout <= 8'b00011111; // 1697 :  31 - 0x1f
      13'h6A2: dout <= 8'b01111111; // 1698 : 127 - 0x7f
      13'h6A3: dout <= 8'b00111111; // 1699 :  63 - 0x3f
      13'h6A4: dout <= 8'b00001111; // 1700 :  15 - 0xf
      13'h6A5: dout <= 8'b00000111; // 1701 :   7 - 0x7
      13'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      13'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      13'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0
      13'h6A9: dout <= 8'b00011111; // 1705 :  31 - 0x1f
      13'h6AA: dout <= 8'b01111111; // 1706 : 127 - 0x7f
      13'h6AB: dout <= 8'b00111111; // 1707 :  63 - 0x3f
      13'h6AC: dout <= 8'b00001111; // 1708 :  15 - 0xf
      13'h6AD: dout <= 8'b00000111; // 1709 :   7 - 0x7
      13'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      13'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      13'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0x6b
      13'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      13'h6B2: dout <= 8'b11000000; // 1714 : 192 - 0xc0
      13'h6B3: dout <= 8'b11110000; // 1715 : 240 - 0xf0
      13'h6B4: dout <= 8'b11111000; // 1716 : 248 - 0xf8
      13'h6B5: dout <= 8'b11111000; // 1717 : 248 - 0xf8
      13'h6B6: dout <= 8'b11100000; // 1718 : 224 - 0xe0
      13'h6B7: dout <= 8'b00000000; // 1719 :   0 - 0x0
      13'h6B8: dout <= 8'b00000000; // 1720 :   0 - 0x0
      13'h6B9: dout <= 8'b00000000; // 1721 :   0 - 0x0
      13'h6BA: dout <= 8'b11000000; // 1722 : 192 - 0xc0
      13'h6BB: dout <= 8'b11110000; // 1723 : 240 - 0xf0
      13'h6BC: dout <= 8'b11111000; // 1724 : 248 - 0xf8
      13'h6BD: dout <= 8'b11111000; // 1725 : 248 - 0xf8
      13'h6BE: dout <= 8'b11100000; // 1726 : 224 - 0xe0
      13'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      13'h6C0: dout <= 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0x6c
      13'h6C1: dout <= 8'b00000000; // 1729 :   0 - 0x0
      13'h6C2: dout <= 8'b00000000; // 1730 :   0 - 0x0
      13'h6C3: dout <= 8'b00000000; // 1731 :   0 - 0x0
      13'h6C4: dout <= 8'b00000000; // 1732 :   0 - 0x0
      13'h6C5: dout <= 8'b00000000; // 1733 :   0 - 0x0
      13'h6C6: dout <= 8'b00000000; // 1734 :   0 - 0x0
      13'h6C7: dout <= 8'b00000000; // 1735 :   0 - 0x0
      13'h6C8: dout <= 8'b00000000; // 1736 :   0 - 0x0
      13'h6C9: dout <= 8'b00000000; // 1737 :   0 - 0x0
      13'h6CA: dout <= 8'b00000000; // 1738 :   0 - 0x0
      13'h6CB: dout <= 8'b00000000; // 1739 :   0 - 0x0
      13'h6CC: dout <= 8'b00000000; // 1740 :   0 - 0x0
      13'h6CD: dout <= 8'b00000000; // 1741 :   0 - 0x0
      13'h6CE: dout <= 8'b00000000; // 1742 :   0 - 0x0
      13'h6CF: dout <= 8'b00000000; // 1743 :   0 - 0x0
      13'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0x6d
      13'h6D1: dout <= 8'b00000000; // 1745 :   0 - 0x0
      13'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      13'h6D3: dout <= 8'b00000000; // 1747 :   0 - 0x0
      13'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      13'h6D5: dout <= 8'b00000000; // 1749 :   0 - 0x0
      13'h6D6: dout <= 8'b00000000; // 1750 :   0 - 0x0
      13'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      13'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0
      13'h6D9: dout <= 8'b00000000; // 1753 :   0 - 0x0
      13'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      13'h6DB: dout <= 8'b00000000; // 1755 :   0 - 0x0
      13'h6DC: dout <= 8'b00000000; // 1756 :   0 - 0x0
      13'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      13'h6DE: dout <= 8'b00000000; // 1758 :   0 - 0x0
      13'h6DF: dout <= 8'b00000000; // 1759 :   0 - 0x0
      13'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0x6e
      13'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      13'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      13'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      13'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      13'h6E5: dout <= 8'b00000000; // 1765 :   0 - 0x0
      13'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      13'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      13'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0
      13'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      13'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      13'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      13'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      13'h6ED: dout <= 8'b00000000; // 1773 :   0 - 0x0
      13'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      13'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      13'h6F0: dout <= 8'b00000000; // 1776 :   0 - 0x0 -- Sprite 0x6f
      13'h6F1: dout <= 8'b00000000; // 1777 :   0 - 0x0
      13'h6F2: dout <= 8'b00000000; // 1778 :   0 - 0x0
      13'h6F3: dout <= 8'b00000000; // 1779 :   0 - 0x0
      13'h6F4: dout <= 8'b00000000; // 1780 :   0 - 0x0
      13'h6F5: dout <= 8'b00000000; // 1781 :   0 - 0x0
      13'h6F6: dout <= 8'b00000000; // 1782 :   0 - 0x0
      13'h6F7: dout <= 8'b00000000; // 1783 :   0 - 0x0
      13'h6F8: dout <= 8'b00000000; // 1784 :   0 - 0x0
      13'h6F9: dout <= 8'b00000000; // 1785 :   0 - 0x0
      13'h6FA: dout <= 8'b00000000; // 1786 :   0 - 0x0
      13'h6FB: dout <= 8'b00000000; // 1787 :   0 - 0x0
      13'h6FC: dout <= 8'b00000000; // 1788 :   0 - 0x0
      13'h6FD: dout <= 8'b00000000; // 1789 :   0 - 0x0
      13'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      13'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      13'h700: dout <= 8'b11111111; // 1792 : 255 - 0xff -- Sprite 0x70
      13'h701: dout <= 8'b11111111; // 1793 : 255 - 0xff
      13'h702: dout <= 8'b11111111; // 1794 : 255 - 0xff
      13'h703: dout <= 8'b11111111; // 1795 : 255 - 0xff
      13'h704: dout <= 8'b11111111; // 1796 : 255 - 0xff
      13'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      13'h706: dout <= 8'b11111111; // 1798 : 255 - 0xff
      13'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      13'h708: dout <= 8'b11111111; // 1800 : 255 - 0xff
      13'h709: dout <= 8'b11111111; // 1801 : 255 - 0xff
      13'h70A: dout <= 8'b11111111; // 1802 : 255 - 0xff
      13'h70B: dout <= 8'b11111111; // 1803 : 255 - 0xff
      13'h70C: dout <= 8'b11111111; // 1804 : 255 - 0xff
      13'h70D: dout <= 8'b11111111; // 1805 : 255 - 0xff
      13'h70E: dout <= 8'b11111111; // 1806 : 255 - 0xff
      13'h70F: dout <= 8'b11111111; // 1807 : 255 - 0xff
      13'h710: dout <= 8'b11111111; // 1808 : 255 - 0xff -- Sprite 0x71
      13'h711: dout <= 8'b11111111; // 1809 : 255 - 0xff
      13'h712: dout <= 8'b11111111; // 1810 : 255 - 0xff
      13'h713: dout <= 8'b11111111; // 1811 : 255 - 0xff
      13'h714: dout <= 8'b11111111; // 1812 : 255 - 0xff
      13'h715: dout <= 8'b11111111; // 1813 : 255 - 0xff
      13'h716: dout <= 8'b11111111; // 1814 : 255 - 0xff
      13'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      13'h718: dout <= 8'b11111111; // 1816 : 255 - 0xff
      13'h719: dout <= 8'b11111111; // 1817 : 255 - 0xff
      13'h71A: dout <= 8'b11111111; // 1818 : 255 - 0xff
      13'h71B: dout <= 8'b11111111; // 1819 : 255 - 0xff
      13'h71C: dout <= 8'b11111111; // 1820 : 255 - 0xff
      13'h71D: dout <= 8'b11111111; // 1821 : 255 - 0xff
      13'h71E: dout <= 8'b11111111; // 1822 : 255 - 0xff
      13'h71F: dout <= 8'b11111111; // 1823 : 255 - 0xff
      13'h720: dout <= 8'b11111111; // 1824 : 255 - 0xff -- Sprite 0x72
      13'h721: dout <= 8'b11111111; // 1825 : 255 - 0xff
      13'h722: dout <= 8'b11111111; // 1826 : 255 - 0xff
      13'h723: dout <= 8'b11111111; // 1827 : 255 - 0xff
      13'h724: dout <= 8'b11111111; // 1828 : 255 - 0xff
      13'h725: dout <= 8'b11111111; // 1829 : 255 - 0xff
      13'h726: dout <= 8'b11111111; // 1830 : 255 - 0xff
      13'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      13'h728: dout <= 8'b11111111; // 1832 : 255 - 0xff
      13'h729: dout <= 8'b11111111; // 1833 : 255 - 0xff
      13'h72A: dout <= 8'b11111111; // 1834 : 255 - 0xff
      13'h72B: dout <= 8'b11111111; // 1835 : 255 - 0xff
      13'h72C: dout <= 8'b11111111; // 1836 : 255 - 0xff
      13'h72D: dout <= 8'b11111111; // 1837 : 255 - 0xff
      13'h72E: dout <= 8'b11111111; // 1838 : 255 - 0xff
      13'h72F: dout <= 8'b11111111; // 1839 : 255 - 0xff
      13'h730: dout <= 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0x73
      13'h731: dout <= 8'b11111111; // 1841 : 255 - 0xff
      13'h732: dout <= 8'b11111111; // 1842 : 255 - 0xff
      13'h733: dout <= 8'b11111111; // 1843 : 255 - 0xff
      13'h734: dout <= 8'b11111111; // 1844 : 255 - 0xff
      13'h735: dout <= 8'b11111111; // 1845 : 255 - 0xff
      13'h736: dout <= 8'b11111111; // 1846 : 255 - 0xff
      13'h737: dout <= 8'b11111111; // 1847 : 255 - 0xff
      13'h738: dout <= 8'b11111111; // 1848 : 255 - 0xff
      13'h739: dout <= 8'b11111111; // 1849 : 255 - 0xff
      13'h73A: dout <= 8'b11111111; // 1850 : 255 - 0xff
      13'h73B: dout <= 8'b11111111; // 1851 : 255 - 0xff
      13'h73C: dout <= 8'b11111111; // 1852 : 255 - 0xff
      13'h73D: dout <= 8'b11111111; // 1853 : 255 - 0xff
      13'h73E: dout <= 8'b11111111; // 1854 : 255 - 0xff
      13'h73F: dout <= 8'b11111111; // 1855 : 255 - 0xff
      13'h740: dout <= 8'b11111111; // 1856 : 255 - 0xff -- Sprite 0x74
      13'h741: dout <= 8'b11111111; // 1857 : 255 - 0xff
      13'h742: dout <= 8'b11111111; // 1858 : 255 - 0xff
      13'h743: dout <= 8'b11111111; // 1859 : 255 - 0xff
      13'h744: dout <= 8'b11111111; // 1860 : 255 - 0xff
      13'h745: dout <= 8'b11111111; // 1861 : 255 - 0xff
      13'h746: dout <= 8'b11111111; // 1862 : 255 - 0xff
      13'h747: dout <= 8'b11111111; // 1863 : 255 - 0xff
      13'h748: dout <= 8'b11111111; // 1864 : 255 - 0xff
      13'h749: dout <= 8'b11111111; // 1865 : 255 - 0xff
      13'h74A: dout <= 8'b11111111; // 1866 : 255 - 0xff
      13'h74B: dout <= 8'b11111111; // 1867 : 255 - 0xff
      13'h74C: dout <= 8'b11111111; // 1868 : 255 - 0xff
      13'h74D: dout <= 8'b11111111; // 1869 : 255 - 0xff
      13'h74E: dout <= 8'b11111111; // 1870 : 255 - 0xff
      13'h74F: dout <= 8'b11111111; // 1871 : 255 - 0xff
      13'h750: dout <= 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0x75
      13'h751: dout <= 8'b11111111; // 1873 : 255 - 0xff
      13'h752: dout <= 8'b11111111; // 1874 : 255 - 0xff
      13'h753: dout <= 8'b11111111; // 1875 : 255 - 0xff
      13'h754: dout <= 8'b11111111; // 1876 : 255 - 0xff
      13'h755: dout <= 8'b11111111; // 1877 : 255 - 0xff
      13'h756: dout <= 8'b11111111; // 1878 : 255 - 0xff
      13'h757: dout <= 8'b11111111; // 1879 : 255 - 0xff
      13'h758: dout <= 8'b11111111; // 1880 : 255 - 0xff
      13'h759: dout <= 8'b11111111; // 1881 : 255 - 0xff
      13'h75A: dout <= 8'b11111111; // 1882 : 255 - 0xff
      13'h75B: dout <= 8'b11111111; // 1883 : 255 - 0xff
      13'h75C: dout <= 8'b11111111; // 1884 : 255 - 0xff
      13'h75D: dout <= 8'b11111111; // 1885 : 255 - 0xff
      13'h75E: dout <= 8'b11111111; // 1886 : 255 - 0xff
      13'h75F: dout <= 8'b11111111; // 1887 : 255 - 0xff
      13'h760: dout <= 8'b11111111; // 1888 : 255 - 0xff -- Sprite 0x76
      13'h761: dout <= 8'b11111111; // 1889 : 255 - 0xff
      13'h762: dout <= 8'b11111111; // 1890 : 255 - 0xff
      13'h763: dout <= 8'b11111111; // 1891 : 255 - 0xff
      13'h764: dout <= 8'b11111111; // 1892 : 255 - 0xff
      13'h765: dout <= 8'b11111111; // 1893 : 255 - 0xff
      13'h766: dout <= 8'b11111111; // 1894 : 255 - 0xff
      13'h767: dout <= 8'b11111111; // 1895 : 255 - 0xff
      13'h768: dout <= 8'b11111111; // 1896 : 255 - 0xff
      13'h769: dout <= 8'b11111111; // 1897 : 255 - 0xff
      13'h76A: dout <= 8'b11111111; // 1898 : 255 - 0xff
      13'h76B: dout <= 8'b11111111; // 1899 : 255 - 0xff
      13'h76C: dout <= 8'b11111111; // 1900 : 255 - 0xff
      13'h76D: dout <= 8'b11111111; // 1901 : 255 - 0xff
      13'h76E: dout <= 8'b11111111; // 1902 : 255 - 0xff
      13'h76F: dout <= 8'b11111111; // 1903 : 255 - 0xff
      13'h770: dout <= 8'b11111111; // 1904 : 255 - 0xff -- Sprite 0x77
      13'h771: dout <= 8'b11111111; // 1905 : 255 - 0xff
      13'h772: dout <= 8'b11111111; // 1906 : 255 - 0xff
      13'h773: dout <= 8'b11111111; // 1907 : 255 - 0xff
      13'h774: dout <= 8'b11111111; // 1908 : 255 - 0xff
      13'h775: dout <= 8'b11111111; // 1909 : 255 - 0xff
      13'h776: dout <= 8'b11111111; // 1910 : 255 - 0xff
      13'h777: dout <= 8'b11111111; // 1911 : 255 - 0xff
      13'h778: dout <= 8'b11111111; // 1912 : 255 - 0xff
      13'h779: dout <= 8'b11111111; // 1913 : 255 - 0xff
      13'h77A: dout <= 8'b11111111; // 1914 : 255 - 0xff
      13'h77B: dout <= 8'b11111111; // 1915 : 255 - 0xff
      13'h77C: dout <= 8'b11111111; // 1916 : 255 - 0xff
      13'h77D: dout <= 8'b11111111; // 1917 : 255 - 0xff
      13'h77E: dout <= 8'b11111111; // 1918 : 255 - 0xff
      13'h77F: dout <= 8'b11111111; // 1919 : 255 - 0xff
      13'h780: dout <= 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0x78
      13'h781: dout <= 8'b11111111; // 1921 : 255 - 0xff
      13'h782: dout <= 8'b11111111; // 1922 : 255 - 0xff
      13'h783: dout <= 8'b11111111; // 1923 : 255 - 0xff
      13'h784: dout <= 8'b11111111; // 1924 : 255 - 0xff
      13'h785: dout <= 8'b11111111; // 1925 : 255 - 0xff
      13'h786: dout <= 8'b11111111; // 1926 : 255 - 0xff
      13'h787: dout <= 8'b11111111; // 1927 : 255 - 0xff
      13'h788: dout <= 8'b11111111; // 1928 : 255 - 0xff
      13'h789: dout <= 8'b11111111; // 1929 : 255 - 0xff
      13'h78A: dout <= 8'b11111111; // 1930 : 255 - 0xff
      13'h78B: dout <= 8'b11111111; // 1931 : 255 - 0xff
      13'h78C: dout <= 8'b11111111; // 1932 : 255 - 0xff
      13'h78D: dout <= 8'b11111111; // 1933 : 255 - 0xff
      13'h78E: dout <= 8'b11111111; // 1934 : 255 - 0xff
      13'h78F: dout <= 8'b11111111; // 1935 : 255 - 0xff
      13'h790: dout <= 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0x79
      13'h791: dout <= 8'b11111111; // 1937 : 255 - 0xff
      13'h792: dout <= 8'b11111111; // 1938 : 255 - 0xff
      13'h793: dout <= 8'b11111111; // 1939 : 255 - 0xff
      13'h794: dout <= 8'b11111111; // 1940 : 255 - 0xff
      13'h795: dout <= 8'b11111111; // 1941 : 255 - 0xff
      13'h796: dout <= 8'b11111111; // 1942 : 255 - 0xff
      13'h797: dout <= 8'b11111111; // 1943 : 255 - 0xff
      13'h798: dout <= 8'b11111111; // 1944 : 255 - 0xff
      13'h799: dout <= 8'b11111111; // 1945 : 255 - 0xff
      13'h79A: dout <= 8'b11111111; // 1946 : 255 - 0xff
      13'h79B: dout <= 8'b11111111; // 1947 : 255 - 0xff
      13'h79C: dout <= 8'b11111111; // 1948 : 255 - 0xff
      13'h79D: dout <= 8'b11111111; // 1949 : 255 - 0xff
      13'h79E: dout <= 8'b11111111; // 1950 : 255 - 0xff
      13'h79F: dout <= 8'b11111111; // 1951 : 255 - 0xff
      13'h7A0: dout <= 8'b11111111; // 1952 : 255 - 0xff -- Sprite 0x7a
      13'h7A1: dout <= 8'b11111111; // 1953 : 255 - 0xff
      13'h7A2: dout <= 8'b11111111; // 1954 : 255 - 0xff
      13'h7A3: dout <= 8'b11111111; // 1955 : 255 - 0xff
      13'h7A4: dout <= 8'b11111111; // 1956 : 255 - 0xff
      13'h7A5: dout <= 8'b11111111; // 1957 : 255 - 0xff
      13'h7A6: dout <= 8'b11111111; // 1958 : 255 - 0xff
      13'h7A7: dout <= 8'b11111111; // 1959 : 255 - 0xff
      13'h7A8: dout <= 8'b11111111; // 1960 : 255 - 0xff
      13'h7A9: dout <= 8'b11111111; // 1961 : 255 - 0xff
      13'h7AA: dout <= 8'b11111111; // 1962 : 255 - 0xff
      13'h7AB: dout <= 8'b11111111; // 1963 : 255 - 0xff
      13'h7AC: dout <= 8'b11111111; // 1964 : 255 - 0xff
      13'h7AD: dout <= 8'b11111111; // 1965 : 255 - 0xff
      13'h7AE: dout <= 8'b11111111; // 1966 : 255 - 0xff
      13'h7AF: dout <= 8'b11111111; // 1967 : 255 - 0xff
      13'h7B0: dout <= 8'b11111111; // 1968 : 255 - 0xff -- Sprite 0x7b
      13'h7B1: dout <= 8'b11111111; // 1969 : 255 - 0xff
      13'h7B2: dout <= 8'b11111111; // 1970 : 255 - 0xff
      13'h7B3: dout <= 8'b11111111; // 1971 : 255 - 0xff
      13'h7B4: dout <= 8'b11111111; // 1972 : 255 - 0xff
      13'h7B5: dout <= 8'b11111111; // 1973 : 255 - 0xff
      13'h7B6: dout <= 8'b11111111; // 1974 : 255 - 0xff
      13'h7B7: dout <= 8'b11111111; // 1975 : 255 - 0xff
      13'h7B8: dout <= 8'b11111111; // 1976 : 255 - 0xff
      13'h7B9: dout <= 8'b11111111; // 1977 : 255 - 0xff
      13'h7BA: dout <= 8'b11111111; // 1978 : 255 - 0xff
      13'h7BB: dout <= 8'b11111111; // 1979 : 255 - 0xff
      13'h7BC: dout <= 8'b11111111; // 1980 : 255 - 0xff
      13'h7BD: dout <= 8'b11111111; // 1981 : 255 - 0xff
      13'h7BE: dout <= 8'b11111111; // 1982 : 255 - 0xff
      13'h7BF: dout <= 8'b11111111; // 1983 : 255 - 0xff
      13'h7C0: dout <= 8'b11111111; // 1984 : 255 - 0xff -- Sprite 0x7c
      13'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      13'h7C2: dout <= 8'b11111111; // 1986 : 255 - 0xff
      13'h7C3: dout <= 8'b11111111; // 1987 : 255 - 0xff
      13'h7C4: dout <= 8'b11111111; // 1988 : 255 - 0xff
      13'h7C5: dout <= 8'b11111111; // 1989 : 255 - 0xff
      13'h7C6: dout <= 8'b11111111; // 1990 : 255 - 0xff
      13'h7C7: dout <= 8'b11111111; // 1991 : 255 - 0xff
      13'h7C8: dout <= 8'b11111111; // 1992 : 255 - 0xff
      13'h7C9: dout <= 8'b11111111; // 1993 : 255 - 0xff
      13'h7CA: dout <= 8'b11111111; // 1994 : 255 - 0xff
      13'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      13'h7CC: dout <= 8'b11111111; // 1996 : 255 - 0xff
      13'h7CD: dout <= 8'b11111111; // 1997 : 255 - 0xff
      13'h7CE: dout <= 8'b11111111; // 1998 : 255 - 0xff
      13'h7CF: dout <= 8'b11111111; // 1999 : 255 - 0xff
      13'h7D0: dout <= 8'b11111111; // 2000 : 255 - 0xff -- Sprite 0x7d
      13'h7D1: dout <= 8'b11111111; // 2001 : 255 - 0xff
      13'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      13'h7D3: dout <= 8'b11111111; // 2003 : 255 - 0xff
      13'h7D4: dout <= 8'b11111111; // 2004 : 255 - 0xff
      13'h7D5: dout <= 8'b11111111; // 2005 : 255 - 0xff
      13'h7D6: dout <= 8'b11111111; // 2006 : 255 - 0xff
      13'h7D7: dout <= 8'b11111111; // 2007 : 255 - 0xff
      13'h7D8: dout <= 8'b11111111; // 2008 : 255 - 0xff
      13'h7D9: dout <= 8'b11111111; // 2009 : 255 - 0xff
      13'h7DA: dout <= 8'b11111111; // 2010 : 255 - 0xff
      13'h7DB: dout <= 8'b11111111; // 2011 : 255 - 0xff
      13'h7DC: dout <= 8'b11111111; // 2012 : 255 - 0xff
      13'h7DD: dout <= 8'b11111111; // 2013 : 255 - 0xff
      13'h7DE: dout <= 8'b11111111; // 2014 : 255 - 0xff
      13'h7DF: dout <= 8'b11111111; // 2015 : 255 - 0xff
      13'h7E0: dout <= 8'b11111111; // 2016 : 255 - 0xff -- Sprite 0x7e
      13'h7E1: dout <= 8'b11111111; // 2017 : 255 - 0xff
      13'h7E2: dout <= 8'b11111111; // 2018 : 255 - 0xff
      13'h7E3: dout <= 8'b11111111; // 2019 : 255 - 0xff
      13'h7E4: dout <= 8'b11111111; // 2020 : 255 - 0xff
      13'h7E5: dout <= 8'b11111111; // 2021 : 255 - 0xff
      13'h7E6: dout <= 8'b11111111; // 2022 : 255 - 0xff
      13'h7E7: dout <= 8'b11111111; // 2023 : 255 - 0xff
      13'h7E8: dout <= 8'b11111111; // 2024 : 255 - 0xff
      13'h7E9: dout <= 8'b11111111; // 2025 : 255 - 0xff
      13'h7EA: dout <= 8'b11111111; // 2026 : 255 - 0xff
      13'h7EB: dout <= 8'b11111111; // 2027 : 255 - 0xff
      13'h7EC: dout <= 8'b11111111; // 2028 : 255 - 0xff
      13'h7ED: dout <= 8'b11111111; // 2029 : 255 - 0xff
      13'h7EE: dout <= 8'b11111111; // 2030 : 255 - 0xff
      13'h7EF: dout <= 8'b11111111; // 2031 : 255 - 0xff
      13'h7F0: dout <= 8'b11111111; // 2032 : 255 - 0xff -- Sprite 0x7f
      13'h7F1: dout <= 8'b11111111; // 2033 : 255 - 0xff
      13'h7F2: dout <= 8'b11111111; // 2034 : 255 - 0xff
      13'h7F3: dout <= 8'b11111111; // 2035 : 255 - 0xff
      13'h7F4: dout <= 8'b11111111; // 2036 : 255 - 0xff
      13'h7F5: dout <= 8'b11111111; // 2037 : 255 - 0xff
      13'h7F6: dout <= 8'b11111111; // 2038 : 255 - 0xff
      13'h7F7: dout <= 8'b11111111; // 2039 : 255 - 0xff
      13'h7F8: dout <= 8'b11111111; // 2040 : 255 - 0xff
      13'h7F9: dout <= 8'b11111111; // 2041 : 255 - 0xff
      13'h7FA: dout <= 8'b11111111; // 2042 : 255 - 0xff
      13'h7FB: dout <= 8'b11111111; // 2043 : 255 - 0xff
      13'h7FC: dout <= 8'b11111111; // 2044 : 255 - 0xff
      13'h7FD: dout <= 8'b11111111; // 2045 : 255 - 0xff
      13'h7FE: dout <= 8'b11111111; // 2046 : 255 - 0xff
      13'h7FF: dout <= 8'b11111111; // 2047 : 255 - 0xff
      13'h800: dout <= 8'b11111111; // 2048 : 255 - 0xff -- Sprite 0x80
      13'h801: dout <= 8'b11111111; // 2049 : 255 - 0xff
      13'h802: dout <= 8'b11111111; // 2050 : 255 - 0xff
      13'h803: dout <= 8'b11111111; // 2051 : 255 - 0xff
      13'h804: dout <= 8'b11111111; // 2052 : 255 - 0xff
      13'h805: dout <= 8'b11111111; // 2053 : 255 - 0xff
      13'h806: dout <= 8'b11111111; // 2054 : 255 - 0xff
      13'h807: dout <= 8'b11111111; // 2055 : 255 - 0xff
      13'h808: dout <= 8'b11111111; // 2056 : 255 - 0xff
      13'h809: dout <= 8'b11111111; // 2057 : 255 - 0xff
      13'h80A: dout <= 8'b11111111; // 2058 : 255 - 0xff
      13'h80B: dout <= 8'b11111111; // 2059 : 255 - 0xff
      13'h80C: dout <= 8'b11111111; // 2060 : 255 - 0xff
      13'h80D: dout <= 8'b11111111; // 2061 : 255 - 0xff
      13'h80E: dout <= 8'b11111111; // 2062 : 255 - 0xff
      13'h80F: dout <= 8'b11111111; // 2063 : 255 - 0xff
      13'h810: dout <= 8'b11111111; // 2064 : 255 - 0xff -- Sprite 0x81
      13'h811: dout <= 8'b11111111; // 2065 : 255 - 0xff
      13'h812: dout <= 8'b11111111; // 2066 : 255 - 0xff
      13'h813: dout <= 8'b11111111; // 2067 : 255 - 0xff
      13'h814: dout <= 8'b11111111; // 2068 : 255 - 0xff
      13'h815: dout <= 8'b11111111; // 2069 : 255 - 0xff
      13'h816: dout <= 8'b11111111; // 2070 : 255 - 0xff
      13'h817: dout <= 8'b11111111; // 2071 : 255 - 0xff
      13'h818: dout <= 8'b11111111; // 2072 : 255 - 0xff
      13'h819: dout <= 8'b11111111; // 2073 : 255 - 0xff
      13'h81A: dout <= 8'b11111111; // 2074 : 255 - 0xff
      13'h81B: dout <= 8'b11111111; // 2075 : 255 - 0xff
      13'h81C: dout <= 8'b11111111; // 2076 : 255 - 0xff
      13'h81D: dout <= 8'b11111111; // 2077 : 255 - 0xff
      13'h81E: dout <= 8'b11111111; // 2078 : 255 - 0xff
      13'h81F: dout <= 8'b11111111; // 2079 : 255 - 0xff
      13'h820: dout <= 8'b11111111; // 2080 : 255 - 0xff -- Sprite 0x82
      13'h821: dout <= 8'b11111111; // 2081 : 255 - 0xff
      13'h822: dout <= 8'b11111111; // 2082 : 255 - 0xff
      13'h823: dout <= 8'b11111111; // 2083 : 255 - 0xff
      13'h824: dout <= 8'b11111111; // 2084 : 255 - 0xff
      13'h825: dout <= 8'b11111111; // 2085 : 255 - 0xff
      13'h826: dout <= 8'b11111111; // 2086 : 255 - 0xff
      13'h827: dout <= 8'b11111111; // 2087 : 255 - 0xff
      13'h828: dout <= 8'b11111111; // 2088 : 255 - 0xff
      13'h829: dout <= 8'b11111111; // 2089 : 255 - 0xff
      13'h82A: dout <= 8'b11111111; // 2090 : 255 - 0xff
      13'h82B: dout <= 8'b11111111; // 2091 : 255 - 0xff
      13'h82C: dout <= 8'b11111111; // 2092 : 255 - 0xff
      13'h82D: dout <= 8'b11111111; // 2093 : 255 - 0xff
      13'h82E: dout <= 8'b11111111; // 2094 : 255 - 0xff
      13'h82F: dout <= 8'b11111111; // 2095 : 255 - 0xff
      13'h830: dout <= 8'b11111111; // 2096 : 255 - 0xff -- Sprite 0x83
      13'h831: dout <= 8'b11111111; // 2097 : 255 - 0xff
      13'h832: dout <= 8'b11111111; // 2098 : 255 - 0xff
      13'h833: dout <= 8'b11111111; // 2099 : 255 - 0xff
      13'h834: dout <= 8'b11111111; // 2100 : 255 - 0xff
      13'h835: dout <= 8'b11111111; // 2101 : 255 - 0xff
      13'h836: dout <= 8'b11111111; // 2102 : 255 - 0xff
      13'h837: dout <= 8'b11111111; // 2103 : 255 - 0xff
      13'h838: dout <= 8'b11111111; // 2104 : 255 - 0xff
      13'h839: dout <= 8'b11111111; // 2105 : 255 - 0xff
      13'h83A: dout <= 8'b11111111; // 2106 : 255 - 0xff
      13'h83B: dout <= 8'b11111111; // 2107 : 255 - 0xff
      13'h83C: dout <= 8'b11111111; // 2108 : 255 - 0xff
      13'h83D: dout <= 8'b11111111; // 2109 : 255 - 0xff
      13'h83E: dout <= 8'b11111111; // 2110 : 255 - 0xff
      13'h83F: dout <= 8'b11111111; // 2111 : 255 - 0xff
      13'h840: dout <= 8'b11111111; // 2112 : 255 - 0xff -- Sprite 0x84
      13'h841: dout <= 8'b11111111; // 2113 : 255 - 0xff
      13'h842: dout <= 8'b11111111; // 2114 : 255 - 0xff
      13'h843: dout <= 8'b11111111; // 2115 : 255 - 0xff
      13'h844: dout <= 8'b11111111; // 2116 : 255 - 0xff
      13'h845: dout <= 8'b11111111; // 2117 : 255 - 0xff
      13'h846: dout <= 8'b11111111; // 2118 : 255 - 0xff
      13'h847: dout <= 8'b11111111; // 2119 : 255 - 0xff
      13'h848: dout <= 8'b11111111; // 2120 : 255 - 0xff
      13'h849: dout <= 8'b11111111; // 2121 : 255 - 0xff
      13'h84A: dout <= 8'b11111111; // 2122 : 255 - 0xff
      13'h84B: dout <= 8'b11111111; // 2123 : 255 - 0xff
      13'h84C: dout <= 8'b11111111; // 2124 : 255 - 0xff
      13'h84D: dout <= 8'b11111111; // 2125 : 255 - 0xff
      13'h84E: dout <= 8'b11111111; // 2126 : 255 - 0xff
      13'h84F: dout <= 8'b11111111; // 2127 : 255 - 0xff
      13'h850: dout <= 8'b11111111; // 2128 : 255 - 0xff -- Sprite 0x85
      13'h851: dout <= 8'b11111111; // 2129 : 255 - 0xff
      13'h852: dout <= 8'b11111111; // 2130 : 255 - 0xff
      13'h853: dout <= 8'b11111111; // 2131 : 255 - 0xff
      13'h854: dout <= 8'b11111111; // 2132 : 255 - 0xff
      13'h855: dout <= 8'b11111111; // 2133 : 255 - 0xff
      13'h856: dout <= 8'b11111111; // 2134 : 255 - 0xff
      13'h857: dout <= 8'b11111111; // 2135 : 255 - 0xff
      13'h858: dout <= 8'b11111111; // 2136 : 255 - 0xff
      13'h859: dout <= 8'b11111111; // 2137 : 255 - 0xff
      13'h85A: dout <= 8'b11111111; // 2138 : 255 - 0xff
      13'h85B: dout <= 8'b11111111; // 2139 : 255 - 0xff
      13'h85C: dout <= 8'b11111111; // 2140 : 255 - 0xff
      13'h85D: dout <= 8'b11111111; // 2141 : 255 - 0xff
      13'h85E: dout <= 8'b11111111; // 2142 : 255 - 0xff
      13'h85F: dout <= 8'b11111111; // 2143 : 255 - 0xff
      13'h860: dout <= 8'b11111111; // 2144 : 255 - 0xff -- Sprite 0x86
      13'h861: dout <= 8'b11111111; // 2145 : 255 - 0xff
      13'h862: dout <= 8'b11111111; // 2146 : 255 - 0xff
      13'h863: dout <= 8'b11111111; // 2147 : 255 - 0xff
      13'h864: dout <= 8'b11111111; // 2148 : 255 - 0xff
      13'h865: dout <= 8'b11111111; // 2149 : 255 - 0xff
      13'h866: dout <= 8'b11111111; // 2150 : 255 - 0xff
      13'h867: dout <= 8'b11111111; // 2151 : 255 - 0xff
      13'h868: dout <= 8'b11111111; // 2152 : 255 - 0xff
      13'h869: dout <= 8'b11111111; // 2153 : 255 - 0xff
      13'h86A: dout <= 8'b11111111; // 2154 : 255 - 0xff
      13'h86B: dout <= 8'b11111111; // 2155 : 255 - 0xff
      13'h86C: dout <= 8'b11111111; // 2156 : 255 - 0xff
      13'h86D: dout <= 8'b11111111; // 2157 : 255 - 0xff
      13'h86E: dout <= 8'b11111111; // 2158 : 255 - 0xff
      13'h86F: dout <= 8'b11111111; // 2159 : 255 - 0xff
      13'h870: dout <= 8'b11111111; // 2160 : 255 - 0xff -- Sprite 0x87
      13'h871: dout <= 8'b11111111; // 2161 : 255 - 0xff
      13'h872: dout <= 8'b11111111; // 2162 : 255 - 0xff
      13'h873: dout <= 8'b11111111; // 2163 : 255 - 0xff
      13'h874: dout <= 8'b11111111; // 2164 : 255 - 0xff
      13'h875: dout <= 8'b11111111; // 2165 : 255 - 0xff
      13'h876: dout <= 8'b11111111; // 2166 : 255 - 0xff
      13'h877: dout <= 8'b11111111; // 2167 : 255 - 0xff
      13'h878: dout <= 8'b11111111; // 2168 : 255 - 0xff
      13'h879: dout <= 8'b11111111; // 2169 : 255 - 0xff
      13'h87A: dout <= 8'b11111111; // 2170 : 255 - 0xff
      13'h87B: dout <= 8'b11111111; // 2171 : 255 - 0xff
      13'h87C: dout <= 8'b11111111; // 2172 : 255 - 0xff
      13'h87D: dout <= 8'b11111111; // 2173 : 255 - 0xff
      13'h87E: dout <= 8'b11111111; // 2174 : 255 - 0xff
      13'h87F: dout <= 8'b11111111; // 2175 : 255 - 0xff
      13'h880: dout <= 8'b11111111; // 2176 : 255 - 0xff -- Sprite 0x88
      13'h881: dout <= 8'b11111111; // 2177 : 255 - 0xff
      13'h882: dout <= 8'b11111111; // 2178 : 255 - 0xff
      13'h883: dout <= 8'b11111111; // 2179 : 255 - 0xff
      13'h884: dout <= 8'b11111111; // 2180 : 255 - 0xff
      13'h885: dout <= 8'b11111111; // 2181 : 255 - 0xff
      13'h886: dout <= 8'b11111111; // 2182 : 255 - 0xff
      13'h887: dout <= 8'b11111111; // 2183 : 255 - 0xff
      13'h888: dout <= 8'b11111111; // 2184 : 255 - 0xff
      13'h889: dout <= 8'b11111111; // 2185 : 255 - 0xff
      13'h88A: dout <= 8'b11111111; // 2186 : 255 - 0xff
      13'h88B: dout <= 8'b11111111; // 2187 : 255 - 0xff
      13'h88C: dout <= 8'b11111111; // 2188 : 255 - 0xff
      13'h88D: dout <= 8'b11111111; // 2189 : 255 - 0xff
      13'h88E: dout <= 8'b11111111; // 2190 : 255 - 0xff
      13'h88F: dout <= 8'b11111111; // 2191 : 255 - 0xff
      13'h890: dout <= 8'b11111111; // 2192 : 255 - 0xff -- Sprite 0x89
      13'h891: dout <= 8'b11111111; // 2193 : 255 - 0xff
      13'h892: dout <= 8'b11111111; // 2194 : 255 - 0xff
      13'h893: dout <= 8'b11111111; // 2195 : 255 - 0xff
      13'h894: dout <= 8'b11111111; // 2196 : 255 - 0xff
      13'h895: dout <= 8'b11111111; // 2197 : 255 - 0xff
      13'h896: dout <= 8'b11111111; // 2198 : 255 - 0xff
      13'h897: dout <= 8'b11111111; // 2199 : 255 - 0xff
      13'h898: dout <= 8'b11111111; // 2200 : 255 - 0xff
      13'h899: dout <= 8'b11111111; // 2201 : 255 - 0xff
      13'h89A: dout <= 8'b11111111; // 2202 : 255 - 0xff
      13'h89B: dout <= 8'b11111111; // 2203 : 255 - 0xff
      13'h89C: dout <= 8'b11111111; // 2204 : 255 - 0xff
      13'h89D: dout <= 8'b11111111; // 2205 : 255 - 0xff
      13'h89E: dout <= 8'b11111111; // 2206 : 255 - 0xff
      13'h89F: dout <= 8'b11111111; // 2207 : 255 - 0xff
      13'h8A0: dout <= 8'b11111111; // 2208 : 255 - 0xff -- Sprite 0x8a
      13'h8A1: dout <= 8'b11111111; // 2209 : 255 - 0xff
      13'h8A2: dout <= 8'b11111111; // 2210 : 255 - 0xff
      13'h8A3: dout <= 8'b11111111; // 2211 : 255 - 0xff
      13'h8A4: dout <= 8'b11111111; // 2212 : 255 - 0xff
      13'h8A5: dout <= 8'b11111111; // 2213 : 255 - 0xff
      13'h8A6: dout <= 8'b11111111; // 2214 : 255 - 0xff
      13'h8A7: dout <= 8'b11111111; // 2215 : 255 - 0xff
      13'h8A8: dout <= 8'b11111111; // 2216 : 255 - 0xff
      13'h8A9: dout <= 8'b11111111; // 2217 : 255 - 0xff
      13'h8AA: dout <= 8'b11111111; // 2218 : 255 - 0xff
      13'h8AB: dout <= 8'b11111111; // 2219 : 255 - 0xff
      13'h8AC: dout <= 8'b11111111; // 2220 : 255 - 0xff
      13'h8AD: dout <= 8'b11111111; // 2221 : 255 - 0xff
      13'h8AE: dout <= 8'b11111111; // 2222 : 255 - 0xff
      13'h8AF: dout <= 8'b11111111; // 2223 : 255 - 0xff
      13'h8B0: dout <= 8'b11111111; // 2224 : 255 - 0xff -- Sprite 0x8b
      13'h8B1: dout <= 8'b11111111; // 2225 : 255 - 0xff
      13'h8B2: dout <= 8'b11111111; // 2226 : 255 - 0xff
      13'h8B3: dout <= 8'b11111111; // 2227 : 255 - 0xff
      13'h8B4: dout <= 8'b11111111; // 2228 : 255 - 0xff
      13'h8B5: dout <= 8'b11111111; // 2229 : 255 - 0xff
      13'h8B6: dout <= 8'b11111111; // 2230 : 255 - 0xff
      13'h8B7: dout <= 8'b11111111; // 2231 : 255 - 0xff
      13'h8B8: dout <= 8'b11111111; // 2232 : 255 - 0xff
      13'h8B9: dout <= 8'b11111111; // 2233 : 255 - 0xff
      13'h8BA: dout <= 8'b11111111; // 2234 : 255 - 0xff
      13'h8BB: dout <= 8'b11111111; // 2235 : 255 - 0xff
      13'h8BC: dout <= 8'b11111111; // 2236 : 255 - 0xff
      13'h8BD: dout <= 8'b11111111; // 2237 : 255 - 0xff
      13'h8BE: dout <= 8'b11111111; // 2238 : 255 - 0xff
      13'h8BF: dout <= 8'b11111111; // 2239 : 255 - 0xff
      13'h8C0: dout <= 8'b11111111; // 2240 : 255 - 0xff -- Sprite 0x8c
      13'h8C1: dout <= 8'b11111111; // 2241 : 255 - 0xff
      13'h8C2: dout <= 8'b11111111; // 2242 : 255 - 0xff
      13'h8C3: dout <= 8'b11111111; // 2243 : 255 - 0xff
      13'h8C4: dout <= 8'b11111111; // 2244 : 255 - 0xff
      13'h8C5: dout <= 8'b11111111; // 2245 : 255 - 0xff
      13'h8C6: dout <= 8'b11111111; // 2246 : 255 - 0xff
      13'h8C7: dout <= 8'b11111111; // 2247 : 255 - 0xff
      13'h8C8: dout <= 8'b11111111; // 2248 : 255 - 0xff
      13'h8C9: dout <= 8'b11111111; // 2249 : 255 - 0xff
      13'h8CA: dout <= 8'b11111111; // 2250 : 255 - 0xff
      13'h8CB: dout <= 8'b11111111; // 2251 : 255 - 0xff
      13'h8CC: dout <= 8'b11111111; // 2252 : 255 - 0xff
      13'h8CD: dout <= 8'b11111111; // 2253 : 255 - 0xff
      13'h8CE: dout <= 8'b11111111; // 2254 : 255 - 0xff
      13'h8CF: dout <= 8'b11111111; // 2255 : 255 - 0xff
      13'h8D0: dout <= 8'b11111111; // 2256 : 255 - 0xff -- Sprite 0x8d
      13'h8D1: dout <= 8'b11111111; // 2257 : 255 - 0xff
      13'h8D2: dout <= 8'b11111111; // 2258 : 255 - 0xff
      13'h8D3: dout <= 8'b11111111; // 2259 : 255 - 0xff
      13'h8D4: dout <= 8'b11111111; // 2260 : 255 - 0xff
      13'h8D5: dout <= 8'b11111111; // 2261 : 255 - 0xff
      13'h8D6: dout <= 8'b11111111; // 2262 : 255 - 0xff
      13'h8D7: dout <= 8'b11111111; // 2263 : 255 - 0xff
      13'h8D8: dout <= 8'b11111111; // 2264 : 255 - 0xff
      13'h8D9: dout <= 8'b11111111; // 2265 : 255 - 0xff
      13'h8DA: dout <= 8'b11111111; // 2266 : 255 - 0xff
      13'h8DB: dout <= 8'b11111111; // 2267 : 255 - 0xff
      13'h8DC: dout <= 8'b11111111; // 2268 : 255 - 0xff
      13'h8DD: dout <= 8'b11111111; // 2269 : 255 - 0xff
      13'h8DE: dout <= 8'b11111111; // 2270 : 255 - 0xff
      13'h8DF: dout <= 8'b11111111; // 2271 : 255 - 0xff
      13'h8E0: dout <= 8'b11111111; // 2272 : 255 - 0xff -- Sprite 0x8e
      13'h8E1: dout <= 8'b11111111; // 2273 : 255 - 0xff
      13'h8E2: dout <= 8'b11111111; // 2274 : 255 - 0xff
      13'h8E3: dout <= 8'b11111111; // 2275 : 255 - 0xff
      13'h8E4: dout <= 8'b11111111; // 2276 : 255 - 0xff
      13'h8E5: dout <= 8'b11111111; // 2277 : 255 - 0xff
      13'h8E6: dout <= 8'b11111111; // 2278 : 255 - 0xff
      13'h8E7: dout <= 8'b11111111; // 2279 : 255 - 0xff
      13'h8E8: dout <= 8'b11111111; // 2280 : 255 - 0xff
      13'h8E9: dout <= 8'b11111111; // 2281 : 255 - 0xff
      13'h8EA: dout <= 8'b11111111; // 2282 : 255 - 0xff
      13'h8EB: dout <= 8'b11111111; // 2283 : 255 - 0xff
      13'h8EC: dout <= 8'b11111111; // 2284 : 255 - 0xff
      13'h8ED: dout <= 8'b11111111; // 2285 : 255 - 0xff
      13'h8EE: dout <= 8'b11111111; // 2286 : 255 - 0xff
      13'h8EF: dout <= 8'b11111111; // 2287 : 255 - 0xff
      13'h8F0: dout <= 8'b11111111; // 2288 : 255 - 0xff -- Sprite 0x8f
      13'h8F1: dout <= 8'b11111111; // 2289 : 255 - 0xff
      13'h8F2: dout <= 8'b11111111; // 2290 : 255 - 0xff
      13'h8F3: dout <= 8'b11111111; // 2291 : 255 - 0xff
      13'h8F4: dout <= 8'b11111111; // 2292 : 255 - 0xff
      13'h8F5: dout <= 8'b11111111; // 2293 : 255 - 0xff
      13'h8F6: dout <= 8'b11111111; // 2294 : 255 - 0xff
      13'h8F7: dout <= 8'b11111111; // 2295 : 255 - 0xff
      13'h8F8: dout <= 8'b11111111; // 2296 : 255 - 0xff
      13'h8F9: dout <= 8'b11111111; // 2297 : 255 - 0xff
      13'h8FA: dout <= 8'b11111111; // 2298 : 255 - 0xff
      13'h8FB: dout <= 8'b11111111; // 2299 : 255 - 0xff
      13'h8FC: dout <= 8'b11111111; // 2300 : 255 - 0xff
      13'h8FD: dout <= 8'b11111111; // 2301 : 255 - 0xff
      13'h8FE: dout <= 8'b11111111; // 2302 : 255 - 0xff
      13'h8FF: dout <= 8'b11111111; // 2303 : 255 - 0xff
      13'h900: dout <= 8'b00000000; // 2304 :   0 - 0x0 -- Sprite 0x90
      13'h901: dout <= 8'b00000000; // 2305 :   0 - 0x0
      13'h902: dout <= 8'b00000000; // 2306 :   0 - 0x0
      13'h903: dout <= 8'b00000000; // 2307 :   0 - 0x0
      13'h904: dout <= 8'b00000000; // 2308 :   0 - 0x0
      13'h905: dout <= 8'b00000001; // 2309 :   1 - 0x1
      13'h906: dout <= 8'b00011110; // 2310 :  30 - 0x1e
      13'h907: dout <= 8'b00111011; // 2311 :  59 - 0x3b
      13'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0
      13'h909: dout <= 8'b00000000; // 2313 :   0 - 0x0
      13'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      13'h90B: dout <= 8'b00000000; // 2315 :   0 - 0x0
      13'h90C: dout <= 8'b00000000; // 2316 :   0 - 0x0
      13'h90D: dout <= 8'b00000000; // 2317 :   0 - 0x0
      13'h90E: dout <= 8'b00000000; // 2318 :   0 - 0x0
      13'h90F: dout <= 8'b00000000; // 2319 :   0 - 0x0
      13'h910: dout <= 8'b00000000; // 2320 :   0 - 0x0 -- Sprite 0x91
      13'h911: dout <= 8'b00000000; // 2321 :   0 - 0x0
      13'h912: dout <= 8'b00001100; // 2322 :  12 - 0xc
      13'h913: dout <= 8'b00111100; // 2323 :  60 - 0x3c
      13'h914: dout <= 8'b11010000; // 2324 : 208 - 0xd0
      13'h915: dout <= 8'b00010000; // 2325 :  16 - 0x10
      13'h916: dout <= 8'b00100000; // 2326 :  32 - 0x20
      13'h917: dout <= 8'b01000000; // 2327 :  64 - 0x40
      13'h918: dout <= 8'b00000000; // 2328 :   0 - 0x0
      13'h919: dout <= 8'b00000000; // 2329 :   0 - 0x0
      13'h91A: dout <= 8'b00000000; // 2330 :   0 - 0x0
      13'h91B: dout <= 8'b00000000; // 2331 :   0 - 0x0
      13'h91C: dout <= 8'b00000000; // 2332 :   0 - 0x0
      13'h91D: dout <= 8'b00000000; // 2333 :   0 - 0x0
      13'h91E: dout <= 8'b00000000; // 2334 :   0 - 0x0
      13'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      13'h920: dout <= 8'b00111110; // 2336 :  62 - 0x3e -- Sprite 0x92
      13'h921: dout <= 8'b00101101; // 2337 :  45 - 0x2d
      13'h922: dout <= 8'b00110101; // 2338 :  53 - 0x35
      13'h923: dout <= 8'b00011101; // 2339 :  29 - 0x1d
      13'h924: dout <= 8'b00000001; // 2340 :   1 - 0x1
      13'h925: dout <= 8'b00000000; // 2341 :   0 - 0x0
      13'h926: dout <= 8'b00000000; // 2342 :   0 - 0x0
      13'h927: dout <= 8'b00000000; // 2343 :   0 - 0x0
      13'h928: dout <= 8'b00000000; // 2344 :   0 - 0x0
      13'h929: dout <= 8'b00000000; // 2345 :   0 - 0x0
      13'h92A: dout <= 8'b00000000; // 2346 :   0 - 0x0
      13'h92B: dout <= 8'b00000000; // 2347 :   0 - 0x0
      13'h92C: dout <= 8'b00000000; // 2348 :   0 - 0x0
      13'h92D: dout <= 8'b00000000; // 2349 :   0 - 0x0
      13'h92E: dout <= 8'b00000000; // 2350 :   0 - 0x0
      13'h92F: dout <= 8'b00000000; // 2351 :   0 - 0x0
      13'h930: dout <= 8'b10110000; // 2352 : 176 - 0xb0 -- Sprite 0x93
      13'h931: dout <= 8'b10111000; // 2353 : 184 - 0xb8
      13'h932: dout <= 8'b11111000; // 2354 : 248 - 0xf8
      13'h933: dout <= 8'b01111000; // 2355 : 120 - 0x78
      13'h934: dout <= 8'b10011000; // 2356 : 152 - 0x98
      13'h935: dout <= 8'b11110000; // 2357 : 240 - 0xf0
      13'h936: dout <= 8'b00000000; // 2358 :   0 - 0x0
      13'h937: dout <= 8'b00000000; // 2359 :   0 - 0x0
      13'h938: dout <= 8'b00000000; // 2360 :   0 - 0x0
      13'h939: dout <= 8'b00000000; // 2361 :   0 - 0x0
      13'h93A: dout <= 8'b00000000; // 2362 :   0 - 0x0
      13'h93B: dout <= 8'b00000000; // 2363 :   0 - 0x0
      13'h93C: dout <= 8'b00000000; // 2364 :   0 - 0x0
      13'h93D: dout <= 8'b00000000; // 2365 :   0 - 0x0
      13'h93E: dout <= 8'b00000000; // 2366 :   0 - 0x0
      13'h93F: dout <= 8'b00000000; // 2367 :   0 - 0x0
      13'h940: dout <= 8'b00000000; // 2368 :   0 - 0x0 -- Sprite 0x94
      13'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      13'h942: dout <= 8'b00000111; // 2370 :   7 - 0x7
      13'h943: dout <= 8'b00000011; // 2371 :   3 - 0x3
      13'h944: dout <= 8'b00001101; // 2372 :  13 - 0xd
      13'h945: dout <= 8'b00011110; // 2373 :  30 - 0x1e
      13'h946: dout <= 8'b00010111; // 2374 :  23 - 0x17
      13'h947: dout <= 8'b00011101; // 2375 :  29 - 0x1d
      13'h948: dout <= 8'b00000000; // 2376 :   0 - 0x0
      13'h949: dout <= 8'b00000000; // 2377 :   0 - 0x0
      13'h94A: dout <= 8'b00000000; // 2378 :   0 - 0x0
      13'h94B: dout <= 8'b00000000; // 2379 :   0 - 0x0
      13'h94C: dout <= 8'b00000000; // 2380 :   0 - 0x0
      13'h94D: dout <= 8'b00000000; // 2381 :   0 - 0x0
      13'h94E: dout <= 8'b00000000; // 2382 :   0 - 0x0
      13'h94F: dout <= 8'b00000000; // 2383 :   0 - 0x0
      13'h950: dout <= 8'b00000000; // 2384 :   0 - 0x0 -- Sprite 0x95
      13'h951: dout <= 8'b10000000; // 2385 : 128 - 0x80
      13'h952: dout <= 8'b01110000; // 2386 : 112 - 0x70
      13'h953: dout <= 8'b11100000; // 2387 : 224 - 0xe0
      13'h954: dout <= 8'b11011000; // 2388 : 216 - 0xd8
      13'h955: dout <= 8'b10111100; // 2389 : 188 - 0xbc
      13'h956: dout <= 8'b01110100; // 2390 : 116 - 0x74
      13'h957: dout <= 8'b11011100; // 2391 : 220 - 0xdc
      13'h958: dout <= 8'b00000000; // 2392 :   0 - 0x0
      13'h959: dout <= 8'b00000000; // 2393 :   0 - 0x0
      13'h95A: dout <= 8'b00000000; // 2394 :   0 - 0x0
      13'h95B: dout <= 8'b00000000; // 2395 :   0 - 0x0
      13'h95C: dout <= 8'b00000000; // 2396 :   0 - 0x0
      13'h95D: dout <= 8'b00000000; // 2397 :   0 - 0x0
      13'h95E: dout <= 8'b00000000; // 2398 :   0 - 0x0
      13'h95F: dout <= 8'b00000000; // 2399 :   0 - 0x0
      13'h960: dout <= 8'b00011111; // 2400 :  31 - 0x1f -- Sprite 0x96
      13'h961: dout <= 8'b00001011; // 2401 :  11 - 0xb
      13'h962: dout <= 8'b00001111; // 2402 :  15 - 0xf
      13'h963: dout <= 8'b00000101; // 2403 :   5 - 0x5
      13'h964: dout <= 8'b00000011; // 2404 :   3 - 0x3
      13'h965: dout <= 8'b00000001; // 2405 :   1 - 0x1
      13'h966: dout <= 8'b00000000; // 2406 :   0 - 0x0
      13'h967: dout <= 8'b00000000; // 2407 :   0 - 0x0
      13'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0
      13'h969: dout <= 8'b00000000; // 2409 :   0 - 0x0
      13'h96A: dout <= 8'b00000000; // 2410 :   0 - 0x0
      13'h96B: dout <= 8'b00000000; // 2411 :   0 - 0x0
      13'h96C: dout <= 8'b00000000; // 2412 :   0 - 0x0
      13'h96D: dout <= 8'b00000000; // 2413 :   0 - 0x0
      13'h96E: dout <= 8'b00000000; // 2414 :   0 - 0x0
      13'h96F: dout <= 8'b00000000; // 2415 :   0 - 0x0
      13'h970: dout <= 8'b11111100; // 2416 : 252 - 0xfc -- Sprite 0x97
      13'h971: dout <= 8'b01101000; // 2417 : 104 - 0x68
      13'h972: dout <= 8'b11111000; // 2418 : 248 - 0xf8
      13'h973: dout <= 8'b10110000; // 2419 : 176 - 0xb0
      13'h974: dout <= 8'b11100000; // 2420 : 224 - 0xe0
      13'h975: dout <= 8'b10000000; // 2421 : 128 - 0x80
      13'h976: dout <= 8'b00000000; // 2422 :   0 - 0x0
      13'h977: dout <= 8'b00000000; // 2423 :   0 - 0x0
      13'h978: dout <= 8'b00000000; // 2424 :   0 - 0x0
      13'h979: dout <= 8'b00000000; // 2425 :   0 - 0x0
      13'h97A: dout <= 8'b00000000; // 2426 :   0 - 0x0
      13'h97B: dout <= 8'b00000000; // 2427 :   0 - 0x0
      13'h97C: dout <= 8'b00000000; // 2428 :   0 - 0x0
      13'h97D: dout <= 8'b00000000; // 2429 :   0 - 0x0
      13'h97E: dout <= 8'b00000000; // 2430 :   0 - 0x0
      13'h97F: dout <= 8'b00000000; // 2431 :   0 - 0x0
      13'h980: dout <= 8'b00000000; // 2432 :   0 - 0x0 -- Sprite 0x98
      13'h981: dout <= 8'b00000000; // 2433 :   0 - 0x0
      13'h982: dout <= 8'b00000000; // 2434 :   0 - 0x0
      13'h983: dout <= 8'b00000001; // 2435 :   1 - 0x1
      13'h984: dout <= 8'b00000001; // 2436 :   1 - 0x1
      13'h985: dout <= 8'b00001011; // 2437 :  11 - 0xb
      13'h986: dout <= 8'b00011100; // 2438 :  28 - 0x1c
      13'h987: dout <= 8'b00111111; // 2439 :  63 - 0x3f
      13'h988: dout <= 8'b00000000; // 2440 :   0 - 0x0
      13'h989: dout <= 8'b00000000; // 2441 :   0 - 0x0
      13'h98A: dout <= 8'b00000000; // 2442 :   0 - 0x0
      13'h98B: dout <= 8'b00000000; // 2443 :   0 - 0x0
      13'h98C: dout <= 8'b00000000; // 2444 :   0 - 0x0
      13'h98D: dout <= 8'b00000000; // 2445 :   0 - 0x0
      13'h98E: dout <= 8'b00000000; // 2446 :   0 - 0x0
      13'h98F: dout <= 8'b00000000; // 2447 :   0 - 0x0
      13'h990: dout <= 8'b00000000; // 2448 :   0 - 0x0 -- Sprite 0x99
      13'h991: dout <= 8'b00000000; // 2449 :   0 - 0x0
      13'h992: dout <= 8'b00110000; // 2450 :  48 - 0x30
      13'h993: dout <= 8'b01111000; // 2451 : 120 - 0x78
      13'h994: dout <= 8'b10000000; // 2452 : 128 - 0x80
      13'h995: dout <= 8'b11110000; // 2453 : 240 - 0xf0
      13'h996: dout <= 8'b11111000; // 2454 : 248 - 0xf8
      13'h997: dout <= 8'b11111100; // 2455 : 252 - 0xfc
      13'h998: dout <= 8'b00000000; // 2456 :   0 - 0x0
      13'h999: dout <= 8'b00000000; // 2457 :   0 - 0x0
      13'h99A: dout <= 8'b00000000; // 2458 :   0 - 0x0
      13'h99B: dout <= 8'b00000000; // 2459 :   0 - 0x0
      13'h99C: dout <= 8'b00000000; // 2460 :   0 - 0x0
      13'h99D: dout <= 8'b00000000; // 2461 :   0 - 0x0
      13'h99E: dout <= 8'b00000000; // 2462 :   0 - 0x0
      13'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      13'h9A0: dout <= 8'b00111111; // 2464 :  63 - 0x3f -- Sprite 0x9a
      13'h9A1: dout <= 8'b00111111; // 2465 :  63 - 0x3f
      13'h9A2: dout <= 8'b00111111; // 2466 :  63 - 0x3f
      13'h9A3: dout <= 8'b00011111; // 2467 :  31 - 0x1f
      13'h9A4: dout <= 8'b00011111; // 2468 :  31 - 0x1f
      13'h9A5: dout <= 8'b00000111; // 2469 :   7 - 0x7
      13'h9A6: dout <= 8'b00000000; // 2470 :   0 - 0x0
      13'h9A7: dout <= 8'b00000000; // 2471 :   0 - 0x0
      13'h9A8: dout <= 8'b00000000; // 2472 :   0 - 0x0
      13'h9A9: dout <= 8'b00000000; // 2473 :   0 - 0x0
      13'h9AA: dout <= 8'b00000000; // 2474 :   0 - 0x0
      13'h9AB: dout <= 8'b00000000; // 2475 :   0 - 0x0
      13'h9AC: dout <= 8'b00000000; // 2476 :   0 - 0x0
      13'h9AD: dout <= 8'b00000000; // 2477 :   0 - 0x0
      13'h9AE: dout <= 8'b00000000; // 2478 :   0 - 0x0
      13'h9AF: dout <= 8'b00000000; // 2479 :   0 - 0x0
      13'h9B0: dout <= 8'b11111100; // 2480 : 252 - 0xfc -- Sprite 0x9b
      13'h9B1: dout <= 8'b11101100; // 2481 : 236 - 0xec
      13'h9B2: dout <= 8'b11101100; // 2482 : 236 - 0xec
      13'h9B3: dout <= 8'b11011000; // 2483 : 216 - 0xd8
      13'h9B4: dout <= 8'b11111000; // 2484 : 248 - 0xf8
      13'h9B5: dout <= 8'b11100000; // 2485 : 224 - 0xe0
      13'h9B6: dout <= 8'b00000000; // 2486 :   0 - 0x0
      13'h9B7: dout <= 8'b00000000; // 2487 :   0 - 0x0
      13'h9B8: dout <= 8'b00000000; // 2488 :   0 - 0x0
      13'h9B9: dout <= 8'b00000000; // 2489 :   0 - 0x0
      13'h9BA: dout <= 8'b00000000; // 2490 :   0 - 0x0
      13'h9BB: dout <= 8'b00000000; // 2491 :   0 - 0x0
      13'h9BC: dout <= 8'b00000000; // 2492 :   0 - 0x0
      13'h9BD: dout <= 8'b00000000; // 2493 :   0 - 0x0
      13'h9BE: dout <= 8'b00000000; // 2494 :   0 - 0x0
      13'h9BF: dout <= 8'b00000000; // 2495 :   0 - 0x0
      13'h9C0: dout <= 8'b00000000; // 2496 :   0 - 0x0 -- Sprite 0x9c
      13'h9C1: dout <= 8'b00000000; // 2497 :   0 - 0x0
      13'h9C2: dout <= 8'b00000001; // 2498 :   1 - 0x1
      13'h9C3: dout <= 8'b00011101; // 2499 :  29 - 0x1d
      13'h9C4: dout <= 8'b00111110; // 2500 :  62 - 0x3e
      13'h9C5: dout <= 8'b00111111; // 2501 :  63 - 0x3f
      13'h9C6: dout <= 8'b00111111; // 2502 :  63 - 0x3f
      13'h9C7: dout <= 8'b00111111; // 2503 :  63 - 0x3f
      13'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0
      13'h9C9: dout <= 8'b00000000; // 2505 :   0 - 0x0
      13'h9CA: dout <= 8'b00000000; // 2506 :   0 - 0x0
      13'h9CB: dout <= 8'b00000000; // 2507 :   0 - 0x0
      13'h9CC: dout <= 8'b00000000; // 2508 :   0 - 0x0
      13'h9CD: dout <= 8'b00000000; // 2509 :   0 - 0x0
      13'h9CE: dout <= 8'b00000000; // 2510 :   0 - 0x0
      13'h9CF: dout <= 8'b00000000; // 2511 :   0 - 0x0
      13'h9D0: dout <= 8'b00000000; // 2512 :   0 - 0x0 -- Sprite 0x9d
      13'h9D1: dout <= 8'b10000000; // 2513 : 128 - 0x80
      13'h9D2: dout <= 8'b00000000; // 2514 :   0 - 0x0
      13'h9D3: dout <= 8'b01110000; // 2515 : 112 - 0x70
      13'h9D4: dout <= 8'b11111000; // 2516 : 248 - 0xf8
      13'h9D5: dout <= 8'b11111100; // 2517 : 252 - 0xfc
      13'h9D6: dout <= 8'b11111100; // 2518 : 252 - 0xfc
      13'h9D7: dout <= 8'b11111100; // 2519 : 252 - 0xfc
      13'h9D8: dout <= 8'b00000000; // 2520 :   0 - 0x0
      13'h9D9: dout <= 8'b00000000; // 2521 :   0 - 0x0
      13'h9DA: dout <= 8'b00000000; // 2522 :   0 - 0x0
      13'h9DB: dout <= 8'b00000000; // 2523 :   0 - 0x0
      13'h9DC: dout <= 8'b00000000; // 2524 :   0 - 0x0
      13'h9DD: dout <= 8'b00000000; // 2525 :   0 - 0x0
      13'h9DE: dout <= 8'b00000000; // 2526 :   0 - 0x0
      13'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      13'h9E0: dout <= 8'b00111111; // 2528 :  63 - 0x3f -- Sprite 0x9e
      13'h9E1: dout <= 8'b00111111; // 2529 :  63 - 0x3f
      13'h9E2: dout <= 8'b00011111; // 2530 :  31 - 0x1f
      13'h9E3: dout <= 8'b00011111; // 2531 :  31 - 0x1f
      13'h9E4: dout <= 8'b00001111; // 2532 :  15 - 0xf
      13'h9E5: dout <= 8'b00000110; // 2533 :   6 - 0x6
      13'h9E6: dout <= 8'b00000000; // 2534 :   0 - 0x0
      13'h9E7: dout <= 8'b00000000; // 2535 :   0 - 0x0
      13'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0
      13'h9E9: dout <= 8'b00000000; // 2537 :   0 - 0x0
      13'h9EA: dout <= 8'b00000000; // 2538 :   0 - 0x0
      13'h9EB: dout <= 8'b00000000; // 2539 :   0 - 0x0
      13'h9EC: dout <= 8'b00000000; // 2540 :   0 - 0x0
      13'h9ED: dout <= 8'b00000000; // 2541 :   0 - 0x0
      13'h9EE: dout <= 8'b00000000; // 2542 :   0 - 0x0
      13'h9EF: dout <= 8'b00000000; // 2543 :   0 - 0x0
      13'h9F0: dout <= 8'b11101100; // 2544 : 236 - 0xec -- Sprite 0x9f
      13'h9F1: dout <= 8'b11101100; // 2545 : 236 - 0xec
      13'h9F2: dout <= 8'b11011000; // 2546 : 216 - 0xd8
      13'h9F3: dout <= 8'b11111000; // 2547 : 248 - 0xf8
      13'h9F4: dout <= 8'b11110000; // 2548 : 240 - 0xf0
      13'h9F5: dout <= 8'b11100000; // 2549 : 224 - 0xe0
      13'h9F6: dout <= 8'b00000000; // 2550 :   0 - 0x0
      13'h9F7: dout <= 8'b00000000; // 2551 :   0 - 0x0
      13'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0
      13'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      13'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      13'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      13'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      13'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      13'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      13'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      13'hA00: dout <= 8'b00000000; // 2560 :   0 - 0x0 -- Sprite 0xa0
      13'hA01: dout <= 8'b00000100; // 2561 :   4 - 0x4
      13'hA02: dout <= 8'b00000011; // 2562 :   3 - 0x3
      13'hA03: dout <= 8'b00000000; // 2563 :   0 - 0x0
      13'hA04: dout <= 8'b00000001; // 2564 :   1 - 0x1
      13'hA05: dout <= 8'b00000111; // 2565 :   7 - 0x7
      13'hA06: dout <= 8'b00001111; // 2566 :  15 - 0xf
      13'hA07: dout <= 8'b00001100; // 2567 :  12 - 0xc
      13'hA08: dout <= 8'b00000000; // 2568 :   0 - 0x0
      13'hA09: dout <= 8'b00000000; // 2569 :   0 - 0x0
      13'hA0A: dout <= 8'b00000000; // 2570 :   0 - 0x0
      13'hA0B: dout <= 8'b00000000; // 2571 :   0 - 0x0
      13'hA0C: dout <= 8'b00000000; // 2572 :   0 - 0x0
      13'hA0D: dout <= 8'b00000000; // 2573 :   0 - 0x0
      13'hA0E: dout <= 8'b00000000; // 2574 :   0 - 0x0
      13'hA0F: dout <= 8'b00000000; // 2575 :   0 - 0x0
      13'hA10: dout <= 8'b00000000; // 2576 :   0 - 0x0 -- Sprite 0xa1
      13'hA11: dout <= 8'b00000000; // 2577 :   0 - 0x0
      13'hA12: dout <= 8'b11100000; // 2578 : 224 - 0xe0
      13'hA13: dout <= 8'b10000000; // 2579 : 128 - 0x80
      13'hA14: dout <= 8'b01000000; // 2580 :  64 - 0x40
      13'hA15: dout <= 8'b11110000; // 2581 : 240 - 0xf0
      13'hA16: dout <= 8'b10011000; // 2582 : 152 - 0x98
      13'hA17: dout <= 8'b11111000; // 2583 : 248 - 0xf8
      13'hA18: dout <= 8'b00000000; // 2584 :   0 - 0x0
      13'hA19: dout <= 8'b00000000; // 2585 :   0 - 0x0
      13'hA1A: dout <= 8'b00000000; // 2586 :   0 - 0x0
      13'hA1B: dout <= 8'b00000000; // 2587 :   0 - 0x0
      13'hA1C: dout <= 8'b00000000; // 2588 :   0 - 0x0
      13'hA1D: dout <= 8'b00000000; // 2589 :   0 - 0x0
      13'hA1E: dout <= 8'b00000000; // 2590 :   0 - 0x0
      13'hA1F: dout <= 8'b00000000; // 2591 :   0 - 0x0
      13'hA20: dout <= 8'b00011111; // 2592 :  31 - 0x1f -- Sprite 0xa2
      13'hA21: dout <= 8'b00010011; // 2593 :  19 - 0x13
      13'hA22: dout <= 8'b00011111; // 2594 :  31 - 0x1f
      13'hA23: dout <= 8'b00001111; // 2595 :  15 - 0xf
      13'hA24: dout <= 8'b00001001; // 2596 :   9 - 0x9
      13'hA25: dout <= 8'b00000111; // 2597 :   7 - 0x7
      13'hA26: dout <= 8'b00000001; // 2598 :   1 - 0x1
      13'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      13'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0
      13'hA29: dout <= 8'b00000000; // 2601 :   0 - 0x0
      13'hA2A: dout <= 8'b00000000; // 2602 :   0 - 0x0
      13'hA2B: dout <= 8'b00000000; // 2603 :   0 - 0x0
      13'hA2C: dout <= 8'b00000000; // 2604 :   0 - 0x0
      13'hA2D: dout <= 8'b00000000; // 2605 :   0 - 0x0
      13'hA2E: dout <= 8'b00000000; // 2606 :   0 - 0x0
      13'hA2F: dout <= 8'b00000000; // 2607 :   0 - 0x0
      13'hA30: dout <= 8'b11100100; // 2608 : 228 - 0xe4 -- Sprite 0xa3
      13'hA31: dout <= 8'b00111100; // 2609 :  60 - 0x3c
      13'hA32: dout <= 8'b11100100; // 2610 : 228 - 0xe4
      13'hA33: dout <= 8'b00111000; // 2611 :  56 - 0x38
      13'hA34: dout <= 8'b11111000; // 2612 : 248 - 0xf8
      13'hA35: dout <= 8'b11110000; // 2613 : 240 - 0xf0
      13'hA36: dout <= 8'b11000000; // 2614 : 192 - 0xc0
      13'hA37: dout <= 8'b00000000; // 2615 :   0 - 0x0
      13'hA38: dout <= 8'b00000000; // 2616 :   0 - 0x0
      13'hA39: dout <= 8'b00000000; // 2617 :   0 - 0x0
      13'hA3A: dout <= 8'b00000000; // 2618 :   0 - 0x0
      13'hA3B: dout <= 8'b00000000; // 2619 :   0 - 0x0
      13'hA3C: dout <= 8'b00000000; // 2620 :   0 - 0x0
      13'hA3D: dout <= 8'b00000000; // 2621 :   0 - 0x0
      13'hA3E: dout <= 8'b00000000; // 2622 :   0 - 0x0
      13'hA3F: dout <= 8'b00000000; // 2623 :   0 - 0x0
      13'hA40: dout <= 8'b00000000; // 2624 :   0 - 0x0 -- Sprite 0xa4
      13'hA41: dout <= 8'b00000000; // 2625 :   0 - 0x0
      13'hA42: dout <= 8'b00000000; // 2626 :   0 - 0x0
      13'hA43: dout <= 8'b00000000; // 2627 :   0 - 0x0
      13'hA44: dout <= 8'b00010001; // 2628 :  17 - 0x11
      13'hA45: dout <= 8'b00010011; // 2629 :  19 - 0x13
      13'hA46: dout <= 8'b00011111; // 2630 :  31 - 0x1f
      13'hA47: dout <= 8'b00011111; // 2631 :  31 - 0x1f
      13'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0
      13'hA49: dout <= 8'b00000000; // 2633 :   0 - 0x0
      13'hA4A: dout <= 8'b00000000; // 2634 :   0 - 0x0
      13'hA4B: dout <= 8'b00000000; // 2635 :   0 - 0x0
      13'hA4C: dout <= 8'b00000000; // 2636 :   0 - 0x0
      13'hA4D: dout <= 8'b00000000; // 2637 :   0 - 0x0
      13'hA4E: dout <= 8'b00000000; // 2638 :   0 - 0x0
      13'hA4F: dout <= 8'b00000000; // 2639 :   0 - 0x0
      13'hA50: dout <= 8'b00000000; // 2640 :   0 - 0x0 -- Sprite 0xa5
      13'hA51: dout <= 8'b00000000; // 2641 :   0 - 0x0
      13'hA52: dout <= 8'b00000000; // 2642 :   0 - 0x0
      13'hA53: dout <= 8'b10000000; // 2643 : 128 - 0x80
      13'hA54: dout <= 8'b11000100; // 2644 : 196 - 0xc4
      13'hA55: dout <= 8'b11100100; // 2645 : 228 - 0xe4
      13'hA56: dout <= 8'b11111100; // 2646 : 252 - 0xfc
      13'hA57: dout <= 8'b11111100; // 2647 : 252 - 0xfc
      13'hA58: dout <= 8'b00000000; // 2648 :   0 - 0x0
      13'hA59: dout <= 8'b00000000; // 2649 :   0 - 0x0
      13'hA5A: dout <= 8'b00000000; // 2650 :   0 - 0x0
      13'hA5B: dout <= 8'b00000000; // 2651 :   0 - 0x0
      13'hA5C: dout <= 8'b00000000; // 2652 :   0 - 0x0
      13'hA5D: dout <= 8'b00000000; // 2653 :   0 - 0x0
      13'hA5E: dout <= 8'b00000000; // 2654 :   0 - 0x0
      13'hA5F: dout <= 8'b00000000; // 2655 :   0 - 0x0
      13'hA60: dout <= 8'b00011111; // 2656 :  31 - 0x1f -- Sprite 0xa6
      13'hA61: dout <= 8'b00001110; // 2657 :  14 - 0xe
      13'hA62: dout <= 8'b00000110; // 2658 :   6 - 0x6
      13'hA63: dout <= 8'b00000010; // 2659 :   2 - 0x2
      13'hA64: dout <= 8'b00000000; // 2660 :   0 - 0x0
      13'hA65: dout <= 8'b00000000; // 2661 :   0 - 0x0
      13'hA66: dout <= 8'b00000000; // 2662 :   0 - 0x0
      13'hA67: dout <= 8'b00000000; // 2663 :   0 - 0x0
      13'hA68: dout <= 8'b00000000; // 2664 :   0 - 0x0
      13'hA69: dout <= 8'b00000000; // 2665 :   0 - 0x0
      13'hA6A: dout <= 8'b00000000; // 2666 :   0 - 0x0
      13'hA6B: dout <= 8'b00000000; // 2667 :   0 - 0x0
      13'hA6C: dout <= 8'b00000000; // 2668 :   0 - 0x0
      13'hA6D: dout <= 8'b00000000; // 2669 :   0 - 0x0
      13'hA6E: dout <= 8'b00000000; // 2670 :   0 - 0x0
      13'hA6F: dout <= 8'b00000000; // 2671 :   0 - 0x0
      13'hA70: dout <= 8'b11111100; // 2672 : 252 - 0xfc -- Sprite 0xa7
      13'hA71: dout <= 8'b10111000; // 2673 : 184 - 0xb8
      13'hA72: dout <= 8'b10110000; // 2674 : 176 - 0xb0
      13'hA73: dout <= 8'b10100000; // 2675 : 160 - 0xa0
      13'hA74: dout <= 8'b10000000; // 2676 : 128 - 0x80
      13'hA75: dout <= 8'b00000000; // 2677 :   0 - 0x0
      13'hA76: dout <= 8'b00000000; // 2678 :   0 - 0x0
      13'hA77: dout <= 8'b00000000; // 2679 :   0 - 0x0
      13'hA78: dout <= 8'b00000000; // 2680 :   0 - 0x0
      13'hA79: dout <= 8'b00000000; // 2681 :   0 - 0x0
      13'hA7A: dout <= 8'b00000000; // 2682 :   0 - 0x0
      13'hA7B: dout <= 8'b00000000; // 2683 :   0 - 0x0
      13'hA7C: dout <= 8'b00000000; // 2684 :   0 - 0x0
      13'hA7D: dout <= 8'b00000000; // 2685 :   0 - 0x0
      13'hA7E: dout <= 8'b00000000; // 2686 :   0 - 0x0
      13'hA7F: dout <= 8'b00000000; // 2687 :   0 - 0x0
      13'hA80: dout <= 8'b00000000; // 2688 :   0 - 0x0 -- Sprite 0xa8
      13'hA81: dout <= 8'b00000000; // 2689 :   0 - 0x0
      13'hA82: dout <= 8'b00000000; // 2690 :   0 - 0x0
      13'hA83: dout <= 8'b00000001; // 2691 :   1 - 0x1
      13'hA84: dout <= 8'b00000011; // 2692 :   3 - 0x3
      13'hA85: dout <= 8'b00000110; // 2693 :   6 - 0x6
      13'hA86: dout <= 8'b00000110; // 2694 :   6 - 0x6
      13'hA87: dout <= 8'b00001111; // 2695 :  15 - 0xf
      13'hA88: dout <= 8'b00000000; // 2696 :   0 - 0x0
      13'hA89: dout <= 8'b00000000; // 2697 :   0 - 0x0
      13'hA8A: dout <= 8'b00000000; // 2698 :   0 - 0x0
      13'hA8B: dout <= 8'b00000000; // 2699 :   0 - 0x0
      13'hA8C: dout <= 8'b00000000; // 2700 :   0 - 0x0
      13'hA8D: dout <= 8'b00000000; // 2701 :   0 - 0x0
      13'hA8E: dout <= 8'b00000000; // 2702 :   0 - 0x0
      13'hA8F: dout <= 8'b00000000; // 2703 :   0 - 0x0
      13'hA90: dout <= 8'b00000000; // 2704 :   0 - 0x0 -- Sprite 0xa9
      13'hA91: dout <= 8'b00011000; // 2705 :  24 - 0x18
      13'hA92: dout <= 8'b11110100; // 2706 : 244 - 0xf4
      13'hA93: dout <= 8'b11111000; // 2707 : 248 - 0xf8
      13'hA94: dout <= 8'b00111000; // 2708 :  56 - 0x38
      13'hA95: dout <= 8'b01111100; // 2709 : 124 - 0x7c
      13'hA96: dout <= 8'b11111100; // 2710 : 252 - 0xfc
      13'hA97: dout <= 8'b11111100; // 2711 : 252 - 0xfc
      13'hA98: dout <= 8'b00000000; // 2712 :   0 - 0x0
      13'hA99: dout <= 8'b00000000; // 2713 :   0 - 0x0
      13'hA9A: dout <= 8'b00000000; // 2714 :   0 - 0x0
      13'hA9B: dout <= 8'b00000000; // 2715 :   0 - 0x0
      13'hA9C: dout <= 8'b00000000; // 2716 :   0 - 0x0
      13'hA9D: dout <= 8'b00000000; // 2717 :   0 - 0x0
      13'hA9E: dout <= 8'b00000000; // 2718 :   0 - 0x0
      13'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      13'hAA0: dout <= 8'b00001111; // 2720 :  15 - 0xf -- Sprite 0xaa
      13'hAA1: dout <= 8'b00011111; // 2721 :  31 - 0x1f
      13'hAA2: dout <= 8'b00110000; // 2722 :  48 - 0x30
      13'hAA3: dout <= 8'b00111000; // 2723 :  56 - 0x38
      13'hAA4: dout <= 8'b00011101; // 2724 :  29 - 0x1d
      13'hAA5: dout <= 8'b00000011; // 2725 :   3 - 0x3
      13'hAA6: dout <= 8'b00000011; // 2726 :   3 - 0x3
      13'hAA7: dout <= 8'b00000000; // 2727 :   0 - 0x0
      13'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0
      13'hAA9: dout <= 8'b00000000; // 2729 :   0 - 0x0
      13'hAAA: dout <= 8'b00000000; // 2730 :   0 - 0x0
      13'hAAB: dout <= 8'b00000000; // 2731 :   0 - 0x0
      13'hAAC: dout <= 8'b00000000; // 2732 :   0 - 0x0
      13'hAAD: dout <= 8'b00000000; // 2733 :   0 - 0x0
      13'hAAE: dout <= 8'b00000000; // 2734 :   0 - 0x0
      13'hAAF: dout <= 8'b00000000; // 2735 :   0 - 0x0
      13'hAB0: dout <= 8'b11111100; // 2736 : 252 - 0xfc -- Sprite 0xab
      13'hAB1: dout <= 8'b11111100; // 2737 : 252 - 0xfc
      13'hAB2: dout <= 8'b01111100; // 2738 : 124 - 0x7c
      13'hAB3: dout <= 8'b10001110; // 2739 : 142 - 0x8e
      13'hAB4: dout <= 8'b10000110; // 2740 : 134 - 0x86
      13'hAB5: dout <= 8'b10011100; // 2741 : 156 - 0x9c
      13'hAB6: dout <= 8'b01111000; // 2742 : 120 - 0x78
      13'hAB7: dout <= 8'b00000000; // 2743 :   0 - 0x0
      13'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0
      13'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      13'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      13'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      13'hABC: dout <= 8'b00000000; // 2748 :   0 - 0x0
      13'hABD: dout <= 8'b00000000; // 2749 :   0 - 0x0
      13'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      13'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      13'hAC0: dout <= 8'b00000000; // 2752 :   0 - 0x0 -- Sprite 0xac
      13'hAC1: dout <= 8'b00000001; // 2753 :   1 - 0x1
      13'hAC2: dout <= 8'b00000110; // 2754 :   6 - 0x6
      13'hAC3: dout <= 8'b00000111; // 2755 :   7 - 0x7
      13'hAC4: dout <= 8'b00000111; // 2756 :   7 - 0x7
      13'hAC5: dout <= 8'b00000111; // 2757 :   7 - 0x7
      13'hAC6: dout <= 8'b00000001; // 2758 :   1 - 0x1
      13'hAC7: dout <= 8'b00000011; // 2759 :   3 - 0x3
      13'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0
      13'hAC9: dout <= 8'b00000000; // 2761 :   0 - 0x0
      13'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      13'hACB: dout <= 8'b00000000; // 2763 :   0 - 0x0
      13'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      13'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      13'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      13'hACF: dout <= 8'b00000000; // 2767 :   0 - 0x0
      13'hAD0: dout <= 8'b00000000; // 2768 :   0 - 0x0 -- Sprite 0xad
      13'hAD1: dout <= 8'b11000000; // 2769 : 192 - 0xc0
      13'hAD2: dout <= 8'b00110000; // 2770 :  48 - 0x30
      13'hAD3: dout <= 8'b11110000; // 2771 : 240 - 0xf0
      13'hAD4: dout <= 8'b11110000; // 2772 : 240 - 0xf0
      13'hAD5: dout <= 8'b11110000; // 2773 : 240 - 0xf0
      13'hAD6: dout <= 8'b01000000; // 2774 :  64 - 0x40
      13'hAD7: dout <= 8'b01000000; // 2775 :  64 - 0x40
      13'hAD8: dout <= 8'b00000000; // 2776 :   0 - 0x0
      13'hAD9: dout <= 8'b00000000; // 2777 :   0 - 0x0
      13'hADA: dout <= 8'b00000000; // 2778 :   0 - 0x0
      13'hADB: dout <= 8'b00000000; // 2779 :   0 - 0x0
      13'hADC: dout <= 8'b00000000; // 2780 :   0 - 0x0
      13'hADD: dout <= 8'b00000000; // 2781 :   0 - 0x0
      13'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      13'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      13'hAE0: dout <= 8'b00000001; // 2784 :   1 - 0x1 -- Sprite 0xae
      13'hAE1: dout <= 8'b00000000; // 2785 :   0 - 0x0
      13'hAE2: dout <= 8'b00000001; // 2786 :   1 - 0x1
      13'hAE3: dout <= 8'b00000011; // 2787 :   3 - 0x3
      13'hAE4: dout <= 8'b00000001; // 2788 :   1 - 0x1
      13'hAE5: dout <= 8'b00000000; // 2789 :   0 - 0x0
      13'hAE6: dout <= 8'b00000000; // 2790 :   0 - 0x0
      13'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      13'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0
      13'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      13'hAEA: dout <= 8'b00000000; // 2794 :   0 - 0x0
      13'hAEB: dout <= 8'b00000000; // 2795 :   0 - 0x0
      13'hAEC: dout <= 8'b00000000; // 2796 :   0 - 0x0
      13'hAED: dout <= 8'b00000000; // 2797 :   0 - 0x0
      13'hAEE: dout <= 8'b00000000; // 2798 :   0 - 0x0
      13'hAEF: dout <= 8'b00000000; // 2799 :   0 - 0x0
      13'hAF0: dout <= 8'b01000000; // 2800 :  64 - 0x40 -- Sprite 0xaf
      13'hAF1: dout <= 8'b01000000; // 2801 :  64 - 0x40
      13'hAF2: dout <= 8'b01000000; // 2802 :  64 - 0x40
      13'hAF3: dout <= 8'b01000000; // 2803 :  64 - 0x40
      13'hAF4: dout <= 8'b01000000; // 2804 :  64 - 0x40
      13'hAF5: dout <= 8'b10000000; // 2805 : 128 - 0x80
      13'hAF6: dout <= 8'b00000000; // 2806 :   0 - 0x0
      13'hAF7: dout <= 8'b00000000; // 2807 :   0 - 0x0
      13'hAF8: dout <= 8'b00000000; // 2808 :   0 - 0x0
      13'hAF9: dout <= 8'b00000000; // 2809 :   0 - 0x0
      13'hAFA: dout <= 8'b00000000; // 2810 :   0 - 0x0
      13'hAFB: dout <= 8'b00000000; // 2811 :   0 - 0x0
      13'hAFC: dout <= 8'b00000000; // 2812 :   0 - 0x0
      13'hAFD: dout <= 8'b00000000; // 2813 :   0 - 0x0
      13'hAFE: dout <= 8'b00000000; // 2814 :   0 - 0x0
      13'hAFF: dout <= 8'b00000000; // 2815 :   0 - 0x0
      13'hB00: dout <= 8'b01111110; // 2816 : 126 - 0x7e -- Sprite 0xb0
      13'hB01: dout <= 8'b01100011; // 2817 :  99 - 0x63
      13'hB02: dout <= 8'b01100011; // 2818 :  99 - 0x63
      13'hB03: dout <= 8'b01100011; // 2819 :  99 - 0x63
      13'hB04: dout <= 8'b01111110; // 2820 : 126 - 0x7e
      13'hB05: dout <= 8'b01100000; // 2821 :  96 - 0x60
      13'hB06: dout <= 8'b01100000; // 2822 :  96 - 0x60
      13'hB07: dout <= 8'b00000000; // 2823 :   0 - 0x0
      13'hB08: dout <= 8'b01111110; // 2824 : 126 - 0x7e
      13'hB09: dout <= 8'b01100011; // 2825 :  99 - 0x63
      13'hB0A: dout <= 8'b01100011; // 2826 :  99 - 0x63
      13'hB0B: dout <= 8'b01100011; // 2827 :  99 - 0x63
      13'hB0C: dout <= 8'b01111110; // 2828 : 126 - 0x7e
      13'hB0D: dout <= 8'b01100000; // 2829 :  96 - 0x60
      13'hB0E: dout <= 8'b01100000; // 2830 :  96 - 0x60
      13'hB0F: dout <= 8'b00000000; // 2831 :   0 - 0x0
      13'hB10: dout <= 8'b01100000; // 2832 :  96 - 0x60 -- Sprite 0xb1
      13'hB11: dout <= 8'b01100000; // 2833 :  96 - 0x60
      13'hB12: dout <= 8'b01100000; // 2834 :  96 - 0x60
      13'hB13: dout <= 8'b01100000; // 2835 :  96 - 0x60
      13'hB14: dout <= 8'b01100000; // 2836 :  96 - 0x60
      13'hB15: dout <= 8'b01100000; // 2837 :  96 - 0x60
      13'hB16: dout <= 8'b01111111; // 2838 : 127 - 0x7f
      13'hB17: dout <= 8'b00000000; // 2839 :   0 - 0x0
      13'hB18: dout <= 8'b01100000; // 2840 :  96 - 0x60
      13'hB19: dout <= 8'b01100000; // 2841 :  96 - 0x60
      13'hB1A: dout <= 8'b01100000; // 2842 :  96 - 0x60
      13'hB1B: dout <= 8'b01100000; // 2843 :  96 - 0x60
      13'hB1C: dout <= 8'b01100000; // 2844 :  96 - 0x60
      13'hB1D: dout <= 8'b01100000; // 2845 :  96 - 0x60
      13'hB1E: dout <= 8'b01111111; // 2846 : 127 - 0x7f
      13'hB1F: dout <= 8'b00000000; // 2847 :   0 - 0x0
      13'hB20: dout <= 8'b00011100; // 2848 :  28 - 0x1c -- Sprite 0xb2
      13'hB21: dout <= 8'b00110110; // 2849 :  54 - 0x36
      13'hB22: dout <= 8'b01100011; // 2850 :  99 - 0x63
      13'hB23: dout <= 8'b01100011; // 2851 :  99 - 0x63
      13'hB24: dout <= 8'b01111111; // 2852 : 127 - 0x7f
      13'hB25: dout <= 8'b01100011; // 2853 :  99 - 0x63
      13'hB26: dout <= 8'b01100011; // 2854 :  99 - 0x63
      13'hB27: dout <= 8'b00000000; // 2855 :   0 - 0x0
      13'hB28: dout <= 8'b00011100; // 2856 :  28 - 0x1c
      13'hB29: dout <= 8'b00110110; // 2857 :  54 - 0x36
      13'hB2A: dout <= 8'b01100011; // 2858 :  99 - 0x63
      13'hB2B: dout <= 8'b01100011; // 2859 :  99 - 0x63
      13'hB2C: dout <= 8'b01111111; // 2860 : 127 - 0x7f
      13'hB2D: dout <= 8'b01100011; // 2861 :  99 - 0x63
      13'hB2E: dout <= 8'b01100011; // 2862 :  99 - 0x63
      13'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      13'hB30: dout <= 8'b00110011; // 2864 :  51 - 0x33 -- Sprite 0xb3
      13'hB31: dout <= 8'b00110011; // 2865 :  51 - 0x33
      13'hB32: dout <= 8'b00110011; // 2866 :  51 - 0x33
      13'hB33: dout <= 8'b00011110; // 2867 :  30 - 0x1e
      13'hB34: dout <= 8'b00001100; // 2868 :  12 - 0xc
      13'hB35: dout <= 8'b00001100; // 2869 :  12 - 0xc
      13'hB36: dout <= 8'b00001100; // 2870 :  12 - 0xc
      13'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      13'hB38: dout <= 8'b00110011; // 2872 :  51 - 0x33
      13'hB39: dout <= 8'b00110011; // 2873 :  51 - 0x33
      13'hB3A: dout <= 8'b00110011; // 2874 :  51 - 0x33
      13'hB3B: dout <= 8'b00011110; // 2875 :  30 - 0x1e
      13'hB3C: dout <= 8'b00001100; // 2876 :  12 - 0xc
      13'hB3D: dout <= 8'b00001100; // 2877 :  12 - 0xc
      13'hB3E: dout <= 8'b00001100; // 2878 :  12 - 0xc
      13'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      13'hB40: dout <= 8'b01111111; // 2880 : 127 - 0x7f -- Sprite 0xb4
      13'hB41: dout <= 8'b01100000; // 2881 :  96 - 0x60
      13'hB42: dout <= 8'b01100000; // 2882 :  96 - 0x60
      13'hB43: dout <= 8'b01111110; // 2883 : 126 - 0x7e
      13'hB44: dout <= 8'b01100000; // 2884 :  96 - 0x60
      13'hB45: dout <= 8'b01100000; // 2885 :  96 - 0x60
      13'hB46: dout <= 8'b01111111; // 2886 : 127 - 0x7f
      13'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      13'hB48: dout <= 8'b01111111; // 2888 : 127 - 0x7f
      13'hB49: dout <= 8'b01100000; // 2889 :  96 - 0x60
      13'hB4A: dout <= 8'b01100000; // 2890 :  96 - 0x60
      13'hB4B: dout <= 8'b01111110; // 2891 : 126 - 0x7e
      13'hB4C: dout <= 8'b01100000; // 2892 :  96 - 0x60
      13'hB4D: dout <= 8'b01100000; // 2893 :  96 - 0x60
      13'hB4E: dout <= 8'b01111111; // 2894 : 127 - 0x7f
      13'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      13'hB50: dout <= 8'b01111110; // 2896 : 126 - 0x7e -- Sprite 0xb5
      13'hB51: dout <= 8'b01100011; // 2897 :  99 - 0x63
      13'hB52: dout <= 8'b01100011; // 2898 :  99 - 0x63
      13'hB53: dout <= 8'b01100111; // 2899 : 103 - 0x67
      13'hB54: dout <= 8'b01111100; // 2900 : 124 - 0x7c
      13'hB55: dout <= 8'b01101110; // 2901 : 110 - 0x6e
      13'hB56: dout <= 8'b01100111; // 2902 : 103 - 0x67
      13'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      13'hB58: dout <= 8'b01111110; // 2904 : 126 - 0x7e
      13'hB59: dout <= 8'b01100011; // 2905 :  99 - 0x63
      13'hB5A: dout <= 8'b01100011; // 2906 :  99 - 0x63
      13'hB5B: dout <= 8'b01100111; // 2907 : 103 - 0x67
      13'hB5C: dout <= 8'b01111100; // 2908 : 124 - 0x7c
      13'hB5D: dout <= 8'b01101110; // 2909 : 110 - 0x6e
      13'hB5E: dout <= 8'b01100111; // 2910 : 103 - 0x67
      13'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      13'hB60: dout <= 8'b00111110; // 2912 :  62 - 0x3e -- Sprite 0xb6
      13'hB61: dout <= 8'b01100011; // 2913 :  99 - 0x63
      13'hB62: dout <= 8'b01100011; // 2914 :  99 - 0x63
      13'hB63: dout <= 8'b01100011; // 2915 :  99 - 0x63
      13'hB64: dout <= 8'b01100011; // 2916 :  99 - 0x63
      13'hB65: dout <= 8'b01100011; // 2917 :  99 - 0x63
      13'hB66: dout <= 8'b00111110; // 2918 :  62 - 0x3e
      13'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      13'hB68: dout <= 8'b00111110; // 2920 :  62 - 0x3e
      13'hB69: dout <= 8'b01100011; // 2921 :  99 - 0x63
      13'hB6A: dout <= 8'b01100011; // 2922 :  99 - 0x63
      13'hB6B: dout <= 8'b01100011; // 2923 :  99 - 0x63
      13'hB6C: dout <= 8'b01100011; // 2924 :  99 - 0x63
      13'hB6D: dout <= 8'b01100011; // 2925 :  99 - 0x63
      13'hB6E: dout <= 8'b00111110; // 2926 :  62 - 0x3e
      13'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      13'hB70: dout <= 8'b01100011; // 2928 :  99 - 0x63 -- Sprite 0xb7
      13'hB71: dout <= 8'b01110011; // 2929 : 115 - 0x73
      13'hB72: dout <= 8'b01111011; // 2930 : 123 - 0x7b
      13'hB73: dout <= 8'b01111111; // 2931 : 127 - 0x7f
      13'hB74: dout <= 8'b01101111; // 2932 : 111 - 0x6f
      13'hB75: dout <= 8'b01100111; // 2933 : 103 - 0x67
      13'hB76: dout <= 8'b01100011; // 2934 :  99 - 0x63
      13'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      13'hB78: dout <= 8'b01100011; // 2936 :  99 - 0x63
      13'hB79: dout <= 8'b01110011; // 2937 : 115 - 0x73
      13'hB7A: dout <= 8'b01111011; // 2938 : 123 - 0x7b
      13'hB7B: dout <= 8'b01111111; // 2939 : 127 - 0x7f
      13'hB7C: dout <= 8'b01101111; // 2940 : 111 - 0x6f
      13'hB7D: dout <= 8'b01100111; // 2941 : 103 - 0x67
      13'hB7E: dout <= 8'b01100011; // 2942 :  99 - 0x63
      13'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      13'hB80: dout <= 8'b00111111; // 2944 :  63 - 0x3f -- Sprite 0xb8
      13'hB81: dout <= 8'b00001100; // 2945 :  12 - 0xc
      13'hB82: dout <= 8'b00001100; // 2946 :  12 - 0xc
      13'hB83: dout <= 8'b00001100; // 2947 :  12 - 0xc
      13'hB84: dout <= 8'b00001100; // 2948 :  12 - 0xc
      13'hB85: dout <= 8'b00001100; // 2949 :  12 - 0xc
      13'hB86: dout <= 8'b00001100; // 2950 :  12 - 0xc
      13'hB87: dout <= 8'b00000000; // 2951 :   0 - 0x0
      13'hB88: dout <= 8'b00111111; // 2952 :  63 - 0x3f
      13'hB89: dout <= 8'b00001100; // 2953 :  12 - 0xc
      13'hB8A: dout <= 8'b00001100; // 2954 :  12 - 0xc
      13'hB8B: dout <= 8'b00001100; // 2955 :  12 - 0xc
      13'hB8C: dout <= 8'b00001100; // 2956 :  12 - 0xc
      13'hB8D: dout <= 8'b00001100; // 2957 :  12 - 0xc
      13'hB8E: dout <= 8'b00001100; // 2958 :  12 - 0xc
      13'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      13'hB90: dout <= 8'b01100011; // 2960 :  99 - 0x63 -- Sprite 0xb9
      13'hB91: dout <= 8'b01100011; // 2961 :  99 - 0x63
      13'hB92: dout <= 8'b01101011; // 2962 : 107 - 0x6b
      13'hB93: dout <= 8'b01111111; // 2963 : 127 - 0x7f
      13'hB94: dout <= 8'b01111111; // 2964 : 127 - 0x7f
      13'hB95: dout <= 8'b01110111; // 2965 : 119 - 0x77
      13'hB96: dout <= 8'b01100011; // 2966 :  99 - 0x63
      13'hB97: dout <= 8'b00000000; // 2967 :   0 - 0x0
      13'hB98: dout <= 8'b01100011; // 2968 :  99 - 0x63
      13'hB99: dout <= 8'b01100011; // 2969 :  99 - 0x63
      13'hB9A: dout <= 8'b01101011; // 2970 : 107 - 0x6b
      13'hB9B: dout <= 8'b01111111; // 2971 : 127 - 0x7f
      13'hB9C: dout <= 8'b01111111; // 2972 : 127 - 0x7f
      13'hB9D: dout <= 8'b01110111; // 2973 : 119 - 0x77
      13'hB9E: dout <= 8'b01100011; // 2974 :  99 - 0x63
      13'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      13'hBA0: dout <= 8'b01111100; // 2976 : 124 - 0x7c -- Sprite 0xba
      13'hBA1: dout <= 8'b01100110; // 2977 : 102 - 0x66
      13'hBA2: dout <= 8'b01100011; // 2978 :  99 - 0x63
      13'hBA3: dout <= 8'b01100011; // 2979 :  99 - 0x63
      13'hBA4: dout <= 8'b01100011; // 2980 :  99 - 0x63
      13'hBA5: dout <= 8'b01100110; // 2981 : 102 - 0x66
      13'hBA6: dout <= 8'b01111100; // 2982 : 124 - 0x7c
      13'hBA7: dout <= 8'b00000000; // 2983 :   0 - 0x0
      13'hBA8: dout <= 8'b00000000; // 2984 :   0 - 0x0
      13'hBA9: dout <= 8'b00000000; // 2985 :   0 - 0x0
      13'hBAA: dout <= 8'b00000000; // 2986 :   0 - 0x0
      13'hBAB: dout <= 8'b00000000; // 2987 :   0 - 0x0
      13'hBAC: dout <= 8'b00000000; // 2988 :   0 - 0x0
      13'hBAD: dout <= 8'b00000000; // 2989 :   0 - 0x0
      13'hBAE: dout <= 8'b00000000; // 2990 :   0 - 0x0
      13'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      13'hBB0: dout <= 8'b00011100; // 2992 :  28 - 0x1c -- Sprite 0xbb
      13'hBB1: dout <= 8'b00011100; // 2993 :  28 - 0x1c
      13'hBB2: dout <= 8'b00011100; // 2994 :  28 - 0x1c
      13'hBB3: dout <= 8'b00011000; // 2995 :  24 - 0x18
      13'hBB4: dout <= 8'b00011000; // 2996 :  24 - 0x18
      13'hBB5: dout <= 8'b00000000; // 2997 :   0 - 0x0
      13'hBB6: dout <= 8'b00011000; // 2998 :  24 - 0x18
      13'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      13'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0
      13'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      13'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      13'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      13'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      13'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      13'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      13'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      13'hBC0: dout <= 8'b00011111; // 3008 :  31 - 0x1f -- Sprite 0xbc
      13'hBC1: dout <= 8'b00110000; // 3009 :  48 - 0x30
      13'hBC2: dout <= 8'b01100000; // 3010 :  96 - 0x60
      13'hBC3: dout <= 8'b01100111; // 3011 : 103 - 0x67
      13'hBC4: dout <= 8'b01100011; // 3012 :  99 - 0x63
      13'hBC5: dout <= 8'b00110011; // 3013 :  51 - 0x33
      13'hBC6: dout <= 8'b00011111; // 3014 :  31 - 0x1f
      13'hBC7: dout <= 8'b00000000; // 3015 :   0 - 0x0
      13'hBC8: dout <= 8'b00011111; // 3016 :  31 - 0x1f
      13'hBC9: dout <= 8'b00110000; // 3017 :  48 - 0x30
      13'hBCA: dout <= 8'b01100000; // 3018 :  96 - 0x60
      13'hBCB: dout <= 8'b01100111; // 3019 : 103 - 0x67
      13'hBCC: dout <= 8'b01100011; // 3020 :  99 - 0x63
      13'hBCD: dout <= 8'b00110011; // 3021 :  51 - 0x33
      13'hBCE: dout <= 8'b00011111; // 3022 :  31 - 0x1f
      13'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      13'hBD0: dout <= 8'b01100011; // 3024 :  99 - 0x63 -- Sprite 0xbd
      13'hBD1: dout <= 8'b01110111; // 3025 : 119 - 0x77
      13'hBD2: dout <= 8'b01111111; // 3026 : 127 - 0x7f
      13'hBD3: dout <= 8'b01111111; // 3027 : 127 - 0x7f
      13'hBD4: dout <= 8'b01101011; // 3028 : 107 - 0x6b
      13'hBD5: dout <= 8'b01100011; // 3029 :  99 - 0x63
      13'hBD6: dout <= 8'b01100011; // 3030 :  99 - 0x63
      13'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      13'hBD8: dout <= 8'b01100011; // 3032 :  99 - 0x63
      13'hBD9: dout <= 8'b01110111; // 3033 : 119 - 0x77
      13'hBDA: dout <= 8'b01111111; // 3034 : 127 - 0x7f
      13'hBDB: dout <= 8'b01111111; // 3035 : 127 - 0x7f
      13'hBDC: dout <= 8'b01101011; // 3036 : 107 - 0x6b
      13'hBDD: dout <= 8'b01100011; // 3037 :  99 - 0x63
      13'hBDE: dout <= 8'b01100011; // 3038 :  99 - 0x63
      13'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      13'hBE0: dout <= 8'b01100011; // 3040 :  99 - 0x63 -- Sprite 0xbe
      13'hBE1: dout <= 8'b01100011; // 3041 :  99 - 0x63
      13'hBE2: dout <= 8'b01100011; // 3042 :  99 - 0x63
      13'hBE3: dout <= 8'b01110111; // 3043 : 119 - 0x77
      13'hBE4: dout <= 8'b00111110; // 3044 :  62 - 0x3e
      13'hBE5: dout <= 8'b00011100; // 3045 :  28 - 0x1c
      13'hBE6: dout <= 8'b00001000; // 3046 :   8 - 0x8
      13'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      13'hBE8: dout <= 8'b01100011; // 3048 :  99 - 0x63
      13'hBE9: dout <= 8'b01100011; // 3049 :  99 - 0x63
      13'hBEA: dout <= 8'b01100011; // 3050 :  99 - 0x63
      13'hBEB: dout <= 8'b01110111; // 3051 : 119 - 0x77
      13'hBEC: dout <= 8'b00111110; // 3052 :  62 - 0x3e
      13'hBED: dout <= 8'b00011100; // 3053 :  28 - 0x1c
      13'hBEE: dout <= 8'b00001000; // 3054 :   8 - 0x8
      13'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      13'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Sprite 0xbf
      13'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      13'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      13'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      13'hBF4: dout <= 8'b00000000; // 3060 :   0 - 0x0
      13'hBF5: dout <= 8'b00000000; // 3061 :   0 - 0x0
      13'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      13'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      13'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0
      13'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      13'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      13'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      13'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      13'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      13'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      13'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      13'hC00: dout <= 8'b00011111; // 3072 :  31 - 0x1f -- Sprite 0xc0
      13'hC01: dout <= 8'b00110000; // 3073 :  48 - 0x30
      13'hC02: dout <= 8'b01100000; // 3074 :  96 - 0x60
      13'hC03: dout <= 8'b01100111; // 3075 : 103 - 0x67
      13'hC04: dout <= 8'b01100011; // 3076 :  99 - 0x63
      13'hC05: dout <= 8'b00110011; // 3077 :  51 - 0x33
      13'hC06: dout <= 8'b00011111; // 3078 :  31 - 0x1f
      13'hC07: dout <= 8'b00000000; // 3079 :   0 - 0x0
      13'hC08: dout <= 8'b00000000; // 3080 :   0 - 0x0
      13'hC09: dout <= 8'b00000000; // 3081 :   0 - 0x0
      13'hC0A: dout <= 8'b00000000; // 3082 :   0 - 0x0
      13'hC0B: dout <= 8'b00000000; // 3083 :   0 - 0x0
      13'hC0C: dout <= 8'b00000000; // 3084 :   0 - 0x0
      13'hC0D: dout <= 8'b00000000; // 3085 :   0 - 0x0
      13'hC0E: dout <= 8'b00000000; // 3086 :   0 - 0x0
      13'hC0F: dout <= 8'b00000000; // 3087 :   0 - 0x0
      13'hC10: dout <= 8'b00011100; // 3088 :  28 - 0x1c -- Sprite 0xc1
      13'hC11: dout <= 8'b00110110; // 3089 :  54 - 0x36
      13'hC12: dout <= 8'b01100011; // 3090 :  99 - 0x63
      13'hC13: dout <= 8'b01100011; // 3091 :  99 - 0x63
      13'hC14: dout <= 8'b01111111; // 3092 : 127 - 0x7f
      13'hC15: dout <= 8'b01100011; // 3093 :  99 - 0x63
      13'hC16: dout <= 8'b01100011; // 3094 :  99 - 0x63
      13'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      13'hC18: dout <= 8'b00000000; // 3096 :   0 - 0x0
      13'hC19: dout <= 8'b00000000; // 3097 :   0 - 0x0
      13'hC1A: dout <= 8'b00000000; // 3098 :   0 - 0x0
      13'hC1B: dout <= 8'b00000000; // 3099 :   0 - 0x0
      13'hC1C: dout <= 8'b00000000; // 3100 :   0 - 0x0
      13'hC1D: dout <= 8'b00000000; // 3101 :   0 - 0x0
      13'hC1E: dout <= 8'b00000000; // 3102 :   0 - 0x0
      13'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      13'hC20: dout <= 8'b01100011; // 3104 :  99 - 0x63 -- Sprite 0xc2
      13'hC21: dout <= 8'b01110111; // 3105 : 119 - 0x77
      13'hC22: dout <= 8'b01111111; // 3106 : 127 - 0x7f
      13'hC23: dout <= 8'b01111111; // 3107 : 127 - 0x7f
      13'hC24: dout <= 8'b01101011; // 3108 : 107 - 0x6b
      13'hC25: dout <= 8'b01100011; // 3109 :  99 - 0x63
      13'hC26: dout <= 8'b01100011; // 3110 :  99 - 0x63
      13'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      13'hC28: dout <= 8'b00000000; // 3112 :   0 - 0x0
      13'hC29: dout <= 8'b00000000; // 3113 :   0 - 0x0
      13'hC2A: dout <= 8'b00000000; // 3114 :   0 - 0x0
      13'hC2B: dout <= 8'b00000000; // 3115 :   0 - 0x0
      13'hC2C: dout <= 8'b00000000; // 3116 :   0 - 0x0
      13'hC2D: dout <= 8'b00000000; // 3117 :   0 - 0x0
      13'hC2E: dout <= 8'b00000000; // 3118 :   0 - 0x0
      13'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      13'hC30: dout <= 8'b01111111; // 3120 : 127 - 0x7f -- Sprite 0xc3
      13'hC31: dout <= 8'b01100000; // 3121 :  96 - 0x60
      13'hC32: dout <= 8'b01100000; // 3122 :  96 - 0x60
      13'hC33: dout <= 8'b01111110; // 3123 : 126 - 0x7e
      13'hC34: dout <= 8'b01100000; // 3124 :  96 - 0x60
      13'hC35: dout <= 8'b01100000; // 3125 :  96 - 0x60
      13'hC36: dout <= 8'b01111111; // 3126 : 127 - 0x7f
      13'hC37: dout <= 8'b00000000; // 3127 :   0 - 0x0
      13'hC38: dout <= 8'b00000000; // 3128 :   0 - 0x0
      13'hC39: dout <= 8'b00000000; // 3129 :   0 - 0x0
      13'hC3A: dout <= 8'b00000000; // 3130 :   0 - 0x0
      13'hC3B: dout <= 8'b00000000; // 3131 :   0 - 0x0
      13'hC3C: dout <= 8'b00000000; // 3132 :   0 - 0x0
      13'hC3D: dout <= 8'b00000000; // 3133 :   0 - 0x0
      13'hC3E: dout <= 8'b00000000; // 3134 :   0 - 0x0
      13'hC3F: dout <= 8'b00000000; // 3135 :   0 - 0x0
      13'hC40: dout <= 8'b00111110; // 3136 :  62 - 0x3e -- Sprite 0xc4
      13'hC41: dout <= 8'b01100011; // 3137 :  99 - 0x63
      13'hC42: dout <= 8'b01100011; // 3138 :  99 - 0x63
      13'hC43: dout <= 8'b01100011; // 3139 :  99 - 0x63
      13'hC44: dout <= 8'b01100011; // 3140 :  99 - 0x63
      13'hC45: dout <= 8'b01100011; // 3141 :  99 - 0x63
      13'hC46: dout <= 8'b00111110; // 3142 :  62 - 0x3e
      13'hC47: dout <= 8'b00000000; // 3143 :   0 - 0x0
      13'hC48: dout <= 8'b00000000; // 3144 :   0 - 0x0
      13'hC49: dout <= 8'b00000000; // 3145 :   0 - 0x0
      13'hC4A: dout <= 8'b00000000; // 3146 :   0 - 0x0
      13'hC4B: dout <= 8'b00000000; // 3147 :   0 - 0x0
      13'hC4C: dout <= 8'b00000000; // 3148 :   0 - 0x0
      13'hC4D: dout <= 8'b00000000; // 3149 :   0 - 0x0
      13'hC4E: dout <= 8'b00000000; // 3150 :   0 - 0x0
      13'hC4F: dout <= 8'b00000000; // 3151 :   0 - 0x0
      13'hC50: dout <= 8'b01100011; // 3152 :  99 - 0x63 -- Sprite 0xc5
      13'hC51: dout <= 8'b01100011; // 3153 :  99 - 0x63
      13'hC52: dout <= 8'b01100011; // 3154 :  99 - 0x63
      13'hC53: dout <= 8'b01110111; // 3155 : 119 - 0x77
      13'hC54: dout <= 8'b00111110; // 3156 :  62 - 0x3e
      13'hC55: dout <= 8'b00011100; // 3157 :  28 - 0x1c
      13'hC56: dout <= 8'b00001000; // 3158 :   8 - 0x8
      13'hC57: dout <= 8'b00000000; // 3159 :   0 - 0x0
      13'hC58: dout <= 8'b00000000; // 3160 :   0 - 0x0
      13'hC59: dout <= 8'b00000000; // 3161 :   0 - 0x0
      13'hC5A: dout <= 8'b00000000; // 3162 :   0 - 0x0
      13'hC5B: dout <= 8'b00000000; // 3163 :   0 - 0x0
      13'hC5C: dout <= 8'b00000000; // 3164 :   0 - 0x0
      13'hC5D: dout <= 8'b00000000; // 3165 :   0 - 0x0
      13'hC5E: dout <= 8'b00000000; // 3166 :   0 - 0x0
      13'hC5F: dout <= 8'b00000000; // 3167 :   0 - 0x0
      13'hC60: dout <= 8'b01111110; // 3168 : 126 - 0x7e -- Sprite 0xc6
      13'hC61: dout <= 8'b01100011; // 3169 :  99 - 0x63
      13'hC62: dout <= 8'b01100011; // 3170 :  99 - 0x63
      13'hC63: dout <= 8'b01100111; // 3171 : 103 - 0x67
      13'hC64: dout <= 8'b01111100; // 3172 : 124 - 0x7c
      13'hC65: dout <= 8'b01101110; // 3173 : 110 - 0x6e
      13'hC66: dout <= 8'b01100111; // 3174 : 103 - 0x67
      13'hC67: dout <= 8'b00000000; // 3175 :   0 - 0x0
      13'hC68: dout <= 8'b00000000; // 3176 :   0 - 0x0
      13'hC69: dout <= 8'b00000000; // 3177 :   0 - 0x0
      13'hC6A: dout <= 8'b00000000; // 3178 :   0 - 0x0
      13'hC6B: dout <= 8'b00000000; // 3179 :   0 - 0x0
      13'hC6C: dout <= 8'b00000000; // 3180 :   0 - 0x0
      13'hC6D: dout <= 8'b00000000; // 3181 :   0 - 0x0
      13'hC6E: dout <= 8'b00000000; // 3182 :   0 - 0x0
      13'hC6F: dout <= 8'b00000000; // 3183 :   0 - 0x0
      13'hC70: dout <= 8'b00110011; // 3184 :  51 - 0x33 -- Sprite 0xc7
      13'hC71: dout <= 8'b00110011; // 3185 :  51 - 0x33
      13'hC72: dout <= 8'b00110011; // 3186 :  51 - 0x33
      13'hC73: dout <= 8'b00011110; // 3187 :  30 - 0x1e
      13'hC74: dout <= 8'b00001100; // 3188 :  12 - 0xc
      13'hC75: dout <= 8'b00001100; // 3189 :  12 - 0xc
      13'hC76: dout <= 8'b00001100; // 3190 :  12 - 0xc
      13'hC77: dout <= 8'b00000000; // 3191 :   0 - 0x0
      13'hC78: dout <= 8'b00000000; // 3192 :   0 - 0x0
      13'hC79: dout <= 8'b00000000; // 3193 :   0 - 0x0
      13'hC7A: dout <= 8'b00000000; // 3194 :   0 - 0x0
      13'hC7B: dout <= 8'b00000000; // 3195 :   0 - 0x0
      13'hC7C: dout <= 8'b00000000; // 3196 :   0 - 0x0
      13'hC7D: dout <= 8'b00000000; // 3197 :   0 - 0x0
      13'hC7E: dout <= 8'b00000000; // 3198 :   0 - 0x0
      13'hC7F: dout <= 8'b00000000; // 3199 :   0 - 0x0
      13'hC80: dout <= 8'b00000000; // 3200 :   0 - 0x0 -- Sprite 0xc8
      13'hC81: dout <= 8'b00000000; // 3201 :   0 - 0x0
      13'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      13'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      13'hC84: dout <= 8'b00000000; // 3204 :   0 - 0x0
      13'hC85: dout <= 8'b00000000; // 3205 :   0 - 0x0
      13'hC86: dout <= 8'b00000000; // 3206 :   0 - 0x0
      13'hC87: dout <= 8'b00000000; // 3207 :   0 - 0x0
      13'hC88: dout <= 8'b00000000; // 3208 :   0 - 0x0
      13'hC89: dout <= 8'b00000000; // 3209 :   0 - 0x0
      13'hC8A: dout <= 8'b00000000; // 3210 :   0 - 0x0
      13'hC8B: dout <= 8'b00000000; // 3211 :   0 - 0x0
      13'hC8C: dout <= 8'b00000000; // 3212 :   0 - 0x0
      13'hC8D: dout <= 8'b00000000; // 3213 :   0 - 0x0
      13'hC8E: dout <= 8'b00000000; // 3214 :   0 - 0x0
      13'hC8F: dout <= 8'b00000000; // 3215 :   0 - 0x0
      13'hC90: dout <= 8'b00000000; // 3216 :   0 - 0x0 -- Sprite 0xc9
      13'hC91: dout <= 8'b00000000; // 3217 :   0 - 0x0
      13'hC92: dout <= 8'b00000000; // 3218 :   0 - 0x0
      13'hC93: dout <= 8'b00000000; // 3219 :   0 - 0x0
      13'hC94: dout <= 8'b00000000; // 3220 :   0 - 0x0
      13'hC95: dout <= 8'b00000000; // 3221 :   0 - 0x0
      13'hC96: dout <= 8'b00000000; // 3222 :   0 - 0x0
      13'hC97: dout <= 8'b00000000; // 3223 :   0 - 0x0
      13'hC98: dout <= 8'b00000000; // 3224 :   0 - 0x0
      13'hC99: dout <= 8'b00000000; // 3225 :   0 - 0x0
      13'hC9A: dout <= 8'b00000000; // 3226 :   0 - 0x0
      13'hC9B: dout <= 8'b00000000; // 3227 :   0 - 0x0
      13'hC9C: dout <= 8'b00000000; // 3228 :   0 - 0x0
      13'hC9D: dout <= 8'b00000000; // 3229 :   0 - 0x0
      13'hC9E: dout <= 8'b00000000; // 3230 :   0 - 0x0
      13'hC9F: dout <= 8'b00000000; // 3231 :   0 - 0x0
      13'hCA0: dout <= 8'b00000000; // 3232 :   0 - 0x0 -- Sprite 0xca
      13'hCA1: dout <= 8'b00000000; // 3233 :   0 - 0x0
      13'hCA2: dout <= 8'b00000000; // 3234 :   0 - 0x0
      13'hCA3: dout <= 8'b00000000; // 3235 :   0 - 0x0
      13'hCA4: dout <= 8'b00000000; // 3236 :   0 - 0x0
      13'hCA5: dout <= 8'b00000000; // 3237 :   0 - 0x0
      13'hCA6: dout <= 8'b00000000; // 3238 :   0 - 0x0
      13'hCA7: dout <= 8'b00000000; // 3239 :   0 - 0x0
      13'hCA8: dout <= 8'b00000000; // 3240 :   0 - 0x0
      13'hCA9: dout <= 8'b00000000; // 3241 :   0 - 0x0
      13'hCAA: dout <= 8'b00000000; // 3242 :   0 - 0x0
      13'hCAB: dout <= 8'b00000000; // 3243 :   0 - 0x0
      13'hCAC: dout <= 8'b00000000; // 3244 :   0 - 0x0
      13'hCAD: dout <= 8'b00000000; // 3245 :   0 - 0x0
      13'hCAE: dout <= 8'b00000000; // 3246 :   0 - 0x0
      13'hCAF: dout <= 8'b00000000; // 3247 :   0 - 0x0
      13'hCB0: dout <= 8'b00000000; // 3248 :   0 - 0x0 -- Sprite 0xcb
      13'hCB1: dout <= 8'b00000000; // 3249 :   0 - 0x0
      13'hCB2: dout <= 8'b00000000; // 3250 :   0 - 0x0
      13'hCB3: dout <= 8'b00000000; // 3251 :   0 - 0x0
      13'hCB4: dout <= 8'b00000000; // 3252 :   0 - 0x0
      13'hCB5: dout <= 8'b00000000; // 3253 :   0 - 0x0
      13'hCB6: dout <= 8'b00000000; // 3254 :   0 - 0x0
      13'hCB7: dout <= 8'b00000000; // 3255 :   0 - 0x0
      13'hCB8: dout <= 8'b00000000; // 3256 :   0 - 0x0
      13'hCB9: dout <= 8'b00000000; // 3257 :   0 - 0x0
      13'hCBA: dout <= 8'b00000000; // 3258 :   0 - 0x0
      13'hCBB: dout <= 8'b00000000; // 3259 :   0 - 0x0
      13'hCBC: dout <= 8'b00000000; // 3260 :   0 - 0x0
      13'hCBD: dout <= 8'b00000000; // 3261 :   0 - 0x0
      13'hCBE: dout <= 8'b00000000; // 3262 :   0 - 0x0
      13'hCBF: dout <= 8'b00000000; // 3263 :   0 - 0x0
      13'hCC0: dout <= 8'b00000000; // 3264 :   0 - 0x0 -- Sprite 0xcc
      13'hCC1: dout <= 8'b00000000; // 3265 :   0 - 0x0
      13'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      13'hCC3: dout <= 8'b00000000; // 3267 :   0 - 0x0
      13'hCC4: dout <= 8'b00000000; // 3268 :   0 - 0x0
      13'hCC5: dout <= 8'b00000000; // 3269 :   0 - 0x0
      13'hCC6: dout <= 8'b00000000; // 3270 :   0 - 0x0
      13'hCC7: dout <= 8'b00000000; // 3271 :   0 - 0x0
      13'hCC8: dout <= 8'b00000000; // 3272 :   0 - 0x0
      13'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      13'hCCA: dout <= 8'b00000000; // 3274 :   0 - 0x0
      13'hCCB: dout <= 8'b00000000; // 3275 :   0 - 0x0
      13'hCCC: dout <= 8'b00000000; // 3276 :   0 - 0x0
      13'hCCD: dout <= 8'b00000000; // 3277 :   0 - 0x0
      13'hCCE: dout <= 8'b00000000; // 3278 :   0 - 0x0
      13'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      13'hCD0: dout <= 8'b00000000; // 3280 :   0 - 0x0 -- Sprite 0xcd
      13'hCD1: dout <= 8'b00000000; // 3281 :   0 - 0x0
      13'hCD2: dout <= 8'b00000000; // 3282 :   0 - 0x0
      13'hCD3: dout <= 8'b00000000; // 3283 :   0 - 0x0
      13'hCD4: dout <= 8'b00000000; // 3284 :   0 - 0x0
      13'hCD5: dout <= 8'b00000000; // 3285 :   0 - 0x0
      13'hCD6: dout <= 8'b00000000; // 3286 :   0 - 0x0
      13'hCD7: dout <= 8'b00000000; // 3287 :   0 - 0x0
      13'hCD8: dout <= 8'b00000000; // 3288 :   0 - 0x0
      13'hCD9: dout <= 8'b00000000; // 3289 :   0 - 0x0
      13'hCDA: dout <= 8'b00000000; // 3290 :   0 - 0x0
      13'hCDB: dout <= 8'b00000000; // 3291 :   0 - 0x0
      13'hCDC: dout <= 8'b00000000; // 3292 :   0 - 0x0
      13'hCDD: dout <= 8'b00000000; // 3293 :   0 - 0x0
      13'hCDE: dout <= 8'b00000000; // 3294 :   0 - 0x0
      13'hCDF: dout <= 8'b00000000; // 3295 :   0 - 0x0
      13'hCE0: dout <= 8'b00000000; // 3296 :   0 - 0x0 -- Sprite 0xce
      13'hCE1: dout <= 8'b00000000; // 3297 :   0 - 0x0
      13'hCE2: dout <= 8'b00000000; // 3298 :   0 - 0x0
      13'hCE3: dout <= 8'b00000000; // 3299 :   0 - 0x0
      13'hCE4: dout <= 8'b00000000; // 3300 :   0 - 0x0
      13'hCE5: dout <= 8'b00000000; // 3301 :   0 - 0x0
      13'hCE6: dout <= 8'b00000000; // 3302 :   0 - 0x0
      13'hCE7: dout <= 8'b00000000; // 3303 :   0 - 0x0
      13'hCE8: dout <= 8'b00000000; // 3304 :   0 - 0x0
      13'hCE9: dout <= 8'b00000000; // 3305 :   0 - 0x0
      13'hCEA: dout <= 8'b00000000; // 3306 :   0 - 0x0
      13'hCEB: dout <= 8'b00000000; // 3307 :   0 - 0x0
      13'hCEC: dout <= 8'b00000000; // 3308 :   0 - 0x0
      13'hCED: dout <= 8'b00000000; // 3309 :   0 - 0x0
      13'hCEE: dout <= 8'b00000000; // 3310 :   0 - 0x0
      13'hCEF: dout <= 8'b00000000; // 3311 :   0 - 0x0
      13'hCF0: dout <= 8'b00000000; // 3312 :   0 - 0x0 -- Sprite 0xcf
      13'hCF1: dout <= 8'b00000000; // 3313 :   0 - 0x0
      13'hCF2: dout <= 8'b00000000; // 3314 :   0 - 0x0
      13'hCF3: dout <= 8'b00000000; // 3315 :   0 - 0x0
      13'hCF4: dout <= 8'b00000000; // 3316 :   0 - 0x0
      13'hCF5: dout <= 8'b00000000; // 3317 :   0 - 0x0
      13'hCF6: dout <= 8'b00000000; // 3318 :   0 - 0x0
      13'hCF7: dout <= 8'b00000000; // 3319 :   0 - 0x0
      13'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0
      13'hCF9: dout <= 8'b00000000; // 3321 :   0 - 0x0
      13'hCFA: dout <= 8'b00000000; // 3322 :   0 - 0x0
      13'hCFB: dout <= 8'b00000000; // 3323 :   0 - 0x0
      13'hCFC: dout <= 8'b00000000; // 3324 :   0 - 0x0
      13'hCFD: dout <= 8'b00000000; // 3325 :   0 - 0x0
      13'hCFE: dout <= 8'b00000000; // 3326 :   0 - 0x0
      13'hCFF: dout <= 8'b00000000; // 3327 :   0 - 0x0
      13'hD00: dout <= 8'b11111111; // 3328 : 255 - 0xff -- Sprite 0xd0
      13'hD01: dout <= 8'b11111111; // 3329 : 255 - 0xff
      13'hD02: dout <= 8'b11111111; // 3330 : 255 - 0xff
      13'hD03: dout <= 8'b11111111; // 3331 : 255 - 0xff
      13'hD04: dout <= 8'b11111111; // 3332 : 255 - 0xff
      13'hD05: dout <= 8'b11111111; // 3333 : 255 - 0xff
      13'hD06: dout <= 8'b11111111; // 3334 : 255 - 0xff
      13'hD07: dout <= 8'b11111111; // 3335 : 255 - 0xff
      13'hD08: dout <= 8'b11111111; // 3336 : 255 - 0xff
      13'hD09: dout <= 8'b11111111; // 3337 : 255 - 0xff
      13'hD0A: dout <= 8'b11111111; // 3338 : 255 - 0xff
      13'hD0B: dout <= 8'b11111111; // 3339 : 255 - 0xff
      13'hD0C: dout <= 8'b11111111; // 3340 : 255 - 0xff
      13'hD0D: dout <= 8'b11111111; // 3341 : 255 - 0xff
      13'hD0E: dout <= 8'b11111111; // 3342 : 255 - 0xff
      13'hD0F: dout <= 8'b11111111; // 3343 : 255 - 0xff
      13'hD10: dout <= 8'b11111111; // 3344 : 255 - 0xff -- Sprite 0xd1
      13'hD11: dout <= 8'b11111111; // 3345 : 255 - 0xff
      13'hD12: dout <= 8'b11111111; // 3346 : 255 - 0xff
      13'hD13: dout <= 8'b11111111; // 3347 : 255 - 0xff
      13'hD14: dout <= 8'b11111111; // 3348 : 255 - 0xff
      13'hD15: dout <= 8'b11111111; // 3349 : 255 - 0xff
      13'hD16: dout <= 8'b11111111; // 3350 : 255 - 0xff
      13'hD17: dout <= 8'b11111111; // 3351 : 255 - 0xff
      13'hD18: dout <= 8'b11111111; // 3352 : 255 - 0xff
      13'hD19: dout <= 8'b11111111; // 3353 : 255 - 0xff
      13'hD1A: dout <= 8'b11111111; // 3354 : 255 - 0xff
      13'hD1B: dout <= 8'b11111111; // 3355 : 255 - 0xff
      13'hD1C: dout <= 8'b11111111; // 3356 : 255 - 0xff
      13'hD1D: dout <= 8'b11111111; // 3357 : 255 - 0xff
      13'hD1E: dout <= 8'b11111111; // 3358 : 255 - 0xff
      13'hD1F: dout <= 8'b11111111; // 3359 : 255 - 0xff
      13'hD20: dout <= 8'b11111111; // 3360 : 255 - 0xff -- Sprite 0xd2
      13'hD21: dout <= 8'b11111111; // 3361 : 255 - 0xff
      13'hD22: dout <= 8'b11111111; // 3362 : 255 - 0xff
      13'hD23: dout <= 8'b11111111; // 3363 : 255 - 0xff
      13'hD24: dout <= 8'b11111111; // 3364 : 255 - 0xff
      13'hD25: dout <= 8'b11111111; // 3365 : 255 - 0xff
      13'hD26: dout <= 8'b11111111; // 3366 : 255 - 0xff
      13'hD27: dout <= 8'b11111111; // 3367 : 255 - 0xff
      13'hD28: dout <= 8'b11111111; // 3368 : 255 - 0xff
      13'hD29: dout <= 8'b11111111; // 3369 : 255 - 0xff
      13'hD2A: dout <= 8'b11111111; // 3370 : 255 - 0xff
      13'hD2B: dout <= 8'b11111111; // 3371 : 255 - 0xff
      13'hD2C: dout <= 8'b11111111; // 3372 : 255 - 0xff
      13'hD2D: dout <= 8'b11111111; // 3373 : 255 - 0xff
      13'hD2E: dout <= 8'b11111111; // 3374 : 255 - 0xff
      13'hD2F: dout <= 8'b11111111; // 3375 : 255 - 0xff
      13'hD30: dout <= 8'b11111111; // 3376 : 255 - 0xff -- Sprite 0xd3
      13'hD31: dout <= 8'b11111111; // 3377 : 255 - 0xff
      13'hD32: dout <= 8'b11111111; // 3378 : 255 - 0xff
      13'hD33: dout <= 8'b11111111; // 3379 : 255 - 0xff
      13'hD34: dout <= 8'b11111111; // 3380 : 255 - 0xff
      13'hD35: dout <= 8'b11111111; // 3381 : 255 - 0xff
      13'hD36: dout <= 8'b11111111; // 3382 : 255 - 0xff
      13'hD37: dout <= 8'b11111111; // 3383 : 255 - 0xff
      13'hD38: dout <= 8'b11111111; // 3384 : 255 - 0xff
      13'hD39: dout <= 8'b11111111; // 3385 : 255 - 0xff
      13'hD3A: dout <= 8'b11111111; // 3386 : 255 - 0xff
      13'hD3B: dout <= 8'b11111111; // 3387 : 255 - 0xff
      13'hD3C: dout <= 8'b11111111; // 3388 : 255 - 0xff
      13'hD3D: dout <= 8'b11111111; // 3389 : 255 - 0xff
      13'hD3E: dout <= 8'b11111111; // 3390 : 255 - 0xff
      13'hD3F: dout <= 8'b11111111; // 3391 : 255 - 0xff
      13'hD40: dout <= 8'b11111111; // 3392 : 255 - 0xff -- Sprite 0xd4
      13'hD41: dout <= 8'b11111111; // 3393 : 255 - 0xff
      13'hD42: dout <= 8'b11111111; // 3394 : 255 - 0xff
      13'hD43: dout <= 8'b11111111; // 3395 : 255 - 0xff
      13'hD44: dout <= 8'b11111111; // 3396 : 255 - 0xff
      13'hD45: dout <= 8'b11111111; // 3397 : 255 - 0xff
      13'hD46: dout <= 8'b11111111; // 3398 : 255 - 0xff
      13'hD47: dout <= 8'b11111111; // 3399 : 255 - 0xff
      13'hD48: dout <= 8'b11111111; // 3400 : 255 - 0xff
      13'hD49: dout <= 8'b11111111; // 3401 : 255 - 0xff
      13'hD4A: dout <= 8'b11111111; // 3402 : 255 - 0xff
      13'hD4B: dout <= 8'b11111111; // 3403 : 255 - 0xff
      13'hD4C: dout <= 8'b11111111; // 3404 : 255 - 0xff
      13'hD4D: dout <= 8'b11111111; // 3405 : 255 - 0xff
      13'hD4E: dout <= 8'b11111111; // 3406 : 255 - 0xff
      13'hD4F: dout <= 8'b11111111; // 3407 : 255 - 0xff
      13'hD50: dout <= 8'b11111111; // 3408 : 255 - 0xff -- Sprite 0xd5
      13'hD51: dout <= 8'b11111111; // 3409 : 255 - 0xff
      13'hD52: dout <= 8'b11111111; // 3410 : 255 - 0xff
      13'hD53: dout <= 8'b11111111; // 3411 : 255 - 0xff
      13'hD54: dout <= 8'b11111111; // 3412 : 255 - 0xff
      13'hD55: dout <= 8'b11111111; // 3413 : 255 - 0xff
      13'hD56: dout <= 8'b11111111; // 3414 : 255 - 0xff
      13'hD57: dout <= 8'b11111111; // 3415 : 255 - 0xff
      13'hD58: dout <= 8'b11111111; // 3416 : 255 - 0xff
      13'hD59: dout <= 8'b11111111; // 3417 : 255 - 0xff
      13'hD5A: dout <= 8'b11111111; // 3418 : 255 - 0xff
      13'hD5B: dout <= 8'b11111111; // 3419 : 255 - 0xff
      13'hD5C: dout <= 8'b11111111; // 3420 : 255 - 0xff
      13'hD5D: dout <= 8'b11111111; // 3421 : 255 - 0xff
      13'hD5E: dout <= 8'b11111111; // 3422 : 255 - 0xff
      13'hD5F: dout <= 8'b11111111; // 3423 : 255 - 0xff
      13'hD60: dout <= 8'b11111111; // 3424 : 255 - 0xff -- Sprite 0xd6
      13'hD61: dout <= 8'b11111111; // 3425 : 255 - 0xff
      13'hD62: dout <= 8'b11111111; // 3426 : 255 - 0xff
      13'hD63: dout <= 8'b11111111; // 3427 : 255 - 0xff
      13'hD64: dout <= 8'b11111111; // 3428 : 255 - 0xff
      13'hD65: dout <= 8'b11111111; // 3429 : 255 - 0xff
      13'hD66: dout <= 8'b11111111; // 3430 : 255 - 0xff
      13'hD67: dout <= 8'b11111111; // 3431 : 255 - 0xff
      13'hD68: dout <= 8'b11111111; // 3432 : 255 - 0xff
      13'hD69: dout <= 8'b11111111; // 3433 : 255 - 0xff
      13'hD6A: dout <= 8'b11111111; // 3434 : 255 - 0xff
      13'hD6B: dout <= 8'b11111111; // 3435 : 255 - 0xff
      13'hD6C: dout <= 8'b11111111; // 3436 : 255 - 0xff
      13'hD6D: dout <= 8'b11111111; // 3437 : 255 - 0xff
      13'hD6E: dout <= 8'b11111111; // 3438 : 255 - 0xff
      13'hD6F: dout <= 8'b11111111; // 3439 : 255 - 0xff
      13'hD70: dout <= 8'b11111111; // 3440 : 255 - 0xff -- Sprite 0xd7
      13'hD71: dout <= 8'b11111111; // 3441 : 255 - 0xff
      13'hD72: dout <= 8'b11111111; // 3442 : 255 - 0xff
      13'hD73: dout <= 8'b11111111; // 3443 : 255 - 0xff
      13'hD74: dout <= 8'b11111111; // 3444 : 255 - 0xff
      13'hD75: dout <= 8'b11111111; // 3445 : 255 - 0xff
      13'hD76: dout <= 8'b11111111; // 3446 : 255 - 0xff
      13'hD77: dout <= 8'b11111111; // 3447 : 255 - 0xff
      13'hD78: dout <= 8'b11111111; // 3448 : 255 - 0xff
      13'hD79: dout <= 8'b11111111; // 3449 : 255 - 0xff
      13'hD7A: dout <= 8'b11111111; // 3450 : 255 - 0xff
      13'hD7B: dout <= 8'b11111111; // 3451 : 255 - 0xff
      13'hD7C: dout <= 8'b11111111; // 3452 : 255 - 0xff
      13'hD7D: dout <= 8'b11111111; // 3453 : 255 - 0xff
      13'hD7E: dout <= 8'b11111111; // 3454 : 255 - 0xff
      13'hD7F: dout <= 8'b11111111; // 3455 : 255 - 0xff
      13'hD80: dout <= 8'b11111111; // 3456 : 255 - 0xff -- Sprite 0xd8
      13'hD81: dout <= 8'b11111111; // 3457 : 255 - 0xff
      13'hD82: dout <= 8'b11111111; // 3458 : 255 - 0xff
      13'hD83: dout <= 8'b11111111; // 3459 : 255 - 0xff
      13'hD84: dout <= 8'b11111111; // 3460 : 255 - 0xff
      13'hD85: dout <= 8'b11111111; // 3461 : 255 - 0xff
      13'hD86: dout <= 8'b11111111; // 3462 : 255 - 0xff
      13'hD87: dout <= 8'b11111111; // 3463 : 255 - 0xff
      13'hD88: dout <= 8'b11111111; // 3464 : 255 - 0xff
      13'hD89: dout <= 8'b11111111; // 3465 : 255 - 0xff
      13'hD8A: dout <= 8'b11111111; // 3466 : 255 - 0xff
      13'hD8B: dout <= 8'b11111111; // 3467 : 255 - 0xff
      13'hD8C: dout <= 8'b11111111; // 3468 : 255 - 0xff
      13'hD8D: dout <= 8'b11111111; // 3469 : 255 - 0xff
      13'hD8E: dout <= 8'b11111111; // 3470 : 255 - 0xff
      13'hD8F: dout <= 8'b11111111; // 3471 : 255 - 0xff
      13'hD90: dout <= 8'b11111111; // 3472 : 255 - 0xff -- Sprite 0xd9
      13'hD91: dout <= 8'b11111111; // 3473 : 255 - 0xff
      13'hD92: dout <= 8'b11111111; // 3474 : 255 - 0xff
      13'hD93: dout <= 8'b11111111; // 3475 : 255 - 0xff
      13'hD94: dout <= 8'b11111111; // 3476 : 255 - 0xff
      13'hD95: dout <= 8'b11111111; // 3477 : 255 - 0xff
      13'hD96: dout <= 8'b11111111; // 3478 : 255 - 0xff
      13'hD97: dout <= 8'b11111111; // 3479 : 255 - 0xff
      13'hD98: dout <= 8'b11111111; // 3480 : 255 - 0xff
      13'hD99: dout <= 8'b11111111; // 3481 : 255 - 0xff
      13'hD9A: dout <= 8'b11111111; // 3482 : 255 - 0xff
      13'hD9B: dout <= 8'b11111111; // 3483 : 255 - 0xff
      13'hD9C: dout <= 8'b11111111; // 3484 : 255 - 0xff
      13'hD9D: dout <= 8'b11111111; // 3485 : 255 - 0xff
      13'hD9E: dout <= 8'b11111111; // 3486 : 255 - 0xff
      13'hD9F: dout <= 8'b11111111; // 3487 : 255 - 0xff
      13'hDA0: dout <= 8'b11111111; // 3488 : 255 - 0xff -- Sprite 0xda
      13'hDA1: dout <= 8'b11111111; // 3489 : 255 - 0xff
      13'hDA2: dout <= 8'b11111111; // 3490 : 255 - 0xff
      13'hDA3: dout <= 8'b11111111; // 3491 : 255 - 0xff
      13'hDA4: dout <= 8'b11111111; // 3492 : 255 - 0xff
      13'hDA5: dout <= 8'b11111111; // 3493 : 255 - 0xff
      13'hDA6: dout <= 8'b11111111; // 3494 : 255 - 0xff
      13'hDA7: dout <= 8'b11111111; // 3495 : 255 - 0xff
      13'hDA8: dout <= 8'b11111111; // 3496 : 255 - 0xff
      13'hDA9: dout <= 8'b11111111; // 3497 : 255 - 0xff
      13'hDAA: dout <= 8'b11111111; // 3498 : 255 - 0xff
      13'hDAB: dout <= 8'b11111111; // 3499 : 255 - 0xff
      13'hDAC: dout <= 8'b11111111; // 3500 : 255 - 0xff
      13'hDAD: dout <= 8'b11111111; // 3501 : 255 - 0xff
      13'hDAE: dout <= 8'b11111111; // 3502 : 255 - 0xff
      13'hDAF: dout <= 8'b11111111; // 3503 : 255 - 0xff
      13'hDB0: dout <= 8'b11111111; // 3504 : 255 - 0xff -- Sprite 0xdb
      13'hDB1: dout <= 8'b11111111; // 3505 : 255 - 0xff
      13'hDB2: dout <= 8'b11111111; // 3506 : 255 - 0xff
      13'hDB3: dout <= 8'b11111111; // 3507 : 255 - 0xff
      13'hDB4: dout <= 8'b11111111; // 3508 : 255 - 0xff
      13'hDB5: dout <= 8'b11111111; // 3509 : 255 - 0xff
      13'hDB6: dout <= 8'b11111111; // 3510 : 255 - 0xff
      13'hDB7: dout <= 8'b11111111; // 3511 : 255 - 0xff
      13'hDB8: dout <= 8'b11111111; // 3512 : 255 - 0xff
      13'hDB9: dout <= 8'b11111111; // 3513 : 255 - 0xff
      13'hDBA: dout <= 8'b11111111; // 3514 : 255 - 0xff
      13'hDBB: dout <= 8'b11111111; // 3515 : 255 - 0xff
      13'hDBC: dout <= 8'b11111111; // 3516 : 255 - 0xff
      13'hDBD: dout <= 8'b11111111; // 3517 : 255 - 0xff
      13'hDBE: dout <= 8'b11111111; // 3518 : 255 - 0xff
      13'hDBF: dout <= 8'b11111111; // 3519 : 255 - 0xff
      13'hDC0: dout <= 8'b11111111; // 3520 : 255 - 0xff -- Sprite 0xdc
      13'hDC1: dout <= 8'b11111111; // 3521 : 255 - 0xff
      13'hDC2: dout <= 8'b11111111; // 3522 : 255 - 0xff
      13'hDC3: dout <= 8'b11111111; // 3523 : 255 - 0xff
      13'hDC4: dout <= 8'b11111111; // 3524 : 255 - 0xff
      13'hDC5: dout <= 8'b11111111; // 3525 : 255 - 0xff
      13'hDC6: dout <= 8'b11111111; // 3526 : 255 - 0xff
      13'hDC7: dout <= 8'b11111111; // 3527 : 255 - 0xff
      13'hDC8: dout <= 8'b11111111; // 3528 : 255 - 0xff
      13'hDC9: dout <= 8'b11111111; // 3529 : 255 - 0xff
      13'hDCA: dout <= 8'b11111111; // 3530 : 255 - 0xff
      13'hDCB: dout <= 8'b11111111; // 3531 : 255 - 0xff
      13'hDCC: dout <= 8'b11111111; // 3532 : 255 - 0xff
      13'hDCD: dout <= 8'b11111111; // 3533 : 255 - 0xff
      13'hDCE: dout <= 8'b11111111; // 3534 : 255 - 0xff
      13'hDCF: dout <= 8'b11111111; // 3535 : 255 - 0xff
      13'hDD0: dout <= 8'b11111111; // 3536 : 255 - 0xff -- Sprite 0xdd
      13'hDD1: dout <= 8'b11111111; // 3537 : 255 - 0xff
      13'hDD2: dout <= 8'b11111111; // 3538 : 255 - 0xff
      13'hDD3: dout <= 8'b11111111; // 3539 : 255 - 0xff
      13'hDD4: dout <= 8'b11111111; // 3540 : 255 - 0xff
      13'hDD5: dout <= 8'b11111111; // 3541 : 255 - 0xff
      13'hDD6: dout <= 8'b11111111; // 3542 : 255 - 0xff
      13'hDD7: dout <= 8'b11111111; // 3543 : 255 - 0xff
      13'hDD8: dout <= 8'b11111111; // 3544 : 255 - 0xff
      13'hDD9: dout <= 8'b11111111; // 3545 : 255 - 0xff
      13'hDDA: dout <= 8'b11111111; // 3546 : 255 - 0xff
      13'hDDB: dout <= 8'b11111111; // 3547 : 255 - 0xff
      13'hDDC: dout <= 8'b11111111; // 3548 : 255 - 0xff
      13'hDDD: dout <= 8'b11111111; // 3549 : 255 - 0xff
      13'hDDE: dout <= 8'b11111111; // 3550 : 255 - 0xff
      13'hDDF: dout <= 8'b11111111; // 3551 : 255 - 0xff
      13'hDE0: dout <= 8'b11111111; // 3552 : 255 - 0xff -- Sprite 0xde
      13'hDE1: dout <= 8'b11111111; // 3553 : 255 - 0xff
      13'hDE2: dout <= 8'b11111111; // 3554 : 255 - 0xff
      13'hDE3: dout <= 8'b11111111; // 3555 : 255 - 0xff
      13'hDE4: dout <= 8'b11111111; // 3556 : 255 - 0xff
      13'hDE5: dout <= 8'b11111111; // 3557 : 255 - 0xff
      13'hDE6: dout <= 8'b11111111; // 3558 : 255 - 0xff
      13'hDE7: dout <= 8'b11111111; // 3559 : 255 - 0xff
      13'hDE8: dout <= 8'b11111111; // 3560 : 255 - 0xff
      13'hDE9: dout <= 8'b11111111; // 3561 : 255 - 0xff
      13'hDEA: dout <= 8'b11111111; // 3562 : 255 - 0xff
      13'hDEB: dout <= 8'b11111111; // 3563 : 255 - 0xff
      13'hDEC: dout <= 8'b11111111; // 3564 : 255 - 0xff
      13'hDED: dout <= 8'b11111111; // 3565 : 255 - 0xff
      13'hDEE: dout <= 8'b11111111; // 3566 : 255 - 0xff
      13'hDEF: dout <= 8'b11111111; // 3567 : 255 - 0xff
      13'hDF0: dout <= 8'b11111111; // 3568 : 255 - 0xff -- Sprite 0xdf
      13'hDF1: dout <= 8'b11111111; // 3569 : 255 - 0xff
      13'hDF2: dout <= 8'b11111111; // 3570 : 255 - 0xff
      13'hDF3: dout <= 8'b11111111; // 3571 : 255 - 0xff
      13'hDF4: dout <= 8'b11111111; // 3572 : 255 - 0xff
      13'hDF5: dout <= 8'b11111111; // 3573 : 255 - 0xff
      13'hDF6: dout <= 8'b11111111; // 3574 : 255 - 0xff
      13'hDF7: dout <= 8'b11111111; // 3575 : 255 - 0xff
      13'hDF8: dout <= 8'b11111111; // 3576 : 255 - 0xff
      13'hDF9: dout <= 8'b11111111; // 3577 : 255 - 0xff
      13'hDFA: dout <= 8'b11111111; // 3578 : 255 - 0xff
      13'hDFB: dout <= 8'b11111111; // 3579 : 255 - 0xff
      13'hDFC: dout <= 8'b11111111; // 3580 : 255 - 0xff
      13'hDFD: dout <= 8'b11111111; // 3581 : 255 - 0xff
      13'hDFE: dout <= 8'b11111111; // 3582 : 255 - 0xff
      13'hDFF: dout <= 8'b11111111; // 3583 : 255 - 0xff
      13'hE00: dout <= 8'b11111111; // 3584 : 255 - 0xff -- Sprite 0xe0
      13'hE01: dout <= 8'b11111111; // 3585 : 255 - 0xff
      13'hE02: dout <= 8'b11111111; // 3586 : 255 - 0xff
      13'hE03: dout <= 8'b11111111; // 3587 : 255 - 0xff
      13'hE04: dout <= 8'b11111111; // 3588 : 255 - 0xff
      13'hE05: dout <= 8'b11111111; // 3589 : 255 - 0xff
      13'hE06: dout <= 8'b11111111; // 3590 : 255 - 0xff
      13'hE07: dout <= 8'b11111111; // 3591 : 255 - 0xff
      13'hE08: dout <= 8'b11111111; // 3592 : 255 - 0xff
      13'hE09: dout <= 8'b11111111; // 3593 : 255 - 0xff
      13'hE0A: dout <= 8'b11111111; // 3594 : 255 - 0xff
      13'hE0B: dout <= 8'b11111111; // 3595 : 255 - 0xff
      13'hE0C: dout <= 8'b11111111; // 3596 : 255 - 0xff
      13'hE0D: dout <= 8'b11111111; // 3597 : 255 - 0xff
      13'hE0E: dout <= 8'b11111111; // 3598 : 255 - 0xff
      13'hE0F: dout <= 8'b11111111; // 3599 : 255 - 0xff
      13'hE10: dout <= 8'b11111111; // 3600 : 255 - 0xff -- Sprite 0xe1
      13'hE11: dout <= 8'b11111111; // 3601 : 255 - 0xff
      13'hE12: dout <= 8'b11111111; // 3602 : 255 - 0xff
      13'hE13: dout <= 8'b11111111; // 3603 : 255 - 0xff
      13'hE14: dout <= 8'b11111111; // 3604 : 255 - 0xff
      13'hE15: dout <= 8'b11111111; // 3605 : 255 - 0xff
      13'hE16: dout <= 8'b11111111; // 3606 : 255 - 0xff
      13'hE17: dout <= 8'b11111111; // 3607 : 255 - 0xff
      13'hE18: dout <= 8'b11111111; // 3608 : 255 - 0xff
      13'hE19: dout <= 8'b11111111; // 3609 : 255 - 0xff
      13'hE1A: dout <= 8'b11111111; // 3610 : 255 - 0xff
      13'hE1B: dout <= 8'b11111111; // 3611 : 255 - 0xff
      13'hE1C: dout <= 8'b11111111; // 3612 : 255 - 0xff
      13'hE1D: dout <= 8'b11111111; // 3613 : 255 - 0xff
      13'hE1E: dout <= 8'b11111111; // 3614 : 255 - 0xff
      13'hE1F: dout <= 8'b11111111; // 3615 : 255 - 0xff
      13'hE20: dout <= 8'b11111111; // 3616 : 255 - 0xff -- Sprite 0xe2
      13'hE21: dout <= 8'b11111111; // 3617 : 255 - 0xff
      13'hE22: dout <= 8'b11111111; // 3618 : 255 - 0xff
      13'hE23: dout <= 8'b11111111; // 3619 : 255 - 0xff
      13'hE24: dout <= 8'b11111111; // 3620 : 255 - 0xff
      13'hE25: dout <= 8'b11111111; // 3621 : 255 - 0xff
      13'hE26: dout <= 8'b11111111; // 3622 : 255 - 0xff
      13'hE27: dout <= 8'b11111111; // 3623 : 255 - 0xff
      13'hE28: dout <= 8'b11111111; // 3624 : 255 - 0xff
      13'hE29: dout <= 8'b11111111; // 3625 : 255 - 0xff
      13'hE2A: dout <= 8'b11111111; // 3626 : 255 - 0xff
      13'hE2B: dout <= 8'b11111111; // 3627 : 255 - 0xff
      13'hE2C: dout <= 8'b11111111; // 3628 : 255 - 0xff
      13'hE2D: dout <= 8'b11111111; // 3629 : 255 - 0xff
      13'hE2E: dout <= 8'b11111111; // 3630 : 255 - 0xff
      13'hE2F: dout <= 8'b11111111; // 3631 : 255 - 0xff
      13'hE30: dout <= 8'b11111111; // 3632 : 255 - 0xff -- Sprite 0xe3
      13'hE31: dout <= 8'b11111111; // 3633 : 255 - 0xff
      13'hE32: dout <= 8'b11111111; // 3634 : 255 - 0xff
      13'hE33: dout <= 8'b11111111; // 3635 : 255 - 0xff
      13'hE34: dout <= 8'b11111111; // 3636 : 255 - 0xff
      13'hE35: dout <= 8'b11111111; // 3637 : 255 - 0xff
      13'hE36: dout <= 8'b11111111; // 3638 : 255 - 0xff
      13'hE37: dout <= 8'b11111111; // 3639 : 255 - 0xff
      13'hE38: dout <= 8'b11111111; // 3640 : 255 - 0xff
      13'hE39: dout <= 8'b11111111; // 3641 : 255 - 0xff
      13'hE3A: dout <= 8'b11111111; // 3642 : 255 - 0xff
      13'hE3B: dout <= 8'b11111111; // 3643 : 255 - 0xff
      13'hE3C: dout <= 8'b11111111; // 3644 : 255 - 0xff
      13'hE3D: dout <= 8'b11111111; // 3645 : 255 - 0xff
      13'hE3E: dout <= 8'b11111111; // 3646 : 255 - 0xff
      13'hE3F: dout <= 8'b11111111; // 3647 : 255 - 0xff
      13'hE40: dout <= 8'b11111111; // 3648 : 255 - 0xff -- Sprite 0xe4
      13'hE41: dout <= 8'b11111111; // 3649 : 255 - 0xff
      13'hE42: dout <= 8'b11111111; // 3650 : 255 - 0xff
      13'hE43: dout <= 8'b11111111; // 3651 : 255 - 0xff
      13'hE44: dout <= 8'b11111111; // 3652 : 255 - 0xff
      13'hE45: dout <= 8'b11111111; // 3653 : 255 - 0xff
      13'hE46: dout <= 8'b11111111; // 3654 : 255 - 0xff
      13'hE47: dout <= 8'b11111111; // 3655 : 255 - 0xff
      13'hE48: dout <= 8'b11111111; // 3656 : 255 - 0xff
      13'hE49: dout <= 8'b11111111; // 3657 : 255 - 0xff
      13'hE4A: dout <= 8'b11111111; // 3658 : 255 - 0xff
      13'hE4B: dout <= 8'b11111111; // 3659 : 255 - 0xff
      13'hE4C: dout <= 8'b11111111; // 3660 : 255 - 0xff
      13'hE4D: dout <= 8'b11111111; // 3661 : 255 - 0xff
      13'hE4E: dout <= 8'b11111111; // 3662 : 255 - 0xff
      13'hE4F: dout <= 8'b11111111; // 3663 : 255 - 0xff
      13'hE50: dout <= 8'b11111111; // 3664 : 255 - 0xff -- Sprite 0xe5
      13'hE51: dout <= 8'b11111111; // 3665 : 255 - 0xff
      13'hE52: dout <= 8'b11111111; // 3666 : 255 - 0xff
      13'hE53: dout <= 8'b11111111; // 3667 : 255 - 0xff
      13'hE54: dout <= 8'b11111111; // 3668 : 255 - 0xff
      13'hE55: dout <= 8'b11111111; // 3669 : 255 - 0xff
      13'hE56: dout <= 8'b11111111; // 3670 : 255 - 0xff
      13'hE57: dout <= 8'b11111111; // 3671 : 255 - 0xff
      13'hE58: dout <= 8'b11111111; // 3672 : 255 - 0xff
      13'hE59: dout <= 8'b11111111; // 3673 : 255 - 0xff
      13'hE5A: dout <= 8'b11111111; // 3674 : 255 - 0xff
      13'hE5B: dout <= 8'b11111111; // 3675 : 255 - 0xff
      13'hE5C: dout <= 8'b11111111; // 3676 : 255 - 0xff
      13'hE5D: dout <= 8'b11111111; // 3677 : 255 - 0xff
      13'hE5E: dout <= 8'b11111111; // 3678 : 255 - 0xff
      13'hE5F: dout <= 8'b11111111; // 3679 : 255 - 0xff
      13'hE60: dout <= 8'b11111111; // 3680 : 255 - 0xff -- Sprite 0xe6
      13'hE61: dout <= 8'b11111111; // 3681 : 255 - 0xff
      13'hE62: dout <= 8'b11111111; // 3682 : 255 - 0xff
      13'hE63: dout <= 8'b11111111; // 3683 : 255 - 0xff
      13'hE64: dout <= 8'b11111111; // 3684 : 255 - 0xff
      13'hE65: dout <= 8'b11111111; // 3685 : 255 - 0xff
      13'hE66: dout <= 8'b11111111; // 3686 : 255 - 0xff
      13'hE67: dout <= 8'b11111111; // 3687 : 255 - 0xff
      13'hE68: dout <= 8'b11111111; // 3688 : 255 - 0xff
      13'hE69: dout <= 8'b11111111; // 3689 : 255 - 0xff
      13'hE6A: dout <= 8'b11111111; // 3690 : 255 - 0xff
      13'hE6B: dout <= 8'b11111111; // 3691 : 255 - 0xff
      13'hE6C: dout <= 8'b11111111; // 3692 : 255 - 0xff
      13'hE6D: dout <= 8'b11111111; // 3693 : 255 - 0xff
      13'hE6E: dout <= 8'b11111111; // 3694 : 255 - 0xff
      13'hE6F: dout <= 8'b11111111; // 3695 : 255 - 0xff
      13'hE70: dout <= 8'b11111111; // 3696 : 255 - 0xff -- Sprite 0xe7
      13'hE71: dout <= 8'b11111111; // 3697 : 255 - 0xff
      13'hE72: dout <= 8'b11111111; // 3698 : 255 - 0xff
      13'hE73: dout <= 8'b11111111; // 3699 : 255 - 0xff
      13'hE74: dout <= 8'b11111111; // 3700 : 255 - 0xff
      13'hE75: dout <= 8'b11111111; // 3701 : 255 - 0xff
      13'hE76: dout <= 8'b11111111; // 3702 : 255 - 0xff
      13'hE77: dout <= 8'b11111111; // 3703 : 255 - 0xff
      13'hE78: dout <= 8'b11111111; // 3704 : 255 - 0xff
      13'hE79: dout <= 8'b11111111; // 3705 : 255 - 0xff
      13'hE7A: dout <= 8'b11111111; // 3706 : 255 - 0xff
      13'hE7B: dout <= 8'b11111111; // 3707 : 255 - 0xff
      13'hE7C: dout <= 8'b11111111; // 3708 : 255 - 0xff
      13'hE7D: dout <= 8'b11111111; // 3709 : 255 - 0xff
      13'hE7E: dout <= 8'b11111111; // 3710 : 255 - 0xff
      13'hE7F: dout <= 8'b11111111; // 3711 : 255 - 0xff
      13'hE80: dout <= 8'b11111111; // 3712 : 255 - 0xff -- Sprite 0xe8
      13'hE81: dout <= 8'b11111111; // 3713 : 255 - 0xff
      13'hE82: dout <= 8'b11111111; // 3714 : 255 - 0xff
      13'hE83: dout <= 8'b11111111; // 3715 : 255 - 0xff
      13'hE84: dout <= 8'b11111111; // 3716 : 255 - 0xff
      13'hE85: dout <= 8'b11111111; // 3717 : 255 - 0xff
      13'hE86: dout <= 8'b11111111; // 3718 : 255 - 0xff
      13'hE87: dout <= 8'b11111111; // 3719 : 255 - 0xff
      13'hE88: dout <= 8'b11111111; // 3720 : 255 - 0xff
      13'hE89: dout <= 8'b11111111; // 3721 : 255 - 0xff
      13'hE8A: dout <= 8'b11111111; // 3722 : 255 - 0xff
      13'hE8B: dout <= 8'b11111111; // 3723 : 255 - 0xff
      13'hE8C: dout <= 8'b11111111; // 3724 : 255 - 0xff
      13'hE8D: dout <= 8'b11111111; // 3725 : 255 - 0xff
      13'hE8E: dout <= 8'b11111111; // 3726 : 255 - 0xff
      13'hE8F: dout <= 8'b11111111; // 3727 : 255 - 0xff
      13'hE90: dout <= 8'b11111111; // 3728 : 255 - 0xff -- Sprite 0xe9
      13'hE91: dout <= 8'b11111111; // 3729 : 255 - 0xff
      13'hE92: dout <= 8'b11111111; // 3730 : 255 - 0xff
      13'hE93: dout <= 8'b11111111; // 3731 : 255 - 0xff
      13'hE94: dout <= 8'b11111111; // 3732 : 255 - 0xff
      13'hE95: dout <= 8'b11111111; // 3733 : 255 - 0xff
      13'hE96: dout <= 8'b11111111; // 3734 : 255 - 0xff
      13'hE97: dout <= 8'b11111111; // 3735 : 255 - 0xff
      13'hE98: dout <= 8'b11111111; // 3736 : 255 - 0xff
      13'hE99: dout <= 8'b11111111; // 3737 : 255 - 0xff
      13'hE9A: dout <= 8'b11111111; // 3738 : 255 - 0xff
      13'hE9B: dout <= 8'b11111111; // 3739 : 255 - 0xff
      13'hE9C: dout <= 8'b11111111; // 3740 : 255 - 0xff
      13'hE9D: dout <= 8'b11111111; // 3741 : 255 - 0xff
      13'hE9E: dout <= 8'b11111111; // 3742 : 255 - 0xff
      13'hE9F: dout <= 8'b11111111; // 3743 : 255 - 0xff
      13'hEA0: dout <= 8'b11111111; // 3744 : 255 - 0xff -- Sprite 0xea
      13'hEA1: dout <= 8'b11111111; // 3745 : 255 - 0xff
      13'hEA2: dout <= 8'b11111111; // 3746 : 255 - 0xff
      13'hEA3: dout <= 8'b11111111; // 3747 : 255 - 0xff
      13'hEA4: dout <= 8'b11111111; // 3748 : 255 - 0xff
      13'hEA5: dout <= 8'b11111111; // 3749 : 255 - 0xff
      13'hEA6: dout <= 8'b11111111; // 3750 : 255 - 0xff
      13'hEA7: dout <= 8'b11111111; // 3751 : 255 - 0xff
      13'hEA8: dout <= 8'b11111111; // 3752 : 255 - 0xff
      13'hEA9: dout <= 8'b11111111; // 3753 : 255 - 0xff
      13'hEAA: dout <= 8'b11111111; // 3754 : 255 - 0xff
      13'hEAB: dout <= 8'b11111111; // 3755 : 255 - 0xff
      13'hEAC: dout <= 8'b11111111; // 3756 : 255 - 0xff
      13'hEAD: dout <= 8'b11111111; // 3757 : 255 - 0xff
      13'hEAE: dout <= 8'b11111111; // 3758 : 255 - 0xff
      13'hEAF: dout <= 8'b11111111; // 3759 : 255 - 0xff
      13'hEB0: dout <= 8'b11111111; // 3760 : 255 - 0xff -- Sprite 0xeb
      13'hEB1: dout <= 8'b11111111; // 3761 : 255 - 0xff
      13'hEB2: dout <= 8'b11111111; // 3762 : 255 - 0xff
      13'hEB3: dout <= 8'b11111111; // 3763 : 255 - 0xff
      13'hEB4: dout <= 8'b11111111; // 3764 : 255 - 0xff
      13'hEB5: dout <= 8'b11111111; // 3765 : 255 - 0xff
      13'hEB6: dout <= 8'b11111111; // 3766 : 255 - 0xff
      13'hEB7: dout <= 8'b11111111; // 3767 : 255 - 0xff
      13'hEB8: dout <= 8'b11111111; // 3768 : 255 - 0xff
      13'hEB9: dout <= 8'b11111111; // 3769 : 255 - 0xff
      13'hEBA: dout <= 8'b11111111; // 3770 : 255 - 0xff
      13'hEBB: dout <= 8'b11111111; // 3771 : 255 - 0xff
      13'hEBC: dout <= 8'b11111111; // 3772 : 255 - 0xff
      13'hEBD: dout <= 8'b11111111; // 3773 : 255 - 0xff
      13'hEBE: dout <= 8'b11111111; // 3774 : 255 - 0xff
      13'hEBF: dout <= 8'b11111111; // 3775 : 255 - 0xff
      13'hEC0: dout <= 8'b11111111; // 3776 : 255 - 0xff -- Sprite 0xec
      13'hEC1: dout <= 8'b11111111; // 3777 : 255 - 0xff
      13'hEC2: dout <= 8'b11111111; // 3778 : 255 - 0xff
      13'hEC3: dout <= 8'b11111111; // 3779 : 255 - 0xff
      13'hEC4: dout <= 8'b11111111; // 3780 : 255 - 0xff
      13'hEC5: dout <= 8'b11111111; // 3781 : 255 - 0xff
      13'hEC6: dout <= 8'b11111111; // 3782 : 255 - 0xff
      13'hEC7: dout <= 8'b11111111; // 3783 : 255 - 0xff
      13'hEC8: dout <= 8'b11111111; // 3784 : 255 - 0xff
      13'hEC9: dout <= 8'b11111111; // 3785 : 255 - 0xff
      13'hECA: dout <= 8'b11111111; // 3786 : 255 - 0xff
      13'hECB: dout <= 8'b11111111; // 3787 : 255 - 0xff
      13'hECC: dout <= 8'b11111111; // 3788 : 255 - 0xff
      13'hECD: dout <= 8'b11111111; // 3789 : 255 - 0xff
      13'hECE: dout <= 8'b11111111; // 3790 : 255 - 0xff
      13'hECF: dout <= 8'b11111111; // 3791 : 255 - 0xff
      13'hED0: dout <= 8'b11111111; // 3792 : 255 - 0xff -- Sprite 0xed
      13'hED1: dout <= 8'b11111111; // 3793 : 255 - 0xff
      13'hED2: dout <= 8'b11111111; // 3794 : 255 - 0xff
      13'hED3: dout <= 8'b11111111; // 3795 : 255 - 0xff
      13'hED4: dout <= 8'b11111111; // 3796 : 255 - 0xff
      13'hED5: dout <= 8'b11111111; // 3797 : 255 - 0xff
      13'hED6: dout <= 8'b11111111; // 3798 : 255 - 0xff
      13'hED7: dout <= 8'b11111111; // 3799 : 255 - 0xff
      13'hED8: dout <= 8'b11111111; // 3800 : 255 - 0xff
      13'hED9: dout <= 8'b11111111; // 3801 : 255 - 0xff
      13'hEDA: dout <= 8'b11111111; // 3802 : 255 - 0xff
      13'hEDB: dout <= 8'b11111111; // 3803 : 255 - 0xff
      13'hEDC: dout <= 8'b11111111; // 3804 : 255 - 0xff
      13'hEDD: dout <= 8'b11111111; // 3805 : 255 - 0xff
      13'hEDE: dout <= 8'b11111111; // 3806 : 255 - 0xff
      13'hEDF: dout <= 8'b11111111; // 3807 : 255 - 0xff
      13'hEE0: dout <= 8'b11111111; // 3808 : 255 - 0xff -- Sprite 0xee
      13'hEE1: dout <= 8'b11111111; // 3809 : 255 - 0xff
      13'hEE2: dout <= 8'b11111111; // 3810 : 255 - 0xff
      13'hEE3: dout <= 8'b11111111; // 3811 : 255 - 0xff
      13'hEE4: dout <= 8'b11111111; // 3812 : 255 - 0xff
      13'hEE5: dout <= 8'b11111111; // 3813 : 255 - 0xff
      13'hEE6: dout <= 8'b11111111; // 3814 : 255 - 0xff
      13'hEE7: dout <= 8'b11111111; // 3815 : 255 - 0xff
      13'hEE8: dout <= 8'b11111111; // 3816 : 255 - 0xff
      13'hEE9: dout <= 8'b11111111; // 3817 : 255 - 0xff
      13'hEEA: dout <= 8'b11111111; // 3818 : 255 - 0xff
      13'hEEB: dout <= 8'b11111111; // 3819 : 255 - 0xff
      13'hEEC: dout <= 8'b11111111; // 3820 : 255 - 0xff
      13'hEED: dout <= 8'b11111111; // 3821 : 255 - 0xff
      13'hEEE: dout <= 8'b11111111; // 3822 : 255 - 0xff
      13'hEEF: dout <= 8'b11111111; // 3823 : 255 - 0xff
      13'hEF0: dout <= 8'b11111111; // 3824 : 255 - 0xff -- Sprite 0xef
      13'hEF1: dout <= 8'b11111111; // 3825 : 255 - 0xff
      13'hEF2: dout <= 8'b11111111; // 3826 : 255 - 0xff
      13'hEF3: dout <= 8'b11111111; // 3827 : 255 - 0xff
      13'hEF4: dout <= 8'b11111111; // 3828 : 255 - 0xff
      13'hEF5: dout <= 8'b11111111; // 3829 : 255 - 0xff
      13'hEF6: dout <= 8'b11111111; // 3830 : 255 - 0xff
      13'hEF7: dout <= 8'b11111111; // 3831 : 255 - 0xff
      13'hEF8: dout <= 8'b11111111; // 3832 : 255 - 0xff
      13'hEF9: dout <= 8'b11111111; // 3833 : 255 - 0xff
      13'hEFA: dout <= 8'b11111111; // 3834 : 255 - 0xff
      13'hEFB: dout <= 8'b11111111; // 3835 : 255 - 0xff
      13'hEFC: dout <= 8'b11111111; // 3836 : 255 - 0xff
      13'hEFD: dout <= 8'b11111111; // 3837 : 255 - 0xff
      13'hEFE: dout <= 8'b11111111; // 3838 : 255 - 0xff
      13'hEFF: dout <= 8'b11111111; // 3839 : 255 - 0xff
      13'hF00: dout <= 8'b11111111; // 3840 : 255 - 0xff -- Sprite 0xf0
      13'hF01: dout <= 8'b11111111; // 3841 : 255 - 0xff
      13'hF02: dout <= 8'b11111111; // 3842 : 255 - 0xff
      13'hF03: dout <= 8'b11111111; // 3843 : 255 - 0xff
      13'hF04: dout <= 8'b11111111; // 3844 : 255 - 0xff
      13'hF05: dout <= 8'b11111111; // 3845 : 255 - 0xff
      13'hF06: dout <= 8'b11111111; // 3846 : 255 - 0xff
      13'hF07: dout <= 8'b11111111; // 3847 : 255 - 0xff
      13'hF08: dout <= 8'b11111111; // 3848 : 255 - 0xff
      13'hF09: dout <= 8'b11111111; // 3849 : 255 - 0xff
      13'hF0A: dout <= 8'b11111111; // 3850 : 255 - 0xff
      13'hF0B: dout <= 8'b11111111; // 3851 : 255 - 0xff
      13'hF0C: dout <= 8'b11111111; // 3852 : 255 - 0xff
      13'hF0D: dout <= 8'b11111111; // 3853 : 255 - 0xff
      13'hF0E: dout <= 8'b11111111; // 3854 : 255 - 0xff
      13'hF0F: dout <= 8'b11111111; // 3855 : 255 - 0xff
      13'hF10: dout <= 8'b11111111; // 3856 : 255 - 0xff -- Sprite 0xf1
      13'hF11: dout <= 8'b11111111; // 3857 : 255 - 0xff
      13'hF12: dout <= 8'b11111111; // 3858 : 255 - 0xff
      13'hF13: dout <= 8'b11111111; // 3859 : 255 - 0xff
      13'hF14: dout <= 8'b11111111; // 3860 : 255 - 0xff
      13'hF15: dout <= 8'b11111111; // 3861 : 255 - 0xff
      13'hF16: dout <= 8'b11111111; // 3862 : 255 - 0xff
      13'hF17: dout <= 8'b11111111; // 3863 : 255 - 0xff
      13'hF18: dout <= 8'b11111111; // 3864 : 255 - 0xff
      13'hF19: dout <= 8'b11111111; // 3865 : 255 - 0xff
      13'hF1A: dout <= 8'b11111111; // 3866 : 255 - 0xff
      13'hF1B: dout <= 8'b11111111; // 3867 : 255 - 0xff
      13'hF1C: dout <= 8'b11111111; // 3868 : 255 - 0xff
      13'hF1D: dout <= 8'b11111111; // 3869 : 255 - 0xff
      13'hF1E: dout <= 8'b11111111; // 3870 : 255 - 0xff
      13'hF1F: dout <= 8'b11111111; // 3871 : 255 - 0xff
      13'hF20: dout <= 8'b11111111; // 3872 : 255 - 0xff -- Sprite 0xf2
      13'hF21: dout <= 8'b11111111; // 3873 : 255 - 0xff
      13'hF22: dout <= 8'b11111111; // 3874 : 255 - 0xff
      13'hF23: dout <= 8'b11111111; // 3875 : 255 - 0xff
      13'hF24: dout <= 8'b11111111; // 3876 : 255 - 0xff
      13'hF25: dout <= 8'b11111111; // 3877 : 255 - 0xff
      13'hF26: dout <= 8'b11111111; // 3878 : 255 - 0xff
      13'hF27: dout <= 8'b11111111; // 3879 : 255 - 0xff
      13'hF28: dout <= 8'b11111111; // 3880 : 255 - 0xff
      13'hF29: dout <= 8'b11111111; // 3881 : 255 - 0xff
      13'hF2A: dout <= 8'b11111111; // 3882 : 255 - 0xff
      13'hF2B: dout <= 8'b11111111; // 3883 : 255 - 0xff
      13'hF2C: dout <= 8'b11111111; // 3884 : 255 - 0xff
      13'hF2D: dout <= 8'b11111111; // 3885 : 255 - 0xff
      13'hF2E: dout <= 8'b11111111; // 3886 : 255 - 0xff
      13'hF2F: dout <= 8'b11111111; // 3887 : 255 - 0xff
      13'hF30: dout <= 8'b11111111; // 3888 : 255 - 0xff -- Sprite 0xf3
      13'hF31: dout <= 8'b11111111; // 3889 : 255 - 0xff
      13'hF32: dout <= 8'b11111111; // 3890 : 255 - 0xff
      13'hF33: dout <= 8'b11111111; // 3891 : 255 - 0xff
      13'hF34: dout <= 8'b11111111; // 3892 : 255 - 0xff
      13'hF35: dout <= 8'b11111111; // 3893 : 255 - 0xff
      13'hF36: dout <= 8'b11111111; // 3894 : 255 - 0xff
      13'hF37: dout <= 8'b11111111; // 3895 : 255 - 0xff
      13'hF38: dout <= 8'b11111111; // 3896 : 255 - 0xff
      13'hF39: dout <= 8'b11111111; // 3897 : 255 - 0xff
      13'hF3A: dout <= 8'b11111111; // 3898 : 255 - 0xff
      13'hF3B: dout <= 8'b11111111; // 3899 : 255 - 0xff
      13'hF3C: dout <= 8'b11111111; // 3900 : 255 - 0xff
      13'hF3D: dout <= 8'b11111111; // 3901 : 255 - 0xff
      13'hF3E: dout <= 8'b11111111; // 3902 : 255 - 0xff
      13'hF3F: dout <= 8'b11111111; // 3903 : 255 - 0xff
      13'hF40: dout <= 8'b11111111; // 3904 : 255 - 0xff -- Sprite 0xf4
      13'hF41: dout <= 8'b11111111; // 3905 : 255 - 0xff
      13'hF42: dout <= 8'b11111111; // 3906 : 255 - 0xff
      13'hF43: dout <= 8'b11111111; // 3907 : 255 - 0xff
      13'hF44: dout <= 8'b11111111; // 3908 : 255 - 0xff
      13'hF45: dout <= 8'b11111111; // 3909 : 255 - 0xff
      13'hF46: dout <= 8'b11111111; // 3910 : 255 - 0xff
      13'hF47: dout <= 8'b11111111; // 3911 : 255 - 0xff
      13'hF48: dout <= 8'b11111111; // 3912 : 255 - 0xff
      13'hF49: dout <= 8'b11111111; // 3913 : 255 - 0xff
      13'hF4A: dout <= 8'b11111111; // 3914 : 255 - 0xff
      13'hF4B: dout <= 8'b11111111; // 3915 : 255 - 0xff
      13'hF4C: dout <= 8'b11111111; // 3916 : 255 - 0xff
      13'hF4D: dout <= 8'b11111111; // 3917 : 255 - 0xff
      13'hF4E: dout <= 8'b11111111; // 3918 : 255 - 0xff
      13'hF4F: dout <= 8'b11111111; // 3919 : 255 - 0xff
      13'hF50: dout <= 8'b11111111; // 3920 : 255 - 0xff -- Sprite 0xf5
      13'hF51: dout <= 8'b11111111; // 3921 : 255 - 0xff
      13'hF52: dout <= 8'b11111111; // 3922 : 255 - 0xff
      13'hF53: dout <= 8'b11111111; // 3923 : 255 - 0xff
      13'hF54: dout <= 8'b11111111; // 3924 : 255 - 0xff
      13'hF55: dout <= 8'b11111111; // 3925 : 255 - 0xff
      13'hF56: dout <= 8'b11111111; // 3926 : 255 - 0xff
      13'hF57: dout <= 8'b11111111; // 3927 : 255 - 0xff
      13'hF58: dout <= 8'b11111111; // 3928 : 255 - 0xff
      13'hF59: dout <= 8'b11111111; // 3929 : 255 - 0xff
      13'hF5A: dout <= 8'b11111111; // 3930 : 255 - 0xff
      13'hF5B: dout <= 8'b11111111; // 3931 : 255 - 0xff
      13'hF5C: dout <= 8'b11111111; // 3932 : 255 - 0xff
      13'hF5D: dout <= 8'b11111111; // 3933 : 255 - 0xff
      13'hF5E: dout <= 8'b11111111; // 3934 : 255 - 0xff
      13'hF5F: dout <= 8'b11111111; // 3935 : 255 - 0xff
      13'hF60: dout <= 8'b11111111; // 3936 : 255 - 0xff -- Sprite 0xf6
      13'hF61: dout <= 8'b11111111; // 3937 : 255 - 0xff
      13'hF62: dout <= 8'b11111111; // 3938 : 255 - 0xff
      13'hF63: dout <= 8'b11111111; // 3939 : 255 - 0xff
      13'hF64: dout <= 8'b11111111; // 3940 : 255 - 0xff
      13'hF65: dout <= 8'b11111111; // 3941 : 255 - 0xff
      13'hF66: dout <= 8'b11111111; // 3942 : 255 - 0xff
      13'hF67: dout <= 8'b11111111; // 3943 : 255 - 0xff
      13'hF68: dout <= 8'b11111111; // 3944 : 255 - 0xff
      13'hF69: dout <= 8'b11111111; // 3945 : 255 - 0xff
      13'hF6A: dout <= 8'b11111111; // 3946 : 255 - 0xff
      13'hF6B: dout <= 8'b11111111; // 3947 : 255 - 0xff
      13'hF6C: dout <= 8'b11111111; // 3948 : 255 - 0xff
      13'hF6D: dout <= 8'b11111111; // 3949 : 255 - 0xff
      13'hF6E: dout <= 8'b11111111; // 3950 : 255 - 0xff
      13'hF6F: dout <= 8'b11111111; // 3951 : 255 - 0xff
      13'hF70: dout <= 8'b11111111; // 3952 : 255 - 0xff -- Sprite 0xf7
      13'hF71: dout <= 8'b11111111; // 3953 : 255 - 0xff
      13'hF72: dout <= 8'b11111111; // 3954 : 255 - 0xff
      13'hF73: dout <= 8'b11111111; // 3955 : 255 - 0xff
      13'hF74: dout <= 8'b11111111; // 3956 : 255 - 0xff
      13'hF75: dout <= 8'b11111111; // 3957 : 255 - 0xff
      13'hF76: dout <= 8'b11111111; // 3958 : 255 - 0xff
      13'hF77: dout <= 8'b11111111; // 3959 : 255 - 0xff
      13'hF78: dout <= 8'b11111111; // 3960 : 255 - 0xff
      13'hF79: dout <= 8'b11111111; // 3961 : 255 - 0xff
      13'hF7A: dout <= 8'b11111111; // 3962 : 255 - 0xff
      13'hF7B: dout <= 8'b11111111; // 3963 : 255 - 0xff
      13'hF7C: dout <= 8'b11111111; // 3964 : 255 - 0xff
      13'hF7D: dout <= 8'b11111111; // 3965 : 255 - 0xff
      13'hF7E: dout <= 8'b11111111; // 3966 : 255 - 0xff
      13'hF7F: dout <= 8'b11111111; // 3967 : 255 - 0xff
      13'hF80: dout <= 8'b11111111; // 3968 : 255 - 0xff -- Sprite 0xf8
      13'hF81: dout <= 8'b11111111; // 3969 : 255 - 0xff
      13'hF82: dout <= 8'b11111111; // 3970 : 255 - 0xff
      13'hF83: dout <= 8'b11111111; // 3971 : 255 - 0xff
      13'hF84: dout <= 8'b11111111; // 3972 : 255 - 0xff
      13'hF85: dout <= 8'b11111111; // 3973 : 255 - 0xff
      13'hF86: dout <= 8'b11111111; // 3974 : 255 - 0xff
      13'hF87: dout <= 8'b11111111; // 3975 : 255 - 0xff
      13'hF88: dout <= 8'b11111111; // 3976 : 255 - 0xff
      13'hF89: dout <= 8'b11111111; // 3977 : 255 - 0xff
      13'hF8A: dout <= 8'b11111111; // 3978 : 255 - 0xff
      13'hF8B: dout <= 8'b11111111; // 3979 : 255 - 0xff
      13'hF8C: dout <= 8'b11111111; // 3980 : 255 - 0xff
      13'hF8D: dout <= 8'b11111111; // 3981 : 255 - 0xff
      13'hF8E: dout <= 8'b11111111; // 3982 : 255 - 0xff
      13'hF8F: dout <= 8'b11111111; // 3983 : 255 - 0xff
      13'hF90: dout <= 8'b11111111; // 3984 : 255 - 0xff -- Sprite 0xf9
      13'hF91: dout <= 8'b11111111; // 3985 : 255 - 0xff
      13'hF92: dout <= 8'b11111111; // 3986 : 255 - 0xff
      13'hF93: dout <= 8'b11111111; // 3987 : 255 - 0xff
      13'hF94: dout <= 8'b11111111; // 3988 : 255 - 0xff
      13'hF95: dout <= 8'b11111111; // 3989 : 255 - 0xff
      13'hF96: dout <= 8'b11111111; // 3990 : 255 - 0xff
      13'hF97: dout <= 8'b11111111; // 3991 : 255 - 0xff
      13'hF98: dout <= 8'b11111111; // 3992 : 255 - 0xff
      13'hF99: dout <= 8'b11111111; // 3993 : 255 - 0xff
      13'hF9A: dout <= 8'b11111111; // 3994 : 255 - 0xff
      13'hF9B: dout <= 8'b11111111; // 3995 : 255 - 0xff
      13'hF9C: dout <= 8'b11111111; // 3996 : 255 - 0xff
      13'hF9D: dout <= 8'b11111111; // 3997 : 255 - 0xff
      13'hF9E: dout <= 8'b11111111; // 3998 : 255 - 0xff
      13'hF9F: dout <= 8'b11111111; // 3999 : 255 - 0xff
      13'hFA0: dout <= 8'b11111111; // 4000 : 255 - 0xff -- Sprite 0xfa
      13'hFA1: dout <= 8'b11111111; // 4001 : 255 - 0xff
      13'hFA2: dout <= 8'b11111111; // 4002 : 255 - 0xff
      13'hFA3: dout <= 8'b11111111; // 4003 : 255 - 0xff
      13'hFA4: dout <= 8'b11111111; // 4004 : 255 - 0xff
      13'hFA5: dout <= 8'b11111111; // 4005 : 255 - 0xff
      13'hFA6: dout <= 8'b11111111; // 4006 : 255 - 0xff
      13'hFA7: dout <= 8'b11111111; // 4007 : 255 - 0xff
      13'hFA8: dout <= 8'b11111111; // 4008 : 255 - 0xff
      13'hFA9: dout <= 8'b11111111; // 4009 : 255 - 0xff
      13'hFAA: dout <= 8'b11111111; // 4010 : 255 - 0xff
      13'hFAB: dout <= 8'b11111111; // 4011 : 255 - 0xff
      13'hFAC: dout <= 8'b11111111; // 4012 : 255 - 0xff
      13'hFAD: dout <= 8'b11111111; // 4013 : 255 - 0xff
      13'hFAE: dout <= 8'b11111111; // 4014 : 255 - 0xff
      13'hFAF: dout <= 8'b11111111; // 4015 : 255 - 0xff
      13'hFB0: dout <= 8'b11111111; // 4016 : 255 - 0xff -- Sprite 0xfb
      13'hFB1: dout <= 8'b11111111; // 4017 : 255 - 0xff
      13'hFB2: dout <= 8'b11111111; // 4018 : 255 - 0xff
      13'hFB3: dout <= 8'b11111111; // 4019 : 255 - 0xff
      13'hFB4: dout <= 8'b11111111; // 4020 : 255 - 0xff
      13'hFB5: dout <= 8'b11111111; // 4021 : 255 - 0xff
      13'hFB6: dout <= 8'b11111111; // 4022 : 255 - 0xff
      13'hFB7: dout <= 8'b11111111; // 4023 : 255 - 0xff
      13'hFB8: dout <= 8'b11111111; // 4024 : 255 - 0xff
      13'hFB9: dout <= 8'b11111111; // 4025 : 255 - 0xff
      13'hFBA: dout <= 8'b11111111; // 4026 : 255 - 0xff
      13'hFBB: dout <= 8'b11111111; // 4027 : 255 - 0xff
      13'hFBC: dout <= 8'b11111111; // 4028 : 255 - 0xff
      13'hFBD: dout <= 8'b11111111; // 4029 : 255 - 0xff
      13'hFBE: dout <= 8'b11111111; // 4030 : 255 - 0xff
      13'hFBF: dout <= 8'b11111111; // 4031 : 255 - 0xff
      13'hFC0: dout <= 8'b11111111; // 4032 : 255 - 0xff -- Sprite 0xfc
      13'hFC1: dout <= 8'b11111111; // 4033 : 255 - 0xff
      13'hFC2: dout <= 8'b11111111; // 4034 : 255 - 0xff
      13'hFC3: dout <= 8'b11111111; // 4035 : 255 - 0xff
      13'hFC4: dout <= 8'b11111111; // 4036 : 255 - 0xff
      13'hFC5: dout <= 8'b11111111; // 4037 : 255 - 0xff
      13'hFC6: dout <= 8'b11111111; // 4038 : 255 - 0xff
      13'hFC7: dout <= 8'b11111111; // 4039 : 255 - 0xff
      13'hFC8: dout <= 8'b11111111; // 4040 : 255 - 0xff
      13'hFC9: dout <= 8'b11111111; // 4041 : 255 - 0xff
      13'hFCA: dout <= 8'b11111111; // 4042 : 255 - 0xff
      13'hFCB: dout <= 8'b11111111; // 4043 : 255 - 0xff
      13'hFCC: dout <= 8'b11111111; // 4044 : 255 - 0xff
      13'hFCD: dout <= 8'b11111111; // 4045 : 255 - 0xff
      13'hFCE: dout <= 8'b11111111; // 4046 : 255 - 0xff
      13'hFCF: dout <= 8'b11111111; // 4047 : 255 - 0xff
      13'hFD0: dout <= 8'b11111111; // 4048 : 255 - 0xff -- Sprite 0xfd
      13'hFD1: dout <= 8'b11111111; // 4049 : 255 - 0xff
      13'hFD2: dout <= 8'b11111111; // 4050 : 255 - 0xff
      13'hFD3: dout <= 8'b11111111; // 4051 : 255 - 0xff
      13'hFD4: dout <= 8'b11111111; // 4052 : 255 - 0xff
      13'hFD5: dout <= 8'b11111111; // 4053 : 255 - 0xff
      13'hFD6: dout <= 8'b11111111; // 4054 : 255 - 0xff
      13'hFD7: dout <= 8'b11111111; // 4055 : 255 - 0xff
      13'hFD8: dout <= 8'b11111111; // 4056 : 255 - 0xff
      13'hFD9: dout <= 8'b11111111; // 4057 : 255 - 0xff
      13'hFDA: dout <= 8'b11111111; // 4058 : 255 - 0xff
      13'hFDB: dout <= 8'b11111111; // 4059 : 255 - 0xff
      13'hFDC: dout <= 8'b11111111; // 4060 : 255 - 0xff
      13'hFDD: dout <= 8'b11111111; // 4061 : 255 - 0xff
      13'hFDE: dout <= 8'b11111111; // 4062 : 255 - 0xff
      13'hFDF: dout <= 8'b11111111; // 4063 : 255 - 0xff
      13'hFE0: dout <= 8'b11111111; // 4064 : 255 - 0xff -- Sprite 0xfe
      13'hFE1: dout <= 8'b11111111; // 4065 : 255 - 0xff
      13'hFE2: dout <= 8'b11111111; // 4066 : 255 - 0xff
      13'hFE3: dout <= 8'b11111111; // 4067 : 255 - 0xff
      13'hFE4: dout <= 8'b11111111; // 4068 : 255 - 0xff
      13'hFE5: dout <= 8'b11111111; // 4069 : 255 - 0xff
      13'hFE6: dout <= 8'b11111111; // 4070 : 255 - 0xff
      13'hFE7: dout <= 8'b11111111; // 4071 : 255 - 0xff
      13'hFE8: dout <= 8'b11111111; // 4072 : 255 - 0xff
      13'hFE9: dout <= 8'b11111111; // 4073 : 255 - 0xff
      13'hFEA: dout <= 8'b11111111; // 4074 : 255 - 0xff
      13'hFEB: dout <= 8'b11111111; // 4075 : 255 - 0xff
      13'hFEC: dout <= 8'b11111111; // 4076 : 255 - 0xff
      13'hFED: dout <= 8'b11111111; // 4077 : 255 - 0xff
      13'hFEE: dout <= 8'b11111111; // 4078 : 255 - 0xff
      13'hFEF: dout <= 8'b11111111; // 4079 : 255 - 0xff
      13'hFF0: dout <= 8'b11111111; // 4080 : 255 - 0xff -- Sprite 0xff
      13'hFF1: dout <= 8'b11111111; // 4081 : 255 - 0xff
      13'hFF2: dout <= 8'b11111111; // 4082 : 255 - 0xff
      13'hFF3: dout <= 8'b11111111; // 4083 : 255 - 0xff
      13'hFF4: dout <= 8'b11111111; // 4084 : 255 - 0xff
      13'hFF5: dout <= 8'b11111111; // 4085 : 255 - 0xff
      13'hFF6: dout <= 8'b11111111; // 4086 : 255 - 0xff
      13'hFF7: dout <= 8'b11111111; // 4087 : 255 - 0xff
      13'hFF8: dout <= 8'b11111111; // 4088 : 255 - 0xff
      13'hFF9: dout <= 8'b11111111; // 4089 : 255 - 0xff
      13'hFFA: dout <= 8'b11111111; // 4090 : 255 - 0xff
      13'hFFB: dout <= 8'b11111111; // 4091 : 255 - 0xff
      13'hFFC: dout <= 8'b11111111; // 4092 : 255 - 0xff
      13'hFFD: dout <= 8'b11111111; // 4093 : 255 - 0xff
      13'hFFE: dout <= 8'b11111111; // 4094 : 255 - 0xff
      13'hFFF: dout <= 8'b11111111; // 4095 : 255 - 0xff
          // Pattern Table 1---------
      13'h1000: dout <= 8'b00000000; // 4096 :   0 - 0x0 -- Background 0x0
      13'h1001: dout <= 8'b00000000; // 4097 :   0 - 0x0
      13'h1002: dout <= 8'b00000000; // 4098 :   0 - 0x0
      13'h1003: dout <= 8'b00000000; // 4099 :   0 - 0x0
      13'h1004: dout <= 8'b00000000; // 4100 :   0 - 0x0
      13'h1005: dout <= 8'b00000000; // 4101 :   0 - 0x0
      13'h1006: dout <= 8'b00000000; // 4102 :   0 - 0x0
      13'h1007: dout <= 8'b00000000; // 4103 :   0 - 0x0
      13'h1008: dout <= 8'b00000000; // 4104 :   0 - 0x0
      13'h1009: dout <= 8'b00000000; // 4105 :   0 - 0x0
      13'h100A: dout <= 8'b00000000; // 4106 :   0 - 0x0
      13'h100B: dout <= 8'b00000000; // 4107 :   0 - 0x0
      13'h100C: dout <= 8'b00000000; // 4108 :   0 - 0x0
      13'h100D: dout <= 8'b00000000; // 4109 :   0 - 0x0
      13'h100E: dout <= 8'b00000000; // 4110 :   0 - 0x0
      13'h100F: dout <= 8'b00000000; // 4111 :   0 - 0x0
      13'h1010: dout <= 8'b00000000; // 4112 :   0 - 0x0 -- Background 0x1
      13'h1011: dout <= 8'b00111000; // 4113 :  56 - 0x38
      13'h1012: dout <= 8'b01111100; // 4114 : 124 - 0x7c
      13'h1013: dout <= 8'b11111110; // 4115 : 254 - 0xfe
      13'h1014: dout <= 8'b11111110; // 4116 : 254 - 0xfe
      13'h1015: dout <= 8'b11111110; // 4117 : 254 - 0xfe
      13'h1016: dout <= 8'b01111100; // 4118 : 124 - 0x7c
      13'h1017: dout <= 8'b00111000; // 4119 :  56 - 0x38
      13'h1018: dout <= 8'b00000000; // 4120 :   0 - 0x0
      13'h1019: dout <= 8'b00111000; // 4121 :  56 - 0x38
      13'h101A: dout <= 8'b01111100; // 4122 : 124 - 0x7c
      13'h101B: dout <= 8'b11111110; // 4123 : 254 - 0xfe
      13'h101C: dout <= 8'b11111110; // 4124 : 254 - 0xfe
      13'h101D: dout <= 8'b11111110; // 4125 : 254 - 0xfe
      13'h101E: dout <= 8'b01111100; // 4126 : 124 - 0x7c
      13'h101F: dout <= 8'b00111000; // 4127 :  56 - 0x38
      13'h1020: dout <= 8'b00000000; // 4128 :   0 - 0x0 -- Background 0x2
      13'h1021: dout <= 8'b00000000; // 4129 :   0 - 0x0
      13'h1022: dout <= 8'b00000000; // 4130 :   0 - 0x0
      13'h1023: dout <= 8'b00000000; // 4131 :   0 - 0x0
      13'h1024: dout <= 8'b00000000; // 4132 :   0 - 0x0
      13'h1025: dout <= 8'b00000000; // 4133 :   0 - 0x0
      13'h1026: dout <= 8'b00000000; // 4134 :   0 - 0x0
      13'h1027: dout <= 8'b00000000; // 4135 :   0 - 0x0
      13'h1028: dout <= 8'b00000000; // 4136 :   0 - 0x0
      13'h1029: dout <= 8'b00000000; // 4137 :   0 - 0x0
      13'h102A: dout <= 8'b00000000; // 4138 :   0 - 0x0
      13'h102B: dout <= 8'b00000000; // 4139 :   0 - 0x0
      13'h102C: dout <= 8'b00000000; // 4140 :   0 - 0x0
      13'h102D: dout <= 8'b00000000; // 4141 :   0 - 0x0
      13'h102E: dout <= 8'b00000000; // 4142 :   0 - 0x0
      13'h102F: dout <= 8'b00000000; // 4143 :   0 - 0x0
      13'h1030: dout <= 8'b00000000; // 4144 :   0 - 0x0 -- Background 0x3
      13'h1031: dout <= 8'b00000000; // 4145 :   0 - 0x0
      13'h1032: dout <= 8'b00000000; // 4146 :   0 - 0x0
      13'h1033: dout <= 8'b00011000; // 4147 :  24 - 0x18
      13'h1034: dout <= 8'b00011000; // 4148 :  24 - 0x18
      13'h1035: dout <= 8'b00000000; // 4149 :   0 - 0x0
      13'h1036: dout <= 8'b00000000; // 4150 :   0 - 0x0
      13'h1037: dout <= 8'b00000000; // 4151 :   0 - 0x0
      13'h1038: dout <= 8'b00000000; // 4152 :   0 - 0x0
      13'h1039: dout <= 8'b00000000; // 4153 :   0 - 0x0
      13'h103A: dout <= 8'b00000000; // 4154 :   0 - 0x0
      13'h103B: dout <= 8'b00011000; // 4155 :  24 - 0x18
      13'h103C: dout <= 8'b00011000; // 4156 :  24 - 0x18
      13'h103D: dout <= 8'b00000000; // 4157 :   0 - 0x0
      13'h103E: dout <= 8'b00000000; // 4158 :   0 - 0x0
      13'h103F: dout <= 8'b00000000; // 4159 :   0 - 0x0
      13'h1040: dout <= 8'b00000000; // 4160 :   0 - 0x0 -- Background 0x4
      13'h1041: dout <= 8'b00000000; // 4161 :   0 - 0x0
      13'h1042: dout <= 8'b00000000; // 4162 :   0 - 0x0
      13'h1043: dout <= 8'b00000000; // 4163 :   0 - 0x0
      13'h1044: dout <= 8'b00000000; // 4164 :   0 - 0x0
      13'h1045: dout <= 8'b00000000; // 4165 :   0 - 0x0
      13'h1046: dout <= 8'b00000000; // 4166 :   0 - 0x0
      13'h1047: dout <= 8'b00000000; // 4167 :   0 - 0x0
      13'h1048: dout <= 8'b11111111; // 4168 : 255 - 0xff
      13'h1049: dout <= 8'b11111111; // 4169 : 255 - 0xff
      13'h104A: dout <= 8'b11111111; // 4170 : 255 - 0xff
      13'h104B: dout <= 8'b11111111; // 4171 : 255 - 0xff
      13'h104C: dout <= 8'b11111111; // 4172 : 255 - 0xff
      13'h104D: dout <= 8'b11111111; // 4173 : 255 - 0xff
      13'h104E: dout <= 8'b11111111; // 4174 : 255 - 0xff
      13'h104F: dout <= 8'b11111111; // 4175 : 255 - 0xff
      13'h1050: dout <= 8'b00000000; // 4176 :   0 - 0x0 -- Background 0x5
      13'h1051: dout <= 8'b00000000; // 4177 :   0 - 0x0
      13'h1052: dout <= 8'b00000000; // 4178 :   0 - 0x0
      13'h1053: dout <= 8'b00000000; // 4179 :   0 - 0x0
      13'h1054: dout <= 8'b00000000; // 4180 :   0 - 0x0
      13'h1055: dout <= 8'b00000000; // 4181 :   0 - 0x0
      13'h1056: dout <= 8'b00000000; // 4182 :   0 - 0x0
      13'h1057: dout <= 8'b00000000; // 4183 :   0 - 0x0
      13'h1058: dout <= 8'b00001111; // 4184 :  15 - 0xf
      13'h1059: dout <= 8'b00001111; // 4185 :  15 - 0xf
      13'h105A: dout <= 8'b00001111; // 4186 :  15 - 0xf
      13'h105B: dout <= 8'b00001111; // 4187 :  15 - 0xf
      13'h105C: dout <= 8'b00001111; // 4188 :  15 - 0xf
      13'h105D: dout <= 8'b00001111; // 4189 :  15 - 0xf
      13'h105E: dout <= 8'b00001111; // 4190 :  15 - 0xf
      13'h105F: dout <= 8'b00001111; // 4191 :  15 - 0xf
      13'h1060: dout <= 8'b00000000; // 4192 :   0 - 0x0 -- Background 0x6
      13'h1061: dout <= 8'b00000000; // 4193 :   0 - 0x0
      13'h1062: dout <= 8'b00000000; // 4194 :   0 - 0x0
      13'h1063: dout <= 8'b00000000; // 4195 :   0 - 0x0
      13'h1064: dout <= 8'b00000000; // 4196 :   0 - 0x0
      13'h1065: dout <= 8'b00000000; // 4197 :   0 - 0x0
      13'h1066: dout <= 8'b00000000; // 4198 :   0 - 0x0
      13'h1067: dout <= 8'b00000000; // 4199 :   0 - 0x0
      13'h1068: dout <= 8'b11110000; // 4200 : 240 - 0xf0
      13'h1069: dout <= 8'b11110000; // 4201 : 240 - 0xf0
      13'h106A: dout <= 8'b11110000; // 4202 : 240 - 0xf0
      13'h106B: dout <= 8'b11110000; // 4203 : 240 - 0xf0
      13'h106C: dout <= 8'b11110000; // 4204 : 240 - 0xf0
      13'h106D: dout <= 8'b11110000; // 4205 : 240 - 0xf0
      13'h106E: dout <= 8'b11110000; // 4206 : 240 - 0xf0
      13'h106F: dout <= 8'b11110000; // 4207 : 240 - 0xf0
      13'h1070: dout <= 8'b00000000; // 4208 :   0 - 0x0 -- Background 0x7
      13'h1071: dout <= 8'b00000000; // 4209 :   0 - 0x0
      13'h1072: dout <= 8'b00000000; // 4210 :   0 - 0x0
      13'h1073: dout <= 8'b00000000; // 4211 :   0 - 0x0
      13'h1074: dout <= 8'b00000000; // 4212 :   0 - 0x0
      13'h1075: dout <= 8'b00000000; // 4213 :   0 - 0x0
      13'h1076: dout <= 8'b00000000; // 4214 :   0 - 0x0
      13'h1077: dout <= 8'b00000000; // 4215 :   0 - 0x0
      13'h1078: dout <= 8'b00000000; // 4216 :   0 - 0x0
      13'h1079: dout <= 8'b00000000; // 4217 :   0 - 0x0
      13'h107A: dout <= 8'b00000000; // 4218 :   0 - 0x0
      13'h107B: dout <= 8'b00000000; // 4219 :   0 - 0x0
      13'h107C: dout <= 8'b00000000; // 4220 :   0 - 0x0
      13'h107D: dout <= 8'b00000000; // 4221 :   0 - 0x0
      13'h107E: dout <= 8'b00000000; // 4222 :   0 - 0x0
      13'h107F: dout <= 8'b00000000; // 4223 :   0 - 0x0
      13'h1080: dout <= 8'b00000000; // 4224 :   0 - 0x0 -- Background 0x8
      13'h1081: dout <= 8'b00000000; // 4225 :   0 - 0x0
      13'h1082: dout <= 8'b00000000; // 4226 :   0 - 0x0
      13'h1083: dout <= 8'b00000000; // 4227 :   0 - 0x0
      13'h1084: dout <= 8'b00000000; // 4228 :   0 - 0x0
      13'h1085: dout <= 8'b00000000; // 4229 :   0 - 0x0
      13'h1086: dout <= 8'b00000000; // 4230 :   0 - 0x0
      13'h1087: dout <= 8'b00000000; // 4231 :   0 - 0x0
      13'h1088: dout <= 8'b00000000; // 4232 :   0 - 0x0
      13'h1089: dout <= 8'b00000000; // 4233 :   0 - 0x0
      13'h108A: dout <= 8'b00000000; // 4234 :   0 - 0x0
      13'h108B: dout <= 8'b00000000; // 4235 :   0 - 0x0
      13'h108C: dout <= 8'b00000000; // 4236 :   0 - 0x0
      13'h108D: dout <= 8'b00000000; // 4237 :   0 - 0x0
      13'h108E: dout <= 8'b00000000; // 4238 :   0 - 0x0
      13'h108F: dout <= 8'b00000000; // 4239 :   0 - 0x0
      13'h1090: dout <= 8'b00000000; // 4240 :   0 - 0x0 -- Background 0x9
      13'h1091: dout <= 8'b00000000; // 4241 :   0 - 0x0
      13'h1092: dout <= 8'b00000000; // 4242 :   0 - 0x0
      13'h1093: dout <= 8'b00011000; // 4243 :  24 - 0x18
      13'h1094: dout <= 8'b00011000; // 4244 :  24 - 0x18
      13'h1095: dout <= 8'b00000000; // 4245 :   0 - 0x0
      13'h1096: dout <= 8'b00000000; // 4246 :   0 - 0x0
      13'h1097: dout <= 8'b00000000; // 4247 :   0 - 0x0
      13'h1098: dout <= 8'b00000000; // 4248 :   0 - 0x0
      13'h1099: dout <= 8'b00000000; // 4249 :   0 - 0x0
      13'h109A: dout <= 8'b00000000; // 4250 :   0 - 0x0
      13'h109B: dout <= 8'b00011000; // 4251 :  24 - 0x18
      13'h109C: dout <= 8'b00011000; // 4252 :  24 - 0x18
      13'h109D: dout <= 8'b00000000; // 4253 :   0 - 0x0
      13'h109E: dout <= 8'b00000000; // 4254 :   0 - 0x0
      13'h109F: dout <= 8'b00000000; // 4255 :   0 - 0x0
      13'h10A0: dout <= 8'b00000000; // 4256 :   0 - 0x0 -- Background 0xa
      13'h10A1: dout <= 8'b00000000; // 4257 :   0 - 0x0
      13'h10A2: dout <= 8'b00000000; // 4258 :   0 - 0x0
      13'h10A3: dout <= 8'b00000000; // 4259 :   0 - 0x0
      13'h10A4: dout <= 8'b00000000; // 4260 :   0 - 0x0
      13'h10A5: dout <= 8'b00000000; // 4261 :   0 - 0x0
      13'h10A6: dout <= 8'b00000000; // 4262 :   0 - 0x0
      13'h10A7: dout <= 8'b00000000; // 4263 :   0 - 0x0
      13'h10A8: dout <= 8'b00000000; // 4264 :   0 - 0x0
      13'h10A9: dout <= 8'b00000000; // 4265 :   0 - 0x0
      13'h10AA: dout <= 8'b00000000; // 4266 :   0 - 0x0
      13'h10AB: dout <= 8'b00000000; // 4267 :   0 - 0x0
      13'h10AC: dout <= 8'b00000000; // 4268 :   0 - 0x0
      13'h10AD: dout <= 8'b00000000; // 4269 :   0 - 0x0
      13'h10AE: dout <= 8'b00000000; // 4270 :   0 - 0x0
      13'h10AF: dout <= 8'b00000000; // 4271 :   0 - 0x0
      13'h10B0: dout <= 8'b00000000; // 4272 :   0 - 0x0 -- Background 0xb
      13'h10B1: dout <= 8'b00000000; // 4273 :   0 - 0x0
      13'h10B2: dout <= 8'b00000000; // 4274 :   0 - 0x0
      13'h10B3: dout <= 8'b00000000; // 4275 :   0 - 0x0
      13'h10B4: dout <= 8'b00000000; // 4276 :   0 - 0x0
      13'h10B5: dout <= 8'b00000000; // 4277 :   0 - 0x0
      13'h10B6: dout <= 8'b00000000; // 4278 :   0 - 0x0
      13'h10B7: dout <= 8'b00000000; // 4279 :   0 - 0x0
      13'h10B8: dout <= 8'b00000000; // 4280 :   0 - 0x0
      13'h10B9: dout <= 8'b00000000; // 4281 :   0 - 0x0
      13'h10BA: dout <= 8'b00000000; // 4282 :   0 - 0x0
      13'h10BB: dout <= 8'b00000000; // 4283 :   0 - 0x0
      13'h10BC: dout <= 8'b00000000; // 4284 :   0 - 0x0
      13'h10BD: dout <= 8'b00000000; // 4285 :   0 - 0x0
      13'h10BE: dout <= 8'b00000000; // 4286 :   0 - 0x0
      13'h10BF: dout <= 8'b00000000; // 4287 :   0 - 0x0
      13'h10C0: dout <= 8'b00000000; // 4288 :   0 - 0x0 -- Background 0xc
      13'h10C1: dout <= 8'b00000000; // 4289 :   0 - 0x0
      13'h10C2: dout <= 8'b00000000; // 4290 :   0 - 0x0
      13'h10C3: dout <= 8'b00000000; // 4291 :   0 - 0x0
      13'h10C4: dout <= 8'b00000000; // 4292 :   0 - 0x0
      13'h10C5: dout <= 8'b00000000; // 4293 :   0 - 0x0
      13'h10C6: dout <= 8'b00000000; // 4294 :   0 - 0x0
      13'h10C7: dout <= 8'b00000000; // 4295 :   0 - 0x0
      13'h10C8: dout <= 8'b00000000; // 4296 :   0 - 0x0
      13'h10C9: dout <= 8'b00000000; // 4297 :   0 - 0x0
      13'h10CA: dout <= 8'b00000000; // 4298 :   0 - 0x0
      13'h10CB: dout <= 8'b00000000; // 4299 :   0 - 0x0
      13'h10CC: dout <= 8'b00000000; // 4300 :   0 - 0x0
      13'h10CD: dout <= 8'b00000000; // 4301 :   0 - 0x0
      13'h10CE: dout <= 8'b00000000; // 4302 :   0 - 0x0
      13'h10CF: dout <= 8'b00000000; // 4303 :   0 - 0x0
      13'h10D0: dout <= 8'b00000000; // 4304 :   0 - 0x0 -- Background 0xd
      13'h10D1: dout <= 8'b00000000; // 4305 :   0 - 0x0
      13'h10D2: dout <= 8'b00000000; // 4306 :   0 - 0x0
      13'h10D3: dout <= 8'b00000000; // 4307 :   0 - 0x0
      13'h10D4: dout <= 8'b00000000; // 4308 :   0 - 0x0
      13'h10D5: dout <= 8'b00000000; // 4309 :   0 - 0x0
      13'h10D6: dout <= 8'b00000000; // 4310 :   0 - 0x0
      13'h10D7: dout <= 8'b00000000; // 4311 :   0 - 0x0
      13'h10D8: dout <= 8'b00000000; // 4312 :   0 - 0x0
      13'h10D9: dout <= 8'b00000000; // 4313 :   0 - 0x0
      13'h10DA: dout <= 8'b00000000; // 4314 :   0 - 0x0
      13'h10DB: dout <= 8'b00000000; // 4315 :   0 - 0x0
      13'h10DC: dout <= 8'b00000000; // 4316 :   0 - 0x0
      13'h10DD: dout <= 8'b00000000; // 4317 :   0 - 0x0
      13'h10DE: dout <= 8'b00000000; // 4318 :   0 - 0x0
      13'h10DF: dout <= 8'b00000000; // 4319 :   0 - 0x0
      13'h10E0: dout <= 8'b00000000; // 4320 :   0 - 0x0 -- Background 0xe
      13'h10E1: dout <= 8'b00000000; // 4321 :   0 - 0x0
      13'h10E2: dout <= 8'b00000000; // 4322 :   0 - 0x0
      13'h10E3: dout <= 8'b00000000; // 4323 :   0 - 0x0
      13'h10E4: dout <= 8'b00000000; // 4324 :   0 - 0x0
      13'h10E5: dout <= 8'b00000000; // 4325 :   0 - 0x0
      13'h10E6: dout <= 8'b00000000; // 4326 :   0 - 0x0
      13'h10E7: dout <= 8'b00000000; // 4327 :   0 - 0x0
      13'h10E8: dout <= 8'b00000000; // 4328 :   0 - 0x0
      13'h10E9: dout <= 8'b00000000; // 4329 :   0 - 0x0
      13'h10EA: dout <= 8'b00000000; // 4330 :   0 - 0x0
      13'h10EB: dout <= 8'b00000000; // 4331 :   0 - 0x0
      13'h10EC: dout <= 8'b00000000; // 4332 :   0 - 0x0
      13'h10ED: dout <= 8'b00000000; // 4333 :   0 - 0x0
      13'h10EE: dout <= 8'b00000000; // 4334 :   0 - 0x0
      13'h10EF: dout <= 8'b00000000; // 4335 :   0 - 0x0
      13'h10F0: dout <= 8'b00000000; // 4336 :   0 - 0x0 -- Background 0xf
      13'h10F1: dout <= 8'b00000000; // 4337 :   0 - 0x0
      13'h10F2: dout <= 8'b00000000; // 4338 :   0 - 0x0
      13'h10F3: dout <= 8'b00000000; // 4339 :   0 - 0x0
      13'h10F4: dout <= 8'b00000000; // 4340 :   0 - 0x0
      13'h10F5: dout <= 8'b00000000; // 4341 :   0 - 0x0
      13'h10F6: dout <= 8'b00000000; // 4342 :   0 - 0x0
      13'h10F7: dout <= 8'b00000000; // 4343 :   0 - 0x0
      13'h10F8: dout <= 8'b00000000; // 4344 :   0 - 0x0
      13'h10F9: dout <= 8'b00000000; // 4345 :   0 - 0x0
      13'h10FA: dout <= 8'b00000000; // 4346 :   0 - 0x0
      13'h10FB: dout <= 8'b00000000; // 4347 :   0 - 0x0
      13'h10FC: dout <= 8'b00000000; // 4348 :   0 - 0x0
      13'h10FD: dout <= 8'b00000000; // 4349 :   0 - 0x0
      13'h10FE: dout <= 8'b00000000; // 4350 :   0 - 0x0
      13'h10FF: dout <= 8'b00000000; // 4351 :   0 - 0x0
      13'h1100: dout <= 8'b00000000; // 4352 :   0 - 0x0 -- Background 0x10
      13'h1101: dout <= 8'b00000000; // 4353 :   0 - 0x0
      13'h1102: dout <= 8'b11111111; // 4354 : 255 - 0xff
      13'h1103: dout <= 8'b00000000; // 4355 :   0 - 0x0
      13'h1104: dout <= 8'b00000000; // 4356 :   0 - 0x0
      13'h1105: dout <= 8'b11111111; // 4357 : 255 - 0xff
      13'h1106: dout <= 8'b00000000; // 4358 :   0 - 0x0
      13'h1107: dout <= 8'b00000000; // 4359 :   0 - 0x0
      13'h1108: dout <= 8'b00000000; // 4360 :   0 - 0x0
      13'h1109: dout <= 8'b00000000; // 4361 :   0 - 0x0
      13'h110A: dout <= 8'b00000000; // 4362 :   0 - 0x0
      13'h110B: dout <= 8'b00000000; // 4363 :   0 - 0x0
      13'h110C: dout <= 8'b00000000; // 4364 :   0 - 0x0
      13'h110D: dout <= 8'b00000000; // 4365 :   0 - 0x0
      13'h110E: dout <= 8'b00000000; // 4366 :   0 - 0x0
      13'h110F: dout <= 8'b00000000; // 4367 :   0 - 0x0
      13'h1110: dout <= 8'b00100100; // 4368 :  36 - 0x24 -- Background 0x11
      13'h1111: dout <= 8'b00100100; // 4369 :  36 - 0x24
      13'h1112: dout <= 8'b00100100; // 4370 :  36 - 0x24
      13'h1113: dout <= 8'b00100100; // 4371 :  36 - 0x24
      13'h1114: dout <= 8'b00100100; // 4372 :  36 - 0x24
      13'h1115: dout <= 8'b00100100; // 4373 :  36 - 0x24
      13'h1116: dout <= 8'b00100100; // 4374 :  36 - 0x24
      13'h1117: dout <= 8'b00100100; // 4375 :  36 - 0x24
      13'h1118: dout <= 8'b00000000; // 4376 :   0 - 0x0
      13'h1119: dout <= 8'b00000000; // 4377 :   0 - 0x0
      13'h111A: dout <= 8'b00000000; // 4378 :   0 - 0x0
      13'h111B: dout <= 8'b00000000; // 4379 :   0 - 0x0
      13'h111C: dout <= 8'b00000000; // 4380 :   0 - 0x0
      13'h111D: dout <= 8'b00000000; // 4381 :   0 - 0x0
      13'h111E: dout <= 8'b00000000; // 4382 :   0 - 0x0
      13'h111F: dout <= 8'b00000000; // 4383 :   0 - 0x0
      13'h1120: dout <= 8'b00100100; // 4384 :  36 - 0x24 -- Background 0x12
      13'h1121: dout <= 8'b00100100; // 4385 :  36 - 0x24
      13'h1122: dout <= 8'b11000011; // 4386 : 195 - 0xc3
      13'h1123: dout <= 8'b00000000; // 4387 :   0 - 0x0
      13'h1124: dout <= 8'b00000000; // 4388 :   0 - 0x0
      13'h1125: dout <= 8'b11111111; // 4389 : 255 - 0xff
      13'h1126: dout <= 8'b00000000; // 4390 :   0 - 0x0
      13'h1127: dout <= 8'b00000000; // 4391 :   0 - 0x0
      13'h1128: dout <= 8'b00000000; // 4392 :   0 - 0x0
      13'h1129: dout <= 8'b00000000; // 4393 :   0 - 0x0
      13'h112A: dout <= 8'b00000000; // 4394 :   0 - 0x0
      13'h112B: dout <= 8'b00000000; // 4395 :   0 - 0x0
      13'h112C: dout <= 8'b00000000; // 4396 :   0 - 0x0
      13'h112D: dout <= 8'b00000000; // 4397 :   0 - 0x0
      13'h112E: dout <= 8'b00000000; // 4398 :   0 - 0x0
      13'h112F: dout <= 8'b00000000; // 4399 :   0 - 0x0
      13'h1130: dout <= 8'b00000000; // 4400 :   0 - 0x0 -- Background 0x13
      13'h1131: dout <= 8'b00000000; // 4401 :   0 - 0x0
      13'h1132: dout <= 8'b11111111; // 4402 : 255 - 0xff
      13'h1133: dout <= 8'b00000000; // 4403 :   0 - 0x0
      13'h1134: dout <= 8'b00000000; // 4404 :   0 - 0x0
      13'h1135: dout <= 8'b11000011; // 4405 : 195 - 0xc3
      13'h1136: dout <= 8'b00100100; // 4406 :  36 - 0x24
      13'h1137: dout <= 8'b00100100; // 4407 :  36 - 0x24
      13'h1138: dout <= 8'b00000000; // 4408 :   0 - 0x0
      13'h1139: dout <= 8'b00000000; // 4409 :   0 - 0x0
      13'h113A: dout <= 8'b00000000; // 4410 :   0 - 0x0
      13'h113B: dout <= 8'b00000000; // 4411 :   0 - 0x0
      13'h113C: dout <= 8'b00000000; // 4412 :   0 - 0x0
      13'h113D: dout <= 8'b00000000; // 4413 :   0 - 0x0
      13'h113E: dout <= 8'b00000000; // 4414 :   0 - 0x0
      13'h113F: dout <= 8'b00000000; // 4415 :   0 - 0x0
      13'h1140: dout <= 8'b00100100; // 4416 :  36 - 0x24 -- Background 0x14
      13'h1141: dout <= 8'b00100100; // 4417 :  36 - 0x24
      13'h1142: dout <= 8'b11000100; // 4418 : 196 - 0xc4
      13'h1143: dout <= 8'b00000100; // 4419 :   4 - 0x4
      13'h1144: dout <= 8'b00000100; // 4420 :   4 - 0x4
      13'h1145: dout <= 8'b11000100; // 4421 : 196 - 0xc4
      13'h1146: dout <= 8'b00100100; // 4422 :  36 - 0x24
      13'h1147: dout <= 8'b00100100; // 4423 :  36 - 0x24
      13'h1148: dout <= 8'b00000000; // 4424 :   0 - 0x0
      13'h1149: dout <= 8'b00000000; // 4425 :   0 - 0x0
      13'h114A: dout <= 8'b00000000; // 4426 :   0 - 0x0
      13'h114B: dout <= 8'b00000000; // 4427 :   0 - 0x0
      13'h114C: dout <= 8'b00000000; // 4428 :   0 - 0x0
      13'h114D: dout <= 8'b00000000; // 4429 :   0 - 0x0
      13'h114E: dout <= 8'b00000000; // 4430 :   0 - 0x0
      13'h114F: dout <= 8'b00000000; // 4431 :   0 - 0x0
      13'h1150: dout <= 8'b00100100; // 4432 :  36 - 0x24 -- Background 0x15
      13'h1151: dout <= 8'b00100100; // 4433 :  36 - 0x24
      13'h1152: dout <= 8'b00100011; // 4434 :  35 - 0x23
      13'h1153: dout <= 8'b00100000; // 4435 :  32 - 0x20
      13'h1154: dout <= 8'b00100000; // 4436 :  32 - 0x20
      13'h1155: dout <= 8'b00100011; // 4437 :  35 - 0x23
      13'h1156: dout <= 8'b00100100; // 4438 :  36 - 0x24
      13'h1157: dout <= 8'b00100100; // 4439 :  36 - 0x24
      13'h1158: dout <= 8'b00000000; // 4440 :   0 - 0x0
      13'h1159: dout <= 8'b00000000; // 4441 :   0 - 0x0
      13'h115A: dout <= 8'b00000000; // 4442 :   0 - 0x0
      13'h115B: dout <= 8'b00000000; // 4443 :   0 - 0x0
      13'h115C: dout <= 8'b00000000; // 4444 :   0 - 0x0
      13'h115D: dout <= 8'b00000000; // 4445 :   0 - 0x0
      13'h115E: dout <= 8'b00000000; // 4446 :   0 - 0x0
      13'h115F: dout <= 8'b00000000; // 4447 :   0 - 0x0
      13'h1160: dout <= 8'b00000000; // 4448 :   0 - 0x0 -- Background 0x16
      13'h1161: dout <= 8'b00000000; // 4449 :   0 - 0x0
      13'h1162: dout <= 8'b00001111; // 4450 :  15 - 0xf
      13'h1163: dout <= 8'b00010000; // 4451 :  16 - 0x10
      13'h1164: dout <= 8'b11110000; // 4452 : 240 - 0xf0
      13'h1165: dout <= 8'b00001111; // 4453 :  15 - 0xf
      13'h1166: dout <= 8'b00000000; // 4454 :   0 - 0x0
      13'h1167: dout <= 8'b00000000; // 4455 :   0 - 0x0
      13'h1168: dout <= 8'b00000000; // 4456 :   0 - 0x0
      13'h1169: dout <= 8'b00000000; // 4457 :   0 - 0x0
      13'h116A: dout <= 8'b00000000; // 4458 :   0 - 0x0
      13'h116B: dout <= 8'b00000000; // 4459 :   0 - 0x0
      13'h116C: dout <= 8'b00000000; // 4460 :   0 - 0x0
      13'h116D: dout <= 8'b00000000; // 4461 :   0 - 0x0
      13'h116E: dout <= 8'b00000000; // 4462 :   0 - 0x0
      13'h116F: dout <= 8'b00000000; // 4463 :   0 - 0x0
      13'h1170: dout <= 8'b00000000; // 4464 :   0 - 0x0 -- Background 0x17
      13'h1171: dout <= 8'b00000000; // 4465 :   0 - 0x0
      13'h1172: dout <= 8'b11110000; // 4466 : 240 - 0xf0
      13'h1173: dout <= 8'b00001000; // 4467 :   8 - 0x8
      13'h1174: dout <= 8'b00001111; // 4468 :  15 - 0xf
      13'h1175: dout <= 8'b11110000; // 4469 : 240 - 0xf0
      13'h1176: dout <= 8'b00000000; // 4470 :   0 - 0x0
      13'h1177: dout <= 8'b00000000; // 4471 :   0 - 0x0
      13'h1178: dout <= 8'b00000000; // 4472 :   0 - 0x0
      13'h1179: dout <= 8'b00000000; // 4473 :   0 - 0x0
      13'h117A: dout <= 8'b00000000; // 4474 :   0 - 0x0
      13'h117B: dout <= 8'b00000000; // 4475 :   0 - 0x0
      13'h117C: dout <= 8'b00000000; // 4476 :   0 - 0x0
      13'h117D: dout <= 8'b00000000; // 4477 :   0 - 0x0
      13'h117E: dout <= 8'b00000000; // 4478 :   0 - 0x0
      13'h117F: dout <= 8'b00000000; // 4479 :   0 - 0x0
      13'h1180: dout <= 8'b00000000; // 4480 :   0 - 0x0 -- Background 0x18
      13'h1181: dout <= 8'b00000000; // 4481 :   0 - 0x0
      13'h1182: dout <= 8'b11110000; // 4482 : 240 - 0xf0
      13'h1183: dout <= 8'b00001000; // 4483 :   8 - 0x8
      13'h1184: dout <= 8'b00001000; // 4484 :   8 - 0x8
      13'h1185: dout <= 8'b11110000; // 4485 : 240 - 0xf0
      13'h1186: dout <= 8'b00000000; // 4486 :   0 - 0x0
      13'h1187: dout <= 8'b00000000; // 4487 :   0 - 0x0
      13'h1188: dout <= 8'b00000000; // 4488 :   0 - 0x0
      13'h1189: dout <= 8'b00000000; // 4489 :   0 - 0x0
      13'h118A: dout <= 8'b00000000; // 4490 :   0 - 0x0
      13'h118B: dout <= 8'b00000000; // 4491 :   0 - 0x0
      13'h118C: dout <= 8'b00000000; // 4492 :   0 - 0x0
      13'h118D: dout <= 8'b00000000; // 4493 :   0 - 0x0
      13'h118E: dout <= 8'b00000000; // 4494 :   0 - 0x0
      13'h118F: dout <= 8'b00000000; // 4495 :   0 - 0x0
      13'h1190: dout <= 8'b00000000; // 4496 :   0 - 0x0 -- Background 0x19
      13'h1191: dout <= 8'b00000000; // 4497 :   0 - 0x0
      13'h1192: dout <= 8'b00001111; // 4498 :  15 - 0xf
      13'h1193: dout <= 8'b00010000; // 4499 :  16 - 0x10
      13'h1194: dout <= 8'b00010000; // 4500 :  16 - 0x10
      13'h1195: dout <= 8'b00001111; // 4501 :  15 - 0xf
      13'h1196: dout <= 8'b00000000; // 4502 :   0 - 0x0
      13'h1197: dout <= 8'b00000000; // 4503 :   0 - 0x0
      13'h1198: dout <= 8'b00000000; // 4504 :   0 - 0x0
      13'h1199: dout <= 8'b00000000; // 4505 :   0 - 0x0
      13'h119A: dout <= 8'b00000000; // 4506 :   0 - 0x0
      13'h119B: dout <= 8'b00000000; // 4507 :   0 - 0x0
      13'h119C: dout <= 8'b00000000; // 4508 :   0 - 0x0
      13'h119D: dout <= 8'b00000000; // 4509 :   0 - 0x0
      13'h119E: dout <= 8'b00000000; // 4510 :   0 - 0x0
      13'h119F: dout <= 8'b00000000; // 4511 :   0 - 0x0
      13'h11A0: dout <= 8'b00100100; // 4512 :  36 - 0x24 -- Background 0x1a
      13'h11A1: dout <= 8'b00100100; // 4513 :  36 - 0x24
      13'h11A2: dout <= 8'b00100100; // 4514 :  36 - 0x24
      13'h11A3: dout <= 8'b00100100; // 4515 :  36 - 0x24
      13'h11A4: dout <= 8'b00011000; // 4516 :  24 - 0x18
      13'h11A5: dout <= 8'b00000000; // 4517 :   0 - 0x0
      13'h11A6: dout <= 8'b00000000; // 4518 :   0 - 0x0
      13'h11A7: dout <= 8'b00000000; // 4519 :   0 - 0x0
      13'h11A8: dout <= 8'b00000000; // 4520 :   0 - 0x0
      13'h11A9: dout <= 8'b00000000; // 4521 :   0 - 0x0
      13'h11AA: dout <= 8'b00000000; // 4522 :   0 - 0x0
      13'h11AB: dout <= 8'b00000000; // 4523 :   0 - 0x0
      13'h11AC: dout <= 8'b00000000; // 4524 :   0 - 0x0
      13'h11AD: dout <= 8'b00000000; // 4525 :   0 - 0x0
      13'h11AE: dout <= 8'b00000000; // 4526 :   0 - 0x0
      13'h11AF: dout <= 8'b00000000; // 4527 :   0 - 0x0
      13'h11B0: dout <= 8'b00000000; // 4528 :   0 - 0x0 -- Background 0x1b
      13'h11B1: dout <= 8'b00000000; // 4529 :   0 - 0x0
      13'h11B2: dout <= 8'b00000000; // 4530 :   0 - 0x0
      13'h11B3: dout <= 8'b00011000; // 4531 :  24 - 0x18
      13'h11B4: dout <= 8'b00100100; // 4532 :  36 - 0x24
      13'h11B5: dout <= 8'b00100100; // 4533 :  36 - 0x24
      13'h11B6: dout <= 8'b00100100; // 4534 :  36 - 0x24
      13'h11B7: dout <= 8'b00100100; // 4535 :  36 - 0x24
      13'h11B8: dout <= 8'b00000000; // 4536 :   0 - 0x0
      13'h11B9: dout <= 8'b00000000; // 4537 :   0 - 0x0
      13'h11BA: dout <= 8'b00000000; // 4538 :   0 - 0x0
      13'h11BB: dout <= 8'b00000000; // 4539 :   0 - 0x0
      13'h11BC: dout <= 8'b00000000; // 4540 :   0 - 0x0
      13'h11BD: dout <= 8'b00000000; // 4541 :   0 - 0x0
      13'h11BE: dout <= 8'b00000000; // 4542 :   0 - 0x0
      13'h11BF: dout <= 8'b00000000; // 4543 :   0 - 0x0
      13'h11C0: dout <= 8'b00100100; // 4544 :  36 - 0x24 -- Background 0x1c
      13'h11C1: dout <= 8'b00100100; // 4545 :  36 - 0x24
      13'h11C2: dout <= 8'b11000100; // 4546 : 196 - 0xc4
      13'h11C3: dout <= 8'b00000100; // 4547 :   4 - 0x4
      13'h11C4: dout <= 8'b00001000; // 4548 :   8 - 0x8
      13'h11C5: dout <= 8'b11110000; // 4549 : 240 - 0xf0
      13'h11C6: dout <= 8'b00000000; // 4550 :   0 - 0x0
      13'h11C7: dout <= 8'b00000000; // 4551 :   0 - 0x0
      13'h11C8: dout <= 8'b00000000; // 4552 :   0 - 0x0
      13'h11C9: dout <= 8'b00000000; // 4553 :   0 - 0x0
      13'h11CA: dout <= 8'b00000000; // 4554 :   0 - 0x0
      13'h11CB: dout <= 8'b00000000; // 4555 :   0 - 0x0
      13'h11CC: dout <= 8'b00000000; // 4556 :   0 - 0x0
      13'h11CD: dout <= 8'b00000000; // 4557 :   0 - 0x0
      13'h11CE: dout <= 8'b00000000; // 4558 :   0 - 0x0
      13'h11CF: dout <= 8'b00000000; // 4559 :   0 - 0x0
      13'h11D0: dout <= 8'b00000000; // 4560 :   0 - 0x0 -- Background 0x1d
      13'h11D1: dout <= 8'b00000000; // 4561 :   0 - 0x0
      13'h11D2: dout <= 8'b11110000; // 4562 : 240 - 0xf0
      13'h11D3: dout <= 8'b00001000; // 4563 :   8 - 0x8
      13'h11D4: dout <= 8'b00000100; // 4564 :   4 - 0x4
      13'h11D5: dout <= 8'b11000100; // 4565 : 196 - 0xc4
      13'h11D6: dout <= 8'b00100100; // 4566 :  36 - 0x24
      13'h11D7: dout <= 8'b00100100; // 4567 :  36 - 0x24
      13'h11D8: dout <= 8'b00000000; // 4568 :   0 - 0x0
      13'h11D9: dout <= 8'b00000000; // 4569 :   0 - 0x0
      13'h11DA: dout <= 8'b00000000; // 4570 :   0 - 0x0
      13'h11DB: dout <= 8'b00000000; // 4571 :   0 - 0x0
      13'h11DC: dout <= 8'b00000000; // 4572 :   0 - 0x0
      13'h11DD: dout <= 8'b00000000; // 4573 :   0 - 0x0
      13'h11DE: dout <= 8'b00000000; // 4574 :   0 - 0x0
      13'h11DF: dout <= 8'b00000000; // 4575 :   0 - 0x0
      13'h11E0: dout <= 8'b00100100; // 4576 :  36 - 0x24 -- Background 0x1e
      13'h11E1: dout <= 8'b00100100; // 4577 :  36 - 0x24
      13'h11E2: dout <= 8'b00100011; // 4578 :  35 - 0x23
      13'h11E3: dout <= 8'b00100000; // 4579 :  32 - 0x20
      13'h11E4: dout <= 8'b00010000; // 4580 :  16 - 0x10
      13'h11E5: dout <= 8'b00001111; // 4581 :  15 - 0xf
      13'h11E6: dout <= 8'b00000000; // 4582 :   0 - 0x0
      13'h11E7: dout <= 8'b00000000; // 4583 :   0 - 0x0
      13'h11E8: dout <= 8'b00000000; // 4584 :   0 - 0x0
      13'h11E9: dout <= 8'b00000000; // 4585 :   0 - 0x0
      13'h11EA: dout <= 8'b00000000; // 4586 :   0 - 0x0
      13'h11EB: dout <= 8'b00000000; // 4587 :   0 - 0x0
      13'h11EC: dout <= 8'b00000000; // 4588 :   0 - 0x0
      13'h11ED: dout <= 8'b00000000; // 4589 :   0 - 0x0
      13'h11EE: dout <= 8'b00000000; // 4590 :   0 - 0x0
      13'h11EF: dout <= 8'b00000000; // 4591 :   0 - 0x0
      13'h11F0: dout <= 8'b00000000; // 4592 :   0 - 0x0 -- Background 0x1f
      13'h11F1: dout <= 8'b00000000; // 4593 :   0 - 0x0
      13'h11F2: dout <= 8'b00001111; // 4594 :  15 - 0xf
      13'h11F3: dout <= 8'b00010000; // 4595 :  16 - 0x10
      13'h11F4: dout <= 8'b00100000; // 4596 :  32 - 0x20
      13'h11F5: dout <= 8'b00100011; // 4597 :  35 - 0x23
      13'h11F6: dout <= 8'b00100100; // 4598 :  36 - 0x24
      13'h11F7: dout <= 8'b00100100; // 4599 :  36 - 0x24
      13'h11F8: dout <= 8'b00000000; // 4600 :   0 - 0x0
      13'h11F9: dout <= 8'b00000000; // 4601 :   0 - 0x0
      13'h11FA: dout <= 8'b00000000; // 4602 :   0 - 0x0
      13'h11FB: dout <= 8'b00000000; // 4603 :   0 - 0x0
      13'h11FC: dout <= 8'b00000000; // 4604 :   0 - 0x0
      13'h11FD: dout <= 8'b00000000; // 4605 :   0 - 0x0
      13'h11FE: dout <= 8'b00000000; // 4606 :   0 - 0x0
      13'h11FF: dout <= 8'b00000000; // 4607 :   0 - 0x0
      13'h1200: dout <= 8'b00000000; // 4608 :   0 - 0x0 -- Background 0x20
      13'h1201: dout <= 8'b00000000; // 4609 :   0 - 0x0
      13'h1202: dout <= 8'b00000000; // 4610 :   0 - 0x0
      13'h1203: dout <= 8'b00000000; // 4611 :   0 - 0x0
      13'h1204: dout <= 8'b00000000; // 4612 :   0 - 0x0
      13'h1205: dout <= 8'b00000000; // 4613 :   0 - 0x0
      13'h1206: dout <= 8'b00000000; // 4614 :   0 - 0x0
      13'h1207: dout <= 8'b00000000; // 4615 :   0 - 0x0
      13'h1208: dout <= 8'b00000000; // 4616 :   0 - 0x0
      13'h1209: dout <= 8'b00000000; // 4617 :   0 - 0x0
      13'h120A: dout <= 8'b00000000; // 4618 :   0 - 0x0
      13'h120B: dout <= 8'b00000000; // 4619 :   0 - 0x0
      13'h120C: dout <= 8'b00000000; // 4620 :   0 - 0x0
      13'h120D: dout <= 8'b00000000; // 4621 :   0 - 0x0
      13'h120E: dout <= 8'b00000000; // 4622 :   0 - 0x0
      13'h120F: dout <= 8'b00000000; // 4623 :   0 - 0x0
      13'h1210: dout <= 8'b00000000; // 4624 :   0 - 0x0 -- Background 0x21
      13'h1211: dout <= 8'b00000000; // 4625 :   0 - 0x0
      13'h1212: dout <= 8'b11110000; // 4626 : 240 - 0xf0
      13'h1213: dout <= 8'b00001000; // 4627 :   8 - 0x8
      13'h1214: dout <= 8'b00001000; // 4628 :   8 - 0x8
      13'h1215: dout <= 8'b11110000; // 4629 : 240 - 0xf0
      13'h1216: dout <= 8'b00000000; // 4630 :   0 - 0x0
      13'h1217: dout <= 8'b00000000; // 4631 :   0 - 0x0
      13'h1218: dout <= 8'b00001111; // 4632 :  15 - 0xf
      13'h1219: dout <= 8'b00001111; // 4633 :  15 - 0xf
      13'h121A: dout <= 8'b00001111; // 4634 :  15 - 0xf
      13'h121B: dout <= 8'b00000111; // 4635 :   7 - 0x7
      13'h121C: dout <= 8'b00000111; // 4636 :   7 - 0x7
      13'h121D: dout <= 8'b00001111; // 4637 :  15 - 0xf
      13'h121E: dout <= 8'b00001111; // 4638 :  15 - 0xf
      13'h121F: dout <= 8'b00001111; // 4639 :  15 - 0xf
      13'h1220: dout <= 8'b00000000; // 4640 :   0 - 0x0 -- Background 0x22
      13'h1221: dout <= 8'b00000000; // 4641 :   0 - 0x0
      13'h1222: dout <= 8'b00001111; // 4642 :  15 - 0xf
      13'h1223: dout <= 8'b00010000; // 4643 :  16 - 0x10
      13'h1224: dout <= 8'b00010000; // 4644 :  16 - 0x10
      13'h1225: dout <= 8'b00001111; // 4645 :  15 - 0xf
      13'h1226: dout <= 8'b00000000; // 4646 :   0 - 0x0
      13'h1227: dout <= 8'b00000000; // 4647 :   0 - 0x0
      13'h1228: dout <= 8'b11110000; // 4648 : 240 - 0xf0
      13'h1229: dout <= 8'b11110000; // 4649 : 240 - 0xf0
      13'h122A: dout <= 8'b11110000; // 4650 : 240 - 0xf0
      13'h122B: dout <= 8'b11100000; // 4651 : 224 - 0xe0
      13'h122C: dout <= 8'b11100000; // 4652 : 224 - 0xe0
      13'h122D: dout <= 8'b11110000; // 4653 : 240 - 0xf0
      13'h122E: dout <= 8'b11110000; // 4654 : 240 - 0xf0
      13'h122F: dout <= 8'b11110000; // 4655 : 240 - 0xf0
      13'h1230: dout <= 8'b11111111; // 4656 : 255 - 0xff -- Background 0x23
      13'h1231: dout <= 8'b11111111; // 4657 : 255 - 0xff
      13'h1232: dout <= 8'b11100001; // 4658 : 225 - 0xe1
      13'h1233: dout <= 8'b11100001; // 4659 : 225 - 0xe1
      13'h1234: dout <= 8'b11100001; // 4660 : 225 - 0xe1
      13'h1235: dout <= 8'b11100001; // 4661 : 225 - 0xe1
      13'h1236: dout <= 8'b11100001; // 4662 : 225 - 0xe1
      13'h1237: dout <= 8'b11100001; // 4663 : 225 - 0xe1
      13'h1238: dout <= 8'b11111111; // 4664 : 255 - 0xff
      13'h1239: dout <= 8'b11111111; // 4665 : 255 - 0xff
      13'h123A: dout <= 8'b11100001; // 4666 : 225 - 0xe1
      13'h123B: dout <= 8'b11100001; // 4667 : 225 - 0xe1
      13'h123C: dout <= 8'b11100001; // 4668 : 225 - 0xe1
      13'h123D: dout <= 8'b11100001; // 4669 : 225 - 0xe1
      13'h123E: dout <= 8'b11100001; // 4670 : 225 - 0xe1
      13'h123F: dout <= 8'b11100001; // 4671 : 225 - 0xe1
      13'h1240: dout <= 8'b10000111; // 4672 : 135 - 0x87 -- Background 0x24
      13'h1241: dout <= 8'b11000111; // 4673 : 199 - 0xc7
      13'h1242: dout <= 8'b11000000; // 4674 : 192 - 0xc0
      13'h1243: dout <= 8'b11000111; // 4675 : 199 - 0xc7
      13'h1244: dout <= 8'b11001111; // 4676 : 207 - 0xcf
      13'h1245: dout <= 8'b11001110; // 4677 : 206 - 0xce
      13'h1246: dout <= 8'b11001111; // 4678 : 207 - 0xcf
      13'h1247: dout <= 8'b11000111; // 4679 : 199 - 0xc7
      13'h1248: dout <= 8'b10000111; // 4680 : 135 - 0x87
      13'h1249: dout <= 8'b11000111; // 4681 : 199 - 0xc7
      13'h124A: dout <= 8'b11000000; // 4682 : 192 - 0xc0
      13'h124B: dout <= 8'b11000111; // 4683 : 199 - 0xc7
      13'h124C: dout <= 8'b11001111; // 4684 : 207 - 0xcf
      13'h124D: dout <= 8'b11001110; // 4685 : 206 - 0xce
      13'h124E: dout <= 8'b11001111; // 4686 : 207 - 0xcf
      13'h124F: dout <= 8'b11000111; // 4687 : 199 - 0xc7
      13'h1250: dout <= 8'b11111000; // 4688 : 248 - 0xf8 -- Background 0x25
      13'h1251: dout <= 8'b11111100; // 4689 : 252 - 0xfc
      13'h1252: dout <= 8'b00011100; // 4690 :  28 - 0x1c
      13'h1253: dout <= 8'b11111100; // 4691 : 252 - 0xfc
      13'h1254: dout <= 8'b11111100; // 4692 : 252 - 0xfc
      13'h1255: dout <= 8'b00011100; // 4693 :  28 - 0x1c
      13'h1256: dout <= 8'b11111100; // 4694 : 252 - 0xfc
      13'h1257: dout <= 8'b11111100; // 4695 : 252 - 0xfc
      13'h1258: dout <= 8'b11111000; // 4696 : 248 - 0xf8
      13'h1259: dout <= 8'b11111100; // 4697 : 252 - 0xfc
      13'h125A: dout <= 8'b00011100; // 4698 :  28 - 0x1c
      13'h125B: dout <= 8'b11111100; // 4699 : 252 - 0xfc
      13'h125C: dout <= 8'b11111100; // 4700 : 252 - 0xfc
      13'h125D: dout <= 8'b00011100; // 4701 :  28 - 0x1c
      13'h125E: dout <= 8'b11111100; // 4702 : 252 - 0xfc
      13'h125F: dout <= 8'b11111100; // 4703 : 252 - 0xfc
      13'h1260: dout <= 8'b11111111; // 4704 : 255 - 0xff -- Background 0x26
      13'h1261: dout <= 8'b11111111; // 4705 : 255 - 0xff
      13'h1262: dout <= 8'b11100111; // 4706 : 231 - 0xe7
      13'h1263: dout <= 8'b11100111; // 4707 : 231 - 0xe7
      13'h1264: dout <= 8'b11100111; // 4708 : 231 - 0xe7
      13'h1265: dout <= 8'b11100111; // 4709 : 231 - 0xe7
      13'h1266: dout <= 8'b11100111; // 4710 : 231 - 0xe7
      13'h1267: dout <= 8'b11100111; // 4711 : 231 - 0xe7
      13'h1268: dout <= 8'b11111111; // 4712 : 255 - 0xff
      13'h1269: dout <= 8'b11111111; // 4713 : 255 - 0xff
      13'h126A: dout <= 8'b11100111; // 4714 : 231 - 0xe7
      13'h126B: dout <= 8'b11100111; // 4715 : 231 - 0xe7
      13'h126C: dout <= 8'b11100111; // 4716 : 231 - 0xe7
      13'h126D: dout <= 8'b11100111; // 4717 : 231 - 0xe7
      13'h126E: dout <= 8'b11100111; // 4718 : 231 - 0xe7
      13'h126F: dout <= 8'b11100111; // 4719 : 231 - 0xe7
      13'h1270: dout <= 8'b11110000; // 4720 : 240 - 0xf0 -- Background 0x27
      13'h1271: dout <= 8'b11111001; // 4721 : 249 - 0xf9
      13'h1272: dout <= 8'b00111001; // 4722 :  57 - 0x39
      13'h1273: dout <= 8'b00111001; // 4723 :  57 - 0x39
      13'h1274: dout <= 8'b00111001; // 4724 :  57 - 0x39
      13'h1275: dout <= 8'b00111001; // 4725 :  57 - 0x39
      13'h1276: dout <= 8'b00111001; // 4726 :  57 - 0x39
      13'h1277: dout <= 8'b00111000; // 4727 :  56 - 0x38
      13'h1278: dout <= 8'b11110000; // 4728 : 240 - 0xf0
      13'h1279: dout <= 8'b11111001; // 4729 : 249 - 0xf9
      13'h127A: dout <= 8'b00111001; // 4730 :  57 - 0x39
      13'h127B: dout <= 8'b00111001; // 4731 :  57 - 0x39
      13'h127C: dout <= 8'b00111001; // 4732 :  57 - 0x39
      13'h127D: dout <= 8'b00111001; // 4733 :  57 - 0x39
      13'h127E: dout <= 8'b00111001; // 4734 :  57 - 0x39
      13'h127F: dout <= 8'b00111000; // 4735 :  56 - 0x38
      13'h1280: dout <= 8'b11111111; // 4736 : 255 - 0xff -- Background 0x28
      13'h1281: dout <= 8'b11111111; // 4737 : 255 - 0xff
      13'h1282: dout <= 8'b11000000; // 4738 : 192 - 0xc0
      13'h1283: dout <= 8'b11000000; // 4739 : 192 - 0xc0
      13'h1284: dout <= 8'b11000000; // 4740 : 192 - 0xc0
      13'h1285: dout <= 8'b11000000; // 4741 : 192 - 0xc0
      13'h1286: dout <= 8'b11111111; // 4742 : 255 - 0xff
      13'h1287: dout <= 8'b11111111; // 4743 : 255 - 0xff
      13'h1288: dout <= 8'b11111111; // 4744 : 255 - 0xff
      13'h1289: dout <= 8'b11111111; // 4745 : 255 - 0xff
      13'h128A: dout <= 8'b11000000; // 4746 : 192 - 0xc0
      13'h128B: dout <= 8'b11000000; // 4747 : 192 - 0xc0
      13'h128C: dout <= 8'b11000000; // 4748 : 192 - 0xc0
      13'h128D: dout <= 8'b11000000; // 4749 : 192 - 0xc0
      13'h128E: dout <= 8'b11111111; // 4750 : 255 - 0xff
      13'h128F: dout <= 8'b11111111; // 4751 : 255 - 0xff
      13'h1290: dout <= 8'b00011111; // 4752 :  31 - 0x1f -- Background 0x29
      13'h1291: dout <= 8'b00111111; // 4753 :  63 - 0x3f
      13'h1292: dout <= 8'b00110000; // 4754 :  48 - 0x30
      13'h1293: dout <= 8'b00110000; // 4755 :  48 - 0x30
      13'h1294: dout <= 8'b00110000; // 4756 :  48 - 0x30
      13'h1295: dout <= 8'b00110000; // 4757 :  48 - 0x30
      13'h1296: dout <= 8'b00111111; // 4758 :  63 - 0x3f
      13'h1297: dout <= 8'b00011111; // 4759 :  31 - 0x1f
      13'h1298: dout <= 8'b00011111; // 4760 :  31 - 0x1f
      13'h1299: dout <= 8'b00111111; // 4761 :  63 - 0x3f
      13'h129A: dout <= 8'b00110000; // 4762 :  48 - 0x30
      13'h129B: dout <= 8'b00110000; // 4763 :  48 - 0x30
      13'h129C: dout <= 8'b00110000; // 4764 :  48 - 0x30
      13'h129D: dout <= 8'b00110000; // 4765 :  48 - 0x30
      13'h129E: dout <= 8'b00111111; // 4766 :  63 - 0x3f
      13'h129F: dout <= 8'b00011111; // 4767 :  31 - 0x1f
      13'h12A0: dout <= 8'b11100011; // 4768 : 227 - 0xe3 -- Background 0x2a
      13'h12A1: dout <= 8'b11110011; // 4769 : 243 - 0xf3
      13'h12A2: dout <= 8'b01110000; // 4770 : 112 - 0x70
      13'h12A3: dout <= 8'b01110000; // 4771 : 112 - 0x70
      13'h12A4: dout <= 8'b01110000; // 4772 : 112 - 0x70
      13'h12A5: dout <= 8'b01110000; // 4773 : 112 - 0x70
      13'h12A6: dout <= 8'b11110000; // 4774 : 240 - 0xf0
      13'h12A7: dout <= 8'b11100000; // 4775 : 224 - 0xe0
      13'h12A8: dout <= 8'b11100011; // 4776 : 227 - 0xe3
      13'h12A9: dout <= 8'b11110011; // 4777 : 243 - 0xf3
      13'h12AA: dout <= 8'b01110000; // 4778 : 112 - 0x70
      13'h12AB: dout <= 8'b01110000; // 4779 : 112 - 0x70
      13'h12AC: dout <= 8'b01110000; // 4780 : 112 - 0x70
      13'h12AD: dout <= 8'b01110000; // 4781 : 112 - 0x70
      13'h12AE: dout <= 8'b11110000; // 4782 : 240 - 0xf0
      13'h12AF: dout <= 8'b11100000; // 4783 : 224 - 0xe0
      13'h12B0: dout <= 8'b11111110; // 4784 : 254 - 0xfe -- Background 0x2b
      13'h12B1: dout <= 8'b11111110; // 4785 : 254 - 0xfe
      13'h12B2: dout <= 8'b01110000; // 4786 : 112 - 0x70
      13'h12B3: dout <= 8'b01110000; // 4787 : 112 - 0x70
      13'h12B4: dout <= 8'b01110000; // 4788 : 112 - 0x70
      13'h12B5: dout <= 8'b01110000; // 4789 : 112 - 0x70
      13'h12B6: dout <= 8'b01110000; // 4790 : 112 - 0x70
      13'h12B7: dout <= 8'b01110000; // 4791 : 112 - 0x70
      13'h12B8: dout <= 8'b11111110; // 4792 : 254 - 0xfe
      13'h12B9: dout <= 8'b11111110; // 4793 : 254 - 0xfe
      13'h12BA: dout <= 8'b01110000; // 4794 : 112 - 0x70
      13'h12BB: dout <= 8'b01110000; // 4795 : 112 - 0x70
      13'h12BC: dout <= 8'b01110000; // 4796 : 112 - 0x70
      13'h12BD: dout <= 8'b01110000; // 4797 : 112 - 0x70
      13'h12BE: dout <= 8'b01110000; // 4798 : 112 - 0x70
      13'h12BF: dout <= 8'b01110000; // 4799 : 112 - 0x70
      13'h12C0: dout <= 8'b00000000; // 4800 :   0 - 0x0 -- Background 0x2c
      13'h12C1: dout <= 8'b00000000; // 4801 :   0 - 0x0
      13'h12C2: dout <= 8'b00000000; // 4802 :   0 - 0x0
      13'h12C3: dout <= 8'b00000000; // 4803 :   0 - 0x0
      13'h12C4: dout <= 8'b11111111; // 4804 : 255 - 0xff
      13'h12C5: dout <= 8'b00000000; // 4805 :   0 - 0x0
      13'h12C6: dout <= 8'b00000000; // 4806 :   0 - 0x0
      13'h12C7: dout <= 8'b00000000; // 4807 :   0 - 0x0
      13'h12C8: dout <= 8'b00000000; // 4808 :   0 - 0x0
      13'h12C9: dout <= 8'b00000000; // 4809 :   0 - 0x0
      13'h12CA: dout <= 8'b00000000; // 4810 :   0 - 0x0
      13'h12CB: dout <= 8'b00000000; // 4811 :   0 - 0x0
      13'h12CC: dout <= 8'b00000000; // 4812 :   0 - 0x0
      13'h12CD: dout <= 8'b00000000; // 4813 :   0 - 0x0
      13'h12CE: dout <= 8'b00000000; // 4814 :   0 - 0x0
      13'h12CF: dout <= 8'b00000000; // 4815 :   0 - 0x0
      13'h12D0: dout <= 8'b00000000; // 4816 :   0 - 0x0 -- Background 0x2d
      13'h12D1: dout <= 8'b00000000; // 4817 :   0 - 0x0
      13'h12D2: dout <= 8'b00000000; // 4818 :   0 - 0x0
      13'h12D3: dout <= 8'b00000000; // 4819 :   0 - 0x0
      13'h12D4: dout <= 8'b00000000; // 4820 :   0 - 0x0
      13'h12D5: dout <= 8'b00000000; // 4821 :   0 - 0x0
      13'h12D6: dout <= 8'b00000000; // 4822 :   0 - 0x0
      13'h12D7: dout <= 8'b00000000; // 4823 :   0 - 0x0
      13'h12D8: dout <= 8'b11111111; // 4824 : 255 - 0xff
      13'h12D9: dout <= 8'b11111111; // 4825 : 255 - 0xff
      13'h12DA: dout <= 8'b11111111; // 4826 : 255 - 0xff
      13'h12DB: dout <= 8'b11111111; // 4827 : 255 - 0xff
      13'h12DC: dout <= 8'b11111111; // 4828 : 255 - 0xff
      13'h12DD: dout <= 8'b11111111; // 4829 : 255 - 0xff
      13'h12DE: dout <= 8'b11111111; // 4830 : 255 - 0xff
      13'h12DF: dout <= 8'b11111111; // 4831 : 255 - 0xff
      13'h12E0: dout <= 8'b00000000; // 4832 :   0 - 0x0 -- Background 0x2e
      13'h12E1: dout <= 8'b00000000; // 4833 :   0 - 0x0
      13'h12E2: dout <= 8'b00000000; // 4834 :   0 - 0x0
      13'h12E3: dout <= 8'b00011000; // 4835 :  24 - 0x18
      13'h12E4: dout <= 8'b00011000; // 4836 :  24 - 0x18
      13'h12E5: dout <= 8'b00000000; // 4837 :   0 - 0x0
      13'h12E6: dout <= 8'b00000000; // 4838 :   0 - 0x0
      13'h12E7: dout <= 8'b00000000; // 4839 :   0 - 0x0
      13'h12E8: dout <= 8'b00000000; // 4840 :   0 - 0x0
      13'h12E9: dout <= 8'b00000000; // 4841 :   0 - 0x0
      13'h12EA: dout <= 8'b00000000; // 4842 :   0 - 0x0
      13'h12EB: dout <= 8'b00000000; // 4843 :   0 - 0x0
      13'h12EC: dout <= 8'b00000000; // 4844 :   0 - 0x0
      13'h12ED: dout <= 8'b00000000; // 4845 :   0 - 0x0
      13'h12EE: dout <= 8'b00000000; // 4846 :   0 - 0x0
      13'h12EF: dout <= 8'b00000000; // 4847 :   0 - 0x0
      13'h12F0: dout <= 8'b00000000; // 4848 :   0 - 0x0 -- Background 0x2f
      13'h12F1: dout <= 8'b00000000; // 4849 :   0 - 0x0
      13'h12F2: dout <= 8'b00000000; // 4850 :   0 - 0x0
      13'h12F3: dout <= 8'b00000000; // 4851 :   0 - 0x0
      13'h12F4: dout <= 8'b00000000; // 4852 :   0 - 0x0
      13'h12F5: dout <= 8'b00000000; // 4853 :   0 - 0x0
      13'h12F6: dout <= 8'b00000000; // 4854 :   0 - 0x0
      13'h12F7: dout <= 8'b00000000; // 4855 :   0 - 0x0
      13'h12F8: dout <= 8'b00000000; // 4856 :   0 - 0x0
      13'h12F9: dout <= 8'b00000000; // 4857 :   0 - 0x0
      13'h12FA: dout <= 8'b00000000; // 4858 :   0 - 0x0
      13'h12FB: dout <= 8'b00011000; // 4859 :  24 - 0x18
      13'h12FC: dout <= 8'b00011000; // 4860 :  24 - 0x18
      13'h12FD: dout <= 8'b00000000; // 4861 :   0 - 0x0
      13'h12FE: dout <= 8'b00000000; // 4862 :   0 - 0x0
      13'h12FF: dout <= 8'b00000000; // 4863 :   0 - 0x0
      13'h1300: dout <= 8'b00011100; // 4864 :  28 - 0x1c -- Background 0x30
      13'h1301: dout <= 8'b00100110; // 4865 :  38 - 0x26
      13'h1302: dout <= 8'b01100011; // 4866 :  99 - 0x63
      13'h1303: dout <= 8'b01100011; // 4867 :  99 - 0x63
      13'h1304: dout <= 8'b01100011; // 4868 :  99 - 0x63
      13'h1305: dout <= 8'b00110010; // 4869 :  50 - 0x32
      13'h1306: dout <= 8'b00011100; // 4870 :  28 - 0x1c
      13'h1307: dout <= 8'b00000000; // 4871 :   0 - 0x0
      13'h1308: dout <= 8'b00000000; // 4872 :   0 - 0x0
      13'h1309: dout <= 8'b00000000; // 4873 :   0 - 0x0
      13'h130A: dout <= 8'b00000000; // 4874 :   0 - 0x0
      13'h130B: dout <= 8'b00000000; // 4875 :   0 - 0x0
      13'h130C: dout <= 8'b00000000; // 4876 :   0 - 0x0
      13'h130D: dout <= 8'b00000000; // 4877 :   0 - 0x0
      13'h130E: dout <= 8'b00000000; // 4878 :   0 - 0x0
      13'h130F: dout <= 8'b00000000; // 4879 :   0 - 0x0
      13'h1310: dout <= 8'b00001100; // 4880 :  12 - 0xc -- Background 0x31
      13'h1311: dout <= 8'b00011100; // 4881 :  28 - 0x1c
      13'h1312: dout <= 8'b00001100; // 4882 :  12 - 0xc
      13'h1313: dout <= 8'b00001100; // 4883 :  12 - 0xc
      13'h1314: dout <= 8'b00001100; // 4884 :  12 - 0xc
      13'h1315: dout <= 8'b00001100; // 4885 :  12 - 0xc
      13'h1316: dout <= 8'b00111111; // 4886 :  63 - 0x3f
      13'h1317: dout <= 8'b00000000; // 4887 :   0 - 0x0
      13'h1318: dout <= 8'b00000000; // 4888 :   0 - 0x0
      13'h1319: dout <= 8'b00000000; // 4889 :   0 - 0x0
      13'h131A: dout <= 8'b00000000; // 4890 :   0 - 0x0
      13'h131B: dout <= 8'b00000000; // 4891 :   0 - 0x0
      13'h131C: dout <= 8'b00000000; // 4892 :   0 - 0x0
      13'h131D: dout <= 8'b00000000; // 4893 :   0 - 0x0
      13'h131E: dout <= 8'b00000000; // 4894 :   0 - 0x0
      13'h131F: dout <= 8'b00000000; // 4895 :   0 - 0x0
      13'h1320: dout <= 8'b00111110; // 4896 :  62 - 0x3e -- Background 0x32
      13'h1321: dout <= 8'b01100011; // 4897 :  99 - 0x63
      13'h1322: dout <= 8'b00000111; // 4898 :   7 - 0x7
      13'h1323: dout <= 8'b00011110; // 4899 :  30 - 0x1e
      13'h1324: dout <= 8'b00111100; // 4900 :  60 - 0x3c
      13'h1325: dout <= 8'b01110000; // 4901 : 112 - 0x70
      13'h1326: dout <= 8'b01111111; // 4902 : 127 - 0x7f
      13'h1327: dout <= 8'b00000000; // 4903 :   0 - 0x0
      13'h1328: dout <= 8'b00000000; // 4904 :   0 - 0x0
      13'h1329: dout <= 8'b00000000; // 4905 :   0 - 0x0
      13'h132A: dout <= 8'b00000000; // 4906 :   0 - 0x0
      13'h132B: dout <= 8'b00000000; // 4907 :   0 - 0x0
      13'h132C: dout <= 8'b00000000; // 4908 :   0 - 0x0
      13'h132D: dout <= 8'b00000000; // 4909 :   0 - 0x0
      13'h132E: dout <= 8'b00000000; // 4910 :   0 - 0x0
      13'h132F: dout <= 8'b00000000; // 4911 :   0 - 0x0
      13'h1330: dout <= 8'b00111111; // 4912 :  63 - 0x3f -- Background 0x33
      13'h1331: dout <= 8'b00000110; // 4913 :   6 - 0x6
      13'h1332: dout <= 8'b00001100; // 4914 :  12 - 0xc
      13'h1333: dout <= 8'b00011110; // 4915 :  30 - 0x1e
      13'h1334: dout <= 8'b00000011; // 4916 :   3 - 0x3
      13'h1335: dout <= 8'b01100011; // 4917 :  99 - 0x63
      13'h1336: dout <= 8'b00111110; // 4918 :  62 - 0x3e
      13'h1337: dout <= 8'b00000000; // 4919 :   0 - 0x0
      13'h1338: dout <= 8'b00000000; // 4920 :   0 - 0x0
      13'h1339: dout <= 8'b00000000; // 4921 :   0 - 0x0
      13'h133A: dout <= 8'b00000000; // 4922 :   0 - 0x0
      13'h133B: dout <= 8'b00000000; // 4923 :   0 - 0x0
      13'h133C: dout <= 8'b00000000; // 4924 :   0 - 0x0
      13'h133D: dout <= 8'b00000000; // 4925 :   0 - 0x0
      13'h133E: dout <= 8'b00000000; // 4926 :   0 - 0x0
      13'h133F: dout <= 8'b00000000; // 4927 :   0 - 0x0
      13'h1340: dout <= 8'b00001110; // 4928 :  14 - 0xe -- Background 0x34
      13'h1341: dout <= 8'b00011110; // 4929 :  30 - 0x1e
      13'h1342: dout <= 8'b00110110; // 4930 :  54 - 0x36
      13'h1343: dout <= 8'b01100110; // 4931 : 102 - 0x66
      13'h1344: dout <= 8'b01111111; // 4932 : 127 - 0x7f
      13'h1345: dout <= 8'b00000110; // 4933 :   6 - 0x6
      13'h1346: dout <= 8'b00000110; // 4934 :   6 - 0x6
      13'h1347: dout <= 8'b00000000; // 4935 :   0 - 0x0
      13'h1348: dout <= 8'b00000000; // 4936 :   0 - 0x0
      13'h1349: dout <= 8'b00000000; // 4937 :   0 - 0x0
      13'h134A: dout <= 8'b00000000; // 4938 :   0 - 0x0
      13'h134B: dout <= 8'b00000000; // 4939 :   0 - 0x0
      13'h134C: dout <= 8'b00000000; // 4940 :   0 - 0x0
      13'h134D: dout <= 8'b00000000; // 4941 :   0 - 0x0
      13'h134E: dout <= 8'b00000000; // 4942 :   0 - 0x0
      13'h134F: dout <= 8'b00000000; // 4943 :   0 - 0x0
      13'h1350: dout <= 8'b01111110; // 4944 : 126 - 0x7e -- Background 0x35
      13'h1351: dout <= 8'b01100000; // 4945 :  96 - 0x60
      13'h1352: dout <= 8'b01111110; // 4946 : 126 - 0x7e
      13'h1353: dout <= 8'b00000011; // 4947 :   3 - 0x3
      13'h1354: dout <= 8'b00000011; // 4948 :   3 - 0x3
      13'h1355: dout <= 8'b01100011; // 4949 :  99 - 0x63
      13'h1356: dout <= 8'b00111110; // 4950 :  62 - 0x3e
      13'h1357: dout <= 8'b00000000; // 4951 :   0 - 0x0
      13'h1358: dout <= 8'b00000000; // 4952 :   0 - 0x0
      13'h1359: dout <= 8'b00000000; // 4953 :   0 - 0x0
      13'h135A: dout <= 8'b00000000; // 4954 :   0 - 0x0
      13'h135B: dout <= 8'b00000000; // 4955 :   0 - 0x0
      13'h135C: dout <= 8'b00000000; // 4956 :   0 - 0x0
      13'h135D: dout <= 8'b00000000; // 4957 :   0 - 0x0
      13'h135E: dout <= 8'b00000000; // 4958 :   0 - 0x0
      13'h135F: dout <= 8'b00000000; // 4959 :   0 - 0x0
      13'h1360: dout <= 8'b00011110; // 4960 :  30 - 0x1e -- Background 0x36
      13'h1361: dout <= 8'b00110000; // 4961 :  48 - 0x30
      13'h1362: dout <= 8'b01100000; // 4962 :  96 - 0x60
      13'h1363: dout <= 8'b01111110; // 4963 : 126 - 0x7e
      13'h1364: dout <= 8'b01100011; // 4964 :  99 - 0x63
      13'h1365: dout <= 8'b01100011; // 4965 :  99 - 0x63
      13'h1366: dout <= 8'b00111110; // 4966 :  62 - 0x3e
      13'h1367: dout <= 8'b00000000; // 4967 :   0 - 0x0
      13'h1368: dout <= 8'b00000000; // 4968 :   0 - 0x0
      13'h1369: dout <= 8'b00000000; // 4969 :   0 - 0x0
      13'h136A: dout <= 8'b00000000; // 4970 :   0 - 0x0
      13'h136B: dout <= 8'b00000000; // 4971 :   0 - 0x0
      13'h136C: dout <= 8'b00000000; // 4972 :   0 - 0x0
      13'h136D: dout <= 8'b00000000; // 4973 :   0 - 0x0
      13'h136E: dout <= 8'b00000000; // 4974 :   0 - 0x0
      13'h136F: dout <= 8'b00000000; // 4975 :   0 - 0x0
      13'h1370: dout <= 8'b01111111; // 4976 : 127 - 0x7f -- Background 0x37
      13'h1371: dout <= 8'b01100011; // 4977 :  99 - 0x63
      13'h1372: dout <= 8'b00000110; // 4978 :   6 - 0x6
      13'h1373: dout <= 8'b00001100; // 4979 :  12 - 0xc
      13'h1374: dout <= 8'b00011000; // 4980 :  24 - 0x18
      13'h1375: dout <= 8'b00011000; // 4981 :  24 - 0x18
      13'h1376: dout <= 8'b00011000; // 4982 :  24 - 0x18
      13'h1377: dout <= 8'b00000000; // 4983 :   0 - 0x0
      13'h1378: dout <= 8'b00000000; // 4984 :   0 - 0x0
      13'h1379: dout <= 8'b00000000; // 4985 :   0 - 0x0
      13'h137A: dout <= 8'b00000000; // 4986 :   0 - 0x0
      13'h137B: dout <= 8'b00000000; // 4987 :   0 - 0x0
      13'h137C: dout <= 8'b00000000; // 4988 :   0 - 0x0
      13'h137D: dout <= 8'b00000000; // 4989 :   0 - 0x0
      13'h137E: dout <= 8'b00000000; // 4990 :   0 - 0x0
      13'h137F: dout <= 8'b00000000; // 4991 :   0 - 0x0
      13'h1380: dout <= 8'b00111100; // 4992 :  60 - 0x3c -- Background 0x38
      13'h1381: dout <= 8'b01100010; // 4993 :  98 - 0x62
      13'h1382: dout <= 8'b01110010; // 4994 : 114 - 0x72
      13'h1383: dout <= 8'b00111100; // 4995 :  60 - 0x3c
      13'h1384: dout <= 8'b01001111; // 4996 :  79 - 0x4f
      13'h1385: dout <= 8'b01000011; // 4997 :  67 - 0x43
      13'h1386: dout <= 8'b00111110; // 4998 :  62 - 0x3e
      13'h1387: dout <= 8'b00000000; // 4999 :   0 - 0x0
      13'h1388: dout <= 8'b00000000; // 5000 :   0 - 0x0
      13'h1389: dout <= 8'b00000000; // 5001 :   0 - 0x0
      13'h138A: dout <= 8'b00000000; // 5002 :   0 - 0x0
      13'h138B: dout <= 8'b00000000; // 5003 :   0 - 0x0
      13'h138C: dout <= 8'b00000000; // 5004 :   0 - 0x0
      13'h138D: dout <= 8'b00000000; // 5005 :   0 - 0x0
      13'h138E: dout <= 8'b00000000; // 5006 :   0 - 0x0
      13'h138F: dout <= 8'b00000000; // 5007 :   0 - 0x0
      13'h1390: dout <= 8'b00111110; // 5008 :  62 - 0x3e -- Background 0x39
      13'h1391: dout <= 8'b01100011; // 5009 :  99 - 0x63
      13'h1392: dout <= 8'b01100011; // 5010 :  99 - 0x63
      13'h1393: dout <= 8'b00111111; // 5011 :  63 - 0x3f
      13'h1394: dout <= 8'b00000011; // 5012 :   3 - 0x3
      13'h1395: dout <= 8'b00000110; // 5013 :   6 - 0x6
      13'h1396: dout <= 8'b00111100; // 5014 :  60 - 0x3c
      13'h1397: dout <= 8'b00000000; // 5015 :   0 - 0x0
      13'h1398: dout <= 8'b00000000; // 5016 :   0 - 0x0
      13'h1399: dout <= 8'b00000000; // 5017 :   0 - 0x0
      13'h139A: dout <= 8'b00000000; // 5018 :   0 - 0x0
      13'h139B: dout <= 8'b00000000; // 5019 :   0 - 0x0
      13'h139C: dout <= 8'b00000000; // 5020 :   0 - 0x0
      13'h139D: dout <= 8'b00000000; // 5021 :   0 - 0x0
      13'h139E: dout <= 8'b00000000; // 5022 :   0 - 0x0
      13'h139F: dout <= 8'b00000000; // 5023 :   0 - 0x0
      13'h13A0: dout <= 8'b00000000; // 5024 :   0 - 0x0 -- Background 0x3a
      13'h13A1: dout <= 8'b00000000; // 5025 :   0 - 0x0
      13'h13A2: dout <= 8'b00000000; // 5026 :   0 - 0x0
      13'h13A3: dout <= 8'b01111110; // 5027 : 126 - 0x7e
      13'h13A4: dout <= 8'b00000000; // 5028 :   0 - 0x0
      13'h13A5: dout <= 8'b00000000; // 5029 :   0 - 0x0
      13'h13A6: dout <= 8'b00000000; // 5030 :   0 - 0x0
      13'h13A7: dout <= 8'b00000000; // 5031 :   0 - 0x0
      13'h13A8: dout <= 8'b00000000; // 5032 :   0 - 0x0
      13'h13A9: dout <= 8'b00000000; // 5033 :   0 - 0x0
      13'h13AA: dout <= 8'b00000000; // 5034 :   0 - 0x0
      13'h13AB: dout <= 8'b00000000; // 5035 :   0 - 0x0
      13'h13AC: dout <= 8'b00000000; // 5036 :   0 - 0x0
      13'h13AD: dout <= 8'b00000000; // 5037 :   0 - 0x0
      13'h13AE: dout <= 8'b00000000; // 5038 :   0 - 0x0
      13'h13AF: dout <= 8'b00000000; // 5039 :   0 - 0x0
      13'h13B0: dout <= 8'b00000000; // 5040 :   0 - 0x0 -- Background 0x3b
      13'h13B1: dout <= 8'b00000010; // 5041 :   2 - 0x2
      13'h13B2: dout <= 8'b00000100; // 5042 :   4 - 0x4
      13'h13B3: dout <= 8'b00001000; // 5043 :   8 - 0x8
      13'h13B4: dout <= 8'b00010000; // 5044 :  16 - 0x10
      13'h13B5: dout <= 8'b00100000; // 5045 :  32 - 0x20
      13'h13B6: dout <= 8'b00000000; // 5046 :   0 - 0x0
      13'h13B7: dout <= 8'b00000000; // 5047 :   0 - 0x0
      13'h13B8: dout <= 8'b00000000; // 5048 :   0 - 0x0
      13'h13B9: dout <= 8'b00000000; // 5049 :   0 - 0x0
      13'h13BA: dout <= 8'b00000000; // 5050 :   0 - 0x0
      13'h13BB: dout <= 8'b00000000; // 5051 :   0 - 0x0
      13'h13BC: dout <= 8'b00000000; // 5052 :   0 - 0x0
      13'h13BD: dout <= 8'b00000000; // 5053 :   0 - 0x0
      13'h13BE: dout <= 8'b00000000; // 5054 :   0 - 0x0
      13'h13BF: dout <= 8'b00000000; // 5055 :   0 - 0x0
      13'h13C0: dout <= 8'b00000000; // 5056 :   0 - 0x0 -- Background 0x3c
      13'h13C1: dout <= 8'b00000111; // 5057 :   7 - 0x7
      13'h13C2: dout <= 8'b00011111; // 5058 :  31 - 0x1f
      13'h13C3: dout <= 8'b00111111; // 5059 :  63 - 0x3f
      13'h13C4: dout <= 8'b00111111; // 5060 :  63 - 0x3f
      13'h13C5: dout <= 8'b00001111; // 5061 :  15 - 0xf
      13'h13C6: dout <= 8'b00000011; // 5062 :   3 - 0x3
      13'h13C7: dout <= 8'b00000000; // 5063 :   0 - 0x0
      13'h13C8: dout <= 8'b00000000; // 5064 :   0 - 0x0
      13'h13C9: dout <= 8'b00000111; // 5065 :   7 - 0x7
      13'h13CA: dout <= 8'b00011111; // 5066 :  31 - 0x1f
      13'h13CB: dout <= 8'b00111111; // 5067 :  63 - 0x3f
      13'h13CC: dout <= 8'b00111111; // 5068 :  63 - 0x3f
      13'h13CD: dout <= 8'b00001111; // 5069 :  15 - 0xf
      13'h13CE: dout <= 8'b00000011; // 5070 :   3 - 0x3
      13'h13CF: dout <= 8'b00000000; // 5071 :   0 - 0x0
      13'h13D0: dout <= 8'b00000000; // 5072 :   0 - 0x0 -- Background 0x3d
      13'h13D1: dout <= 8'b11000000; // 5073 : 192 - 0xc0
      13'h13D2: dout <= 8'b11110000; // 5074 : 240 - 0xf0
      13'h13D3: dout <= 8'b11111000; // 5075 : 248 - 0xf8
      13'h13D4: dout <= 8'b11111000; // 5076 : 248 - 0xf8
      13'h13D5: dout <= 8'b11111100; // 5077 : 252 - 0xfc
      13'h13D6: dout <= 8'b11111100; // 5078 : 252 - 0xfc
      13'h13D7: dout <= 8'b11111100; // 5079 : 252 - 0xfc
      13'h13D8: dout <= 8'b00000000; // 5080 :   0 - 0x0
      13'h13D9: dout <= 8'b11000000; // 5081 : 192 - 0xc0
      13'h13DA: dout <= 8'b11110000; // 5082 : 240 - 0xf0
      13'h13DB: dout <= 8'b11111000; // 5083 : 248 - 0xf8
      13'h13DC: dout <= 8'b11111000; // 5084 : 248 - 0xf8
      13'h13DD: dout <= 8'b11111100; // 5085 : 252 - 0xfc
      13'h13DE: dout <= 8'b11111100; // 5086 : 252 - 0xfc
      13'h13DF: dout <= 8'b11111100; // 5087 : 252 - 0xfc
      13'h13E0: dout <= 8'b00000000; // 5088 :   0 - 0x0 -- Background 0x3e
      13'h13E1: dout <= 8'b00000011; // 5089 :   3 - 0x3
      13'h13E2: dout <= 8'b00001111; // 5090 :  15 - 0xf
      13'h13E3: dout <= 8'b00111111; // 5091 :  63 - 0x3f
      13'h13E4: dout <= 8'b00111111; // 5092 :  63 - 0x3f
      13'h13E5: dout <= 8'b00011111; // 5093 :  31 - 0x1f
      13'h13E6: dout <= 8'b00000111; // 5094 :   7 - 0x7
      13'h13E7: dout <= 8'b00000000; // 5095 :   0 - 0x0
      13'h13E8: dout <= 8'b00000000; // 5096 :   0 - 0x0
      13'h13E9: dout <= 8'b00000011; // 5097 :   3 - 0x3
      13'h13EA: dout <= 8'b00001111; // 5098 :  15 - 0xf
      13'h13EB: dout <= 8'b00111111; // 5099 :  63 - 0x3f
      13'h13EC: dout <= 8'b00111111; // 5100 :  63 - 0x3f
      13'h13ED: dout <= 8'b00011111; // 5101 :  31 - 0x1f
      13'h13EE: dout <= 8'b00000111; // 5102 :   7 - 0x7
      13'h13EF: dout <= 8'b00000000; // 5103 :   0 - 0x0
      13'h13F0: dout <= 8'b11111100; // 5104 : 252 - 0xfc -- Background 0x3f
      13'h13F1: dout <= 8'b11111100; // 5105 : 252 - 0xfc
      13'h13F2: dout <= 8'b11111100; // 5106 : 252 - 0xfc
      13'h13F3: dout <= 8'b11111000; // 5107 : 248 - 0xf8
      13'h13F4: dout <= 8'b11111000; // 5108 : 248 - 0xf8
      13'h13F5: dout <= 8'b11110000; // 5109 : 240 - 0xf0
      13'h13F6: dout <= 8'b11000000; // 5110 : 192 - 0xc0
      13'h13F7: dout <= 8'b00000000; // 5111 :   0 - 0x0
      13'h13F8: dout <= 8'b11111100; // 5112 : 252 - 0xfc
      13'h13F9: dout <= 8'b11111100; // 5113 : 252 - 0xfc
      13'h13FA: dout <= 8'b11111100; // 5114 : 252 - 0xfc
      13'h13FB: dout <= 8'b11111000; // 5115 : 248 - 0xf8
      13'h13FC: dout <= 8'b11111000; // 5116 : 248 - 0xf8
      13'h13FD: dout <= 8'b11110000; // 5117 : 240 - 0xf0
      13'h13FE: dout <= 8'b11000000; // 5118 : 192 - 0xc0
      13'h13FF: dout <= 8'b00000000; // 5119 :   0 - 0x0
      13'h1400: dout <= 8'b00000000; // 5120 :   0 - 0x0 -- Background 0x40
      13'h1401: dout <= 8'b00000000; // 5121 :   0 - 0x0
      13'h1402: dout <= 8'b00000000; // 5122 :   0 - 0x0
      13'h1403: dout <= 8'b00000000; // 5123 :   0 - 0x0
      13'h1404: dout <= 8'b00000000; // 5124 :   0 - 0x0
      13'h1405: dout <= 8'b00000000; // 5125 :   0 - 0x0
      13'h1406: dout <= 8'b00000000; // 5126 :   0 - 0x0
      13'h1407: dout <= 8'b00000000; // 5127 :   0 - 0x0
      13'h1408: dout <= 8'b00000000; // 5128 :   0 - 0x0
      13'h1409: dout <= 8'b00000000; // 5129 :   0 - 0x0
      13'h140A: dout <= 8'b00000000; // 5130 :   0 - 0x0
      13'h140B: dout <= 8'b00000000; // 5131 :   0 - 0x0
      13'h140C: dout <= 8'b00000000; // 5132 :   0 - 0x0
      13'h140D: dout <= 8'b00000000; // 5133 :   0 - 0x0
      13'h140E: dout <= 8'b00000000; // 5134 :   0 - 0x0
      13'h140F: dout <= 8'b00000000; // 5135 :   0 - 0x0
      13'h1410: dout <= 8'b00011100; // 5136 :  28 - 0x1c -- Background 0x41
      13'h1411: dout <= 8'b00110110; // 5137 :  54 - 0x36
      13'h1412: dout <= 8'b01100011; // 5138 :  99 - 0x63
      13'h1413: dout <= 8'b01100011; // 5139 :  99 - 0x63
      13'h1414: dout <= 8'b01111111; // 5140 : 127 - 0x7f
      13'h1415: dout <= 8'b01100011; // 5141 :  99 - 0x63
      13'h1416: dout <= 8'b01100011; // 5142 :  99 - 0x63
      13'h1417: dout <= 8'b00000000; // 5143 :   0 - 0x0
      13'h1418: dout <= 8'b00000000; // 5144 :   0 - 0x0
      13'h1419: dout <= 8'b00000000; // 5145 :   0 - 0x0
      13'h141A: dout <= 8'b00000000; // 5146 :   0 - 0x0
      13'h141B: dout <= 8'b00000000; // 5147 :   0 - 0x0
      13'h141C: dout <= 8'b00000000; // 5148 :   0 - 0x0
      13'h141D: dout <= 8'b00000000; // 5149 :   0 - 0x0
      13'h141E: dout <= 8'b00000000; // 5150 :   0 - 0x0
      13'h141F: dout <= 8'b00000000; // 5151 :   0 - 0x0
      13'h1420: dout <= 8'b01111110; // 5152 : 126 - 0x7e -- Background 0x42
      13'h1421: dout <= 8'b01100011; // 5153 :  99 - 0x63
      13'h1422: dout <= 8'b01100011; // 5154 :  99 - 0x63
      13'h1423: dout <= 8'b01111110; // 5155 : 126 - 0x7e
      13'h1424: dout <= 8'b01100011; // 5156 :  99 - 0x63
      13'h1425: dout <= 8'b01100011; // 5157 :  99 - 0x63
      13'h1426: dout <= 8'b01111110; // 5158 : 126 - 0x7e
      13'h1427: dout <= 8'b00000000; // 5159 :   0 - 0x0
      13'h1428: dout <= 8'b00000000; // 5160 :   0 - 0x0
      13'h1429: dout <= 8'b00000000; // 5161 :   0 - 0x0
      13'h142A: dout <= 8'b00000000; // 5162 :   0 - 0x0
      13'h142B: dout <= 8'b00000000; // 5163 :   0 - 0x0
      13'h142C: dout <= 8'b00000000; // 5164 :   0 - 0x0
      13'h142D: dout <= 8'b00000000; // 5165 :   0 - 0x0
      13'h142E: dout <= 8'b00000000; // 5166 :   0 - 0x0
      13'h142F: dout <= 8'b00000000; // 5167 :   0 - 0x0
      13'h1430: dout <= 8'b00011110; // 5168 :  30 - 0x1e -- Background 0x43
      13'h1431: dout <= 8'b00110011; // 5169 :  51 - 0x33
      13'h1432: dout <= 8'b01100000; // 5170 :  96 - 0x60
      13'h1433: dout <= 8'b01100000; // 5171 :  96 - 0x60
      13'h1434: dout <= 8'b01100000; // 5172 :  96 - 0x60
      13'h1435: dout <= 8'b00110011; // 5173 :  51 - 0x33
      13'h1436: dout <= 8'b00011110; // 5174 :  30 - 0x1e
      13'h1437: dout <= 8'b00000000; // 5175 :   0 - 0x0
      13'h1438: dout <= 8'b00000000; // 5176 :   0 - 0x0
      13'h1439: dout <= 8'b00000000; // 5177 :   0 - 0x0
      13'h143A: dout <= 8'b00000000; // 5178 :   0 - 0x0
      13'h143B: dout <= 8'b00000000; // 5179 :   0 - 0x0
      13'h143C: dout <= 8'b00000000; // 5180 :   0 - 0x0
      13'h143D: dout <= 8'b00000000; // 5181 :   0 - 0x0
      13'h143E: dout <= 8'b00000000; // 5182 :   0 - 0x0
      13'h143F: dout <= 8'b00000000; // 5183 :   0 - 0x0
      13'h1440: dout <= 8'b01111100; // 5184 : 124 - 0x7c -- Background 0x44
      13'h1441: dout <= 8'b01100110; // 5185 : 102 - 0x66
      13'h1442: dout <= 8'b01100011; // 5186 :  99 - 0x63
      13'h1443: dout <= 8'b01100011; // 5187 :  99 - 0x63
      13'h1444: dout <= 8'b01100011; // 5188 :  99 - 0x63
      13'h1445: dout <= 8'b01100110; // 5189 : 102 - 0x66
      13'h1446: dout <= 8'b01111100; // 5190 : 124 - 0x7c
      13'h1447: dout <= 8'b00000000; // 5191 :   0 - 0x0
      13'h1448: dout <= 8'b00000000; // 5192 :   0 - 0x0
      13'h1449: dout <= 8'b00000000; // 5193 :   0 - 0x0
      13'h144A: dout <= 8'b00000000; // 5194 :   0 - 0x0
      13'h144B: dout <= 8'b00000000; // 5195 :   0 - 0x0
      13'h144C: dout <= 8'b00000000; // 5196 :   0 - 0x0
      13'h144D: dout <= 8'b00000000; // 5197 :   0 - 0x0
      13'h144E: dout <= 8'b00000000; // 5198 :   0 - 0x0
      13'h144F: dout <= 8'b00000000; // 5199 :   0 - 0x0
      13'h1450: dout <= 8'b01111111; // 5200 : 127 - 0x7f -- Background 0x45
      13'h1451: dout <= 8'b01100000; // 5201 :  96 - 0x60
      13'h1452: dout <= 8'b01100000; // 5202 :  96 - 0x60
      13'h1453: dout <= 8'b01111110; // 5203 : 126 - 0x7e
      13'h1454: dout <= 8'b01100000; // 5204 :  96 - 0x60
      13'h1455: dout <= 8'b01100000; // 5205 :  96 - 0x60
      13'h1456: dout <= 8'b01111111; // 5206 : 127 - 0x7f
      13'h1457: dout <= 8'b00000000; // 5207 :   0 - 0x0
      13'h1458: dout <= 8'b00000000; // 5208 :   0 - 0x0
      13'h1459: dout <= 8'b00000000; // 5209 :   0 - 0x0
      13'h145A: dout <= 8'b00000000; // 5210 :   0 - 0x0
      13'h145B: dout <= 8'b00000000; // 5211 :   0 - 0x0
      13'h145C: dout <= 8'b00000000; // 5212 :   0 - 0x0
      13'h145D: dout <= 8'b00000000; // 5213 :   0 - 0x0
      13'h145E: dout <= 8'b00000000; // 5214 :   0 - 0x0
      13'h145F: dout <= 8'b00000000; // 5215 :   0 - 0x0
      13'h1460: dout <= 8'b01111111; // 5216 : 127 - 0x7f -- Background 0x46
      13'h1461: dout <= 8'b01100000; // 5217 :  96 - 0x60
      13'h1462: dout <= 8'b01100000; // 5218 :  96 - 0x60
      13'h1463: dout <= 8'b01111110; // 5219 : 126 - 0x7e
      13'h1464: dout <= 8'b01100000; // 5220 :  96 - 0x60
      13'h1465: dout <= 8'b01100000; // 5221 :  96 - 0x60
      13'h1466: dout <= 8'b01100000; // 5222 :  96 - 0x60
      13'h1467: dout <= 8'b00000000; // 5223 :   0 - 0x0
      13'h1468: dout <= 8'b00000000; // 5224 :   0 - 0x0
      13'h1469: dout <= 8'b00000000; // 5225 :   0 - 0x0
      13'h146A: dout <= 8'b00000000; // 5226 :   0 - 0x0
      13'h146B: dout <= 8'b00000000; // 5227 :   0 - 0x0
      13'h146C: dout <= 8'b00000000; // 5228 :   0 - 0x0
      13'h146D: dout <= 8'b00000000; // 5229 :   0 - 0x0
      13'h146E: dout <= 8'b00000000; // 5230 :   0 - 0x0
      13'h146F: dout <= 8'b00000000; // 5231 :   0 - 0x0
      13'h1470: dout <= 8'b00011111; // 5232 :  31 - 0x1f -- Background 0x47
      13'h1471: dout <= 8'b00110000; // 5233 :  48 - 0x30
      13'h1472: dout <= 8'b01100000; // 5234 :  96 - 0x60
      13'h1473: dout <= 8'b01100111; // 5235 : 103 - 0x67
      13'h1474: dout <= 8'b01100011; // 5236 :  99 - 0x63
      13'h1475: dout <= 8'b00110011; // 5237 :  51 - 0x33
      13'h1476: dout <= 8'b00011111; // 5238 :  31 - 0x1f
      13'h1477: dout <= 8'b00000000; // 5239 :   0 - 0x0
      13'h1478: dout <= 8'b00000000; // 5240 :   0 - 0x0
      13'h1479: dout <= 8'b00000000; // 5241 :   0 - 0x0
      13'h147A: dout <= 8'b00000000; // 5242 :   0 - 0x0
      13'h147B: dout <= 8'b00000000; // 5243 :   0 - 0x0
      13'h147C: dout <= 8'b00000000; // 5244 :   0 - 0x0
      13'h147D: dout <= 8'b00000000; // 5245 :   0 - 0x0
      13'h147E: dout <= 8'b00000000; // 5246 :   0 - 0x0
      13'h147F: dout <= 8'b00000000; // 5247 :   0 - 0x0
      13'h1480: dout <= 8'b01100011; // 5248 :  99 - 0x63 -- Background 0x48
      13'h1481: dout <= 8'b01100011; // 5249 :  99 - 0x63
      13'h1482: dout <= 8'b01100011; // 5250 :  99 - 0x63
      13'h1483: dout <= 8'b01111111; // 5251 : 127 - 0x7f
      13'h1484: dout <= 8'b01100011; // 5252 :  99 - 0x63
      13'h1485: dout <= 8'b01100011; // 5253 :  99 - 0x63
      13'h1486: dout <= 8'b01100011; // 5254 :  99 - 0x63
      13'h1487: dout <= 8'b00000000; // 5255 :   0 - 0x0
      13'h1488: dout <= 8'b00000000; // 5256 :   0 - 0x0
      13'h1489: dout <= 8'b00000000; // 5257 :   0 - 0x0
      13'h148A: dout <= 8'b00000000; // 5258 :   0 - 0x0
      13'h148B: dout <= 8'b00000000; // 5259 :   0 - 0x0
      13'h148C: dout <= 8'b00000000; // 5260 :   0 - 0x0
      13'h148D: dout <= 8'b00000000; // 5261 :   0 - 0x0
      13'h148E: dout <= 8'b00000000; // 5262 :   0 - 0x0
      13'h148F: dout <= 8'b00000000; // 5263 :   0 - 0x0
      13'h1490: dout <= 8'b00111111; // 5264 :  63 - 0x3f -- Background 0x49
      13'h1491: dout <= 8'b00001100; // 5265 :  12 - 0xc
      13'h1492: dout <= 8'b00001100; // 5266 :  12 - 0xc
      13'h1493: dout <= 8'b00001100; // 5267 :  12 - 0xc
      13'h1494: dout <= 8'b00001100; // 5268 :  12 - 0xc
      13'h1495: dout <= 8'b00001100; // 5269 :  12 - 0xc
      13'h1496: dout <= 8'b00111111; // 5270 :  63 - 0x3f
      13'h1497: dout <= 8'b00000000; // 5271 :   0 - 0x0
      13'h1498: dout <= 8'b00000000; // 5272 :   0 - 0x0
      13'h1499: dout <= 8'b00000000; // 5273 :   0 - 0x0
      13'h149A: dout <= 8'b00000000; // 5274 :   0 - 0x0
      13'h149B: dout <= 8'b00000000; // 5275 :   0 - 0x0
      13'h149C: dout <= 8'b00000000; // 5276 :   0 - 0x0
      13'h149D: dout <= 8'b00000000; // 5277 :   0 - 0x0
      13'h149E: dout <= 8'b00000000; // 5278 :   0 - 0x0
      13'h149F: dout <= 8'b00000000; // 5279 :   0 - 0x0
      13'h14A0: dout <= 8'b00000011; // 5280 :   3 - 0x3 -- Background 0x4a
      13'h14A1: dout <= 8'b00000011; // 5281 :   3 - 0x3
      13'h14A2: dout <= 8'b00000011; // 5282 :   3 - 0x3
      13'h14A3: dout <= 8'b00000011; // 5283 :   3 - 0x3
      13'h14A4: dout <= 8'b00000011; // 5284 :   3 - 0x3
      13'h14A5: dout <= 8'b01100011; // 5285 :  99 - 0x63
      13'h14A6: dout <= 8'b00111110; // 5286 :  62 - 0x3e
      13'h14A7: dout <= 8'b00000000; // 5287 :   0 - 0x0
      13'h14A8: dout <= 8'b00000000; // 5288 :   0 - 0x0
      13'h14A9: dout <= 8'b00000000; // 5289 :   0 - 0x0
      13'h14AA: dout <= 8'b00000000; // 5290 :   0 - 0x0
      13'h14AB: dout <= 8'b00000000; // 5291 :   0 - 0x0
      13'h14AC: dout <= 8'b00000000; // 5292 :   0 - 0x0
      13'h14AD: dout <= 8'b00000000; // 5293 :   0 - 0x0
      13'h14AE: dout <= 8'b00000000; // 5294 :   0 - 0x0
      13'h14AF: dout <= 8'b00000000; // 5295 :   0 - 0x0
      13'h14B0: dout <= 8'b01100011; // 5296 :  99 - 0x63 -- Background 0x4b
      13'h14B1: dout <= 8'b01100110; // 5297 : 102 - 0x66
      13'h14B2: dout <= 8'b01101100; // 5298 : 108 - 0x6c
      13'h14B3: dout <= 8'b01111000; // 5299 : 120 - 0x78
      13'h14B4: dout <= 8'b01111100; // 5300 : 124 - 0x7c
      13'h14B5: dout <= 8'b01100110; // 5301 : 102 - 0x66
      13'h14B6: dout <= 8'b01100011; // 5302 :  99 - 0x63
      13'h14B7: dout <= 8'b00000000; // 5303 :   0 - 0x0
      13'h14B8: dout <= 8'b00000000; // 5304 :   0 - 0x0
      13'h14B9: dout <= 8'b00000000; // 5305 :   0 - 0x0
      13'h14BA: dout <= 8'b00000000; // 5306 :   0 - 0x0
      13'h14BB: dout <= 8'b00000000; // 5307 :   0 - 0x0
      13'h14BC: dout <= 8'b00000000; // 5308 :   0 - 0x0
      13'h14BD: dout <= 8'b00000000; // 5309 :   0 - 0x0
      13'h14BE: dout <= 8'b00000000; // 5310 :   0 - 0x0
      13'h14BF: dout <= 8'b00000000; // 5311 :   0 - 0x0
      13'h14C0: dout <= 8'b01100000; // 5312 :  96 - 0x60 -- Background 0x4c
      13'h14C1: dout <= 8'b01100000; // 5313 :  96 - 0x60
      13'h14C2: dout <= 8'b01100000; // 5314 :  96 - 0x60
      13'h14C3: dout <= 8'b01100000; // 5315 :  96 - 0x60
      13'h14C4: dout <= 8'b01100000; // 5316 :  96 - 0x60
      13'h14C5: dout <= 8'b01100000; // 5317 :  96 - 0x60
      13'h14C6: dout <= 8'b01111111; // 5318 : 127 - 0x7f
      13'h14C7: dout <= 8'b00000000; // 5319 :   0 - 0x0
      13'h14C8: dout <= 8'b00000000; // 5320 :   0 - 0x0
      13'h14C9: dout <= 8'b00000000; // 5321 :   0 - 0x0
      13'h14CA: dout <= 8'b00000000; // 5322 :   0 - 0x0
      13'h14CB: dout <= 8'b00000000; // 5323 :   0 - 0x0
      13'h14CC: dout <= 8'b00000000; // 5324 :   0 - 0x0
      13'h14CD: dout <= 8'b00000000; // 5325 :   0 - 0x0
      13'h14CE: dout <= 8'b00000000; // 5326 :   0 - 0x0
      13'h14CF: dout <= 8'b00000000; // 5327 :   0 - 0x0
      13'h14D0: dout <= 8'b01100011; // 5328 :  99 - 0x63 -- Background 0x4d
      13'h14D1: dout <= 8'b01110111; // 5329 : 119 - 0x77
      13'h14D2: dout <= 8'b01111111; // 5330 : 127 - 0x7f
      13'h14D3: dout <= 8'b01111111; // 5331 : 127 - 0x7f
      13'h14D4: dout <= 8'b01101011; // 5332 : 107 - 0x6b
      13'h14D5: dout <= 8'b01100011; // 5333 :  99 - 0x63
      13'h14D6: dout <= 8'b01100011; // 5334 :  99 - 0x63
      13'h14D7: dout <= 8'b00000000; // 5335 :   0 - 0x0
      13'h14D8: dout <= 8'b00000000; // 5336 :   0 - 0x0
      13'h14D9: dout <= 8'b00000000; // 5337 :   0 - 0x0
      13'h14DA: dout <= 8'b00000000; // 5338 :   0 - 0x0
      13'h14DB: dout <= 8'b00000000; // 5339 :   0 - 0x0
      13'h14DC: dout <= 8'b00000000; // 5340 :   0 - 0x0
      13'h14DD: dout <= 8'b00000000; // 5341 :   0 - 0x0
      13'h14DE: dout <= 8'b00000000; // 5342 :   0 - 0x0
      13'h14DF: dout <= 8'b00000000; // 5343 :   0 - 0x0
      13'h14E0: dout <= 8'b01100011; // 5344 :  99 - 0x63 -- Background 0x4e
      13'h14E1: dout <= 8'b01110011; // 5345 : 115 - 0x73
      13'h14E2: dout <= 8'b01111011; // 5346 : 123 - 0x7b
      13'h14E3: dout <= 8'b01111111; // 5347 : 127 - 0x7f
      13'h14E4: dout <= 8'b01101111; // 5348 : 111 - 0x6f
      13'h14E5: dout <= 8'b01100111; // 5349 : 103 - 0x67
      13'h14E6: dout <= 8'b01100011; // 5350 :  99 - 0x63
      13'h14E7: dout <= 8'b00000000; // 5351 :   0 - 0x0
      13'h14E8: dout <= 8'b00000000; // 5352 :   0 - 0x0
      13'h14E9: dout <= 8'b00000000; // 5353 :   0 - 0x0
      13'h14EA: dout <= 8'b00000000; // 5354 :   0 - 0x0
      13'h14EB: dout <= 8'b00000000; // 5355 :   0 - 0x0
      13'h14EC: dout <= 8'b00000000; // 5356 :   0 - 0x0
      13'h14ED: dout <= 8'b00000000; // 5357 :   0 - 0x0
      13'h14EE: dout <= 8'b00000000; // 5358 :   0 - 0x0
      13'h14EF: dout <= 8'b00000000; // 5359 :   0 - 0x0
      13'h14F0: dout <= 8'b00111110; // 5360 :  62 - 0x3e -- Background 0x4f
      13'h14F1: dout <= 8'b01100011; // 5361 :  99 - 0x63
      13'h14F2: dout <= 8'b01100011; // 5362 :  99 - 0x63
      13'h14F3: dout <= 8'b01100011; // 5363 :  99 - 0x63
      13'h14F4: dout <= 8'b01100011; // 5364 :  99 - 0x63
      13'h14F5: dout <= 8'b01100011; // 5365 :  99 - 0x63
      13'h14F6: dout <= 8'b00111110; // 5366 :  62 - 0x3e
      13'h14F7: dout <= 8'b00000000; // 5367 :   0 - 0x0
      13'h14F8: dout <= 8'b00000000; // 5368 :   0 - 0x0
      13'h14F9: dout <= 8'b00000000; // 5369 :   0 - 0x0
      13'h14FA: dout <= 8'b00000000; // 5370 :   0 - 0x0
      13'h14FB: dout <= 8'b00000000; // 5371 :   0 - 0x0
      13'h14FC: dout <= 8'b00000000; // 5372 :   0 - 0x0
      13'h14FD: dout <= 8'b00000000; // 5373 :   0 - 0x0
      13'h14FE: dout <= 8'b00000000; // 5374 :   0 - 0x0
      13'h14FF: dout <= 8'b00000000; // 5375 :   0 - 0x0
      13'h1500: dout <= 8'b01111110; // 5376 : 126 - 0x7e -- Background 0x50
      13'h1501: dout <= 8'b01100011; // 5377 :  99 - 0x63
      13'h1502: dout <= 8'b01100011; // 5378 :  99 - 0x63
      13'h1503: dout <= 8'b01100011; // 5379 :  99 - 0x63
      13'h1504: dout <= 8'b01111110; // 5380 : 126 - 0x7e
      13'h1505: dout <= 8'b01100000; // 5381 :  96 - 0x60
      13'h1506: dout <= 8'b01100000; // 5382 :  96 - 0x60
      13'h1507: dout <= 8'b00000000; // 5383 :   0 - 0x0
      13'h1508: dout <= 8'b00000000; // 5384 :   0 - 0x0
      13'h1509: dout <= 8'b00000000; // 5385 :   0 - 0x0
      13'h150A: dout <= 8'b00000000; // 5386 :   0 - 0x0
      13'h150B: dout <= 8'b00000000; // 5387 :   0 - 0x0
      13'h150C: dout <= 8'b00000000; // 5388 :   0 - 0x0
      13'h150D: dout <= 8'b00000000; // 5389 :   0 - 0x0
      13'h150E: dout <= 8'b00000000; // 5390 :   0 - 0x0
      13'h150F: dout <= 8'b00000000; // 5391 :   0 - 0x0
      13'h1510: dout <= 8'b00111110; // 5392 :  62 - 0x3e -- Background 0x51
      13'h1511: dout <= 8'b01100011; // 5393 :  99 - 0x63
      13'h1512: dout <= 8'b01100011; // 5394 :  99 - 0x63
      13'h1513: dout <= 8'b01100011; // 5395 :  99 - 0x63
      13'h1514: dout <= 8'b01101111; // 5396 : 111 - 0x6f
      13'h1515: dout <= 8'b01100110; // 5397 : 102 - 0x66
      13'h1516: dout <= 8'b00111101; // 5398 :  61 - 0x3d
      13'h1517: dout <= 8'b00000000; // 5399 :   0 - 0x0
      13'h1518: dout <= 8'b00000000; // 5400 :   0 - 0x0
      13'h1519: dout <= 8'b00000000; // 5401 :   0 - 0x0
      13'h151A: dout <= 8'b00000000; // 5402 :   0 - 0x0
      13'h151B: dout <= 8'b00000000; // 5403 :   0 - 0x0
      13'h151C: dout <= 8'b00000000; // 5404 :   0 - 0x0
      13'h151D: dout <= 8'b00000000; // 5405 :   0 - 0x0
      13'h151E: dout <= 8'b00000000; // 5406 :   0 - 0x0
      13'h151F: dout <= 8'b00000000; // 5407 :   0 - 0x0
      13'h1520: dout <= 8'b01111110; // 5408 : 126 - 0x7e -- Background 0x52
      13'h1521: dout <= 8'b01100011; // 5409 :  99 - 0x63
      13'h1522: dout <= 8'b01100011; // 5410 :  99 - 0x63
      13'h1523: dout <= 8'b01100111; // 5411 : 103 - 0x67
      13'h1524: dout <= 8'b01111100; // 5412 : 124 - 0x7c
      13'h1525: dout <= 8'b01101110; // 5413 : 110 - 0x6e
      13'h1526: dout <= 8'b01100111; // 5414 : 103 - 0x67
      13'h1527: dout <= 8'b00000000; // 5415 :   0 - 0x0
      13'h1528: dout <= 8'b00000000; // 5416 :   0 - 0x0
      13'h1529: dout <= 8'b00000000; // 5417 :   0 - 0x0
      13'h152A: dout <= 8'b00000000; // 5418 :   0 - 0x0
      13'h152B: dout <= 8'b00000000; // 5419 :   0 - 0x0
      13'h152C: dout <= 8'b00000000; // 5420 :   0 - 0x0
      13'h152D: dout <= 8'b00000000; // 5421 :   0 - 0x0
      13'h152E: dout <= 8'b00000000; // 5422 :   0 - 0x0
      13'h152F: dout <= 8'b00000000; // 5423 :   0 - 0x0
      13'h1530: dout <= 8'b00111100; // 5424 :  60 - 0x3c -- Background 0x53
      13'h1531: dout <= 8'b01100110; // 5425 : 102 - 0x66
      13'h1532: dout <= 8'b01100000; // 5426 :  96 - 0x60
      13'h1533: dout <= 8'b00111110; // 5427 :  62 - 0x3e
      13'h1534: dout <= 8'b00000011; // 5428 :   3 - 0x3
      13'h1535: dout <= 8'b01100011; // 5429 :  99 - 0x63
      13'h1536: dout <= 8'b00111110; // 5430 :  62 - 0x3e
      13'h1537: dout <= 8'b00000000; // 5431 :   0 - 0x0
      13'h1538: dout <= 8'b00000000; // 5432 :   0 - 0x0
      13'h1539: dout <= 8'b00000000; // 5433 :   0 - 0x0
      13'h153A: dout <= 8'b00000000; // 5434 :   0 - 0x0
      13'h153B: dout <= 8'b00000000; // 5435 :   0 - 0x0
      13'h153C: dout <= 8'b00000000; // 5436 :   0 - 0x0
      13'h153D: dout <= 8'b00000000; // 5437 :   0 - 0x0
      13'h153E: dout <= 8'b00000000; // 5438 :   0 - 0x0
      13'h153F: dout <= 8'b00000000; // 5439 :   0 - 0x0
      13'h1540: dout <= 8'b00111111; // 5440 :  63 - 0x3f -- Background 0x54
      13'h1541: dout <= 8'b00001100; // 5441 :  12 - 0xc
      13'h1542: dout <= 8'b00001100; // 5442 :  12 - 0xc
      13'h1543: dout <= 8'b00001100; // 5443 :  12 - 0xc
      13'h1544: dout <= 8'b00001100; // 5444 :  12 - 0xc
      13'h1545: dout <= 8'b00001100; // 5445 :  12 - 0xc
      13'h1546: dout <= 8'b00001100; // 5446 :  12 - 0xc
      13'h1547: dout <= 8'b00000000; // 5447 :   0 - 0x0
      13'h1548: dout <= 8'b00000000; // 5448 :   0 - 0x0
      13'h1549: dout <= 8'b00000000; // 5449 :   0 - 0x0
      13'h154A: dout <= 8'b00000000; // 5450 :   0 - 0x0
      13'h154B: dout <= 8'b00000000; // 5451 :   0 - 0x0
      13'h154C: dout <= 8'b00000000; // 5452 :   0 - 0x0
      13'h154D: dout <= 8'b00000000; // 5453 :   0 - 0x0
      13'h154E: dout <= 8'b00000000; // 5454 :   0 - 0x0
      13'h154F: dout <= 8'b00000000; // 5455 :   0 - 0x0
      13'h1550: dout <= 8'b01100011; // 5456 :  99 - 0x63 -- Background 0x55
      13'h1551: dout <= 8'b01100011; // 5457 :  99 - 0x63
      13'h1552: dout <= 8'b01100011; // 5458 :  99 - 0x63
      13'h1553: dout <= 8'b01100011; // 5459 :  99 - 0x63
      13'h1554: dout <= 8'b01100011; // 5460 :  99 - 0x63
      13'h1555: dout <= 8'b01100011; // 5461 :  99 - 0x63
      13'h1556: dout <= 8'b00111110; // 5462 :  62 - 0x3e
      13'h1557: dout <= 8'b00000000; // 5463 :   0 - 0x0
      13'h1558: dout <= 8'b00000000; // 5464 :   0 - 0x0
      13'h1559: dout <= 8'b00000000; // 5465 :   0 - 0x0
      13'h155A: dout <= 8'b00000000; // 5466 :   0 - 0x0
      13'h155B: dout <= 8'b00000000; // 5467 :   0 - 0x0
      13'h155C: dout <= 8'b00000000; // 5468 :   0 - 0x0
      13'h155D: dout <= 8'b00000000; // 5469 :   0 - 0x0
      13'h155E: dout <= 8'b00000000; // 5470 :   0 - 0x0
      13'h155F: dout <= 8'b00000000; // 5471 :   0 - 0x0
      13'h1560: dout <= 8'b01100011; // 5472 :  99 - 0x63 -- Background 0x56
      13'h1561: dout <= 8'b01100011; // 5473 :  99 - 0x63
      13'h1562: dout <= 8'b01100011; // 5474 :  99 - 0x63
      13'h1563: dout <= 8'b01110111; // 5475 : 119 - 0x77
      13'h1564: dout <= 8'b00111110; // 5476 :  62 - 0x3e
      13'h1565: dout <= 8'b00011100; // 5477 :  28 - 0x1c
      13'h1566: dout <= 8'b00001000; // 5478 :   8 - 0x8
      13'h1567: dout <= 8'b00000000; // 5479 :   0 - 0x0
      13'h1568: dout <= 8'b00000000; // 5480 :   0 - 0x0
      13'h1569: dout <= 8'b00000000; // 5481 :   0 - 0x0
      13'h156A: dout <= 8'b00000000; // 5482 :   0 - 0x0
      13'h156B: dout <= 8'b00000000; // 5483 :   0 - 0x0
      13'h156C: dout <= 8'b00000000; // 5484 :   0 - 0x0
      13'h156D: dout <= 8'b00000000; // 5485 :   0 - 0x0
      13'h156E: dout <= 8'b00000000; // 5486 :   0 - 0x0
      13'h156F: dout <= 8'b00000000; // 5487 :   0 - 0x0
      13'h1570: dout <= 8'b01100011; // 5488 :  99 - 0x63 -- Background 0x57
      13'h1571: dout <= 8'b01100011; // 5489 :  99 - 0x63
      13'h1572: dout <= 8'b01101011; // 5490 : 107 - 0x6b
      13'h1573: dout <= 8'b01111111; // 5491 : 127 - 0x7f
      13'h1574: dout <= 8'b01111111; // 5492 : 127 - 0x7f
      13'h1575: dout <= 8'b01110111; // 5493 : 119 - 0x77
      13'h1576: dout <= 8'b01100011; // 5494 :  99 - 0x63
      13'h1577: dout <= 8'b00000000; // 5495 :   0 - 0x0
      13'h1578: dout <= 8'b00000000; // 5496 :   0 - 0x0
      13'h1579: dout <= 8'b00000000; // 5497 :   0 - 0x0
      13'h157A: dout <= 8'b00000000; // 5498 :   0 - 0x0
      13'h157B: dout <= 8'b00000000; // 5499 :   0 - 0x0
      13'h157C: dout <= 8'b00000000; // 5500 :   0 - 0x0
      13'h157D: dout <= 8'b00000000; // 5501 :   0 - 0x0
      13'h157E: dout <= 8'b00000000; // 5502 :   0 - 0x0
      13'h157F: dout <= 8'b00000000; // 5503 :   0 - 0x0
      13'h1580: dout <= 8'b01100011; // 5504 :  99 - 0x63 -- Background 0x58
      13'h1581: dout <= 8'b01110111; // 5505 : 119 - 0x77
      13'h1582: dout <= 8'b00111110; // 5506 :  62 - 0x3e
      13'h1583: dout <= 8'b00011100; // 5507 :  28 - 0x1c
      13'h1584: dout <= 8'b00111110; // 5508 :  62 - 0x3e
      13'h1585: dout <= 8'b01110111; // 5509 : 119 - 0x77
      13'h1586: dout <= 8'b01100011; // 5510 :  99 - 0x63
      13'h1587: dout <= 8'b00000000; // 5511 :   0 - 0x0
      13'h1588: dout <= 8'b00000000; // 5512 :   0 - 0x0
      13'h1589: dout <= 8'b00000000; // 5513 :   0 - 0x0
      13'h158A: dout <= 8'b00000000; // 5514 :   0 - 0x0
      13'h158B: dout <= 8'b00000000; // 5515 :   0 - 0x0
      13'h158C: dout <= 8'b00000000; // 5516 :   0 - 0x0
      13'h158D: dout <= 8'b00000000; // 5517 :   0 - 0x0
      13'h158E: dout <= 8'b00000000; // 5518 :   0 - 0x0
      13'h158F: dout <= 8'b00000000; // 5519 :   0 - 0x0
      13'h1590: dout <= 8'b00110011; // 5520 :  51 - 0x33 -- Background 0x59
      13'h1591: dout <= 8'b00110011; // 5521 :  51 - 0x33
      13'h1592: dout <= 8'b00110011; // 5522 :  51 - 0x33
      13'h1593: dout <= 8'b00011110; // 5523 :  30 - 0x1e
      13'h1594: dout <= 8'b00001100; // 5524 :  12 - 0xc
      13'h1595: dout <= 8'b00001100; // 5525 :  12 - 0xc
      13'h1596: dout <= 8'b00001100; // 5526 :  12 - 0xc
      13'h1597: dout <= 8'b00000000; // 5527 :   0 - 0x0
      13'h1598: dout <= 8'b00000000; // 5528 :   0 - 0x0
      13'h1599: dout <= 8'b00000000; // 5529 :   0 - 0x0
      13'h159A: dout <= 8'b00000000; // 5530 :   0 - 0x0
      13'h159B: dout <= 8'b00000000; // 5531 :   0 - 0x0
      13'h159C: dout <= 8'b00000000; // 5532 :   0 - 0x0
      13'h159D: dout <= 8'b00000000; // 5533 :   0 - 0x0
      13'h159E: dout <= 8'b00000000; // 5534 :   0 - 0x0
      13'h159F: dout <= 8'b00000000; // 5535 :   0 - 0x0
      13'h15A0: dout <= 8'b01111111; // 5536 : 127 - 0x7f -- Background 0x5a
      13'h15A1: dout <= 8'b00000111; // 5537 :   7 - 0x7
      13'h15A2: dout <= 8'b00001110; // 5538 :  14 - 0xe
      13'h15A3: dout <= 8'b00011100; // 5539 :  28 - 0x1c
      13'h15A4: dout <= 8'b00111000; // 5540 :  56 - 0x38
      13'h15A5: dout <= 8'b01110000; // 5541 : 112 - 0x70
      13'h15A6: dout <= 8'b01111111; // 5542 : 127 - 0x7f
      13'h15A7: dout <= 8'b00000000; // 5543 :   0 - 0x0
      13'h15A8: dout <= 8'b00000000; // 5544 :   0 - 0x0
      13'h15A9: dout <= 8'b00000000; // 5545 :   0 - 0x0
      13'h15AA: dout <= 8'b00000000; // 5546 :   0 - 0x0
      13'h15AB: dout <= 8'b00000000; // 5547 :   0 - 0x0
      13'h15AC: dout <= 8'b00000000; // 5548 :   0 - 0x0
      13'h15AD: dout <= 8'b00000000; // 5549 :   0 - 0x0
      13'h15AE: dout <= 8'b00000000; // 5550 :   0 - 0x0
      13'h15AF: dout <= 8'b00000000; // 5551 :   0 - 0x0
      13'h15B0: dout <= 8'b00000000; // 5552 :   0 - 0x0 -- Background 0x5b
      13'h15B1: dout <= 8'b00000000; // 5553 :   0 - 0x0
      13'h15B2: dout <= 8'b00000000; // 5554 :   0 - 0x0
      13'h15B3: dout <= 8'b00000000; // 5555 :   0 - 0x0
      13'h15B4: dout <= 8'b00000000; // 5556 :   0 - 0x0
      13'h15B5: dout <= 8'b00110000; // 5557 :  48 - 0x30
      13'h15B6: dout <= 8'b00110000; // 5558 :  48 - 0x30
      13'h15B7: dout <= 8'b00000000; // 5559 :   0 - 0x0
      13'h15B8: dout <= 8'b00000000; // 5560 :   0 - 0x0
      13'h15B9: dout <= 8'b00000000; // 5561 :   0 - 0x0
      13'h15BA: dout <= 8'b00000000; // 5562 :   0 - 0x0
      13'h15BB: dout <= 8'b00000000; // 5563 :   0 - 0x0
      13'h15BC: dout <= 8'b00000000; // 5564 :   0 - 0x0
      13'h15BD: dout <= 8'b00000000; // 5565 :   0 - 0x0
      13'h15BE: dout <= 8'b00000000; // 5566 :   0 - 0x0
      13'h15BF: dout <= 8'b00000000; // 5567 :   0 - 0x0
      13'h15C0: dout <= 8'b11000000; // 5568 : 192 - 0xc0 -- Background 0x5c
      13'h15C1: dout <= 8'b11110000; // 5569 : 240 - 0xf0
      13'h15C2: dout <= 8'b11111100; // 5570 : 252 - 0xfc
      13'h15C3: dout <= 8'b11111111; // 5571 : 255 - 0xff
      13'h15C4: dout <= 8'b11111100; // 5572 : 252 - 0xfc
      13'h15C5: dout <= 8'b11110000; // 5573 : 240 - 0xf0
      13'h15C6: dout <= 8'b11000000; // 5574 : 192 - 0xc0
      13'h15C7: dout <= 8'b00000000; // 5575 :   0 - 0x0
      13'h15C8: dout <= 8'b00000000; // 5576 :   0 - 0x0
      13'h15C9: dout <= 8'b00000000; // 5577 :   0 - 0x0
      13'h15CA: dout <= 8'b00000000; // 5578 :   0 - 0x0
      13'h15CB: dout <= 8'b00000000; // 5579 :   0 - 0x0
      13'h15CC: dout <= 8'b00000000; // 5580 :   0 - 0x0
      13'h15CD: dout <= 8'b00000000; // 5581 :   0 - 0x0
      13'h15CE: dout <= 8'b00000000; // 5582 :   0 - 0x0
      13'h15CF: dout <= 8'b00000000; // 5583 :   0 - 0x0
      13'h15D0: dout <= 8'b00111100; // 5584 :  60 - 0x3c -- Background 0x5d
      13'h15D1: dout <= 8'b01000010; // 5585 :  66 - 0x42
      13'h15D2: dout <= 8'b10011001; // 5586 : 153 - 0x99
      13'h15D3: dout <= 8'b10100001; // 5587 : 161 - 0xa1
      13'h15D4: dout <= 8'b10100001; // 5588 : 161 - 0xa1
      13'h15D5: dout <= 8'b10011001; // 5589 : 153 - 0x99
      13'h15D6: dout <= 8'b01000010; // 5590 :  66 - 0x42
      13'h15D7: dout <= 8'b00111100; // 5591 :  60 - 0x3c
      13'h15D8: dout <= 8'b00000000; // 5592 :   0 - 0x0
      13'h15D9: dout <= 8'b00000000; // 5593 :   0 - 0x0
      13'h15DA: dout <= 8'b00000000; // 5594 :   0 - 0x0
      13'h15DB: dout <= 8'b00000000; // 5595 :   0 - 0x0
      13'h15DC: dout <= 8'b00000000; // 5596 :   0 - 0x0
      13'h15DD: dout <= 8'b00000000; // 5597 :   0 - 0x0
      13'h15DE: dout <= 8'b00000000; // 5598 :   0 - 0x0
      13'h15DF: dout <= 8'b00000000; // 5599 :   0 - 0x0
      13'h15E0: dout <= 8'b00000000; // 5600 :   0 - 0x0 -- Background 0x5e
      13'h15E1: dout <= 8'b00000000; // 5601 :   0 - 0x0
      13'h15E2: dout <= 8'b00010000; // 5602 :  16 - 0x10
      13'h15E3: dout <= 8'b00010000; // 5603 :  16 - 0x10
      13'h15E4: dout <= 8'b00010000; // 5604 :  16 - 0x10
      13'h15E5: dout <= 8'b00010000; // 5605 :  16 - 0x10
      13'h15E6: dout <= 8'b00000000; // 5606 :   0 - 0x0
      13'h15E7: dout <= 8'b00000000; // 5607 :   0 - 0x0
      13'h15E8: dout <= 8'b00000000; // 5608 :   0 - 0x0
      13'h15E9: dout <= 8'b00000000; // 5609 :   0 - 0x0
      13'h15EA: dout <= 8'b00010000; // 5610 :  16 - 0x10
      13'h15EB: dout <= 8'b00010000; // 5611 :  16 - 0x10
      13'h15EC: dout <= 8'b00010000; // 5612 :  16 - 0x10
      13'h15ED: dout <= 8'b00010000; // 5613 :  16 - 0x10
      13'h15EE: dout <= 8'b00000000; // 5614 :   0 - 0x0
      13'h15EF: dout <= 8'b00000000; // 5615 :   0 - 0x0
      13'h15F0: dout <= 8'b00110110; // 5616 :  54 - 0x36 -- Background 0x5f
      13'h15F1: dout <= 8'b00110110; // 5617 :  54 - 0x36
      13'h15F2: dout <= 8'b00010010; // 5618 :  18 - 0x12
      13'h15F3: dout <= 8'b00000000; // 5619 :   0 - 0x0
      13'h15F4: dout <= 8'b00000000; // 5620 :   0 - 0x0
      13'h15F5: dout <= 8'b00000000; // 5621 :   0 - 0x0
      13'h15F6: dout <= 8'b00000000; // 5622 :   0 - 0x0
      13'h15F7: dout <= 8'b00000000; // 5623 :   0 - 0x0
      13'h15F8: dout <= 8'b00000000; // 5624 :   0 - 0x0
      13'h15F9: dout <= 8'b00000000; // 5625 :   0 - 0x0
      13'h15FA: dout <= 8'b00000000; // 5626 :   0 - 0x0
      13'h15FB: dout <= 8'b00000000; // 5627 :   0 - 0x0
      13'h15FC: dout <= 8'b00000000; // 5628 :   0 - 0x0
      13'h15FD: dout <= 8'b00000000; // 5629 :   0 - 0x0
      13'h15FE: dout <= 8'b00000000; // 5630 :   0 - 0x0
      13'h15FF: dout <= 8'b00000000; // 5631 :   0 - 0x0
      13'h1600: dout <= 8'b00000000; // 5632 :   0 - 0x0 -- Background 0x60
      13'h1601: dout <= 8'b00000000; // 5633 :   0 - 0x0
      13'h1602: dout <= 8'b00000000; // 5634 :   0 - 0x0
      13'h1603: dout <= 8'b00000000; // 5635 :   0 - 0x0
      13'h1604: dout <= 8'b00000000; // 5636 :   0 - 0x0
      13'h1605: dout <= 8'b00000001; // 5637 :   1 - 0x1
      13'h1606: dout <= 8'b00011110; // 5638 :  30 - 0x1e
      13'h1607: dout <= 8'b00111011; // 5639 :  59 - 0x3b
      13'h1608: dout <= 8'b00000000; // 5640 :   0 - 0x0
      13'h1609: dout <= 8'b00000000; // 5641 :   0 - 0x0
      13'h160A: dout <= 8'b00000000; // 5642 :   0 - 0x0
      13'h160B: dout <= 8'b00000000; // 5643 :   0 - 0x0
      13'h160C: dout <= 8'b00000000; // 5644 :   0 - 0x0
      13'h160D: dout <= 8'b00000000; // 5645 :   0 - 0x0
      13'h160E: dout <= 8'b00000000; // 5646 :   0 - 0x0
      13'h160F: dout <= 8'b00000000; // 5647 :   0 - 0x0
      13'h1610: dout <= 8'b00000000; // 5648 :   0 - 0x0 -- Background 0x61
      13'h1611: dout <= 8'b00000000; // 5649 :   0 - 0x0
      13'h1612: dout <= 8'b00001100; // 5650 :  12 - 0xc
      13'h1613: dout <= 8'b00111100; // 5651 :  60 - 0x3c
      13'h1614: dout <= 8'b11010000; // 5652 : 208 - 0xd0
      13'h1615: dout <= 8'b00010000; // 5653 :  16 - 0x10
      13'h1616: dout <= 8'b00100000; // 5654 :  32 - 0x20
      13'h1617: dout <= 8'b01000000; // 5655 :  64 - 0x40
      13'h1618: dout <= 8'b00000000; // 5656 :   0 - 0x0
      13'h1619: dout <= 8'b00000000; // 5657 :   0 - 0x0
      13'h161A: dout <= 8'b00000000; // 5658 :   0 - 0x0
      13'h161B: dout <= 8'b00000000; // 5659 :   0 - 0x0
      13'h161C: dout <= 8'b00000000; // 5660 :   0 - 0x0
      13'h161D: dout <= 8'b00000000; // 5661 :   0 - 0x0
      13'h161E: dout <= 8'b00000000; // 5662 :   0 - 0x0
      13'h161F: dout <= 8'b00000000; // 5663 :   0 - 0x0
      13'h1620: dout <= 8'b00111110; // 5664 :  62 - 0x3e -- Background 0x62
      13'h1621: dout <= 8'b00101101; // 5665 :  45 - 0x2d
      13'h1622: dout <= 8'b00110101; // 5666 :  53 - 0x35
      13'h1623: dout <= 8'b00011101; // 5667 :  29 - 0x1d
      13'h1624: dout <= 8'b00000001; // 5668 :   1 - 0x1
      13'h1625: dout <= 8'b00000000; // 5669 :   0 - 0x0
      13'h1626: dout <= 8'b00000000; // 5670 :   0 - 0x0
      13'h1627: dout <= 8'b00000000; // 5671 :   0 - 0x0
      13'h1628: dout <= 8'b00000000; // 5672 :   0 - 0x0
      13'h1629: dout <= 8'b00000000; // 5673 :   0 - 0x0
      13'h162A: dout <= 8'b00000000; // 5674 :   0 - 0x0
      13'h162B: dout <= 8'b00000000; // 5675 :   0 - 0x0
      13'h162C: dout <= 8'b00000000; // 5676 :   0 - 0x0
      13'h162D: dout <= 8'b00000000; // 5677 :   0 - 0x0
      13'h162E: dout <= 8'b00000000; // 5678 :   0 - 0x0
      13'h162F: dout <= 8'b00000000; // 5679 :   0 - 0x0
      13'h1630: dout <= 8'b10110000; // 5680 : 176 - 0xb0 -- Background 0x63
      13'h1631: dout <= 8'b10111000; // 5681 : 184 - 0xb8
      13'h1632: dout <= 8'b11111000; // 5682 : 248 - 0xf8
      13'h1633: dout <= 8'b01111000; // 5683 : 120 - 0x78
      13'h1634: dout <= 8'b10011000; // 5684 : 152 - 0x98
      13'h1635: dout <= 8'b11110000; // 5685 : 240 - 0xf0
      13'h1636: dout <= 8'b00000000; // 5686 :   0 - 0x0
      13'h1637: dout <= 8'b00000000; // 5687 :   0 - 0x0
      13'h1638: dout <= 8'b00000000; // 5688 :   0 - 0x0
      13'h1639: dout <= 8'b00000000; // 5689 :   0 - 0x0
      13'h163A: dout <= 8'b00000000; // 5690 :   0 - 0x0
      13'h163B: dout <= 8'b00000000; // 5691 :   0 - 0x0
      13'h163C: dout <= 8'b00000000; // 5692 :   0 - 0x0
      13'h163D: dout <= 8'b00000000; // 5693 :   0 - 0x0
      13'h163E: dout <= 8'b00000000; // 5694 :   0 - 0x0
      13'h163F: dout <= 8'b00000000; // 5695 :   0 - 0x0
      13'h1640: dout <= 8'b00000000; // 5696 :   0 - 0x0 -- Background 0x64
      13'h1641: dout <= 8'b00000000; // 5697 :   0 - 0x0
      13'h1642: dout <= 8'b00000111; // 5698 :   7 - 0x7
      13'h1643: dout <= 8'b00000011; // 5699 :   3 - 0x3
      13'h1644: dout <= 8'b00001101; // 5700 :  13 - 0xd
      13'h1645: dout <= 8'b00011110; // 5701 :  30 - 0x1e
      13'h1646: dout <= 8'b00010111; // 5702 :  23 - 0x17
      13'h1647: dout <= 8'b00011101; // 5703 :  29 - 0x1d
      13'h1648: dout <= 8'b00000000; // 5704 :   0 - 0x0
      13'h1649: dout <= 8'b00000000; // 5705 :   0 - 0x0
      13'h164A: dout <= 8'b00000000; // 5706 :   0 - 0x0
      13'h164B: dout <= 8'b00000000; // 5707 :   0 - 0x0
      13'h164C: dout <= 8'b00000000; // 5708 :   0 - 0x0
      13'h164D: dout <= 8'b00000000; // 5709 :   0 - 0x0
      13'h164E: dout <= 8'b00000000; // 5710 :   0 - 0x0
      13'h164F: dout <= 8'b00000000; // 5711 :   0 - 0x0
      13'h1650: dout <= 8'b00000000; // 5712 :   0 - 0x0 -- Background 0x65
      13'h1651: dout <= 8'b10000000; // 5713 : 128 - 0x80
      13'h1652: dout <= 8'b01110000; // 5714 : 112 - 0x70
      13'h1653: dout <= 8'b11100000; // 5715 : 224 - 0xe0
      13'h1654: dout <= 8'b11011000; // 5716 : 216 - 0xd8
      13'h1655: dout <= 8'b10111100; // 5717 : 188 - 0xbc
      13'h1656: dout <= 8'b01110100; // 5718 : 116 - 0x74
      13'h1657: dout <= 8'b11011100; // 5719 : 220 - 0xdc
      13'h1658: dout <= 8'b00000000; // 5720 :   0 - 0x0
      13'h1659: dout <= 8'b00000000; // 5721 :   0 - 0x0
      13'h165A: dout <= 8'b00000000; // 5722 :   0 - 0x0
      13'h165B: dout <= 8'b00000000; // 5723 :   0 - 0x0
      13'h165C: dout <= 8'b00000000; // 5724 :   0 - 0x0
      13'h165D: dout <= 8'b00000000; // 5725 :   0 - 0x0
      13'h165E: dout <= 8'b00000000; // 5726 :   0 - 0x0
      13'h165F: dout <= 8'b00000000; // 5727 :   0 - 0x0
      13'h1660: dout <= 8'b00011111; // 5728 :  31 - 0x1f -- Background 0x66
      13'h1661: dout <= 8'b00001011; // 5729 :  11 - 0xb
      13'h1662: dout <= 8'b00001111; // 5730 :  15 - 0xf
      13'h1663: dout <= 8'b00000101; // 5731 :   5 - 0x5
      13'h1664: dout <= 8'b00000011; // 5732 :   3 - 0x3
      13'h1665: dout <= 8'b00000001; // 5733 :   1 - 0x1
      13'h1666: dout <= 8'b00000000; // 5734 :   0 - 0x0
      13'h1667: dout <= 8'b00000000; // 5735 :   0 - 0x0
      13'h1668: dout <= 8'b00000000; // 5736 :   0 - 0x0
      13'h1669: dout <= 8'b00000000; // 5737 :   0 - 0x0
      13'h166A: dout <= 8'b00000000; // 5738 :   0 - 0x0
      13'h166B: dout <= 8'b00000000; // 5739 :   0 - 0x0
      13'h166C: dout <= 8'b00000000; // 5740 :   0 - 0x0
      13'h166D: dout <= 8'b00000000; // 5741 :   0 - 0x0
      13'h166E: dout <= 8'b00000000; // 5742 :   0 - 0x0
      13'h166F: dout <= 8'b00000000; // 5743 :   0 - 0x0
      13'h1670: dout <= 8'b11111100; // 5744 : 252 - 0xfc -- Background 0x67
      13'h1671: dout <= 8'b01101000; // 5745 : 104 - 0x68
      13'h1672: dout <= 8'b11111000; // 5746 : 248 - 0xf8
      13'h1673: dout <= 8'b10110000; // 5747 : 176 - 0xb0
      13'h1674: dout <= 8'b11100000; // 5748 : 224 - 0xe0
      13'h1675: dout <= 8'b10000000; // 5749 : 128 - 0x80
      13'h1676: dout <= 8'b00000000; // 5750 :   0 - 0x0
      13'h1677: dout <= 8'b00000000; // 5751 :   0 - 0x0
      13'h1678: dout <= 8'b00000000; // 5752 :   0 - 0x0
      13'h1679: dout <= 8'b00000000; // 5753 :   0 - 0x0
      13'h167A: dout <= 8'b00000000; // 5754 :   0 - 0x0
      13'h167B: dout <= 8'b00000000; // 5755 :   0 - 0x0
      13'h167C: dout <= 8'b00000000; // 5756 :   0 - 0x0
      13'h167D: dout <= 8'b00000000; // 5757 :   0 - 0x0
      13'h167E: dout <= 8'b00000000; // 5758 :   0 - 0x0
      13'h167F: dout <= 8'b00000000; // 5759 :   0 - 0x0
      13'h1680: dout <= 8'b00000000; // 5760 :   0 - 0x0 -- Background 0x68
      13'h1681: dout <= 8'b00000000; // 5761 :   0 - 0x0
      13'h1682: dout <= 8'b00000000; // 5762 :   0 - 0x0
      13'h1683: dout <= 8'b00000000; // 5763 :   0 - 0x0
      13'h1684: dout <= 8'b00000000; // 5764 :   0 - 0x0
      13'h1685: dout <= 8'b00000000; // 5765 :   0 - 0x0
      13'h1686: dout <= 8'b00000000; // 5766 :   0 - 0x0
      13'h1687: dout <= 8'b00000000; // 5767 :   0 - 0x0
      13'h1688: dout <= 8'b00000000; // 5768 :   0 - 0x0
      13'h1689: dout <= 8'b00000000; // 5769 :   0 - 0x0
      13'h168A: dout <= 8'b00000000; // 5770 :   0 - 0x0
      13'h168B: dout <= 8'b00000001; // 5771 :   1 - 0x1
      13'h168C: dout <= 8'b00000001; // 5772 :   1 - 0x1
      13'h168D: dout <= 8'b00001011; // 5773 :  11 - 0xb
      13'h168E: dout <= 8'b00011100; // 5774 :  28 - 0x1c
      13'h168F: dout <= 8'b00111111; // 5775 :  63 - 0x3f
      13'h1690: dout <= 8'b00000000; // 5776 :   0 - 0x0 -- Background 0x69
      13'h1691: dout <= 8'b00000000; // 5777 :   0 - 0x0
      13'h1692: dout <= 8'b00000000; // 5778 :   0 - 0x0
      13'h1693: dout <= 8'b00000000; // 5779 :   0 - 0x0
      13'h1694: dout <= 8'b00000000; // 5780 :   0 - 0x0
      13'h1695: dout <= 8'b00000000; // 5781 :   0 - 0x0
      13'h1696: dout <= 8'b00000000; // 5782 :   0 - 0x0
      13'h1697: dout <= 8'b00000000; // 5783 :   0 - 0x0
      13'h1698: dout <= 8'b00000000; // 5784 :   0 - 0x0
      13'h1699: dout <= 8'b00000000; // 5785 :   0 - 0x0
      13'h169A: dout <= 8'b00110000; // 5786 :  48 - 0x30
      13'h169B: dout <= 8'b01111000; // 5787 : 120 - 0x78
      13'h169C: dout <= 8'b10000000; // 5788 : 128 - 0x80
      13'h169D: dout <= 8'b11110000; // 5789 : 240 - 0xf0
      13'h169E: dout <= 8'b11111000; // 5790 : 248 - 0xf8
      13'h169F: dout <= 8'b11111100; // 5791 : 252 - 0xfc
      13'h16A0: dout <= 8'b00000000; // 5792 :   0 - 0x0 -- Background 0x6a
      13'h16A1: dout <= 8'b00000000; // 5793 :   0 - 0x0
      13'h16A2: dout <= 8'b00000000; // 5794 :   0 - 0x0
      13'h16A3: dout <= 8'b00000000; // 5795 :   0 - 0x0
      13'h16A4: dout <= 8'b00000000; // 5796 :   0 - 0x0
      13'h16A5: dout <= 8'b00000000; // 5797 :   0 - 0x0
      13'h16A6: dout <= 8'b00000000; // 5798 :   0 - 0x0
      13'h16A7: dout <= 8'b00000000; // 5799 :   0 - 0x0
      13'h16A8: dout <= 8'b00111111; // 5800 :  63 - 0x3f
      13'h16A9: dout <= 8'b00111111; // 5801 :  63 - 0x3f
      13'h16AA: dout <= 8'b00111111; // 5802 :  63 - 0x3f
      13'h16AB: dout <= 8'b00011111; // 5803 :  31 - 0x1f
      13'h16AC: dout <= 8'b00011111; // 5804 :  31 - 0x1f
      13'h16AD: dout <= 8'b00000111; // 5805 :   7 - 0x7
      13'h16AE: dout <= 8'b00000000; // 5806 :   0 - 0x0
      13'h16AF: dout <= 8'b00000000; // 5807 :   0 - 0x0
      13'h16B0: dout <= 8'b00000000; // 5808 :   0 - 0x0 -- Background 0x6b
      13'h16B1: dout <= 8'b00000000; // 5809 :   0 - 0x0
      13'h16B2: dout <= 8'b00000000; // 5810 :   0 - 0x0
      13'h16B3: dout <= 8'b00000000; // 5811 :   0 - 0x0
      13'h16B4: dout <= 8'b00000000; // 5812 :   0 - 0x0
      13'h16B5: dout <= 8'b00000000; // 5813 :   0 - 0x0
      13'h16B6: dout <= 8'b00000000; // 5814 :   0 - 0x0
      13'h16B7: dout <= 8'b00000000; // 5815 :   0 - 0x0
      13'h16B8: dout <= 8'b11111100; // 5816 : 252 - 0xfc
      13'h16B9: dout <= 8'b11101100; // 5817 : 236 - 0xec
      13'h16BA: dout <= 8'b11101100; // 5818 : 236 - 0xec
      13'h16BB: dout <= 8'b11011000; // 5819 : 216 - 0xd8
      13'h16BC: dout <= 8'b11111000; // 5820 : 248 - 0xf8
      13'h16BD: dout <= 8'b11100000; // 5821 : 224 - 0xe0
      13'h16BE: dout <= 8'b00000000; // 5822 :   0 - 0x0
      13'h16BF: dout <= 8'b00000000; // 5823 :   0 - 0x0
      13'h16C0: dout <= 8'b00000000; // 5824 :   0 - 0x0 -- Background 0x6c
      13'h16C1: dout <= 8'b00000000; // 5825 :   0 - 0x0
      13'h16C2: dout <= 8'b00000001; // 5826 :   1 - 0x1
      13'h16C3: dout <= 8'b00011101; // 5827 :  29 - 0x1d
      13'h16C4: dout <= 8'b00111110; // 5828 :  62 - 0x3e
      13'h16C5: dout <= 8'b00111111; // 5829 :  63 - 0x3f
      13'h16C6: dout <= 8'b00111111; // 5830 :  63 - 0x3f
      13'h16C7: dout <= 8'b00111111; // 5831 :  63 - 0x3f
      13'h16C8: dout <= 8'b00000000; // 5832 :   0 - 0x0
      13'h16C9: dout <= 8'b00000000; // 5833 :   0 - 0x0
      13'h16CA: dout <= 8'b00000001; // 5834 :   1 - 0x1
      13'h16CB: dout <= 8'b00011101; // 5835 :  29 - 0x1d
      13'h16CC: dout <= 8'b00111110; // 5836 :  62 - 0x3e
      13'h16CD: dout <= 8'b00111111; // 5837 :  63 - 0x3f
      13'h16CE: dout <= 8'b00111111; // 5838 :  63 - 0x3f
      13'h16CF: dout <= 8'b00111111; // 5839 :  63 - 0x3f
      13'h16D0: dout <= 8'b00000000; // 5840 :   0 - 0x0 -- Background 0x6d
      13'h16D1: dout <= 8'b10000000; // 5841 : 128 - 0x80
      13'h16D2: dout <= 8'b00000000; // 5842 :   0 - 0x0
      13'h16D3: dout <= 8'b01110000; // 5843 : 112 - 0x70
      13'h16D4: dout <= 8'b11111000; // 5844 : 248 - 0xf8
      13'h16D5: dout <= 8'b11111100; // 5845 : 252 - 0xfc
      13'h16D6: dout <= 8'b11111100; // 5846 : 252 - 0xfc
      13'h16D7: dout <= 8'b11111100; // 5847 : 252 - 0xfc
      13'h16D8: dout <= 8'b00000000; // 5848 :   0 - 0x0
      13'h16D9: dout <= 8'b10000000; // 5849 : 128 - 0x80
      13'h16DA: dout <= 8'b00000000; // 5850 :   0 - 0x0
      13'h16DB: dout <= 8'b01110000; // 5851 : 112 - 0x70
      13'h16DC: dout <= 8'b11111000; // 5852 : 248 - 0xf8
      13'h16DD: dout <= 8'b11111100; // 5853 : 252 - 0xfc
      13'h16DE: dout <= 8'b11111100; // 5854 : 252 - 0xfc
      13'h16DF: dout <= 8'b11111100; // 5855 : 252 - 0xfc
      13'h16E0: dout <= 8'b00111111; // 5856 :  63 - 0x3f -- Background 0x6e
      13'h16E1: dout <= 8'b00111111; // 5857 :  63 - 0x3f
      13'h16E2: dout <= 8'b00011111; // 5858 :  31 - 0x1f
      13'h16E3: dout <= 8'b00011111; // 5859 :  31 - 0x1f
      13'h16E4: dout <= 8'b00001111; // 5860 :  15 - 0xf
      13'h16E5: dout <= 8'b00000110; // 5861 :   6 - 0x6
      13'h16E6: dout <= 8'b00000000; // 5862 :   0 - 0x0
      13'h16E7: dout <= 8'b00000000; // 5863 :   0 - 0x0
      13'h16E8: dout <= 8'b00111111; // 5864 :  63 - 0x3f
      13'h16E9: dout <= 8'b00111111; // 5865 :  63 - 0x3f
      13'h16EA: dout <= 8'b00011111; // 5866 :  31 - 0x1f
      13'h16EB: dout <= 8'b00011111; // 5867 :  31 - 0x1f
      13'h16EC: dout <= 8'b00001111; // 5868 :  15 - 0xf
      13'h16ED: dout <= 8'b00000110; // 5869 :   6 - 0x6
      13'h16EE: dout <= 8'b00000000; // 5870 :   0 - 0x0
      13'h16EF: dout <= 8'b00000000; // 5871 :   0 - 0x0
      13'h16F0: dout <= 8'b11101100; // 5872 : 236 - 0xec -- Background 0x6f
      13'h16F1: dout <= 8'b11101100; // 5873 : 236 - 0xec
      13'h16F2: dout <= 8'b11011000; // 5874 : 216 - 0xd8
      13'h16F3: dout <= 8'b11111000; // 5875 : 248 - 0xf8
      13'h16F4: dout <= 8'b11110000; // 5876 : 240 - 0xf0
      13'h16F5: dout <= 8'b11100000; // 5877 : 224 - 0xe0
      13'h16F6: dout <= 8'b00000000; // 5878 :   0 - 0x0
      13'h16F7: dout <= 8'b00000000; // 5879 :   0 - 0x0
      13'h16F8: dout <= 8'b11101100; // 5880 : 236 - 0xec
      13'h16F9: dout <= 8'b11101100; // 5881 : 236 - 0xec
      13'h16FA: dout <= 8'b11011000; // 5882 : 216 - 0xd8
      13'h16FB: dout <= 8'b11111000; // 5883 : 248 - 0xf8
      13'h16FC: dout <= 8'b11110000; // 5884 : 240 - 0xf0
      13'h16FD: dout <= 8'b11100000; // 5885 : 224 - 0xe0
      13'h16FE: dout <= 8'b00000000; // 5886 :   0 - 0x0
      13'h16FF: dout <= 8'b00000000; // 5887 :   0 - 0x0
      13'h1700: dout <= 8'b00000000; // 5888 :   0 - 0x0 -- Background 0x70
      13'h1701: dout <= 8'b00000100; // 5889 :   4 - 0x4
      13'h1702: dout <= 8'b00000011; // 5890 :   3 - 0x3
      13'h1703: dout <= 8'b00000000; // 5891 :   0 - 0x0
      13'h1704: dout <= 8'b00000001; // 5892 :   1 - 0x1
      13'h1705: dout <= 8'b00000111; // 5893 :   7 - 0x7
      13'h1706: dout <= 8'b00001111; // 5894 :  15 - 0xf
      13'h1707: dout <= 8'b00001100; // 5895 :  12 - 0xc
      13'h1708: dout <= 8'b00000000; // 5896 :   0 - 0x0
      13'h1709: dout <= 8'b00000000; // 5897 :   0 - 0x0
      13'h170A: dout <= 8'b00000000; // 5898 :   0 - 0x0
      13'h170B: dout <= 8'b00000000; // 5899 :   0 - 0x0
      13'h170C: dout <= 8'b00000000; // 5900 :   0 - 0x0
      13'h170D: dout <= 8'b00000000; // 5901 :   0 - 0x0
      13'h170E: dout <= 8'b00000000; // 5902 :   0 - 0x0
      13'h170F: dout <= 8'b00000000; // 5903 :   0 - 0x0
      13'h1710: dout <= 8'b00000000; // 5904 :   0 - 0x0 -- Background 0x71
      13'h1711: dout <= 8'b00000000; // 5905 :   0 - 0x0
      13'h1712: dout <= 8'b11100000; // 5906 : 224 - 0xe0
      13'h1713: dout <= 8'b10000000; // 5907 : 128 - 0x80
      13'h1714: dout <= 8'b01000000; // 5908 :  64 - 0x40
      13'h1715: dout <= 8'b11110000; // 5909 : 240 - 0xf0
      13'h1716: dout <= 8'b10011000; // 5910 : 152 - 0x98
      13'h1717: dout <= 8'b11111000; // 5911 : 248 - 0xf8
      13'h1718: dout <= 8'b00000000; // 5912 :   0 - 0x0
      13'h1719: dout <= 8'b00000000; // 5913 :   0 - 0x0
      13'h171A: dout <= 8'b00000000; // 5914 :   0 - 0x0
      13'h171B: dout <= 8'b00000000; // 5915 :   0 - 0x0
      13'h171C: dout <= 8'b00000000; // 5916 :   0 - 0x0
      13'h171D: dout <= 8'b00000000; // 5917 :   0 - 0x0
      13'h171E: dout <= 8'b00000000; // 5918 :   0 - 0x0
      13'h171F: dout <= 8'b00000000; // 5919 :   0 - 0x0
      13'h1720: dout <= 8'b00011111; // 5920 :  31 - 0x1f -- Background 0x72
      13'h1721: dout <= 8'b00010011; // 5921 :  19 - 0x13
      13'h1722: dout <= 8'b00011111; // 5922 :  31 - 0x1f
      13'h1723: dout <= 8'b00001111; // 5923 :  15 - 0xf
      13'h1724: dout <= 8'b00001001; // 5924 :   9 - 0x9
      13'h1725: dout <= 8'b00000111; // 5925 :   7 - 0x7
      13'h1726: dout <= 8'b00000001; // 5926 :   1 - 0x1
      13'h1727: dout <= 8'b00000000; // 5927 :   0 - 0x0
      13'h1728: dout <= 8'b00000000; // 5928 :   0 - 0x0
      13'h1729: dout <= 8'b00000000; // 5929 :   0 - 0x0
      13'h172A: dout <= 8'b00000000; // 5930 :   0 - 0x0
      13'h172B: dout <= 8'b00000000; // 5931 :   0 - 0x0
      13'h172C: dout <= 8'b00000000; // 5932 :   0 - 0x0
      13'h172D: dout <= 8'b00000000; // 5933 :   0 - 0x0
      13'h172E: dout <= 8'b00000000; // 5934 :   0 - 0x0
      13'h172F: dout <= 8'b00000000; // 5935 :   0 - 0x0
      13'h1730: dout <= 8'b11100100; // 5936 : 228 - 0xe4 -- Background 0x73
      13'h1731: dout <= 8'b00111100; // 5937 :  60 - 0x3c
      13'h1732: dout <= 8'b11100100; // 5938 : 228 - 0xe4
      13'h1733: dout <= 8'b00111000; // 5939 :  56 - 0x38
      13'h1734: dout <= 8'b11111000; // 5940 : 248 - 0xf8
      13'h1735: dout <= 8'b11110000; // 5941 : 240 - 0xf0
      13'h1736: dout <= 8'b11000000; // 5942 : 192 - 0xc0
      13'h1737: dout <= 8'b00000000; // 5943 :   0 - 0x0
      13'h1738: dout <= 8'b00000000; // 5944 :   0 - 0x0
      13'h1739: dout <= 8'b00000000; // 5945 :   0 - 0x0
      13'h173A: dout <= 8'b00000000; // 5946 :   0 - 0x0
      13'h173B: dout <= 8'b00000000; // 5947 :   0 - 0x0
      13'h173C: dout <= 8'b00000000; // 5948 :   0 - 0x0
      13'h173D: dout <= 8'b00000000; // 5949 :   0 - 0x0
      13'h173E: dout <= 8'b00000000; // 5950 :   0 - 0x0
      13'h173F: dout <= 8'b00000000; // 5951 :   0 - 0x0
      13'h1740: dout <= 8'b00000000; // 5952 :   0 - 0x0 -- Background 0x74
      13'h1741: dout <= 8'b00000000; // 5953 :   0 - 0x0
      13'h1742: dout <= 8'b00000000; // 5954 :   0 - 0x0
      13'h1743: dout <= 8'b00000000; // 5955 :   0 - 0x0
      13'h1744: dout <= 8'b00000000; // 5956 :   0 - 0x0
      13'h1745: dout <= 8'b00000000; // 5957 :   0 - 0x0
      13'h1746: dout <= 8'b00000000; // 5958 :   0 - 0x0
      13'h1747: dout <= 8'b00000000; // 5959 :   0 - 0x0
      13'h1748: dout <= 8'b00000000; // 5960 :   0 - 0x0
      13'h1749: dout <= 8'b00000000; // 5961 :   0 - 0x0
      13'h174A: dout <= 8'b00000000; // 5962 :   0 - 0x0
      13'h174B: dout <= 8'b00000000; // 5963 :   0 - 0x0
      13'h174C: dout <= 8'b00010001; // 5964 :  17 - 0x11
      13'h174D: dout <= 8'b00010011; // 5965 :  19 - 0x13
      13'h174E: dout <= 8'b00011111; // 5966 :  31 - 0x1f
      13'h174F: dout <= 8'b00011111; // 5967 :  31 - 0x1f
      13'h1750: dout <= 8'b00000000; // 5968 :   0 - 0x0 -- Background 0x75
      13'h1751: dout <= 8'b00000000; // 5969 :   0 - 0x0
      13'h1752: dout <= 8'b00000000; // 5970 :   0 - 0x0
      13'h1753: dout <= 8'b00000000; // 5971 :   0 - 0x0
      13'h1754: dout <= 8'b00000000; // 5972 :   0 - 0x0
      13'h1755: dout <= 8'b00000000; // 5973 :   0 - 0x0
      13'h1756: dout <= 8'b00000000; // 5974 :   0 - 0x0
      13'h1757: dout <= 8'b00000000; // 5975 :   0 - 0x0
      13'h1758: dout <= 8'b00000000; // 5976 :   0 - 0x0
      13'h1759: dout <= 8'b00000000; // 5977 :   0 - 0x0
      13'h175A: dout <= 8'b00000000; // 5978 :   0 - 0x0
      13'h175B: dout <= 8'b10000000; // 5979 : 128 - 0x80
      13'h175C: dout <= 8'b11000100; // 5980 : 196 - 0xc4
      13'h175D: dout <= 8'b11100100; // 5981 : 228 - 0xe4
      13'h175E: dout <= 8'b11111100; // 5982 : 252 - 0xfc
      13'h175F: dout <= 8'b11111100; // 5983 : 252 - 0xfc
      13'h1760: dout <= 8'b00000000; // 5984 :   0 - 0x0 -- Background 0x76
      13'h1761: dout <= 8'b00000000; // 5985 :   0 - 0x0
      13'h1762: dout <= 8'b00000000; // 5986 :   0 - 0x0
      13'h1763: dout <= 8'b00000000; // 5987 :   0 - 0x0
      13'h1764: dout <= 8'b00000000; // 5988 :   0 - 0x0
      13'h1765: dout <= 8'b00000000; // 5989 :   0 - 0x0
      13'h1766: dout <= 8'b00000000; // 5990 :   0 - 0x0
      13'h1767: dout <= 8'b00000000; // 5991 :   0 - 0x0
      13'h1768: dout <= 8'b00011111; // 5992 :  31 - 0x1f
      13'h1769: dout <= 8'b00001110; // 5993 :  14 - 0xe
      13'h176A: dout <= 8'b00000110; // 5994 :   6 - 0x6
      13'h176B: dout <= 8'b00000010; // 5995 :   2 - 0x2
      13'h176C: dout <= 8'b00000000; // 5996 :   0 - 0x0
      13'h176D: dout <= 8'b00000000; // 5997 :   0 - 0x0
      13'h176E: dout <= 8'b00000000; // 5998 :   0 - 0x0
      13'h176F: dout <= 8'b00000000; // 5999 :   0 - 0x0
      13'h1770: dout <= 8'b00000000; // 6000 :   0 - 0x0 -- Background 0x77
      13'h1771: dout <= 8'b00000000; // 6001 :   0 - 0x0
      13'h1772: dout <= 8'b00000000; // 6002 :   0 - 0x0
      13'h1773: dout <= 8'b00000000; // 6003 :   0 - 0x0
      13'h1774: dout <= 8'b00000000; // 6004 :   0 - 0x0
      13'h1775: dout <= 8'b00000000; // 6005 :   0 - 0x0
      13'h1776: dout <= 8'b00000000; // 6006 :   0 - 0x0
      13'h1777: dout <= 8'b00000000; // 6007 :   0 - 0x0
      13'h1778: dout <= 8'b11111100; // 6008 : 252 - 0xfc
      13'h1779: dout <= 8'b10111000; // 6009 : 184 - 0xb8
      13'h177A: dout <= 8'b10110000; // 6010 : 176 - 0xb0
      13'h177B: dout <= 8'b10100000; // 6011 : 160 - 0xa0
      13'h177C: dout <= 8'b10000000; // 6012 : 128 - 0x80
      13'h177D: dout <= 8'b00000000; // 6013 :   0 - 0x0
      13'h177E: dout <= 8'b00000000; // 6014 :   0 - 0x0
      13'h177F: dout <= 8'b00000000; // 6015 :   0 - 0x0
      13'h1780: dout <= 8'b00000000; // 6016 :   0 - 0x0 -- Background 0x78
      13'h1781: dout <= 8'b00000000; // 6017 :   0 - 0x0
      13'h1782: dout <= 8'b00000000; // 6018 :   0 - 0x0
      13'h1783: dout <= 8'b00000000; // 6019 :   0 - 0x0
      13'h1784: dout <= 8'b00000000; // 6020 :   0 - 0x0
      13'h1785: dout <= 8'b00000000; // 6021 :   0 - 0x0
      13'h1786: dout <= 8'b00000000; // 6022 :   0 - 0x0
      13'h1787: dout <= 8'b00000000; // 6023 :   0 - 0x0
      13'h1788: dout <= 8'b00000000; // 6024 :   0 - 0x0
      13'h1789: dout <= 8'b00000000; // 6025 :   0 - 0x0
      13'h178A: dout <= 8'b00000000; // 6026 :   0 - 0x0
      13'h178B: dout <= 8'b00000001; // 6027 :   1 - 0x1
      13'h178C: dout <= 8'b00000011; // 6028 :   3 - 0x3
      13'h178D: dout <= 8'b00000110; // 6029 :   6 - 0x6
      13'h178E: dout <= 8'b00000110; // 6030 :   6 - 0x6
      13'h178F: dout <= 8'b00001111; // 6031 :  15 - 0xf
      13'h1790: dout <= 8'b00000000; // 6032 :   0 - 0x0 -- Background 0x79
      13'h1791: dout <= 8'b00000000; // 6033 :   0 - 0x0
      13'h1792: dout <= 8'b00000000; // 6034 :   0 - 0x0
      13'h1793: dout <= 8'b00000000; // 6035 :   0 - 0x0
      13'h1794: dout <= 8'b00000000; // 6036 :   0 - 0x0
      13'h1795: dout <= 8'b00000000; // 6037 :   0 - 0x0
      13'h1796: dout <= 8'b00000000; // 6038 :   0 - 0x0
      13'h1797: dout <= 8'b00000000; // 6039 :   0 - 0x0
      13'h1798: dout <= 8'b00000000; // 6040 :   0 - 0x0
      13'h1799: dout <= 8'b00011000; // 6041 :  24 - 0x18
      13'h179A: dout <= 8'b11110100; // 6042 : 244 - 0xf4
      13'h179B: dout <= 8'b11111000; // 6043 : 248 - 0xf8
      13'h179C: dout <= 8'b00111000; // 6044 :  56 - 0x38
      13'h179D: dout <= 8'b01111100; // 6045 : 124 - 0x7c
      13'h179E: dout <= 8'b11111100; // 6046 : 252 - 0xfc
      13'h179F: dout <= 8'b11111100; // 6047 : 252 - 0xfc
      13'h17A0: dout <= 8'b00000000; // 6048 :   0 - 0x0 -- Background 0x7a
      13'h17A1: dout <= 8'b00000000; // 6049 :   0 - 0x0
      13'h17A2: dout <= 8'b00000000; // 6050 :   0 - 0x0
      13'h17A3: dout <= 8'b00000000; // 6051 :   0 - 0x0
      13'h17A4: dout <= 8'b00000000; // 6052 :   0 - 0x0
      13'h17A5: dout <= 8'b00000000; // 6053 :   0 - 0x0
      13'h17A6: dout <= 8'b00000000; // 6054 :   0 - 0x0
      13'h17A7: dout <= 8'b00000000; // 6055 :   0 - 0x0
      13'h17A8: dout <= 8'b00001111; // 6056 :  15 - 0xf
      13'h17A9: dout <= 8'b00011111; // 6057 :  31 - 0x1f
      13'h17AA: dout <= 8'b00110000; // 6058 :  48 - 0x30
      13'h17AB: dout <= 8'b00111000; // 6059 :  56 - 0x38
      13'h17AC: dout <= 8'b00011101; // 6060 :  29 - 0x1d
      13'h17AD: dout <= 8'b00000011; // 6061 :   3 - 0x3
      13'h17AE: dout <= 8'b00000011; // 6062 :   3 - 0x3
      13'h17AF: dout <= 8'b00000000; // 6063 :   0 - 0x0
      13'h17B0: dout <= 8'b00000000; // 6064 :   0 - 0x0 -- Background 0x7b
      13'h17B1: dout <= 8'b00000000; // 6065 :   0 - 0x0
      13'h17B2: dout <= 8'b00000000; // 6066 :   0 - 0x0
      13'h17B3: dout <= 8'b00000000; // 6067 :   0 - 0x0
      13'h17B4: dout <= 8'b00000000; // 6068 :   0 - 0x0
      13'h17B5: dout <= 8'b00000000; // 6069 :   0 - 0x0
      13'h17B6: dout <= 8'b00000000; // 6070 :   0 - 0x0
      13'h17B7: dout <= 8'b00000000; // 6071 :   0 - 0x0
      13'h17B8: dout <= 8'b11111100; // 6072 : 252 - 0xfc
      13'h17B9: dout <= 8'b11111100; // 6073 : 252 - 0xfc
      13'h17BA: dout <= 8'b01111100; // 6074 : 124 - 0x7c
      13'h17BB: dout <= 8'b10001110; // 6075 : 142 - 0x8e
      13'h17BC: dout <= 8'b10000110; // 6076 : 134 - 0x86
      13'h17BD: dout <= 8'b10011100; // 6077 : 156 - 0x9c
      13'h17BE: dout <= 8'b01111000; // 6078 : 120 - 0x78
      13'h17BF: dout <= 8'b00000000; // 6079 :   0 - 0x0
      13'h17C0: dout <= 8'b00000000; // 6080 :   0 - 0x0 -- Background 0x7c
      13'h17C1: dout <= 8'b00000001; // 6081 :   1 - 0x1
      13'h17C2: dout <= 8'b00000110; // 6082 :   6 - 0x6
      13'h17C3: dout <= 8'b00000111; // 6083 :   7 - 0x7
      13'h17C4: dout <= 8'b00000111; // 6084 :   7 - 0x7
      13'h17C5: dout <= 8'b00000111; // 6085 :   7 - 0x7
      13'h17C6: dout <= 8'b00000001; // 6086 :   1 - 0x1
      13'h17C7: dout <= 8'b00000011; // 6087 :   3 - 0x3
      13'h17C8: dout <= 8'b00000000; // 6088 :   0 - 0x0
      13'h17C9: dout <= 8'b00000001; // 6089 :   1 - 0x1
      13'h17CA: dout <= 8'b00000110; // 6090 :   6 - 0x6
      13'h17CB: dout <= 8'b00000111; // 6091 :   7 - 0x7
      13'h17CC: dout <= 8'b00000111; // 6092 :   7 - 0x7
      13'h17CD: dout <= 8'b00000111; // 6093 :   7 - 0x7
      13'h17CE: dout <= 8'b00000001; // 6094 :   1 - 0x1
      13'h17CF: dout <= 8'b00000011; // 6095 :   3 - 0x3
      13'h17D0: dout <= 8'b00000000; // 6096 :   0 - 0x0 -- Background 0x7d
      13'h17D1: dout <= 8'b11000000; // 6097 : 192 - 0xc0
      13'h17D2: dout <= 8'b00110000; // 6098 :  48 - 0x30
      13'h17D3: dout <= 8'b11110000; // 6099 : 240 - 0xf0
      13'h17D4: dout <= 8'b11110000; // 6100 : 240 - 0xf0
      13'h17D5: dout <= 8'b11110000; // 6101 : 240 - 0xf0
      13'h17D6: dout <= 8'b01000000; // 6102 :  64 - 0x40
      13'h17D7: dout <= 8'b01000000; // 6103 :  64 - 0x40
      13'h17D8: dout <= 8'b00000000; // 6104 :   0 - 0x0
      13'h17D9: dout <= 8'b11000000; // 6105 : 192 - 0xc0
      13'h17DA: dout <= 8'b00110000; // 6106 :  48 - 0x30
      13'h17DB: dout <= 8'b11110000; // 6107 : 240 - 0xf0
      13'h17DC: dout <= 8'b11110000; // 6108 : 240 - 0xf0
      13'h17DD: dout <= 8'b11110000; // 6109 : 240 - 0xf0
      13'h17DE: dout <= 8'b01000000; // 6110 :  64 - 0x40
      13'h17DF: dout <= 8'b01000000; // 6111 :  64 - 0x40
      13'h17E0: dout <= 8'b00000001; // 6112 :   1 - 0x1 -- Background 0x7e
      13'h17E1: dout <= 8'b00000000; // 6113 :   0 - 0x0
      13'h17E2: dout <= 8'b00000001; // 6114 :   1 - 0x1
      13'h17E3: dout <= 8'b00000011; // 6115 :   3 - 0x3
      13'h17E4: dout <= 8'b00000001; // 6116 :   1 - 0x1
      13'h17E5: dout <= 8'b00000000; // 6117 :   0 - 0x0
      13'h17E6: dout <= 8'b00000000; // 6118 :   0 - 0x0
      13'h17E7: dout <= 8'b00000000; // 6119 :   0 - 0x0
      13'h17E8: dout <= 8'b00000001; // 6120 :   1 - 0x1
      13'h17E9: dout <= 8'b00000000; // 6121 :   0 - 0x0
      13'h17EA: dout <= 8'b00000001; // 6122 :   1 - 0x1
      13'h17EB: dout <= 8'b00000011; // 6123 :   3 - 0x3
      13'h17EC: dout <= 8'b00000001; // 6124 :   1 - 0x1
      13'h17ED: dout <= 8'b00000000; // 6125 :   0 - 0x0
      13'h17EE: dout <= 8'b00000000; // 6126 :   0 - 0x0
      13'h17EF: dout <= 8'b00000000; // 6127 :   0 - 0x0
      13'h17F0: dout <= 8'b01000000; // 6128 :  64 - 0x40 -- Background 0x7f
      13'h17F1: dout <= 8'b01000000; // 6129 :  64 - 0x40
      13'h17F2: dout <= 8'b01000000; // 6130 :  64 - 0x40
      13'h17F3: dout <= 8'b01000000; // 6131 :  64 - 0x40
      13'h17F4: dout <= 8'b01000000; // 6132 :  64 - 0x40
      13'h17F5: dout <= 8'b10000000; // 6133 : 128 - 0x80
      13'h17F6: dout <= 8'b00000000; // 6134 :   0 - 0x0
      13'h17F7: dout <= 8'b00000000; // 6135 :   0 - 0x0
      13'h17F8: dout <= 8'b01000000; // 6136 :  64 - 0x40
      13'h17F9: dout <= 8'b01000000; // 6137 :  64 - 0x40
      13'h17FA: dout <= 8'b01000000; // 6138 :  64 - 0x40
      13'h17FB: dout <= 8'b01000000; // 6139 :  64 - 0x40
      13'h17FC: dout <= 8'b01000000; // 6140 :  64 - 0x40
      13'h17FD: dout <= 8'b10000000; // 6141 : 128 - 0x80
      13'h17FE: dout <= 8'b00000000; // 6142 :   0 - 0x0
      13'h17FF: dout <= 8'b00000000; // 6143 :   0 - 0x0
      13'h1800: dout <= 8'b11111111; // 6144 : 255 - 0xff -- Background 0x80
      13'h1801: dout <= 8'b11111111; // 6145 : 255 - 0xff
      13'h1802: dout <= 8'b11111111; // 6146 : 255 - 0xff
      13'h1803: dout <= 8'b11111111; // 6147 : 255 - 0xff
      13'h1804: dout <= 8'b11000000; // 6148 : 192 - 0xc0
      13'h1805: dout <= 8'b11000000; // 6149 : 192 - 0xc0
      13'h1806: dout <= 8'b11000000; // 6150 : 192 - 0xc0
      13'h1807: dout <= 8'b11000111; // 6151 : 199 - 0xc7
      13'h1808: dout <= 8'b00000000; // 6152 :   0 - 0x0
      13'h1809: dout <= 8'b00000000; // 6153 :   0 - 0x0
      13'h180A: dout <= 8'b00000000; // 6154 :   0 - 0x0
      13'h180B: dout <= 8'b00000000; // 6155 :   0 - 0x0
      13'h180C: dout <= 8'b00000000; // 6156 :   0 - 0x0
      13'h180D: dout <= 8'b00011111; // 6157 :  31 - 0x1f
      13'h180E: dout <= 8'b00010000; // 6158 :  16 - 0x10
      13'h180F: dout <= 8'b00010111; // 6159 :  23 - 0x17
      13'h1810: dout <= 8'b11111111; // 6160 : 255 - 0xff -- Background 0x81
      13'h1811: dout <= 8'b11111111; // 6161 : 255 - 0xff
      13'h1812: dout <= 8'b11111111; // 6162 : 255 - 0xff
      13'h1813: dout <= 8'b11111111; // 6163 : 255 - 0xff
      13'h1814: dout <= 8'b00000000; // 6164 :   0 - 0x0
      13'h1815: dout <= 8'b00000000; // 6165 :   0 - 0x0
      13'h1816: dout <= 8'b00000000; // 6166 :   0 - 0x0
      13'h1817: dout <= 8'b11111111; // 6167 : 255 - 0xff
      13'h1818: dout <= 8'b00000000; // 6168 :   0 - 0x0
      13'h1819: dout <= 8'b00000000; // 6169 :   0 - 0x0
      13'h181A: dout <= 8'b00000000; // 6170 :   0 - 0x0
      13'h181B: dout <= 8'b00000000; // 6171 :   0 - 0x0
      13'h181C: dout <= 8'b00000000; // 6172 :   0 - 0x0
      13'h181D: dout <= 8'b11111111; // 6173 : 255 - 0xff
      13'h181E: dout <= 8'b00000000; // 6174 :   0 - 0x0
      13'h181F: dout <= 8'b11111111; // 6175 : 255 - 0xff
      13'h1820: dout <= 8'b11111111; // 6176 : 255 - 0xff -- Background 0x82
      13'h1821: dout <= 8'b11111111; // 6177 : 255 - 0xff
      13'h1822: dout <= 8'b11111111; // 6178 : 255 - 0xff
      13'h1823: dout <= 8'b11111111; // 6179 : 255 - 0xff
      13'h1824: dout <= 8'b01111111; // 6180 : 127 - 0x7f
      13'h1825: dout <= 8'b00111111; // 6181 :  63 - 0x3f
      13'h1826: dout <= 8'b00011111; // 6182 :  31 - 0x1f
      13'h1827: dout <= 8'b11001111; // 6183 : 207 - 0xcf
      13'h1828: dout <= 8'b00000000; // 6184 :   0 - 0x0
      13'h1829: dout <= 8'b00000000; // 6185 :   0 - 0x0
      13'h182A: dout <= 8'b00000000; // 6186 :   0 - 0x0
      13'h182B: dout <= 8'b00000000; // 6187 :   0 - 0x0
      13'h182C: dout <= 8'b00000000; // 6188 :   0 - 0x0
      13'h182D: dout <= 8'b10000000; // 6189 : 128 - 0x80
      13'h182E: dout <= 8'b00000000; // 6190 :   0 - 0x0
      13'h182F: dout <= 8'b11000000; // 6191 : 192 - 0xc0
      13'h1830: dout <= 8'b11111111; // 6192 : 255 - 0xff -- Background 0x83
      13'h1831: dout <= 8'b11111111; // 6193 : 255 - 0xff
      13'h1832: dout <= 8'b11111111; // 6194 : 255 - 0xff
      13'h1833: dout <= 8'b11110111; // 6195 : 247 - 0xf7
      13'h1834: dout <= 8'b11110111; // 6196 : 247 - 0xf7
      13'h1835: dout <= 8'b11100010; // 6197 : 226 - 0xe2
      13'h1836: dout <= 8'b11100000; // 6198 : 224 - 0xe0
      13'h1837: dout <= 8'b11000110; // 6199 : 198 - 0xc6
      13'h1838: dout <= 8'b00000000; // 6200 :   0 - 0x0
      13'h1839: dout <= 8'b00000000; // 6201 :   0 - 0x0
      13'h183A: dout <= 8'b00000000; // 6202 :   0 - 0x0
      13'h183B: dout <= 8'b00000000; // 6203 :   0 - 0x0
      13'h183C: dout <= 8'b00000000; // 6204 :   0 - 0x0
      13'h183D: dout <= 8'b00001000; // 6205 :   8 - 0x8
      13'h183E: dout <= 8'b00001000; // 6206 :   8 - 0x8
      13'h183F: dout <= 8'b00010110; // 6207 :  22 - 0x16
      13'h1840: dout <= 8'b11111111; // 6208 : 255 - 0xff -- Background 0x84
      13'h1841: dout <= 8'b11111111; // 6209 : 255 - 0xff
      13'h1842: dout <= 8'b11111111; // 6210 : 255 - 0xff
      13'h1843: dout <= 8'b11111111; // 6211 : 255 - 0xff
      13'h1844: dout <= 8'b10111111; // 6212 : 191 - 0xbf
      13'h1845: dout <= 8'b10111111; // 6213 : 191 - 0xbf
      13'h1846: dout <= 8'b00011111; // 6214 :  31 - 0x1f
      13'h1847: dout <= 8'b00011111; // 6215 :  31 - 0x1f
      13'h1848: dout <= 8'b00000000; // 6216 :   0 - 0x0
      13'h1849: dout <= 8'b00000000; // 6217 :   0 - 0x0
      13'h184A: dout <= 8'b00000000; // 6218 :   0 - 0x0
      13'h184B: dout <= 8'b00000000; // 6219 :   0 - 0x0
      13'h184C: dout <= 8'b00000000; // 6220 :   0 - 0x0
      13'h184D: dout <= 8'b00000000; // 6221 :   0 - 0x0
      13'h184E: dout <= 8'b01000000; // 6222 :  64 - 0x40
      13'h184F: dout <= 8'b11000000; // 6223 : 192 - 0xc0
      13'h1850: dout <= 8'b11111111; // 6224 : 255 - 0xff -- Background 0x85
      13'h1851: dout <= 8'b11111111; // 6225 : 255 - 0xff
      13'h1852: dout <= 8'b11111111; // 6226 : 255 - 0xff
      13'h1853: dout <= 8'b11111111; // 6227 : 255 - 0xff
      13'h1854: dout <= 8'b11111110; // 6228 : 254 - 0xfe
      13'h1855: dout <= 8'b11111000; // 6229 : 248 - 0xf8
      13'h1856: dout <= 8'b11100000; // 6230 : 224 - 0xe0
      13'h1857: dout <= 8'b11000000; // 6231 : 192 - 0xc0
      13'h1858: dout <= 8'b00000000; // 6232 :   0 - 0x0
      13'h1859: dout <= 8'b00000000; // 6233 :   0 - 0x0
      13'h185A: dout <= 8'b00000000; // 6234 :   0 - 0x0
      13'h185B: dout <= 8'b00000000; // 6235 :   0 - 0x0
      13'h185C: dout <= 8'b00000000; // 6236 :   0 - 0x0
      13'h185D: dout <= 8'b00000001; // 6237 :   1 - 0x1
      13'h185E: dout <= 8'b00000111; // 6238 :   7 - 0x7
      13'h185F: dout <= 8'b00001100; // 6239 :  12 - 0xc
      13'h1860: dout <= 8'b11111111; // 6240 : 255 - 0xff -- Background 0x86
      13'h1861: dout <= 8'b11111111; // 6241 : 255 - 0xff
      13'h1862: dout <= 8'b11111111; // 6242 : 255 - 0xff
      13'h1863: dout <= 8'b11111111; // 6243 : 255 - 0xff
      13'h1864: dout <= 8'b00000111; // 6244 :   7 - 0x7
      13'h1865: dout <= 8'b00000000; // 6245 :   0 - 0x0
      13'h1866: dout <= 8'b00111111; // 6246 :  63 - 0x3f
      13'h1867: dout <= 8'b11111111; // 6247 : 255 - 0xff
      13'h1868: dout <= 8'b00000000; // 6248 :   0 - 0x0
      13'h1869: dout <= 8'b00000000; // 6249 :   0 - 0x0
      13'h186A: dout <= 8'b00000000; // 6250 :   0 - 0x0
      13'h186B: dout <= 8'b00000000; // 6251 :   0 - 0x0
      13'h186C: dout <= 8'b00000000; // 6252 :   0 - 0x0
      13'h186D: dout <= 8'b11000000; // 6253 : 192 - 0xc0
      13'h186E: dout <= 8'b00111111; // 6254 :  63 - 0x3f
      13'h186F: dout <= 8'b11111111; // 6255 : 255 - 0xff
      13'h1870: dout <= 8'b11111111; // 6256 : 255 - 0xff -- Background 0x87
      13'h1871: dout <= 8'b11111111; // 6257 : 255 - 0xff
      13'h1872: dout <= 8'b11111111; // 6258 : 255 - 0xff
      13'h1873: dout <= 8'b11111111; // 6259 : 255 - 0xff
      13'h1874: dout <= 8'b11111111; // 6260 : 255 - 0xff
      13'h1875: dout <= 8'b11111111; // 6261 : 255 - 0xff
      13'h1876: dout <= 8'b00111111; // 6262 :  63 - 0x3f
      13'h1877: dout <= 8'b11001111; // 6263 : 207 - 0xcf
      13'h1878: dout <= 8'b00000000; // 6264 :   0 - 0x0
      13'h1879: dout <= 8'b00000000; // 6265 :   0 - 0x0
      13'h187A: dout <= 8'b00000000; // 6266 :   0 - 0x0
      13'h187B: dout <= 8'b00000000; // 6267 :   0 - 0x0
      13'h187C: dout <= 8'b00000000; // 6268 :   0 - 0x0
      13'h187D: dout <= 8'b00000000; // 6269 :   0 - 0x0
      13'h187E: dout <= 8'b00000000; // 6270 :   0 - 0x0
      13'h187F: dout <= 8'b11000000; // 6271 : 192 - 0xc0
      13'h1880: dout <= 8'b11111111; // 6272 : 255 - 0xff -- Background 0x88
      13'h1881: dout <= 8'b11111111; // 6273 : 255 - 0xff
      13'h1882: dout <= 8'b11111111; // 6274 : 255 - 0xff
      13'h1883: dout <= 8'b11111111; // 6275 : 255 - 0xff
      13'h1884: dout <= 8'b11111111; // 6276 : 255 - 0xff
      13'h1885: dout <= 8'b11111111; // 6277 : 255 - 0xff
      13'h1886: dout <= 8'b11111111; // 6278 : 255 - 0xff
      13'h1887: dout <= 8'b11111111; // 6279 : 255 - 0xff
      13'h1888: dout <= 8'b00000000; // 6280 :   0 - 0x0
      13'h1889: dout <= 8'b00000000; // 6281 :   0 - 0x0
      13'h188A: dout <= 8'b00000000; // 6282 :   0 - 0x0
      13'h188B: dout <= 8'b00000000; // 6283 :   0 - 0x0
      13'h188C: dout <= 8'b00000000; // 6284 :   0 - 0x0
      13'h188D: dout <= 8'b00000000; // 6285 :   0 - 0x0
      13'h188E: dout <= 8'b00000000; // 6286 :   0 - 0x0
      13'h188F: dout <= 8'b00000000; // 6287 :   0 - 0x0
      13'h1890: dout <= 8'b11111111; // 6288 : 255 - 0xff -- Background 0x89
      13'h1891: dout <= 8'b11111111; // 6289 : 255 - 0xff
      13'h1892: dout <= 8'b11111111; // 6290 : 255 - 0xff
      13'h1893: dout <= 8'b01110111; // 6291 : 119 - 0x77
      13'h1894: dout <= 8'b00010011; // 6292 :  19 - 0x13
      13'h1895: dout <= 8'b00000001; // 6293 :   1 - 0x1
      13'h1896: dout <= 8'b00010000; // 6294 :  16 - 0x10
      13'h1897: dout <= 8'b00011000; // 6295 :  24 - 0x18
      13'h1898: dout <= 8'b00000000; // 6296 :   0 - 0x0
      13'h1899: dout <= 8'b00000000; // 6297 :   0 - 0x0
      13'h189A: dout <= 8'b00000000; // 6298 :   0 - 0x0
      13'h189B: dout <= 8'b00000000; // 6299 :   0 - 0x0
      13'h189C: dout <= 8'b00000000; // 6300 :   0 - 0x0
      13'h189D: dout <= 8'b01000100; // 6301 :  68 - 0x44
      13'h189E: dout <= 8'b01010110; // 6302 :  86 - 0x56
      13'h189F: dout <= 8'b01011011; // 6303 :  91 - 0x5b
      13'h18A0: dout <= 8'b11111111; // 6304 : 255 - 0xff -- Background 0x8a
      13'h18A1: dout <= 8'b11111111; // 6305 : 255 - 0xff
      13'h18A2: dout <= 8'b11111111; // 6306 : 255 - 0xff
      13'h18A3: dout <= 8'b11111111; // 6307 : 255 - 0xff
      13'h18A4: dout <= 8'b11111111; // 6308 : 255 - 0xff
      13'h18A5: dout <= 8'b11111111; // 6309 : 255 - 0xff
      13'h18A6: dout <= 8'b11111111; // 6310 : 255 - 0xff
      13'h18A7: dout <= 8'b01111111; // 6311 : 127 - 0x7f
      13'h18A8: dout <= 8'b00000000; // 6312 :   0 - 0x0
      13'h18A9: dout <= 8'b00000000; // 6313 :   0 - 0x0
      13'h18AA: dout <= 8'b00000000; // 6314 :   0 - 0x0
      13'h18AB: dout <= 8'b00000000; // 6315 :   0 - 0x0
      13'h18AC: dout <= 8'b00000000; // 6316 :   0 - 0x0
      13'h18AD: dout <= 8'b00000000; // 6317 :   0 - 0x0
      13'h18AE: dout <= 8'b00000000; // 6318 :   0 - 0x0
      13'h18AF: dout <= 8'b00000000; // 6319 :   0 - 0x0
      13'h18B0: dout <= 8'b11111111; // 6320 : 255 - 0xff -- Background 0x8b
      13'h18B1: dout <= 8'b11111111; // 6321 : 255 - 0xff
      13'h18B2: dout <= 8'b11111111; // 6322 : 255 - 0xff
      13'h18B3: dout <= 8'b11110111; // 6323 : 247 - 0xf7
      13'h18B4: dout <= 8'b11100101; // 6324 : 229 - 0xe5
      13'h18B5: dout <= 8'b11000001; // 6325 : 193 - 0xc1
      13'h18B6: dout <= 8'b10000100; // 6326 : 132 - 0x84
      13'h18B7: dout <= 8'b00001100; // 6327 :  12 - 0xc
      13'h18B8: dout <= 8'b00000000; // 6328 :   0 - 0x0
      13'h18B9: dout <= 8'b00000000; // 6329 :   0 - 0x0
      13'h18BA: dout <= 8'b00000000; // 6330 :   0 - 0x0
      13'h18BB: dout <= 8'b00000000; // 6331 :   0 - 0x0
      13'h18BC: dout <= 8'b00000000; // 6332 :   0 - 0x0
      13'h18BD: dout <= 8'b00010000; // 6333 :  16 - 0x10
      13'h18BE: dout <= 8'b00110100; // 6334 :  52 - 0x34
      13'h18BF: dout <= 8'b01101101; // 6335 : 109 - 0x6d
      13'h18C0: dout <= 8'b11111111; // 6336 : 255 - 0xff -- Background 0x8c
      13'h18C1: dout <= 8'b11111111; // 6337 : 255 - 0xff
      13'h18C2: dout <= 8'b11111111; // 6338 : 255 - 0xff
      13'h18C3: dout <= 8'b11111111; // 6339 : 255 - 0xff
      13'h18C4: dout <= 8'b11111111; // 6340 : 255 - 0xff
      13'h18C5: dout <= 8'b01111111; // 6341 : 127 - 0x7f
      13'h18C6: dout <= 8'b01111110; // 6342 : 126 - 0x7e
      13'h18C7: dout <= 8'b01111110; // 6343 : 126 - 0x7e
      13'h18C8: dout <= 8'b00000000; // 6344 :   0 - 0x0
      13'h18C9: dout <= 8'b00000000; // 6345 :   0 - 0x0
      13'h18CA: dout <= 8'b00000000; // 6346 :   0 - 0x0
      13'h18CB: dout <= 8'b00000000; // 6347 :   0 - 0x0
      13'h18CC: dout <= 8'b00000000; // 6348 :   0 - 0x0
      13'h18CD: dout <= 8'b00000000; // 6349 :   0 - 0x0
      13'h18CE: dout <= 8'b00000000; // 6350 :   0 - 0x0
      13'h18CF: dout <= 8'b00000000; // 6351 :   0 - 0x0
      13'h18D0: dout <= 8'b11111111; // 6352 : 255 - 0xff -- Background 0x8d
      13'h18D1: dout <= 8'b11111111; // 6353 : 255 - 0xff
      13'h18D2: dout <= 8'b10111111; // 6354 : 191 - 0xbf
      13'h18D3: dout <= 8'b10110111; // 6355 : 183 - 0xb7
      13'h18D4: dout <= 8'b00010111; // 6356 :  23 - 0x17
      13'h18D5: dout <= 8'b00000011; // 6357 :   3 - 0x3
      13'h18D6: dout <= 8'b00100011; // 6358 :  35 - 0x23
      13'h18D7: dout <= 8'b00100001; // 6359 :  33 - 0x21
      13'h18D8: dout <= 8'b00000000; // 6360 :   0 - 0x0
      13'h18D9: dout <= 8'b00000000; // 6361 :   0 - 0x0
      13'h18DA: dout <= 8'b00000000; // 6362 :   0 - 0x0
      13'h18DB: dout <= 8'b00000000; // 6363 :   0 - 0x0
      13'h18DC: dout <= 8'b01000000; // 6364 :  64 - 0x40
      13'h18DD: dout <= 8'b01001000; // 6365 :  72 - 0x48
      13'h18DE: dout <= 8'b10101000; // 6366 : 168 - 0xa8
      13'h18DF: dout <= 8'b10101100; // 6367 : 172 - 0xac
      13'h18E0: dout <= 8'b11111111; // 6368 : 255 - 0xff -- Background 0x8e
      13'h18E1: dout <= 8'b11111111; // 6369 : 255 - 0xff
      13'h18E2: dout <= 8'b11111011; // 6370 : 251 - 0xfb
      13'h18E3: dout <= 8'b11111001; // 6371 : 249 - 0xf9
      13'h18E4: dout <= 8'b11111000; // 6372 : 248 - 0xf8
      13'h18E5: dout <= 8'b11111000; // 6373 : 248 - 0xf8
      13'h18E6: dout <= 8'b11111000; // 6374 : 248 - 0xf8
      13'h18E7: dout <= 8'b11111000; // 6375 : 248 - 0xf8
      13'h18E8: dout <= 8'b00000000; // 6376 :   0 - 0x0
      13'h18E9: dout <= 8'b00000000; // 6377 :   0 - 0x0
      13'h18EA: dout <= 8'b00000000; // 6378 :   0 - 0x0
      13'h18EB: dout <= 8'b00000000; // 6379 :   0 - 0x0
      13'h18EC: dout <= 8'b00000010; // 6380 :   2 - 0x2
      13'h18ED: dout <= 8'b00000010; // 6381 :   2 - 0x2
      13'h18EE: dout <= 8'b00000010; // 6382 :   2 - 0x2
      13'h18EF: dout <= 8'b00000010; // 6383 :   2 - 0x2
      13'h18F0: dout <= 8'b11111111; // 6384 : 255 - 0xff -- Background 0x8f
      13'h18F1: dout <= 8'b11111111; // 6385 : 255 - 0xff
      13'h18F2: dout <= 8'b01111000; // 6386 : 120 - 0x78
      13'h18F3: dout <= 8'b00111000; // 6387 :  56 - 0x38
      13'h18F4: dout <= 8'b00011000; // 6388 :  24 - 0x18
      13'h18F5: dout <= 8'b00001000; // 6389 :   8 - 0x8
      13'h18F6: dout <= 8'b10000000; // 6390 : 128 - 0x80
      13'h18F7: dout <= 8'b11000000; // 6391 : 192 - 0xc0
      13'h18F8: dout <= 8'b00000000; // 6392 :   0 - 0x0
      13'h18F9: dout <= 8'b00000000; // 6393 :   0 - 0x0
      13'h18FA: dout <= 8'b00000000; // 6394 :   0 - 0x0
      13'h18FB: dout <= 8'b00000011; // 6395 :   3 - 0x3
      13'h18FC: dout <= 8'b01000011; // 6396 :  67 - 0x43
      13'h18FD: dout <= 8'b01100010; // 6397 :  98 - 0x62
      13'h18FE: dout <= 8'b10110010; // 6398 : 178 - 0xb2
      13'h18FF: dout <= 8'b11011010; // 6399 : 218 - 0xda
      13'h1900: dout <= 8'b11111111; // 6400 : 255 - 0xff -- Background 0x90
      13'h1901: dout <= 8'b11111111; // 6401 : 255 - 0xff
      13'h1902: dout <= 8'b00000001; // 6402 :   1 - 0x1
      13'h1903: dout <= 8'b00000001; // 6403 :   1 - 0x1
      13'h1904: dout <= 8'b00000001; // 6404 :   1 - 0x1
      13'h1905: dout <= 8'b00000000; // 6405 :   0 - 0x0
      13'h1906: dout <= 8'b11111111; // 6406 : 255 - 0xff
      13'h1907: dout <= 8'b11111111; // 6407 : 255 - 0xff
      13'h1908: dout <= 8'b00000000; // 6408 :   0 - 0x0
      13'h1909: dout <= 8'b00000000; // 6409 :   0 - 0x0
      13'h190A: dout <= 8'b00000000; // 6410 :   0 - 0x0
      13'h190B: dout <= 8'b11111100; // 6411 : 252 - 0xfc
      13'h190C: dout <= 8'b11111100; // 6412 : 252 - 0xfc
      13'h190D: dout <= 8'b00000000; // 6413 :   0 - 0x0
      13'h190E: dout <= 8'b11111111; // 6414 : 255 - 0xff
      13'h190F: dout <= 8'b11111111; // 6415 : 255 - 0xff
      13'h1910: dout <= 8'b11111111; // 6416 : 255 - 0xff -- Background 0x91
      13'h1911: dout <= 8'b11111111; // 6417 : 255 - 0xff
      13'h1912: dout <= 8'b11111111; // 6418 : 255 - 0xff
      13'h1913: dout <= 8'b11111111; // 6419 : 255 - 0xff
      13'h1914: dout <= 8'b11111111; // 6420 : 255 - 0xff
      13'h1915: dout <= 8'b11111111; // 6421 : 255 - 0xff
      13'h1916: dout <= 8'b01111111; // 6422 : 127 - 0x7f
      13'h1917: dout <= 8'b00111111; // 6423 :  63 - 0x3f
      13'h1918: dout <= 8'b00000000; // 6424 :   0 - 0x0
      13'h1919: dout <= 8'b00000000; // 6425 :   0 - 0x0
      13'h191A: dout <= 8'b00000000; // 6426 :   0 - 0x0
      13'h191B: dout <= 8'b00000000; // 6427 :   0 - 0x0
      13'h191C: dout <= 8'b00000000; // 6428 :   0 - 0x0
      13'h191D: dout <= 8'b00000000; // 6429 :   0 - 0x0
      13'h191E: dout <= 8'b00000000; // 6430 :   0 - 0x0
      13'h191F: dout <= 8'b00000000; // 6431 :   0 - 0x0
      13'h1920: dout <= 8'b11000111; // 6432 : 199 - 0xc7 -- Background 0x92
      13'h1921: dout <= 8'b11000111; // 6433 : 199 - 0xc7
      13'h1922: dout <= 8'b11000111; // 6434 : 199 - 0xc7
      13'h1923: dout <= 8'b11000111; // 6435 : 199 - 0xc7
      13'h1924: dout <= 8'b11000111; // 6436 : 199 - 0xc7
      13'h1925: dout <= 8'b11000111; // 6437 : 199 - 0xc7
      13'h1926: dout <= 8'b11000111; // 6438 : 199 - 0xc7
      13'h1927: dout <= 8'b11000111; // 6439 : 199 - 0xc7
      13'h1928: dout <= 8'b00010111; // 6440 :  23 - 0x17
      13'h1929: dout <= 8'b00010111; // 6441 :  23 - 0x17
      13'h192A: dout <= 8'b00010111; // 6442 :  23 - 0x17
      13'h192B: dout <= 8'b00010111; // 6443 :  23 - 0x17
      13'h192C: dout <= 8'b00010111; // 6444 :  23 - 0x17
      13'h192D: dout <= 8'b00010111; // 6445 :  23 - 0x17
      13'h192E: dout <= 8'b00010111; // 6446 :  23 - 0x17
      13'h192F: dout <= 8'b00010111; // 6447 :  23 - 0x17
      13'h1930: dout <= 8'b11111111; // 6448 : 255 - 0xff -- Background 0x93
      13'h1931: dout <= 8'b11111111; // 6449 : 255 - 0xff
      13'h1932: dout <= 8'b11111111; // 6450 : 255 - 0xff
      13'h1933: dout <= 8'b11111111; // 6451 : 255 - 0xff
      13'h1934: dout <= 8'b11111001; // 6452 : 249 - 0xf9
      13'h1935: dout <= 8'b11111001; // 6453 : 249 - 0xf9
      13'h1936: dout <= 8'b11111111; // 6454 : 255 - 0xff
      13'h1937: dout <= 8'b11111111; // 6455 : 255 - 0xff
      13'h1938: dout <= 8'b11111111; // 6456 : 255 - 0xff
      13'h1939: dout <= 8'b11111111; // 6457 : 255 - 0xff
      13'h193A: dout <= 8'b11111111; // 6458 : 255 - 0xff
      13'h193B: dout <= 8'b11111111; // 6459 : 255 - 0xff
      13'h193C: dout <= 8'b11111001; // 6460 : 249 - 0xf9
      13'h193D: dout <= 8'b11111001; // 6461 : 249 - 0xf9
      13'h193E: dout <= 8'b11111111; // 6462 : 255 - 0xff
      13'h193F: dout <= 8'b11111111; // 6463 : 255 - 0xff
      13'h1940: dout <= 8'b11110111; // 6464 : 247 - 0xf7 -- Background 0x94
      13'h1941: dout <= 8'b11111011; // 6465 : 251 - 0xfb
      13'h1942: dout <= 8'b11111011; // 6466 : 251 - 0xfb
      13'h1943: dout <= 8'b11111101; // 6467 : 253 - 0xfd
      13'h1944: dout <= 8'b11111100; // 6468 : 252 - 0xfc
      13'h1945: dout <= 8'b11111100; // 6469 : 252 - 0xfc
      13'h1946: dout <= 8'b01111100; // 6470 : 124 - 0x7c
      13'h1947: dout <= 8'b01111100; // 6471 : 124 - 0x7c
      13'h1948: dout <= 8'b11110000; // 6472 : 240 - 0xf0
      13'h1949: dout <= 8'b11111000; // 6473 : 248 - 0xf8
      13'h194A: dout <= 8'b11111000; // 6474 : 248 - 0xf8
      13'h194B: dout <= 8'b11111100; // 6475 : 252 - 0xfc
      13'h194C: dout <= 8'b11111100; // 6476 : 252 - 0xfc
      13'h194D: dout <= 8'b11111100; // 6477 : 252 - 0xfc
      13'h194E: dout <= 8'b01111100; // 6478 : 124 - 0x7c
      13'h194F: dout <= 8'b01111100; // 6479 : 124 - 0x7c
      13'h1950: dout <= 8'b11000111; // 6480 : 199 - 0xc7 -- Background 0x95
      13'h1951: dout <= 8'b10001111; // 6481 : 143 - 0x8f
      13'h1952: dout <= 8'b10001111; // 6482 : 143 - 0x8f
      13'h1953: dout <= 8'b00011111; // 6483 :  31 - 0x1f
      13'h1954: dout <= 8'b00011111; // 6484 :  31 - 0x1f
      13'h1955: dout <= 8'b00111111; // 6485 :  63 - 0x3f
      13'h1956: dout <= 8'b00111111; // 6486 :  63 - 0x3f
      13'h1957: dout <= 8'b01111111; // 6487 : 127 - 0x7f
      13'h1958: dout <= 8'b00010111; // 6488 :  23 - 0x17
      13'h1959: dout <= 8'b00101111; // 6489 :  47 - 0x2f
      13'h195A: dout <= 8'b00101111; // 6490 :  47 - 0x2f
      13'h195B: dout <= 8'b01011111; // 6491 :  95 - 0x5f
      13'h195C: dout <= 8'b01011111; // 6492 :  95 - 0x5f
      13'h195D: dout <= 8'b10111111; // 6493 : 191 - 0xbf
      13'h195E: dout <= 8'b10111111; // 6494 : 191 - 0xbf
      13'h195F: dout <= 8'b01111111; // 6495 : 127 - 0x7f
      13'h1960: dout <= 8'b00001111; // 6496 :  15 - 0xf -- Background 0x96
      13'h1961: dout <= 8'b00001111; // 6497 :  15 - 0xf
      13'h1962: dout <= 8'b10000111; // 6498 : 135 - 0x87
      13'h1963: dout <= 8'b10000111; // 6499 : 135 - 0x87
      13'h1964: dout <= 8'b11000010; // 6500 : 194 - 0xc2
      13'h1965: dout <= 8'b11000010; // 6501 : 194 - 0xc2
      13'h1966: dout <= 8'b11100000; // 6502 : 224 - 0xe0
      13'h1967: dout <= 8'b11100000; // 6503 : 224 - 0xe0
      13'h1968: dout <= 8'b01100000; // 6504 :  96 - 0x60
      13'h1969: dout <= 8'b01100000; // 6505 :  96 - 0x60
      13'h196A: dout <= 8'b10110000; // 6506 : 176 - 0xb0
      13'h196B: dout <= 8'b10110000; // 6507 : 176 - 0xb0
      13'h196C: dout <= 8'b11011000; // 6508 : 216 - 0xd8
      13'h196D: dout <= 8'b11011000; // 6509 : 216 - 0xd8
      13'h196E: dout <= 8'b11101100; // 6510 : 236 - 0xec
      13'h196F: dout <= 8'b11101100; // 6511 : 236 - 0xec
      13'h1970: dout <= 8'b10000011; // 6512 : 131 - 0x83 -- Background 0x97
      13'h1971: dout <= 8'b10001111; // 6513 : 143 - 0x8f
      13'h1972: dout <= 8'b00001111; // 6514 :  15 - 0xf
      13'h1973: dout <= 8'b00011111; // 6515 :  31 - 0x1f
      13'h1974: dout <= 8'b00011111; // 6516 :  31 - 0x1f
      13'h1975: dout <= 8'b00111111; // 6517 :  63 - 0x3f
      13'h1976: dout <= 8'b00111111; // 6518 :  63 - 0x3f
      13'h1977: dout <= 8'b00111111; // 6519 :  63 - 0x3f
      13'h1978: dout <= 8'b00110011; // 6520 :  51 - 0x33
      13'h1979: dout <= 8'b00101111; // 6521 :  47 - 0x2f
      13'h197A: dout <= 8'b01101111; // 6522 : 111 - 0x6f
      13'h197B: dout <= 8'b01011111; // 6523 :  95 - 0x5f
      13'h197C: dout <= 8'b11011111; // 6524 : 223 - 0xdf
      13'h197D: dout <= 8'b10111111; // 6525 : 191 - 0xbf
      13'h197E: dout <= 8'b10111111; // 6526 : 191 - 0xbf
      13'h197F: dout <= 8'b10111111; // 6527 : 191 - 0xbf
      13'h1980: dout <= 8'b11111111; // 6528 : 255 - 0xff -- Background 0x98
      13'h1981: dout <= 8'b11111111; // 6529 : 255 - 0xff
      13'h1982: dout <= 8'b11111111; // 6530 : 255 - 0xff
      13'h1983: dout <= 8'b11111110; // 6531 : 254 - 0xfe
      13'h1984: dout <= 8'b11111001; // 6532 : 249 - 0xf9
      13'h1985: dout <= 8'b11100111; // 6533 : 231 - 0xe7
      13'h1986: dout <= 8'b11111100; // 6534 : 252 - 0xfc
      13'h1987: dout <= 8'b11110000; // 6535 : 240 - 0xf0
      13'h1988: dout <= 8'b11111111; // 6536 : 255 - 0xff
      13'h1989: dout <= 8'b11111111; // 6537 : 255 - 0xff
      13'h198A: dout <= 8'b11111111; // 6538 : 255 - 0xff
      13'h198B: dout <= 8'b11111110; // 6539 : 254 - 0xfe
      13'h198C: dout <= 8'b11111001; // 6540 : 249 - 0xf9
      13'h198D: dout <= 8'b11100111; // 6541 : 231 - 0xe7
      13'h198E: dout <= 8'b11111100; // 6542 : 252 - 0xfc
      13'h198F: dout <= 8'b11110011; // 6543 : 243 - 0xf3
      13'h1990: dout <= 8'b11110111; // 6544 : 247 - 0xf7 -- Background 0x99
      13'h1991: dout <= 8'b11111011; // 6545 : 251 - 0xfb
      13'h1992: dout <= 8'b11111011; // 6546 : 251 - 0xfb
      13'h1993: dout <= 8'b01110011; // 6547 : 115 - 0x73
      13'h1994: dout <= 8'b11000001; // 6548 : 193 - 0xc1
      13'h1995: dout <= 8'b00000011; // 6549 :   3 - 0x3
      13'h1996: dout <= 8'b00001111; // 6550 :  15 - 0xf
      13'h1997: dout <= 8'b00111111; // 6551 :  63 - 0x3f
      13'h1998: dout <= 8'b11110000; // 6552 : 240 - 0xf0
      13'h1999: dout <= 8'b11111000; // 6553 : 248 - 0xf8
      13'h199A: dout <= 8'b11111000; // 6554 : 248 - 0xf8
      13'h199B: dout <= 8'b01110000; // 6555 : 112 - 0x70
      13'h199C: dout <= 8'b11001100; // 6556 : 204 - 0xcc
      13'h199D: dout <= 8'b00110000; // 6557 :  48 - 0x30
      13'h199E: dout <= 8'b11000000; // 6558 : 192 - 0xc0
      13'h199F: dout <= 8'b00000000; // 6559 :   0 - 0x0
      13'h19A0: dout <= 8'b11111111; // 6560 : 255 - 0xff -- Background 0x9a
      13'h19A1: dout <= 8'b11111111; // 6561 : 255 - 0xff
      13'h19A2: dout <= 8'b11111111; // 6562 : 255 - 0xff
      13'h19A3: dout <= 8'b10000000; // 6563 : 128 - 0x80
      13'h19A4: dout <= 8'b10000000; // 6564 : 128 - 0x80
      13'h19A5: dout <= 8'b10000000; // 6565 : 128 - 0x80
      13'h19A6: dout <= 8'b10001111; // 6566 : 143 - 0x8f
      13'h19A7: dout <= 8'b10001111; // 6567 : 143 - 0x8f
      13'h19A8: dout <= 8'b00000000; // 6568 :   0 - 0x0
      13'h19A9: dout <= 8'b00000000; // 6569 :   0 - 0x0
      13'h19AA: dout <= 8'b00000000; // 6570 :   0 - 0x0
      13'h19AB: dout <= 8'b00000000; // 6571 :   0 - 0x0
      13'h19AC: dout <= 8'b00111111; // 6572 :  63 - 0x3f
      13'h19AD: dout <= 8'b00100000; // 6573 :  32 - 0x20
      13'h19AE: dout <= 8'b00101111; // 6574 :  47 - 0x2f
      13'h19AF: dout <= 8'b00101111; // 6575 :  47 - 0x2f
      13'h19B0: dout <= 8'b11111111; // 6576 : 255 - 0xff -- Background 0x9b
      13'h19B1: dout <= 8'b11111111; // 6577 : 255 - 0xff
      13'h19B2: dout <= 8'b11111111; // 6578 : 255 - 0xff
      13'h19B3: dout <= 8'b00001111; // 6579 :  15 - 0xf
      13'h19B4: dout <= 8'b00001111; // 6580 :  15 - 0xf
      13'h19B5: dout <= 8'b00000111; // 6581 :   7 - 0x7
      13'h19B6: dout <= 8'b11110111; // 6582 : 247 - 0xf7
      13'h19B7: dout <= 8'b11110001; // 6583 : 241 - 0xf1
      13'h19B8: dout <= 8'b00000000; // 6584 :   0 - 0x0
      13'h19B9: dout <= 8'b00000000; // 6585 :   0 - 0x0
      13'h19BA: dout <= 8'b00000000; // 6586 :   0 - 0x0
      13'h19BB: dout <= 8'b00000000; // 6587 :   0 - 0x0
      13'h19BC: dout <= 8'b11100000; // 6588 : 224 - 0xe0
      13'h19BD: dout <= 8'b00000000; // 6589 :   0 - 0x0
      13'h19BE: dout <= 8'b11110000; // 6590 : 240 - 0xf0
      13'h19BF: dout <= 8'b11110000; // 6591 : 240 - 0xf0
      13'h19C0: dout <= 8'b00011100; // 6592 :  28 - 0x1c -- Background 0x9c
      13'h19C1: dout <= 8'b00011110; // 6593 :  30 - 0x1e
      13'h19C2: dout <= 8'b00011111; // 6594 :  31 - 0x1f
      13'h19C3: dout <= 8'b00011111; // 6595 :  31 - 0x1f
      13'h19C4: dout <= 8'b00011111; // 6596 :  31 - 0x1f
      13'h19C5: dout <= 8'b00011111; // 6597 :  31 - 0x1f
      13'h19C6: dout <= 8'b00011111; // 6598 :  31 - 0x1f
      13'h19C7: dout <= 8'b00011111; // 6599 :  31 - 0x1f
      13'h19C8: dout <= 8'b01011101; // 6600 :  93 - 0x5d
      13'h19C9: dout <= 8'b01011110; // 6601 :  94 - 0x5e
      13'h19CA: dout <= 8'b01011111; // 6602 :  95 - 0x5f
      13'h19CB: dout <= 8'b01011111; // 6603 :  95 - 0x5f
      13'h19CC: dout <= 8'b01011111; // 6604 :  95 - 0x5f
      13'h19CD: dout <= 8'b01011111; // 6605 :  95 - 0x5f
      13'h19CE: dout <= 8'b01011111; // 6606 :  95 - 0x5f
      13'h19CF: dout <= 8'b01011111; // 6607 :  95 - 0x5f
      13'h19D0: dout <= 8'b00111110; // 6608 :  62 - 0x3e -- Background 0x9d
      13'h19D1: dout <= 8'b00011100; // 6609 :  28 - 0x1c
      13'h19D2: dout <= 8'b00001000; // 6610 :   8 - 0x8
      13'h19D3: dout <= 8'b10000000; // 6611 : 128 - 0x80
      13'h19D4: dout <= 8'b11000001; // 6612 : 193 - 0xc1
      13'h19D5: dout <= 8'b11100011; // 6613 : 227 - 0xe3
      13'h19D6: dout <= 8'b11110111; // 6614 : 247 - 0xf7
      13'h19D7: dout <= 8'b11111111; // 6615 : 255 - 0xff
      13'h19D8: dout <= 8'b10000000; // 6616 : 128 - 0x80
      13'h19D9: dout <= 8'b11000001; // 6617 : 193 - 0xc1
      13'h19DA: dout <= 8'b01100011; // 6618 :  99 - 0x63
      13'h19DB: dout <= 8'b10110110; // 6619 : 182 - 0xb6
      13'h19DC: dout <= 8'b11011001; // 6620 : 217 - 0xd9
      13'h19DD: dout <= 8'b11101011; // 6621 : 235 - 0xeb
      13'h19DE: dout <= 8'b11110111; // 6622 : 247 - 0xf7
      13'h19DF: dout <= 8'b11111111; // 6623 : 255 - 0xff
      13'h19E0: dout <= 8'b00011100; // 6624 :  28 - 0x1c -- Background 0x9e
      13'h19E1: dout <= 8'b00111100; // 6625 :  60 - 0x3c
      13'h19E2: dout <= 8'b01111100; // 6626 : 124 - 0x7c
      13'h19E3: dout <= 8'b11111100; // 6627 : 252 - 0xfc
      13'h19E4: dout <= 8'b11111100; // 6628 : 252 - 0xfc
      13'h19E5: dout <= 8'b11111100; // 6629 : 252 - 0xfc
      13'h19E6: dout <= 8'b11111100; // 6630 : 252 - 0xfc
      13'h19E7: dout <= 8'b11111100; // 6631 : 252 - 0xfc
      13'h19E8: dout <= 8'b11011101; // 6632 : 221 - 0xdd
      13'h19E9: dout <= 8'b10111101; // 6633 : 189 - 0xbd
      13'h19EA: dout <= 8'b01111101; // 6634 : 125 - 0x7d
      13'h19EB: dout <= 8'b11111101; // 6635 : 253 - 0xfd
      13'h19EC: dout <= 8'b11111101; // 6636 : 253 - 0xfd
      13'h19ED: dout <= 8'b11111101; // 6637 : 253 - 0xfd
      13'h19EE: dout <= 8'b11111101; // 6638 : 253 - 0xfd
      13'h19EF: dout <= 8'b11111101; // 6639 : 253 - 0xfd
      13'h19F0: dout <= 8'b01111100; // 6640 : 124 - 0x7c -- Background 0x9f
      13'h19F1: dout <= 8'b01111100; // 6641 : 124 - 0x7c
      13'h19F2: dout <= 8'b01111000; // 6642 : 120 - 0x78
      13'h19F3: dout <= 8'b01111000; // 6643 : 120 - 0x78
      13'h19F4: dout <= 8'b01110001; // 6644 : 113 - 0x71
      13'h19F5: dout <= 8'b01110001; // 6645 : 113 - 0x71
      13'h19F6: dout <= 8'b01100011; // 6646 :  99 - 0x63
      13'h19F7: dout <= 8'b01100011; // 6647 :  99 - 0x63
      13'h19F8: dout <= 8'b00000001; // 6648 :   1 - 0x1
      13'h19F9: dout <= 8'b00000001; // 6649 :   1 - 0x1
      13'h19FA: dout <= 8'b00000010; // 6650 :   2 - 0x2
      13'h19FB: dout <= 8'b00000010; // 6651 :   2 - 0x2
      13'h19FC: dout <= 8'b00000101; // 6652 :   5 - 0x5
      13'h19FD: dout <= 8'b00000101; // 6653 :   5 - 0x5
      13'h19FE: dout <= 8'b00001011; // 6654 :  11 - 0xb
      13'h19FF: dout <= 8'b00001011; // 6655 :  11 - 0xb
      13'h1A00: dout <= 8'b01110001; // 6656 : 113 - 0x71 -- Background 0xa0
      13'h1A01: dout <= 8'b01110000; // 6657 : 112 - 0x70
      13'h1A02: dout <= 8'b11111000; // 6658 : 248 - 0xf8
      13'h1A03: dout <= 8'b11111000; // 6659 : 248 - 0xf8
      13'h1A04: dout <= 8'b11111100; // 6660 : 252 - 0xfc
      13'h1A05: dout <= 8'b11111100; // 6661 : 252 - 0xfc
      13'h1A06: dout <= 8'b11111110; // 6662 : 254 - 0xfe
      13'h1A07: dout <= 8'b11111110; // 6663 : 254 - 0xfe
      13'h1A08: dout <= 8'b01110100; // 6664 : 116 - 0x74
      13'h1A09: dout <= 8'b01110110; // 6665 : 118 - 0x76
      13'h1A0A: dout <= 8'b11111010; // 6666 : 250 - 0xfa
      13'h1A0B: dout <= 8'b11111011; // 6667 : 251 - 0xfb
      13'h1A0C: dout <= 8'b11111101; // 6668 : 253 - 0xfd
      13'h1A0D: dout <= 8'b11111101; // 6669 : 253 - 0xfd
      13'h1A0E: dout <= 8'b11111110; // 6670 : 254 - 0xfe
      13'h1A0F: dout <= 8'b11111110; // 6671 : 254 - 0xfe
      13'h1A10: dout <= 8'b11111000; // 6672 : 248 - 0xf8 -- Background 0xa1
      13'h1A11: dout <= 8'b11111000; // 6673 : 248 - 0xf8
      13'h1A12: dout <= 8'b11111000; // 6674 : 248 - 0xf8
      13'h1A13: dout <= 8'b01111000; // 6675 : 120 - 0x78
      13'h1A14: dout <= 8'b01111000; // 6676 : 120 - 0x78
      13'h1A15: dout <= 8'b00111000; // 6677 :  56 - 0x38
      13'h1A16: dout <= 8'b00111000; // 6678 :  56 - 0x38
      13'h1A17: dout <= 8'b00011000; // 6679 :  24 - 0x18
      13'h1A18: dout <= 8'b00000010; // 6680 :   2 - 0x2
      13'h1A19: dout <= 8'b00000010; // 6681 :   2 - 0x2
      13'h1A1A: dout <= 8'b00000010; // 6682 :   2 - 0x2
      13'h1A1B: dout <= 8'b00000010; // 6683 :   2 - 0x2
      13'h1A1C: dout <= 8'b00000010; // 6684 :   2 - 0x2
      13'h1A1D: dout <= 8'b10000010; // 6685 : 130 - 0x82
      13'h1A1E: dout <= 8'b10000010; // 6686 : 130 - 0x82
      13'h1A1F: dout <= 8'b11000010; // 6687 : 194 - 0xc2
      13'h1A20: dout <= 8'b11100000; // 6688 : 224 - 0xe0 -- Background 0xa2
      13'h1A21: dout <= 8'b11110000; // 6689 : 240 - 0xf0
      13'h1A22: dout <= 8'b11111000; // 6690 : 248 - 0xf8
      13'h1A23: dout <= 8'b11111000; // 6691 : 248 - 0xf8
      13'h1A24: dout <= 8'b11111100; // 6692 : 252 - 0xfc
      13'h1A25: dout <= 8'b11111100; // 6693 : 252 - 0xfc
      13'h1A26: dout <= 8'b11111110; // 6694 : 254 - 0xfe
      13'h1A27: dout <= 8'b11111111; // 6695 : 255 - 0xff
      13'h1A28: dout <= 8'b11101010; // 6696 : 234 - 0xea
      13'h1A29: dout <= 8'b11110110; // 6697 : 246 - 0xf6
      13'h1A2A: dout <= 8'b11111010; // 6698 : 250 - 0xfa
      13'h1A2B: dout <= 8'b11111010; // 6699 : 250 - 0xfa
      13'h1A2C: dout <= 8'b11111100; // 6700 : 252 - 0xfc
      13'h1A2D: dout <= 8'b11111100; // 6701 : 252 - 0xfc
      13'h1A2E: dout <= 8'b11111110; // 6702 : 254 - 0xfe
      13'h1A2F: dout <= 8'b11111111; // 6703 : 255 - 0xff
      13'h1A30: dout <= 8'b11111111; // 6704 : 255 - 0xff -- Background 0xa3
      13'h1A31: dout <= 8'b11111111; // 6705 : 255 - 0xff
      13'h1A32: dout <= 8'b11111111; // 6706 : 255 - 0xff
      13'h1A33: dout <= 8'b11111111; // 6707 : 255 - 0xff
      13'h1A34: dout <= 8'b11111111; // 6708 : 255 - 0xff
      13'h1A35: dout <= 8'b11111111; // 6709 : 255 - 0xff
      13'h1A36: dout <= 8'b11111111; // 6710 : 255 - 0xff
      13'h1A37: dout <= 8'b11111111; // 6711 : 255 - 0xff
      13'h1A38: dout <= 8'b11111111; // 6712 : 255 - 0xff
      13'h1A39: dout <= 8'b11111111; // 6713 : 255 - 0xff
      13'h1A3A: dout <= 8'b11111111; // 6714 : 255 - 0xff
      13'h1A3B: dout <= 8'b11111111; // 6715 : 255 - 0xff
      13'h1A3C: dout <= 8'b11111111; // 6716 : 255 - 0xff
      13'h1A3D: dout <= 8'b11111111; // 6717 : 255 - 0xff
      13'h1A3E: dout <= 8'b11111111; // 6718 : 255 - 0xff
      13'h1A3F: dout <= 8'b11111111; // 6719 : 255 - 0xff
      13'h1A40: dout <= 8'b00011111; // 6720 :  31 - 0x1f -- Background 0xa4
      13'h1A41: dout <= 8'b00011111; // 6721 :  31 - 0x1f
      13'h1A42: dout <= 8'b00011111; // 6722 :  31 - 0x1f
      13'h1A43: dout <= 8'b00011111; // 6723 :  31 - 0x1f
      13'h1A44: dout <= 8'b00011111; // 6724 :  31 - 0x1f
      13'h1A45: dout <= 8'b00011111; // 6725 :  31 - 0x1f
      13'h1A46: dout <= 8'b00011111; // 6726 :  31 - 0x1f
      13'h1A47: dout <= 8'b00011111; // 6727 :  31 - 0x1f
      13'h1A48: dout <= 8'b01000000; // 6728 :  64 - 0x40
      13'h1A49: dout <= 8'b01000000; // 6729 :  64 - 0x40
      13'h1A4A: dout <= 8'b01000000; // 6730 :  64 - 0x40
      13'h1A4B: dout <= 8'b01000000; // 6731 :  64 - 0x40
      13'h1A4C: dout <= 8'b01000000; // 6732 :  64 - 0x40
      13'h1A4D: dout <= 8'b01000000; // 6733 :  64 - 0x40
      13'h1A4E: dout <= 8'b01000000; // 6734 :  64 - 0x40
      13'h1A4F: dout <= 8'b01000000; // 6735 :  64 - 0x40
      13'h1A50: dout <= 8'b11111000; // 6736 : 248 - 0xf8 -- Background 0xa5
      13'h1A51: dout <= 8'b11111111; // 6737 : 255 - 0xff
      13'h1A52: dout <= 8'b11111111; // 6738 : 255 - 0xff
      13'h1A53: dout <= 8'b11111000; // 6739 : 248 - 0xf8
      13'h1A54: dout <= 8'b11111000; // 6740 : 248 - 0xf8
      13'h1A55: dout <= 8'b11111000; // 6741 : 248 - 0xf8
      13'h1A56: dout <= 8'b11111000; // 6742 : 248 - 0xf8
      13'h1A57: dout <= 8'b11111000; // 6743 : 248 - 0xf8
      13'h1A58: dout <= 8'b11111000; // 6744 : 248 - 0xf8
      13'h1A59: dout <= 8'b11111111; // 6745 : 255 - 0xff
      13'h1A5A: dout <= 8'b11111111; // 6746 : 255 - 0xff
      13'h1A5B: dout <= 8'b11111000; // 6747 : 248 - 0xf8
      13'h1A5C: dout <= 8'b11111011; // 6748 : 251 - 0xfb
      13'h1A5D: dout <= 8'b11111010; // 6749 : 250 - 0xfa
      13'h1A5E: dout <= 8'b11111010; // 6750 : 250 - 0xfa
      13'h1A5F: dout <= 8'b11111010; // 6751 : 250 - 0xfa
      13'h1A60: dout <= 8'b11111100; // 6752 : 252 - 0xfc -- Background 0xa6
      13'h1A61: dout <= 8'b11111000; // 6753 : 248 - 0xf8
      13'h1A62: dout <= 8'b11110000; // 6754 : 240 - 0xf0
      13'h1A63: dout <= 8'b00000001; // 6755 :   1 - 0x1
      13'h1A64: dout <= 8'b00000001; // 6756 :   1 - 0x1
      13'h1A65: dout <= 8'b00000011; // 6757 :   3 - 0x3
      13'h1A66: dout <= 8'b11000011; // 6758 : 195 - 0xc3
      13'h1A67: dout <= 8'b10000111; // 6759 : 135 - 0x87
      13'h1A68: dout <= 8'b11111100; // 6760 : 252 - 0xfc
      13'h1A69: dout <= 8'b11111010; // 6761 : 250 - 0xfa
      13'h1A6A: dout <= 8'b11110110; // 6762 : 246 - 0xf6
      13'h1A6B: dout <= 8'b00001101; // 6763 :  13 - 0xd
      13'h1A6C: dout <= 8'b11111001; // 6764 : 249 - 0xf9
      13'h1A6D: dout <= 8'b00000011; // 6765 :   3 - 0x3
      13'h1A6E: dout <= 8'b00010011; // 6766 :  19 - 0x13
      13'h1A6F: dout <= 8'b00110111; // 6767 :  55 - 0x37
      13'h1A70: dout <= 8'b01111111; // 6768 : 127 - 0x7f -- Background 0xa7
      13'h1A71: dout <= 8'b11111001; // 6769 : 249 - 0xf9
      13'h1A72: dout <= 8'b11111001; // 6770 : 249 - 0xf9
      13'h1A73: dout <= 8'b11111111; // 6771 : 255 - 0xff
      13'h1A74: dout <= 8'b11111110; // 6772 : 254 - 0xfe
      13'h1A75: dout <= 8'b11111100; // 6773 : 252 - 0xfc
      13'h1A76: dout <= 8'b11111111; // 6774 : 255 - 0xff
      13'h1A77: dout <= 8'b11111111; // 6775 : 255 - 0xff
      13'h1A78: dout <= 8'b01111111; // 6776 : 127 - 0x7f
      13'h1A79: dout <= 8'b11111001; // 6777 : 249 - 0xf9
      13'h1A7A: dout <= 8'b11111001; // 6778 : 249 - 0xf9
      13'h1A7B: dout <= 8'b11111111; // 6779 : 255 - 0xff
      13'h1A7C: dout <= 8'b11111110; // 6780 : 254 - 0xfe
      13'h1A7D: dout <= 8'b11111100; // 6781 : 252 - 0xfc
      13'h1A7E: dout <= 8'b11111111; // 6782 : 255 - 0xff
      13'h1A7F: dout <= 8'b11111111; // 6783 : 255 - 0xff
      13'h1A80: dout <= 8'b11110000; // 6784 : 240 - 0xf0 -- Background 0xa8
      13'h1A81: dout <= 8'b11110000; // 6785 : 240 - 0xf0
      13'h1A82: dout <= 8'b11111000; // 6786 : 248 - 0xf8
      13'h1A83: dout <= 8'b01111000; // 6787 : 120 - 0x78
      13'h1A84: dout <= 8'b11111100; // 6788 : 252 - 0xfc
      13'h1A85: dout <= 8'b11110100; // 6789 : 244 - 0xf4
      13'h1A86: dout <= 8'b11110110; // 6790 : 246 - 0xf6
      13'h1A87: dout <= 8'b11111010; // 6791 : 250 - 0xfa
      13'h1A88: dout <= 8'b11110110; // 6792 : 246 - 0xf6
      13'h1A89: dout <= 8'b11110110; // 6793 : 246 - 0xf6
      13'h1A8A: dout <= 8'b11111011; // 6794 : 251 - 0xfb
      13'h1A8B: dout <= 8'b01111011; // 6795 : 123 - 0x7b
      13'h1A8C: dout <= 8'b11111101; // 6796 : 253 - 0xfd
      13'h1A8D: dout <= 8'b11110101; // 6797 : 245 - 0xf5
      13'h1A8E: dout <= 8'b11110110; // 6798 : 246 - 0xf6
      13'h1A8F: dout <= 8'b11111010; // 6799 : 250 - 0xfa
      13'h1A90: dout <= 8'b00111111; // 6800 :  63 - 0x3f -- Background 0xa9
      13'h1A91: dout <= 8'b00111111; // 6801 :  63 - 0x3f
      13'h1A92: dout <= 8'b00111111; // 6802 :  63 - 0x3f
      13'h1A93: dout <= 8'b00111111; // 6803 :  63 - 0x3f
      13'h1A94: dout <= 8'b00111111; // 6804 :  63 - 0x3f
      13'h1A95: dout <= 8'b00011111; // 6805 :  31 - 0x1f
      13'h1A96: dout <= 8'b00001111; // 6806 :  15 - 0xf
      13'h1A97: dout <= 8'b00000111; // 6807 :   7 - 0x7
      13'h1A98: dout <= 8'b10111111; // 6808 : 191 - 0xbf
      13'h1A99: dout <= 8'b10111111; // 6809 : 191 - 0xbf
      13'h1A9A: dout <= 8'b00111111; // 6810 :  63 - 0x3f
      13'h1A9B: dout <= 8'b00111111; // 6811 :  63 - 0x3f
      13'h1A9C: dout <= 8'b10111111; // 6812 : 191 - 0xbf
      13'h1A9D: dout <= 8'b10011111; // 6813 : 159 - 0x9f
      13'h1A9E: dout <= 8'b11001111; // 6814 : 207 - 0xcf
      13'h1A9F: dout <= 8'b11010111; // 6815 : 215 - 0xd7
      13'h1AA0: dout <= 8'b11100000; // 6816 : 224 - 0xe0 -- Background 0xaa
      13'h1AA1: dout <= 8'b11111000; // 6817 : 248 - 0xf8
      13'h1AA2: dout <= 8'b11111111; // 6818 : 255 - 0xff
      13'h1AA3: dout <= 8'b11110011; // 6819 : 243 - 0xf3
      13'h1AA4: dout <= 8'b11111100; // 6820 : 252 - 0xfc
      13'h1AA5: dout <= 8'b11111111; // 6821 : 255 - 0xff
      13'h1AA6: dout <= 8'b11111111; // 6822 : 255 - 0xff
      13'h1AA7: dout <= 8'b11111111; // 6823 : 255 - 0xff
      13'h1AA8: dout <= 8'b11100100; // 6824 : 228 - 0xe4
      13'h1AA9: dout <= 8'b11111000; // 6825 : 248 - 0xf8
      13'h1AAA: dout <= 8'b11111111; // 6826 : 255 - 0xff
      13'h1AAB: dout <= 8'b11110011; // 6827 : 243 - 0xf3
      13'h1AAC: dout <= 8'b11111100; // 6828 : 252 - 0xfc
      13'h1AAD: dout <= 8'b11111111; // 6829 : 255 - 0xff
      13'h1AAE: dout <= 8'b11111111; // 6830 : 255 - 0xff
      13'h1AAF: dout <= 8'b11111111; // 6831 : 255 - 0xff
      13'h1AB0: dout <= 8'b11111111; // 6832 : 255 - 0xff -- Background 0xab
      13'h1AB1: dout <= 8'b11111111; // 6833 : 255 - 0xff
      13'h1AB2: dout <= 8'b00111111; // 6834 :  63 - 0x3f
      13'h1AB3: dout <= 8'b11001111; // 6835 : 207 - 0xcf
      13'h1AB4: dout <= 8'b11110011; // 6836 : 243 - 0xf3
      13'h1AB5: dout <= 8'b00111101; // 6837 :  61 - 0x3d
      13'h1AB6: dout <= 8'b11011000; // 6838 : 216 - 0xd8
      13'h1AB7: dout <= 8'b10110000; // 6839 : 176 - 0xb0
      13'h1AB8: dout <= 8'b00000000; // 6840 :   0 - 0x0
      13'h1AB9: dout <= 8'b00000000; // 6841 :   0 - 0x0
      13'h1ABA: dout <= 8'b00000000; // 6842 :   0 - 0x0
      13'h1ABB: dout <= 8'b11000000; // 6843 : 192 - 0xc0
      13'h1ABC: dout <= 8'b11110000; // 6844 : 240 - 0xf0
      13'h1ABD: dout <= 8'b00111100; // 6845 :  60 - 0x3c
      13'h1ABE: dout <= 8'b11011000; // 6846 : 216 - 0xd8
      13'h1ABF: dout <= 8'b10110110; // 6847 : 182 - 0xb6
      13'h1AC0: dout <= 8'b10001111; // 6848 : 143 - 0x8f -- Background 0xac
      13'h1AC1: dout <= 8'b11101111; // 6849 : 239 - 0xef
      13'h1AC2: dout <= 8'b11100000; // 6850 : 224 - 0xe0
      13'h1AC3: dout <= 8'b11111000; // 6851 : 248 - 0xf8
      13'h1AC4: dout <= 8'b11111000; // 6852 : 248 - 0xf8
      13'h1AC5: dout <= 8'b11111111; // 6853 : 255 - 0xff
      13'h1AC6: dout <= 8'b11111111; // 6854 : 255 - 0xff
      13'h1AC7: dout <= 8'b11111111; // 6855 : 255 - 0xff
      13'h1AC8: dout <= 8'b00001111; // 6856 :  15 - 0xf
      13'h1AC9: dout <= 8'b00001111; // 6857 :  15 - 0xf
      13'h1ACA: dout <= 8'b00000000; // 6858 :   0 - 0x0
      13'h1ACB: dout <= 8'b00000011; // 6859 :   3 - 0x3
      13'h1ACC: dout <= 8'b00000000; // 6860 :   0 - 0x0
      13'h1ACD: dout <= 8'b00000000; // 6861 :   0 - 0x0
      13'h1ACE: dout <= 8'b00000000; // 6862 :   0 - 0x0
      13'h1ACF: dout <= 8'b00000000; // 6863 :   0 - 0x0
      13'h1AD0: dout <= 8'b11110001; // 6864 : 241 - 0xf1 -- Background 0xad
      13'h1AD1: dout <= 8'b11110001; // 6865 : 241 - 0xf1
      13'h1AD2: dout <= 8'b00000001; // 6866 :   1 - 0x1
      13'h1AD3: dout <= 8'b00000001; // 6867 :   1 - 0x1
      13'h1AD4: dout <= 8'b00000001; // 6868 :   1 - 0x1
      13'h1AD5: dout <= 8'b11111111; // 6869 : 255 - 0xff
      13'h1AD6: dout <= 8'b11111111; // 6870 : 255 - 0xff
      13'h1AD7: dout <= 8'b11111111; // 6871 : 255 - 0xff
      13'h1AD8: dout <= 8'b11110100; // 6872 : 244 - 0xf4
      13'h1AD9: dout <= 8'b11110100; // 6873 : 244 - 0xf4
      13'h1ADA: dout <= 8'b00000100; // 6874 :   4 - 0x4
      13'h1ADB: dout <= 8'b11111100; // 6875 : 252 - 0xfc
      13'h1ADC: dout <= 8'b00000000; // 6876 :   0 - 0x0
      13'h1ADD: dout <= 8'b00000000; // 6877 :   0 - 0x0
      13'h1ADE: dout <= 8'b00000000; // 6878 :   0 - 0x0
      13'h1ADF: dout <= 8'b00000000; // 6879 :   0 - 0x0
      13'h1AE0: dout <= 8'b00011111; // 6880 :  31 - 0x1f -- Background 0xae
      13'h1AE1: dout <= 8'b00011111; // 6881 :  31 - 0x1f
      13'h1AE2: dout <= 8'b00011111; // 6882 :  31 - 0x1f
      13'h1AE3: dout <= 8'b00011111; // 6883 :  31 - 0x1f
      13'h1AE4: dout <= 8'b00011111; // 6884 :  31 - 0x1f
      13'h1AE5: dout <= 8'b00011111; // 6885 :  31 - 0x1f
      13'h1AE6: dout <= 8'b00011111; // 6886 :  31 - 0x1f
      13'h1AE7: dout <= 8'b00011111; // 6887 :  31 - 0x1f
      13'h1AE8: dout <= 8'b01011111; // 6888 :  95 - 0x5f
      13'h1AE9: dout <= 8'b01011111; // 6889 :  95 - 0x5f
      13'h1AEA: dout <= 8'b01011111; // 6890 :  95 - 0x5f
      13'h1AEB: dout <= 8'b01011111; // 6891 :  95 - 0x5f
      13'h1AEC: dout <= 8'b01011111; // 6892 :  95 - 0x5f
      13'h1AED: dout <= 8'b01011111; // 6893 :  95 - 0x5f
      13'h1AEE: dout <= 8'b01011111; // 6894 :  95 - 0x5f
      13'h1AEF: dout <= 8'b01011111; // 6895 :  95 - 0x5f
      13'h1AF0: dout <= 8'b11111100; // 6896 : 252 - 0xfc -- Background 0xaf
      13'h1AF1: dout <= 8'b11111100; // 6897 : 252 - 0xfc
      13'h1AF2: dout <= 8'b11111100; // 6898 : 252 - 0xfc
      13'h1AF3: dout <= 8'b11111100; // 6899 : 252 - 0xfc
      13'h1AF4: dout <= 8'b11110100; // 6900 : 244 - 0xf4
      13'h1AF5: dout <= 8'b11110100; // 6901 : 244 - 0xf4
      13'h1AF6: dout <= 8'b11110100; // 6902 : 244 - 0xf4
      13'h1AF7: dout <= 8'b11110100; // 6903 : 244 - 0xf4
      13'h1AF8: dout <= 8'b11111101; // 6904 : 253 - 0xfd
      13'h1AF9: dout <= 8'b11111101; // 6905 : 253 - 0xfd
      13'h1AFA: dout <= 8'b11111101; // 6906 : 253 - 0xfd
      13'h1AFB: dout <= 8'b11111101; // 6907 : 253 - 0xfd
      13'h1AFC: dout <= 8'b11110101; // 6908 : 245 - 0xf5
      13'h1AFD: dout <= 8'b11110101; // 6909 : 245 - 0xf5
      13'h1AFE: dout <= 8'b11110101; // 6910 : 245 - 0xf5
      13'h1AFF: dout <= 8'b11110101; // 6911 : 245 - 0xf5
      13'h1B00: dout <= 8'b00001100; // 6912 :  12 - 0xc -- Background 0xb0
      13'h1B01: dout <= 8'b00011100; // 6913 :  28 - 0x1c
      13'h1B02: dout <= 8'b00001100; // 6914 :  12 - 0xc
      13'h1B03: dout <= 8'b00001100; // 6915 :  12 - 0xc
      13'h1B04: dout <= 8'b00001100; // 6916 :  12 - 0xc
      13'h1B05: dout <= 8'b00001100; // 6917 :  12 - 0xc
      13'h1B06: dout <= 8'b00111111; // 6918 :  63 - 0x3f
      13'h1B07: dout <= 8'b00000000; // 6919 :   0 - 0x0
      13'h1B08: dout <= 8'b00001100; // 6920 :  12 - 0xc
      13'h1B09: dout <= 8'b00011100; // 6921 :  28 - 0x1c
      13'h1B0A: dout <= 8'b00001100; // 6922 :  12 - 0xc
      13'h1B0B: dout <= 8'b00001100; // 6923 :  12 - 0xc
      13'h1B0C: dout <= 8'b00001100; // 6924 :  12 - 0xc
      13'h1B0D: dout <= 8'b00001100; // 6925 :  12 - 0xc
      13'h1B0E: dout <= 8'b00111111; // 6926 :  63 - 0x3f
      13'h1B0F: dout <= 8'b00000000; // 6927 :   0 - 0x0
      13'h1B10: dout <= 8'b00111110; // 6928 :  62 - 0x3e -- Background 0xb1
      13'h1B11: dout <= 8'b01100011; // 6929 :  99 - 0x63
      13'h1B12: dout <= 8'b00000111; // 6930 :   7 - 0x7
      13'h1B13: dout <= 8'b00011110; // 6931 :  30 - 0x1e
      13'h1B14: dout <= 8'b00111100; // 6932 :  60 - 0x3c
      13'h1B15: dout <= 8'b01110000; // 6933 : 112 - 0x70
      13'h1B16: dout <= 8'b01111111; // 6934 : 127 - 0x7f
      13'h1B17: dout <= 8'b00000000; // 6935 :   0 - 0x0
      13'h1B18: dout <= 8'b00111110; // 6936 :  62 - 0x3e
      13'h1B19: dout <= 8'b01100011; // 6937 :  99 - 0x63
      13'h1B1A: dout <= 8'b00000111; // 6938 :   7 - 0x7
      13'h1B1B: dout <= 8'b00011110; // 6939 :  30 - 0x1e
      13'h1B1C: dout <= 8'b00111100; // 6940 :  60 - 0x3c
      13'h1B1D: dout <= 8'b01110000; // 6941 : 112 - 0x70
      13'h1B1E: dout <= 8'b01111111; // 6942 : 127 - 0x7f
      13'h1B1F: dout <= 8'b00000000; // 6943 :   0 - 0x0
      13'h1B20: dout <= 8'b01111110; // 6944 : 126 - 0x7e -- Background 0xb2
      13'h1B21: dout <= 8'b01100011; // 6945 :  99 - 0x63
      13'h1B22: dout <= 8'b01100011; // 6946 :  99 - 0x63
      13'h1B23: dout <= 8'b01100011; // 6947 :  99 - 0x63
      13'h1B24: dout <= 8'b01111110; // 6948 : 126 - 0x7e
      13'h1B25: dout <= 8'b01100000; // 6949 :  96 - 0x60
      13'h1B26: dout <= 8'b01100000; // 6950 :  96 - 0x60
      13'h1B27: dout <= 8'b00000000; // 6951 :   0 - 0x0
      13'h1B28: dout <= 8'b01111110; // 6952 : 126 - 0x7e
      13'h1B29: dout <= 8'b01100011; // 6953 :  99 - 0x63
      13'h1B2A: dout <= 8'b01100011; // 6954 :  99 - 0x63
      13'h1B2B: dout <= 8'b01100011; // 6955 :  99 - 0x63
      13'h1B2C: dout <= 8'b01111110; // 6956 : 126 - 0x7e
      13'h1B2D: dout <= 8'b01100000; // 6957 :  96 - 0x60
      13'h1B2E: dout <= 8'b01100000; // 6958 :  96 - 0x60
      13'h1B2F: dout <= 8'b00000000; // 6959 :   0 - 0x0
      13'h1B30: dout <= 8'b01100011; // 6960 :  99 - 0x63 -- Background 0xb3
      13'h1B31: dout <= 8'b01100011; // 6961 :  99 - 0x63
      13'h1B32: dout <= 8'b01100011; // 6962 :  99 - 0x63
      13'h1B33: dout <= 8'b01100011; // 6963 :  99 - 0x63
      13'h1B34: dout <= 8'b01100011; // 6964 :  99 - 0x63
      13'h1B35: dout <= 8'b01100011; // 6965 :  99 - 0x63
      13'h1B36: dout <= 8'b00111110; // 6966 :  62 - 0x3e
      13'h1B37: dout <= 8'b00000000; // 6967 :   0 - 0x0
      13'h1B38: dout <= 8'b01100011; // 6968 :  99 - 0x63
      13'h1B39: dout <= 8'b01100011; // 6969 :  99 - 0x63
      13'h1B3A: dout <= 8'b01100011; // 6970 :  99 - 0x63
      13'h1B3B: dout <= 8'b01100011; // 6971 :  99 - 0x63
      13'h1B3C: dout <= 8'b01100011; // 6972 :  99 - 0x63
      13'h1B3D: dout <= 8'b01100011; // 6973 :  99 - 0x63
      13'h1B3E: dout <= 8'b00111110; // 6974 :  62 - 0x3e
      13'h1B3F: dout <= 8'b00000000; // 6975 :   0 - 0x0
      13'h1B40: dout <= 8'b01100011; // 6976 :  99 - 0x63 -- Background 0xb4
      13'h1B41: dout <= 8'b01100011; // 6977 :  99 - 0x63
      13'h1B42: dout <= 8'b01100011; // 6978 :  99 - 0x63
      13'h1B43: dout <= 8'b01111111; // 6979 : 127 - 0x7f
      13'h1B44: dout <= 8'b01100011; // 6980 :  99 - 0x63
      13'h1B45: dout <= 8'b01100011; // 6981 :  99 - 0x63
      13'h1B46: dout <= 8'b01100011; // 6982 :  99 - 0x63
      13'h1B47: dout <= 8'b00000000; // 6983 :   0 - 0x0
      13'h1B48: dout <= 8'b01100011; // 6984 :  99 - 0x63
      13'h1B49: dout <= 8'b01100011; // 6985 :  99 - 0x63
      13'h1B4A: dout <= 8'b01100011; // 6986 :  99 - 0x63
      13'h1B4B: dout <= 8'b01111111; // 6987 : 127 - 0x7f
      13'h1B4C: dout <= 8'b01100011; // 6988 :  99 - 0x63
      13'h1B4D: dout <= 8'b01100011; // 6989 :  99 - 0x63
      13'h1B4E: dout <= 8'b01100011; // 6990 :  99 - 0x63
      13'h1B4F: dout <= 8'b00000000; // 6991 :   0 - 0x0
      13'h1B50: dout <= 8'b00111111; // 6992 :  63 - 0x3f -- Background 0xb5
      13'h1B51: dout <= 8'b00001100; // 6993 :  12 - 0xc
      13'h1B52: dout <= 8'b00001100; // 6994 :  12 - 0xc
      13'h1B53: dout <= 8'b00001100; // 6995 :  12 - 0xc
      13'h1B54: dout <= 8'b00001100; // 6996 :  12 - 0xc
      13'h1B55: dout <= 8'b00001100; // 6997 :  12 - 0xc
      13'h1B56: dout <= 8'b00111111; // 6998 :  63 - 0x3f
      13'h1B57: dout <= 8'b00000000; // 6999 :   0 - 0x0
      13'h1B58: dout <= 8'b00111111; // 7000 :  63 - 0x3f
      13'h1B59: dout <= 8'b00001100; // 7001 :  12 - 0xc
      13'h1B5A: dout <= 8'b00001100; // 7002 :  12 - 0xc
      13'h1B5B: dout <= 8'b00001100; // 7003 :  12 - 0xc
      13'h1B5C: dout <= 8'b00001100; // 7004 :  12 - 0xc
      13'h1B5D: dout <= 8'b00001100; // 7005 :  12 - 0xc
      13'h1B5E: dout <= 8'b00111111; // 7006 :  63 - 0x3f
      13'h1B5F: dout <= 8'b00000000; // 7007 :   0 - 0x0
      13'h1B60: dout <= 8'b00000000; // 7008 :   0 - 0x0 -- Background 0xb6
      13'h1B61: dout <= 8'b00000000; // 7009 :   0 - 0x0
      13'h1B62: dout <= 8'b00000000; // 7010 :   0 - 0x0
      13'h1B63: dout <= 8'b01111110; // 7011 : 126 - 0x7e
      13'h1B64: dout <= 8'b00000000; // 7012 :   0 - 0x0
      13'h1B65: dout <= 8'b00000000; // 7013 :   0 - 0x0
      13'h1B66: dout <= 8'b00000000; // 7014 :   0 - 0x0
      13'h1B67: dout <= 8'b00000000; // 7015 :   0 - 0x0
      13'h1B68: dout <= 8'b00000000; // 7016 :   0 - 0x0
      13'h1B69: dout <= 8'b00000000; // 7017 :   0 - 0x0
      13'h1B6A: dout <= 8'b00000000; // 7018 :   0 - 0x0
      13'h1B6B: dout <= 8'b01111110; // 7019 : 126 - 0x7e
      13'h1B6C: dout <= 8'b00000000; // 7020 :   0 - 0x0
      13'h1B6D: dout <= 8'b00000000; // 7021 :   0 - 0x0
      13'h1B6E: dout <= 8'b00000000; // 7022 :   0 - 0x0
      13'h1B6F: dout <= 8'b00000000; // 7023 :   0 - 0x0
      13'h1B70: dout <= 8'b00111100; // 7024 :  60 - 0x3c -- Background 0xb7
      13'h1B71: dout <= 8'b01100110; // 7025 : 102 - 0x66
      13'h1B72: dout <= 8'b01100000; // 7026 :  96 - 0x60
      13'h1B73: dout <= 8'b00111110; // 7027 :  62 - 0x3e
      13'h1B74: dout <= 8'b00000011; // 7028 :   3 - 0x3
      13'h1B75: dout <= 8'b01100011; // 7029 :  99 - 0x63
      13'h1B76: dout <= 8'b00111110; // 7030 :  62 - 0x3e
      13'h1B77: dout <= 8'b00000000; // 7031 :   0 - 0x0
      13'h1B78: dout <= 8'b00111100; // 7032 :  60 - 0x3c
      13'h1B79: dout <= 8'b01100110; // 7033 : 102 - 0x66
      13'h1B7A: dout <= 8'b01100000; // 7034 :  96 - 0x60
      13'h1B7B: dout <= 8'b00111110; // 7035 :  62 - 0x3e
      13'h1B7C: dout <= 8'b00000011; // 7036 :   3 - 0x3
      13'h1B7D: dout <= 8'b01100011; // 7037 :  99 - 0x63
      13'h1B7E: dout <= 8'b00111110; // 7038 :  62 - 0x3e
      13'h1B7F: dout <= 8'b00000000; // 7039 :   0 - 0x0
      13'h1B80: dout <= 8'b00011110; // 7040 :  30 - 0x1e -- Background 0xb8
      13'h1B81: dout <= 8'b00110011; // 7041 :  51 - 0x33
      13'h1B82: dout <= 8'b01100000; // 7042 :  96 - 0x60
      13'h1B83: dout <= 8'b01100000; // 7043 :  96 - 0x60
      13'h1B84: dout <= 8'b01100000; // 7044 :  96 - 0x60
      13'h1B85: dout <= 8'b00110011; // 7045 :  51 - 0x33
      13'h1B86: dout <= 8'b00011110; // 7046 :  30 - 0x1e
      13'h1B87: dout <= 8'b00000000; // 7047 :   0 - 0x0
      13'h1B88: dout <= 8'b00011110; // 7048 :  30 - 0x1e
      13'h1B89: dout <= 8'b00110011; // 7049 :  51 - 0x33
      13'h1B8A: dout <= 8'b01100000; // 7050 :  96 - 0x60
      13'h1B8B: dout <= 8'b01100000; // 7051 :  96 - 0x60
      13'h1B8C: dout <= 8'b01100000; // 7052 :  96 - 0x60
      13'h1B8D: dout <= 8'b00110011; // 7053 :  51 - 0x33
      13'h1B8E: dout <= 8'b00011110; // 7054 :  30 - 0x1e
      13'h1B8F: dout <= 8'b00000000; // 7055 :   0 - 0x0
      13'h1B90: dout <= 8'b00111110; // 7056 :  62 - 0x3e -- Background 0xb9
      13'h1B91: dout <= 8'b01100011; // 7057 :  99 - 0x63
      13'h1B92: dout <= 8'b01100011; // 7058 :  99 - 0x63
      13'h1B93: dout <= 8'b01100011; // 7059 :  99 - 0x63
      13'h1B94: dout <= 8'b01100011; // 7060 :  99 - 0x63
      13'h1B95: dout <= 8'b01100011; // 7061 :  99 - 0x63
      13'h1B96: dout <= 8'b00111110; // 7062 :  62 - 0x3e
      13'h1B97: dout <= 8'b00000000; // 7063 :   0 - 0x0
      13'h1B98: dout <= 8'b00111110; // 7064 :  62 - 0x3e
      13'h1B99: dout <= 8'b01100011; // 7065 :  99 - 0x63
      13'h1B9A: dout <= 8'b01100011; // 7066 :  99 - 0x63
      13'h1B9B: dout <= 8'b01100011; // 7067 :  99 - 0x63
      13'h1B9C: dout <= 8'b01100011; // 7068 :  99 - 0x63
      13'h1B9D: dout <= 8'b01100011; // 7069 :  99 - 0x63
      13'h1B9E: dout <= 8'b00111110; // 7070 :  62 - 0x3e
      13'h1B9F: dout <= 8'b00000000; // 7071 :   0 - 0x0
      13'h1BA0: dout <= 8'b01111110; // 7072 : 126 - 0x7e -- Background 0xba
      13'h1BA1: dout <= 8'b01100011; // 7073 :  99 - 0x63
      13'h1BA2: dout <= 8'b01100011; // 7074 :  99 - 0x63
      13'h1BA3: dout <= 8'b01100111; // 7075 : 103 - 0x67
      13'h1BA4: dout <= 8'b01111100; // 7076 : 124 - 0x7c
      13'h1BA5: dout <= 8'b01101110; // 7077 : 110 - 0x6e
      13'h1BA6: dout <= 8'b01100111; // 7078 : 103 - 0x67
      13'h1BA7: dout <= 8'b00000000; // 7079 :   0 - 0x0
      13'h1BA8: dout <= 8'b01111110; // 7080 : 126 - 0x7e
      13'h1BA9: dout <= 8'b01100011; // 7081 :  99 - 0x63
      13'h1BAA: dout <= 8'b01100011; // 7082 :  99 - 0x63
      13'h1BAB: dout <= 8'b01100111; // 7083 : 103 - 0x67
      13'h1BAC: dout <= 8'b01111100; // 7084 : 124 - 0x7c
      13'h1BAD: dout <= 8'b01101110; // 7085 : 110 - 0x6e
      13'h1BAE: dout <= 8'b01100111; // 7086 : 103 - 0x67
      13'h1BAF: dout <= 8'b00000000; // 7087 :   0 - 0x0
      13'h1BB0: dout <= 8'b01111111; // 7088 : 127 - 0x7f -- Background 0xbb
      13'h1BB1: dout <= 8'b01100000; // 7089 :  96 - 0x60
      13'h1BB2: dout <= 8'b01100000; // 7090 :  96 - 0x60
      13'h1BB3: dout <= 8'b01111110; // 7091 : 126 - 0x7e
      13'h1BB4: dout <= 8'b01100000; // 7092 :  96 - 0x60
      13'h1BB5: dout <= 8'b01100000; // 7093 :  96 - 0x60
      13'h1BB6: dout <= 8'b01111111; // 7094 : 127 - 0x7f
      13'h1BB7: dout <= 8'b00000000; // 7095 :   0 - 0x0
      13'h1BB8: dout <= 8'b01111111; // 7096 : 127 - 0x7f
      13'h1BB9: dout <= 8'b01100000; // 7097 :  96 - 0x60
      13'h1BBA: dout <= 8'b01100000; // 7098 :  96 - 0x60
      13'h1BBB: dout <= 8'b01111110; // 7099 : 126 - 0x7e
      13'h1BBC: dout <= 8'b01100000; // 7100 :  96 - 0x60
      13'h1BBD: dout <= 8'b01100000; // 7101 :  96 - 0x60
      13'h1BBE: dout <= 8'b01111111; // 7102 : 127 - 0x7f
      13'h1BBF: dout <= 8'b00000000; // 7103 :   0 - 0x0
      13'h1BC0: dout <= 8'b00000000; // 7104 :   0 - 0x0 -- Background 0xbc
      13'h1BC1: dout <= 8'b00100010; // 7105 :  34 - 0x22
      13'h1BC2: dout <= 8'b01100101; // 7106 : 101 - 0x65
      13'h1BC3: dout <= 8'b00100101; // 7107 :  37 - 0x25
      13'h1BC4: dout <= 8'b00100101; // 7108 :  37 - 0x25
      13'h1BC5: dout <= 8'b01110010; // 7109 : 114 - 0x72
      13'h1BC6: dout <= 8'b00000000; // 7110 :   0 - 0x0
      13'h1BC7: dout <= 8'b00000000; // 7111 :   0 - 0x0
      13'h1BC8: dout <= 8'b00000000; // 7112 :   0 - 0x0
      13'h1BC9: dout <= 8'b00000000; // 7113 :   0 - 0x0
      13'h1BCA: dout <= 8'b00000000; // 7114 :   0 - 0x0
      13'h1BCB: dout <= 8'b00000000; // 7115 :   0 - 0x0
      13'h1BCC: dout <= 8'b00000000; // 7116 :   0 - 0x0
      13'h1BCD: dout <= 8'b00000000; // 7117 :   0 - 0x0
      13'h1BCE: dout <= 8'b00000000; // 7118 :   0 - 0x0
      13'h1BCF: dout <= 8'b00000000; // 7119 :   0 - 0x0
      13'h1BD0: dout <= 8'b00000000; // 7120 :   0 - 0x0 -- Background 0xbd
      13'h1BD1: dout <= 8'b01110010; // 7121 : 114 - 0x72
      13'h1BD2: dout <= 8'b01000101; // 7122 :  69 - 0x45
      13'h1BD3: dout <= 8'b01100101; // 7123 : 101 - 0x65
      13'h1BD4: dout <= 8'b00010101; // 7124 :  21 - 0x15
      13'h1BD5: dout <= 8'b01100010; // 7125 :  98 - 0x62
      13'h1BD6: dout <= 8'b00000000; // 7126 :   0 - 0x0
      13'h1BD7: dout <= 8'b00000000; // 7127 :   0 - 0x0
      13'h1BD8: dout <= 8'b00000000; // 7128 :   0 - 0x0
      13'h1BD9: dout <= 8'b00000000; // 7129 :   0 - 0x0
      13'h1BDA: dout <= 8'b00000000; // 7130 :   0 - 0x0
      13'h1BDB: dout <= 8'b00000000; // 7131 :   0 - 0x0
      13'h1BDC: dout <= 8'b00000000; // 7132 :   0 - 0x0
      13'h1BDD: dout <= 8'b00000000; // 7133 :   0 - 0x0
      13'h1BDE: dout <= 8'b00000000; // 7134 :   0 - 0x0
      13'h1BDF: dout <= 8'b00000000; // 7135 :   0 - 0x0
      13'h1BE0: dout <= 8'b00000000; // 7136 :   0 - 0x0 -- Background 0xbe
      13'h1BE1: dout <= 8'b01100111; // 7137 : 103 - 0x67
      13'h1BE2: dout <= 8'b01010010; // 7138 :  82 - 0x52
      13'h1BE3: dout <= 8'b01100010; // 7139 :  98 - 0x62
      13'h1BE4: dout <= 8'b01000010; // 7140 :  66 - 0x42
      13'h1BE5: dout <= 8'b01000010; // 7141 :  66 - 0x42
      13'h1BE6: dout <= 8'b00000000; // 7142 :   0 - 0x0
      13'h1BE7: dout <= 8'b00000000; // 7143 :   0 - 0x0
      13'h1BE8: dout <= 8'b00000000; // 7144 :   0 - 0x0
      13'h1BE9: dout <= 8'b00000000; // 7145 :   0 - 0x0
      13'h1BEA: dout <= 8'b00000000; // 7146 :   0 - 0x0
      13'h1BEB: dout <= 8'b00000000; // 7147 :   0 - 0x0
      13'h1BEC: dout <= 8'b00000000; // 7148 :   0 - 0x0
      13'h1BED: dout <= 8'b00000000; // 7149 :   0 - 0x0
      13'h1BEE: dout <= 8'b00000000; // 7150 :   0 - 0x0
      13'h1BEF: dout <= 8'b00000000; // 7151 :   0 - 0x0
      13'h1BF0: dout <= 8'b00000000; // 7152 :   0 - 0x0 -- Background 0xbf
      13'h1BF1: dout <= 8'b01100000; // 7153 :  96 - 0x60
      13'h1BF2: dout <= 8'b10000000; // 7154 : 128 - 0x80
      13'h1BF3: dout <= 8'b01000000; // 7155 :  64 - 0x40
      13'h1BF4: dout <= 8'b00100000; // 7156 :  32 - 0x20
      13'h1BF5: dout <= 8'b11000110; // 7157 : 198 - 0xc6
      13'h1BF6: dout <= 8'b00000000; // 7158 :   0 - 0x0
      13'h1BF7: dout <= 8'b00000000; // 7159 :   0 - 0x0
      13'h1BF8: dout <= 8'b00000000; // 7160 :   0 - 0x0
      13'h1BF9: dout <= 8'b00000000; // 7161 :   0 - 0x0
      13'h1BFA: dout <= 8'b00000000; // 7162 :   0 - 0x0
      13'h1BFB: dout <= 8'b00000000; // 7163 :   0 - 0x0
      13'h1BFC: dout <= 8'b00000000; // 7164 :   0 - 0x0
      13'h1BFD: dout <= 8'b00000000; // 7165 :   0 - 0x0
      13'h1BFE: dout <= 8'b00000000; // 7166 :   0 - 0x0
      13'h1BFF: dout <= 8'b00000000; // 7167 :   0 - 0x0
      13'h1C00: dout <= 8'b01100011; // 7168 :  99 - 0x63 -- Background 0xc0
      13'h1C01: dout <= 8'b01100110; // 7169 : 102 - 0x66
      13'h1C02: dout <= 8'b01101100; // 7170 : 108 - 0x6c
      13'h1C03: dout <= 8'b01111000; // 7171 : 120 - 0x78
      13'h1C04: dout <= 8'b01111100; // 7172 : 124 - 0x7c
      13'h1C05: dout <= 8'b01100110; // 7173 : 102 - 0x66
      13'h1C06: dout <= 8'b01100011; // 7174 :  99 - 0x63
      13'h1C07: dout <= 8'b00000000; // 7175 :   0 - 0x0
      13'h1C08: dout <= 8'b01100011; // 7176 :  99 - 0x63
      13'h1C09: dout <= 8'b01100110; // 7177 : 102 - 0x66
      13'h1C0A: dout <= 8'b01101100; // 7178 : 108 - 0x6c
      13'h1C0B: dout <= 8'b01111000; // 7179 : 120 - 0x78
      13'h1C0C: dout <= 8'b01111100; // 7180 : 124 - 0x7c
      13'h1C0D: dout <= 8'b01100110; // 7181 : 102 - 0x66
      13'h1C0E: dout <= 8'b01100011; // 7182 :  99 - 0x63
      13'h1C0F: dout <= 8'b00000000; // 7183 :   0 - 0x0
      13'h1C10: dout <= 8'b00111111; // 7184 :  63 - 0x3f -- Background 0xc1
      13'h1C11: dout <= 8'b00001100; // 7185 :  12 - 0xc
      13'h1C12: dout <= 8'b00001100; // 7186 :  12 - 0xc
      13'h1C13: dout <= 8'b00001100; // 7187 :  12 - 0xc
      13'h1C14: dout <= 8'b00001100; // 7188 :  12 - 0xc
      13'h1C15: dout <= 8'b00001100; // 7189 :  12 - 0xc
      13'h1C16: dout <= 8'b00111111; // 7190 :  63 - 0x3f
      13'h1C17: dout <= 8'b00000000; // 7191 :   0 - 0x0
      13'h1C18: dout <= 8'b00111111; // 7192 :  63 - 0x3f
      13'h1C19: dout <= 8'b00001100; // 7193 :  12 - 0xc
      13'h1C1A: dout <= 8'b00001100; // 7194 :  12 - 0xc
      13'h1C1B: dout <= 8'b00001100; // 7195 :  12 - 0xc
      13'h1C1C: dout <= 8'b00001100; // 7196 :  12 - 0xc
      13'h1C1D: dout <= 8'b00001100; // 7197 :  12 - 0xc
      13'h1C1E: dout <= 8'b00111111; // 7198 :  63 - 0x3f
      13'h1C1F: dout <= 8'b00000000; // 7199 :   0 - 0x0
      13'h1C20: dout <= 8'b01100011; // 7200 :  99 - 0x63 -- Background 0xc2
      13'h1C21: dout <= 8'b01110111; // 7201 : 119 - 0x77
      13'h1C22: dout <= 8'b01111111; // 7202 : 127 - 0x7f
      13'h1C23: dout <= 8'b01111111; // 7203 : 127 - 0x7f
      13'h1C24: dout <= 8'b01101011; // 7204 : 107 - 0x6b
      13'h1C25: dout <= 8'b01100011; // 7205 :  99 - 0x63
      13'h1C26: dout <= 8'b01100011; // 7206 :  99 - 0x63
      13'h1C27: dout <= 8'b00000000; // 7207 :   0 - 0x0
      13'h1C28: dout <= 8'b01100011; // 7208 :  99 - 0x63
      13'h1C29: dout <= 8'b01110111; // 7209 : 119 - 0x77
      13'h1C2A: dout <= 8'b01111111; // 7210 : 127 - 0x7f
      13'h1C2B: dout <= 8'b01111111; // 7211 : 127 - 0x7f
      13'h1C2C: dout <= 8'b01101011; // 7212 : 107 - 0x6b
      13'h1C2D: dout <= 8'b01100011; // 7213 :  99 - 0x63
      13'h1C2E: dout <= 8'b01100011; // 7214 :  99 - 0x63
      13'h1C2F: dout <= 8'b00000000; // 7215 :   0 - 0x0
      13'h1C30: dout <= 8'b00011100; // 7216 :  28 - 0x1c -- Background 0xc3
      13'h1C31: dout <= 8'b00110110; // 7217 :  54 - 0x36
      13'h1C32: dout <= 8'b01100011; // 7218 :  99 - 0x63
      13'h1C33: dout <= 8'b01100011; // 7219 :  99 - 0x63
      13'h1C34: dout <= 8'b01111111; // 7220 : 127 - 0x7f
      13'h1C35: dout <= 8'b01100011; // 7221 :  99 - 0x63
      13'h1C36: dout <= 8'b01100011; // 7222 :  99 - 0x63
      13'h1C37: dout <= 8'b00000000; // 7223 :   0 - 0x0
      13'h1C38: dout <= 8'b00011100; // 7224 :  28 - 0x1c
      13'h1C39: dout <= 8'b00110110; // 7225 :  54 - 0x36
      13'h1C3A: dout <= 8'b01100011; // 7226 :  99 - 0x63
      13'h1C3B: dout <= 8'b01100011; // 7227 :  99 - 0x63
      13'h1C3C: dout <= 8'b01111111; // 7228 : 127 - 0x7f
      13'h1C3D: dout <= 8'b01100011; // 7229 :  99 - 0x63
      13'h1C3E: dout <= 8'b01100011; // 7230 :  99 - 0x63
      13'h1C3F: dout <= 8'b00000000; // 7231 :   0 - 0x0
      13'h1C40: dout <= 8'b00011111; // 7232 :  31 - 0x1f -- Background 0xc4
      13'h1C41: dout <= 8'b00110000; // 7233 :  48 - 0x30
      13'h1C42: dout <= 8'b01100000; // 7234 :  96 - 0x60
      13'h1C43: dout <= 8'b01100111; // 7235 : 103 - 0x67
      13'h1C44: dout <= 8'b01100011; // 7236 :  99 - 0x63
      13'h1C45: dout <= 8'b00110011; // 7237 :  51 - 0x33
      13'h1C46: dout <= 8'b00011111; // 7238 :  31 - 0x1f
      13'h1C47: dout <= 8'b00000000; // 7239 :   0 - 0x0
      13'h1C48: dout <= 8'b00011111; // 7240 :  31 - 0x1f
      13'h1C49: dout <= 8'b00110000; // 7241 :  48 - 0x30
      13'h1C4A: dout <= 8'b01100000; // 7242 :  96 - 0x60
      13'h1C4B: dout <= 8'b01100111; // 7243 : 103 - 0x67
      13'h1C4C: dout <= 8'b01100011; // 7244 :  99 - 0x63
      13'h1C4D: dout <= 8'b00110011; // 7245 :  51 - 0x33
      13'h1C4E: dout <= 8'b00011111; // 7246 :  31 - 0x1f
      13'h1C4F: dout <= 8'b00000000; // 7247 :   0 - 0x0
      13'h1C50: dout <= 8'b01100011; // 7248 :  99 - 0x63 -- Background 0xc5
      13'h1C51: dout <= 8'b01100011; // 7249 :  99 - 0x63
      13'h1C52: dout <= 8'b01100011; // 7250 :  99 - 0x63
      13'h1C53: dout <= 8'b01100011; // 7251 :  99 - 0x63
      13'h1C54: dout <= 8'b01100011; // 7252 :  99 - 0x63
      13'h1C55: dout <= 8'b01100011; // 7253 :  99 - 0x63
      13'h1C56: dout <= 8'b00111110; // 7254 :  62 - 0x3e
      13'h1C57: dout <= 8'b00000000; // 7255 :   0 - 0x0
      13'h1C58: dout <= 8'b01100011; // 7256 :  99 - 0x63
      13'h1C59: dout <= 8'b01100011; // 7257 :  99 - 0x63
      13'h1C5A: dout <= 8'b01100011; // 7258 :  99 - 0x63
      13'h1C5B: dout <= 8'b01100011; // 7259 :  99 - 0x63
      13'h1C5C: dout <= 8'b01100011; // 7260 :  99 - 0x63
      13'h1C5D: dout <= 8'b01100011; // 7261 :  99 - 0x63
      13'h1C5E: dout <= 8'b00111110; // 7262 :  62 - 0x3e
      13'h1C5F: dout <= 8'b00000000; // 7263 :   0 - 0x0
      13'h1C60: dout <= 8'b01111110; // 7264 : 126 - 0x7e -- Background 0xc6
      13'h1C61: dout <= 8'b01100011; // 7265 :  99 - 0x63
      13'h1C62: dout <= 8'b01100011; // 7266 :  99 - 0x63
      13'h1C63: dout <= 8'b01100111; // 7267 : 103 - 0x67
      13'h1C64: dout <= 8'b01111100; // 7268 : 124 - 0x7c
      13'h1C65: dout <= 8'b01101110; // 7269 : 110 - 0x6e
      13'h1C66: dout <= 8'b01100111; // 7270 : 103 - 0x67
      13'h1C67: dout <= 8'b00000000; // 7271 :   0 - 0x0
      13'h1C68: dout <= 8'b01111110; // 7272 : 126 - 0x7e
      13'h1C69: dout <= 8'b01100011; // 7273 :  99 - 0x63
      13'h1C6A: dout <= 8'b01100011; // 7274 :  99 - 0x63
      13'h1C6B: dout <= 8'b01100111; // 7275 : 103 - 0x67
      13'h1C6C: dout <= 8'b01111100; // 7276 : 124 - 0x7c
      13'h1C6D: dout <= 8'b01101110; // 7277 : 110 - 0x6e
      13'h1C6E: dout <= 8'b01100111; // 7278 : 103 - 0x67
      13'h1C6F: dout <= 8'b00000000; // 7279 :   0 - 0x0
      13'h1C70: dout <= 8'b01111111; // 7280 : 127 - 0x7f -- Background 0xc7
      13'h1C71: dout <= 8'b01100000; // 7281 :  96 - 0x60
      13'h1C72: dout <= 8'b01100000; // 7282 :  96 - 0x60
      13'h1C73: dout <= 8'b01111110; // 7283 : 126 - 0x7e
      13'h1C74: dout <= 8'b01100000; // 7284 :  96 - 0x60
      13'h1C75: dout <= 8'b01100000; // 7285 :  96 - 0x60
      13'h1C76: dout <= 8'b01111111; // 7286 : 127 - 0x7f
      13'h1C77: dout <= 8'b00000000; // 7287 :   0 - 0x0
      13'h1C78: dout <= 8'b01111111; // 7288 : 127 - 0x7f
      13'h1C79: dout <= 8'b01100000; // 7289 :  96 - 0x60
      13'h1C7A: dout <= 8'b01100000; // 7290 :  96 - 0x60
      13'h1C7B: dout <= 8'b01111110; // 7291 : 126 - 0x7e
      13'h1C7C: dout <= 8'b01100000; // 7292 :  96 - 0x60
      13'h1C7D: dout <= 8'b01100000; // 7293 :  96 - 0x60
      13'h1C7E: dout <= 8'b01111111; // 7294 : 127 - 0x7f
      13'h1C7F: dout <= 8'b00000000; // 7295 :   0 - 0x0
      13'h1C80: dout <= 8'b00110110; // 7296 :  54 - 0x36 -- Background 0xc8
      13'h1C81: dout <= 8'b00110110; // 7297 :  54 - 0x36
      13'h1C82: dout <= 8'b00010010; // 7298 :  18 - 0x12
      13'h1C83: dout <= 8'b00000000; // 7299 :   0 - 0x0
      13'h1C84: dout <= 8'b00000000; // 7300 :   0 - 0x0
      13'h1C85: dout <= 8'b00000000; // 7301 :   0 - 0x0
      13'h1C86: dout <= 8'b00000000; // 7302 :   0 - 0x0
      13'h1C87: dout <= 8'b00000000; // 7303 :   0 - 0x0
      13'h1C88: dout <= 8'b00110110; // 7304 :  54 - 0x36
      13'h1C89: dout <= 8'b00110110; // 7305 :  54 - 0x36
      13'h1C8A: dout <= 8'b00010010; // 7306 :  18 - 0x12
      13'h1C8B: dout <= 8'b00000000; // 7307 :   0 - 0x0
      13'h1C8C: dout <= 8'b00000000; // 7308 :   0 - 0x0
      13'h1C8D: dout <= 8'b00000000; // 7309 :   0 - 0x0
      13'h1C8E: dout <= 8'b00000000; // 7310 :   0 - 0x0
      13'h1C8F: dout <= 8'b00000000; // 7311 :   0 - 0x0
      13'h1C90: dout <= 8'b00111110; // 7312 :  62 - 0x3e -- Background 0xc9
      13'h1C91: dout <= 8'b01100011; // 7313 :  99 - 0x63
      13'h1C92: dout <= 8'b01100011; // 7314 :  99 - 0x63
      13'h1C93: dout <= 8'b01100011; // 7315 :  99 - 0x63
      13'h1C94: dout <= 8'b01100011; // 7316 :  99 - 0x63
      13'h1C95: dout <= 8'b01100011; // 7317 :  99 - 0x63
      13'h1C96: dout <= 8'b00111110; // 7318 :  62 - 0x3e
      13'h1C97: dout <= 8'b00000000; // 7319 :   0 - 0x0
      13'h1C98: dout <= 8'b00111110; // 7320 :  62 - 0x3e
      13'h1C99: dout <= 8'b01100011; // 7321 :  99 - 0x63
      13'h1C9A: dout <= 8'b01100011; // 7322 :  99 - 0x63
      13'h1C9B: dout <= 8'b01100011; // 7323 :  99 - 0x63
      13'h1C9C: dout <= 8'b01100011; // 7324 :  99 - 0x63
      13'h1C9D: dout <= 8'b01100011; // 7325 :  99 - 0x63
      13'h1C9E: dout <= 8'b00111110; // 7326 :  62 - 0x3e
      13'h1C9F: dout <= 8'b00000000; // 7327 :   0 - 0x0
      13'h1CA0: dout <= 8'b00111100; // 7328 :  60 - 0x3c -- Background 0xca
      13'h1CA1: dout <= 8'b01100110; // 7329 : 102 - 0x66
      13'h1CA2: dout <= 8'b01100000; // 7330 :  96 - 0x60
      13'h1CA3: dout <= 8'b00111110; // 7331 :  62 - 0x3e
      13'h1CA4: dout <= 8'b00000011; // 7332 :   3 - 0x3
      13'h1CA5: dout <= 8'b01100011; // 7333 :  99 - 0x63
      13'h1CA6: dout <= 8'b00111110; // 7334 :  62 - 0x3e
      13'h1CA7: dout <= 8'b00000000; // 7335 :   0 - 0x0
      13'h1CA8: dout <= 8'b00111100; // 7336 :  60 - 0x3c
      13'h1CA9: dout <= 8'b01100110; // 7337 : 102 - 0x66
      13'h1CAA: dout <= 8'b01100000; // 7338 :  96 - 0x60
      13'h1CAB: dout <= 8'b00111110; // 7339 :  62 - 0x3e
      13'h1CAC: dout <= 8'b00000011; // 7340 :   3 - 0x3
      13'h1CAD: dout <= 8'b01100011; // 7341 :  99 - 0x63
      13'h1CAE: dout <= 8'b00111110; // 7342 :  62 - 0x3e
      13'h1CAF: dout <= 8'b00000000; // 7343 :   0 - 0x0
      13'h1CB0: dout <= 8'b00000000; // 7344 :   0 - 0x0 -- Background 0xcb
      13'h1CB1: dout <= 8'b00000000; // 7345 :   0 - 0x0
      13'h1CB2: dout <= 8'b00000000; // 7346 :   0 - 0x0
      13'h1CB3: dout <= 8'b00000000; // 7347 :   0 - 0x0
      13'h1CB4: dout <= 8'b00000000; // 7348 :   0 - 0x0
      13'h1CB5: dout <= 8'b00000000; // 7349 :   0 - 0x0
      13'h1CB6: dout <= 8'b00000000; // 7350 :   0 - 0x0
      13'h1CB7: dout <= 8'b00000000; // 7351 :   0 - 0x0
      13'h1CB8: dout <= 8'b00000000; // 7352 :   0 - 0x0
      13'h1CB9: dout <= 8'b00111000; // 7353 :  56 - 0x38
      13'h1CBA: dout <= 8'b01111100; // 7354 : 124 - 0x7c
      13'h1CBB: dout <= 8'b11111110; // 7355 : 254 - 0xfe
      13'h1CBC: dout <= 8'b11111110; // 7356 : 254 - 0xfe
      13'h1CBD: dout <= 8'b11111110; // 7357 : 254 - 0xfe
      13'h1CBE: dout <= 8'b01111100; // 7358 : 124 - 0x7c
      13'h1CBF: dout <= 8'b00111000; // 7359 :  56 - 0x38
      13'h1CC0: dout <= 8'b00000000; // 7360 :   0 - 0x0 -- Background 0xcc
      13'h1CC1: dout <= 8'b00000000; // 7361 :   0 - 0x0
      13'h1CC2: dout <= 8'b00000000; // 7362 :   0 - 0x0
      13'h1CC3: dout <= 8'b00000000; // 7363 :   0 - 0x0
      13'h1CC4: dout <= 8'b00000000; // 7364 :   0 - 0x0
      13'h1CC5: dout <= 8'b00000000; // 7365 :   0 - 0x0
      13'h1CC6: dout <= 8'b00000000; // 7366 :   0 - 0x0
      13'h1CC7: dout <= 8'b00000000; // 7367 :   0 - 0x0
      13'h1CC8: dout <= 8'b00000000; // 7368 :   0 - 0x0
      13'h1CC9: dout <= 8'b00000000; // 7369 :   0 - 0x0
      13'h1CCA: dout <= 8'b00000000; // 7370 :   0 - 0x0
      13'h1CCB: dout <= 8'b00000000; // 7371 :   0 - 0x0
      13'h1CCC: dout <= 8'b00000000; // 7372 :   0 - 0x0
      13'h1CCD: dout <= 8'b00000000; // 7373 :   0 - 0x0
      13'h1CCE: dout <= 8'b00000000; // 7374 :   0 - 0x0
      13'h1CCF: dout <= 8'b00000000; // 7375 :   0 - 0x0
      13'h1CD0: dout <= 8'b00000000; // 7376 :   0 - 0x0 -- Background 0xcd
      13'h1CD1: dout <= 8'b00000000; // 7377 :   0 - 0x0
      13'h1CD2: dout <= 8'b00000000; // 7378 :   0 - 0x0
      13'h1CD3: dout <= 8'b00000000; // 7379 :   0 - 0x0
      13'h1CD4: dout <= 8'b00000000; // 7380 :   0 - 0x0
      13'h1CD5: dout <= 8'b00000000; // 7381 :   0 - 0x0
      13'h1CD6: dout <= 8'b00000000; // 7382 :   0 - 0x0
      13'h1CD7: dout <= 8'b00000000; // 7383 :   0 - 0x0
      13'h1CD8: dout <= 8'b00000000; // 7384 :   0 - 0x0
      13'h1CD9: dout <= 8'b00000000; // 7385 :   0 - 0x0
      13'h1CDA: dout <= 8'b00000000; // 7386 :   0 - 0x0
      13'h1CDB: dout <= 8'b00000000; // 7387 :   0 - 0x0
      13'h1CDC: dout <= 8'b00000000; // 7388 :   0 - 0x0
      13'h1CDD: dout <= 8'b00000000; // 7389 :   0 - 0x0
      13'h1CDE: dout <= 8'b00000000; // 7390 :   0 - 0x0
      13'h1CDF: dout <= 8'b00000000; // 7391 :   0 - 0x0
      13'h1CE0: dout <= 8'b00000000; // 7392 :   0 - 0x0 -- Background 0xce
      13'h1CE1: dout <= 8'b00000000; // 7393 :   0 - 0x0
      13'h1CE2: dout <= 8'b00000000; // 7394 :   0 - 0x0
      13'h1CE3: dout <= 8'b00000000; // 7395 :   0 - 0x0
      13'h1CE4: dout <= 8'b00000000; // 7396 :   0 - 0x0
      13'h1CE5: dout <= 8'b00000000; // 7397 :   0 - 0x0
      13'h1CE6: dout <= 8'b00000000; // 7398 :   0 - 0x0
      13'h1CE7: dout <= 8'b00000000; // 7399 :   0 - 0x0
      13'h1CE8: dout <= 8'b00000000; // 7400 :   0 - 0x0
      13'h1CE9: dout <= 8'b00000000; // 7401 :   0 - 0x0
      13'h1CEA: dout <= 8'b00000000; // 7402 :   0 - 0x0
      13'h1CEB: dout <= 8'b00000000; // 7403 :   0 - 0x0
      13'h1CEC: dout <= 8'b00000000; // 7404 :   0 - 0x0
      13'h1CED: dout <= 8'b00000000; // 7405 :   0 - 0x0
      13'h1CEE: dout <= 8'b00000000; // 7406 :   0 - 0x0
      13'h1CEF: dout <= 8'b00000000; // 7407 :   0 - 0x0
      13'h1CF0: dout <= 8'b00000000; // 7408 :   0 - 0x0 -- Background 0xcf
      13'h1CF1: dout <= 8'b00000000; // 7409 :   0 - 0x0
      13'h1CF2: dout <= 8'b00000000; // 7410 :   0 - 0x0
      13'h1CF3: dout <= 8'b00000000; // 7411 :   0 - 0x0
      13'h1CF4: dout <= 8'b00000000; // 7412 :   0 - 0x0
      13'h1CF5: dout <= 8'b00000000; // 7413 :   0 - 0x0
      13'h1CF6: dout <= 8'b00000000; // 7414 :   0 - 0x0
      13'h1CF7: dout <= 8'b00000000; // 7415 :   0 - 0x0
      13'h1CF8: dout <= 8'b00000000; // 7416 :   0 - 0x0
      13'h1CF9: dout <= 8'b00000000; // 7417 :   0 - 0x0
      13'h1CFA: dout <= 8'b00000000; // 7418 :   0 - 0x0
      13'h1CFB: dout <= 8'b00000000; // 7419 :   0 - 0x0
      13'h1CFC: dout <= 8'b00000000; // 7420 :   0 - 0x0
      13'h1CFD: dout <= 8'b00000000; // 7421 :   0 - 0x0
      13'h1CFE: dout <= 8'b00000000; // 7422 :   0 - 0x0
      13'h1CFF: dout <= 8'b00000000; // 7423 :   0 - 0x0
      13'h1D00: dout <= 8'b01000111; // 7424 :  71 - 0x47 -- Background 0xd0
      13'h1D01: dout <= 8'b01000111; // 7425 :  71 - 0x47
      13'h1D02: dout <= 8'b00001111; // 7426 :  15 - 0xf
      13'h1D03: dout <= 8'b00001111; // 7427 :  15 - 0xf
      13'h1D04: dout <= 8'b00011111; // 7428 :  31 - 0x1f
      13'h1D05: dout <= 8'b00011111; // 7429 :  31 - 0x1f
      13'h1D06: dout <= 8'b00111111; // 7430 :  63 - 0x3f
      13'h1D07: dout <= 8'b00111111; // 7431 :  63 - 0x3f
      13'h1D08: dout <= 8'b00010111; // 7432 :  23 - 0x17
      13'h1D09: dout <= 8'b00010111; // 7433 :  23 - 0x17
      13'h1D0A: dout <= 8'b00101111; // 7434 :  47 - 0x2f
      13'h1D0B: dout <= 8'b00101111; // 7435 :  47 - 0x2f
      13'h1D0C: dout <= 8'b01011111; // 7436 :  95 - 0x5f
      13'h1D0D: dout <= 8'b01011111; // 7437 :  95 - 0x5f
      13'h1D0E: dout <= 8'b00111111; // 7438 :  63 - 0x3f
      13'h1D0F: dout <= 8'b00111111; // 7439 :  63 - 0x3f
      13'h1D10: dout <= 8'b11111111; // 7440 : 255 - 0xff -- Background 0xd1
      13'h1D11: dout <= 8'b11001111; // 7441 : 207 - 0xcf
      13'h1D12: dout <= 8'b11001111; // 7442 : 207 - 0xcf
      13'h1D13: dout <= 8'b11111011; // 7443 : 251 - 0xfb
      13'h1D14: dout <= 8'b11110111; // 7444 : 247 - 0xf7
      13'h1D15: dout <= 8'b11100111; // 7445 : 231 - 0xe7
      13'h1D16: dout <= 8'b11111111; // 7446 : 255 - 0xff
      13'h1D17: dout <= 8'b11111111; // 7447 : 255 - 0xff
      13'h1D18: dout <= 8'b11111111; // 7448 : 255 - 0xff
      13'h1D19: dout <= 8'b11001111; // 7449 : 207 - 0xcf
      13'h1D1A: dout <= 8'b11001111; // 7450 : 207 - 0xcf
      13'h1D1B: dout <= 8'b11111011; // 7451 : 251 - 0xfb
      13'h1D1C: dout <= 8'b11110111; // 7452 : 247 - 0xf7
      13'h1D1D: dout <= 8'b11100111; // 7453 : 231 - 0xe7
      13'h1D1E: dout <= 8'b11111111; // 7454 : 255 - 0xff
      13'h1D1F: dout <= 8'b11111111; // 7455 : 255 - 0xff
      13'h1D20: dout <= 8'b00011000; // 7456 :  24 - 0x18 -- Background 0xd2
      13'h1D21: dout <= 8'b00001000; // 7457 :   8 - 0x8
      13'h1D22: dout <= 8'b10001000; // 7458 : 136 - 0x88
      13'h1D23: dout <= 8'b10000000; // 7459 : 128 - 0x80
      13'h1D24: dout <= 8'b01000000; // 7460 :  64 - 0x40
      13'h1D25: dout <= 8'b01000000; // 7461 :  64 - 0x40
      13'h1D26: dout <= 8'b10100000; // 7462 : 160 - 0xa0
      13'h1D27: dout <= 8'b10100000; // 7463 : 160 - 0xa0
      13'h1D28: dout <= 8'b01000010; // 7464 :  66 - 0x42
      13'h1D29: dout <= 8'b01100010; // 7465 :  98 - 0x62
      13'h1D2A: dout <= 8'b10100010; // 7466 : 162 - 0xa2
      13'h1D2B: dout <= 8'b10110010; // 7467 : 178 - 0xb2
      13'h1D2C: dout <= 8'b01010010; // 7468 :  82 - 0x52
      13'h1D2D: dout <= 8'b01011010; // 7469 :  90 - 0x5a
      13'h1D2E: dout <= 8'b10101010; // 7470 : 170 - 0xaa
      13'h1D2F: dout <= 8'b10101100; // 7471 : 172 - 0xac
      13'h1D30: dout <= 8'b11111111; // 7472 : 255 - 0xff -- Background 0xd3
      13'h1D31: dout <= 8'b11111111; // 7473 : 255 - 0xff
      13'h1D32: dout <= 8'b11111111; // 7474 : 255 - 0xff
      13'h1D33: dout <= 8'b11111111; // 7475 : 255 - 0xff
      13'h1D34: dout <= 8'b11111101; // 7476 : 253 - 0xfd
      13'h1D35: dout <= 8'b11111101; // 7477 : 253 - 0xfd
      13'h1D36: dout <= 8'b11111101; // 7478 : 253 - 0xfd
      13'h1D37: dout <= 8'b11111101; // 7479 : 253 - 0xfd
      13'h1D38: dout <= 8'b11111111; // 7480 : 255 - 0xff
      13'h1D39: dout <= 8'b11111111; // 7481 : 255 - 0xff
      13'h1D3A: dout <= 8'b11111111; // 7482 : 255 - 0xff
      13'h1D3B: dout <= 8'b11111111; // 7483 : 255 - 0xff
      13'h1D3C: dout <= 8'b11111101; // 7484 : 253 - 0xfd
      13'h1D3D: dout <= 8'b11111101; // 7485 : 253 - 0xfd
      13'h1D3E: dout <= 8'b11111101; // 7486 : 253 - 0xfd
      13'h1D3F: dout <= 8'b11111101; // 7487 : 253 - 0xfd
      13'h1D40: dout <= 8'b11000111; // 7488 : 199 - 0xc7 -- Background 0xd4
      13'h1D41: dout <= 8'b11110111; // 7489 : 247 - 0xf7
      13'h1D42: dout <= 8'b11110000; // 7490 : 240 - 0xf0
      13'h1D43: dout <= 8'b11111000; // 7491 : 248 - 0xf8
      13'h1D44: dout <= 8'b11111000; // 7492 : 248 - 0xf8
      13'h1D45: dout <= 8'b11111111; // 7493 : 255 - 0xff
      13'h1D46: dout <= 8'b11111111; // 7494 : 255 - 0xff
      13'h1D47: dout <= 8'b11111111; // 7495 : 255 - 0xff
      13'h1D48: dout <= 8'b00000111; // 7496 :   7 - 0x7
      13'h1D49: dout <= 8'b00000111; // 7497 :   7 - 0x7
      13'h1D4A: dout <= 8'b00000000; // 7498 :   0 - 0x0
      13'h1D4B: dout <= 8'b00000011; // 7499 :   3 - 0x3
      13'h1D4C: dout <= 8'b00000000; // 7500 :   0 - 0x0
      13'h1D4D: dout <= 8'b00000000; // 7501 :   0 - 0x0
      13'h1D4E: dout <= 8'b00000000; // 7502 :   0 - 0x0
      13'h1D4F: dout <= 8'b00000000; // 7503 :   0 - 0x0
      13'h1D50: dout <= 8'b11111000; // 7504 : 248 - 0xf8 -- Background 0xd5
      13'h1D51: dout <= 8'b11111000; // 7505 : 248 - 0xf8
      13'h1D52: dout <= 8'b00000000; // 7506 :   0 - 0x0
      13'h1D53: dout <= 8'b00000000; // 7507 :   0 - 0x0
      13'h1D54: dout <= 8'b00000000; // 7508 :   0 - 0x0
      13'h1D55: dout <= 8'b11111111; // 7509 : 255 - 0xff
      13'h1D56: dout <= 8'b11111111; // 7510 : 255 - 0xff
      13'h1D57: dout <= 8'b11111111; // 7511 : 255 - 0xff
      13'h1D58: dout <= 8'b11111010; // 7512 : 250 - 0xfa
      13'h1D59: dout <= 8'b11111010; // 7513 : 250 - 0xfa
      13'h1D5A: dout <= 8'b00000010; // 7514 :   2 - 0x2
      13'h1D5B: dout <= 8'b11111110; // 7515 : 254 - 0xfe
      13'h1D5C: dout <= 8'b00000000; // 7516 :   0 - 0x0
      13'h1D5D: dout <= 8'b00000000; // 7517 :   0 - 0x0
      13'h1D5E: dout <= 8'b00000000; // 7518 :   0 - 0x0
      13'h1D5F: dout <= 8'b00000000; // 7519 :   0 - 0x0
      13'h1D60: dout <= 8'b10001111; // 7520 : 143 - 0x8f -- Background 0xd6
      13'h1D61: dout <= 8'b11101111; // 7521 : 239 - 0xef
      13'h1D62: dout <= 8'b11000000; // 7522 : 192 - 0xc0
      13'h1D63: dout <= 8'b11110000; // 7523 : 240 - 0xf0
      13'h1D64: dout <= 8'b11100000; // 7524 : 224 - 0xe0
      13'h1D65: dout <= 8'b11111111; // 7525 : 255 - 0xff
      13'h1D66: dout <= 8'b11111111; // 7526 : 255 - 0xff
      13'h1D67: dout <= 8'b11111111; // 7527 : 255 - 0xff
      13'h1D68: dout <= 8'b00001111; // 7528 :  15 - 0xf
      13'h1D69: dout <= 8'b00001111; // 7529 :  15 - 0xf
      13'h1D6A: dout <= 8'b00000000; // 7530 :   0 - 0x0
      13'h1D6B: dout <= 8'b00000111; // 7531 :   7 - 0x7
      13'h1D6C: dout <= 8'b00000000; // 7532 :   0 - 0x0
      13'h1D6D: dout <= 8'b00000000; // 7533 :   0 - 0x0
      13'h1D6E: dout <= 8'b00000000; // 7534 :   0 - 0x0
      13'h1D6F: dout <= 8'b00000000; // 7535 :   0 - 0x0
      13'h1D70: dout <= 8'b11111111; // 7536 : 255 - 0xff -- Background 0xd7
      13'h1D71: dout <= 8'b11111111; // 7537 : 255 - 0xff
      13'h1D72: dout <= 8'b00000000; // 7538 :   0 - 0x0
      13'h1D73: dout <= 8'b00000000; // 7539 :   0 - 0x0
      13'h1D74: dout <= 8'b00000000; // 7540 :   0 - 0x0
      13'h1D75: dout <= 8'b11111111; // 7541 : 255 - 0xff
      13'h1D76: dout <= 8'b11111111; // 7542 : 255 - 0xff
      13'h1D77: dout <= 8'b11111111; // 7543 : 255 - 0xff
      13'h1D78: dout <= 8'b11111111; // 7544 : 255 - 0xff
      13'h1D79: dout <= 8'b11111111; // 7545 : 255 - 0xff
      13'h1D7A: dout <= 8'b00000000; // 7546 :   0 - 0x0
      13'h1D7B: dout <= 8'b11111111; // 7547 : 255 - 0xff
      13'h1D7C: dout <= 8'b00000000; // 7548 :   0 - 0x0
      13'h1D7D: dout <= 8'b00000000; // 7549 :   0 - 0x0
      13'h1D7E: dout <= 8'b00000000; // 7550 :   0 - 0x0
      13'h1D7F: dout <= 8'b00000000; // 7551 :   0 - 0x0
      13'h1D80: dout <= 8'b11000011; // 7552 : 195 - 0xc3 -- Background 0xd8
      13'h1D81: dout <= 8'b11111111; // 7553 : 255 - 0xff
      13'h1D82: dout <= 8'b00000000; // 7554 :   0 - 0x0
      13'h1D83: dout <= 8'b00000000; // 7555 :   0 - 0x0
      13'h1D84: dout <= 8'b00000000; // 7556 :   0 - 0x0
      13'h1D85: dout <= 8'b11111111; // 7557 : 255 - 0xff
      13'h1D86: dout <= 8'b11111111; // 7558 : 255 - 0xff
      13'h1D87: dout <= 8'b11111111; // 7559 : 255 - 0xff
      13'h1D88: dout <= 8'b11000011; // 7560 : 195 - 0xc3
      13'h1D89: dout <= 8'b11111111; // 7561 : 255 - 0xff
      13'h1D8A: dout <= 8'b00000000; // 7562 :   0 - 0x0
      13'h1D8B: dout <= 8'b11111111; // 7563 : 255 - 0xff
      13'h1D8C: dout <= 8'b00000000; // 7564 :   0 - 0x0
      13'h1D8D: dout <= 8'b00000000; // 7565 :   0 - 0x0
      13'h1D8E: dout <= 8'b00000000; // 7566 :   0 - 0x0
      13'h1D8F: dout <= 8'b00000000; // 7567 :   0 - 0x0
      13'h1D90: dout <= 8'b00000011; // 7568 :   3 - 0x3 -- Background 0xd9
      13'h1D91: dout <= 8'b10000001; // 7569 : 129 - 0x81
      13'h1D92: dout <= 8'b00000000; // 7570 :   0 - 0x0
      13'h1D93: dout <= 8'b00000000; // 7571 :   0 - 0x0
      13'h1D94: dout <= 8'b00000011; // 7572 :   3 - 0x3
      13'h1D95: dout <= 8'b11111111; // 7573 : 255 - 0xff
      13'h1D96: dout <= 8'b11111111; // 7574 : 255 - 0xff
      13'h1D97: dout <= 8'b11111111; // 7575 : 255 - 0xff
      13'h1D98: dout <= 8'b01101011; // 7576 : 107 - 0x6b
      13'h1D99: dout <= 8'b10110101; // 7577 : 181 - 0xb5
      13'h1D9A: dout <= 8'b00110110; // 7578 :  54 - 0x36
      13'h1D9B: dout <= 8'b11111000; // 7579 : 248 - 0xf8
      13'h1D9C: dout <= 8'b00000000; // 7580 :   0 - 0x0
      13'h1D9D: dout <= 8'b00000000; // 7581 :   0 - 0x0
      13'h1D9E: dout <= 8'b00000000; // 7582 :   0 - 0x0
      13'h1D9F: dout <= 8'b00000000; // 7583 :   0 - 0x0
      13'h1DA0: dout <= 8'b11111111; // 7584 : 255 - 0xff -- Background 0xda
      13'h1DA1: dout <= 8'b11111111; // 7585 : 255 - 0xff
      13'h1DA2: dout <= 8'b01111110; // 7586 : 126 - 0x7e
      13'h1DA3: dout <= 8'b00000000; // 7587 :   0 - 0x0
      13'h1DA4: dout <= 8'b00000000; // 7588 :   0 - 0x0
      13'h1DA5: dout <= 8'b11100000; // 7589 : 224 - 0xe0
      13'h1DA6: dout <= 8'b11111111; // 7590 : 255 - 0xff
      13'h1DA7: dout <= 8'b11111111; // 7591 : 255 - 0xff
      13'h1DA8: dout <= 8'b11111111; // 7592 : 255 - 0xff
      13'h1DA9: dout <= 8'b11111111; // 7593 : 255 - 0xff
      13'h1DAA: dout <= 8'b01111110; // 7594 : 126 - 0x7e
      13'h1DAB: dout <= 8'b10000001; // 7595 : 129 - 0x81
      13'h1DAC: dout <= 8'b00011111; // 7596 :  31 - 0x1f
      13'h1DAD: dout <= 8'b00000000; // 7597 :   0 - 0x0
      13'h1DAE: dout <= 8'b00000000; // 7598 :   0 - 0x0
      13'h1DAF: dout <= 8'b00000000; // 7599 :   0 - 0x0
      13'h1DB0: dout <= 8'b01100001; // 7600 :  97 - 0x61 -- Background 0xdb
      13'h1DB1: dout <= 8'b11000011; // 7601 : 195 - 0xc3
      13'h1DB2: dout <= 8'b00000111; // 7602 :   7 - 0x7
      13'h1DB3: dout <= 8'b00001111; // 7603 :  15 - 0xf
      13'h1DB4: dout <= 8'b00011111; // 7604 :  31 - 0x1f
      13'h1DB5: dout <= 8'b01111111; // 7605 : 127 - 0x7f
      13'h1DB6: dout <= 8'b11111111; // 7606 : 255 - 0xff
      13'h1DB7: dout <= 8'b11111111; // 7607 : 255 - 0xff
      13'h1DB8: dout <= 8'b01101100; // 7608 : 108 - 0x6c
      13'h1DB9: dout <= 8'b11011000; // 7609 : 216 - 0xd8
      13'h1DBA: dout <= 8'b00110000; // 7610 :  48 - 0x30
      13'h1DBB: dout <= 8'b11100000; // 7611 : 224 - 0xe0
      13'h1DBC: dout <= 8'b10000000; // 7612 : 128 - 0x80
      13'h1DBD: dout <= 8'b00000000; // 7613 :   0 - 0x0
      13'h1DBE: dout <= 8'b00000000; // 7614 :   0 - 0x0
      13'h1DBF: dout <= 8'b00000000; // 7615 :   0 - 0x0
      13'h1DC0: dout <= 8'b00011111; // 7616 :  31 - 0x1f -- Background 0xdc
      13'h1DC1: dout <= 8'b11011111; // 7617 : 223 - 0xdf
      13'h1DC2: dout <= 8'b11000000; // 7618 : 192 - 0xc0
      13'h1DC3: dout <= 8'b11110000; // 7619 : 240 - 0xf0
      13'h1DC4: dout <= 8'b11110000; // 7620 : 240 - 0xf0
      13'h1DC5: dout <= 8'b11111111; // 7621 : 255 - 0xff
      13'h1DC6: dout <= 8'b11111111; // 7622 : 255 - 0xff
      13'h1DC7: dout <= 8'b11111111; // 7623 : 255 - 0xff
      13'h1DC8: dout <= 8'b00011111; // 7624 :  31 - 0x1f
      13'h1DC9: dout <= 8'b00011111; // 7625 :  31 - 0x1f
      13'h1DCA: dout <= 8'b00000000; // 7626 :   0 - 0x0
      13'h1DCB: dout <= 8'b00000111; // 7627 :   7 - 0x7
      13'h1DCC: dout <= 8'b00000000; // 7628 :   0 - 0x0
      13'h1DCD: dout <= 8'b00000000; // 7629 :   0 - 0x0
      13'h1DCE: dout <= 8'b00000000; // 7630 :   0 - 0x0
      13'h1DCF: dout <= 8'b00000000; // 7631 :   0 - 0x0
      13'h1DD0: dout <= 8'b10000100; // 7632 : 132 - 0x84 -- Background 0xdd
      13'h1DD1: dout <= 8'b11111100; // 7633 : 252 - 0xfc
      13'h1DD2: dout <= 8'b00000000; // 7634 :   0 - 0x0
      13'h1DD3: dout <= 8'b00000000; // 7635 :   0 - 0x0
      13'h1DD4: dout <= 8'b00000000; // 7636 :   0 - 0x0
      13'h1DD5: dout <= 8'b11111111; // 7637 : 255 - 0xff
      13'h1DD6: dout <= 8'b11111111; // 7638 : 255 - 0xff
      13'h1DD7: dout <= 8'b11111111; // 7639 : 255 - 0xff
      13'h1DD8: dout <= 8'b10000101; // 7640 : 133 - 0x85
      13'h1DD9: dout <= 8'b11111101; // 7641 : 253 - 0xfd
      13'h1DDA: dout <= 8'b00000001; // 7642 :   1 - 0x1
      13'h1DDB: dout <= 8'b11111111; // 7643 : 255 - 0xff
      13'h1DDC: dout <= 8'b00000000; // 7644 :   0 - 0x0
      13'h1DDD: dout <= 8'b00000000; // 7645 :   0 - 0x0
      13'h1DDE: dout <= 8'b00000000; // 7646 :   0 - 0x0
      13'h1DDF: dout <= 8'b00000000; // 7647 :   0 - 0x0
      13'h1DE0: dout <= 8'b01111111; // 7648 : 127 - 0x7f -- Background 0xde
      13'h1DE1: dout <= 8'b01111111; // 7649 : 127 - 0x7f
      13'h1DE2: dout <= 8'b00000000; // 7650 :   0 - 0x0
      13'h1DE3: dout <= 8'b00000000; // 7651 :   0 - 0x0
      13'h1DE4: dout <= 8'b00000000; // 7652 :   0 - 0x0
      13'h1DE5: dout <= 8'b11111111; // 7653 : 255 - 0xff
      13'h1DE6: dout <= 8'b11111111; // 7654 : 255 - 0xff
      13'h1DE7: dout <= 8'b11111111; // 7655 : 255 - 0xff
      13'h1DE8: dout <= 8'b01111111; // 7656 : 127 - 0x7f
      13'h1DE9: dout <= 8'b01111111; // 7657 : 127 - 0x7f
      13'h1DEA: dout <= 8'b00000000; // 7658 :   0 - 0x0
      13'h1DEB: dout <= 8'b01011111; // 7659 :  95 - 0x5f
      13'h1DEC: dout <= 8'b00000000; // 7660 :   0 - 0x0
      13'h1DED: dout <= 8'b00000000; // 7661 :   0 - 0x0
      13'h1DEE: dout <= 8'b00000000; // 7662 :   0 - 0x0
      13'h1DEF: dout <= 8'b00000000; // 7663 :   0 - 0x0
      13'h1DF0: dout <= 8'b11111100; // 7664 : 252 - 0xfc -- Background 0xdf
      13'h1DF1: dout <= 8'b11111111; // 7665 : 255 - 0xff
      13'h1DF2: dout <= 8'b00000000; // 7666 :   0 - 0x0
      13'h1DF3: dout <= 8'b00000000; // 7667 :   0 - 0x0
      13'h1DF4: dout <= 8'b00000000; // 7668 :   0 - 0x0
      13'h1DF5: dout <= 8'b11111111; // 7669 : 255 - 0xff
      13'h1DF6: dout <= 8'b11111111; // 7670 : 255 - 0xff
      13'h1DF7: dout <= 8'b11111111; // 7671 : 255 - 0xff
      13'h1DF8: dout <= 8'b11111100; // 7672 : 252 - 0xfc
      13'h1DF9: dout <= 8'b11111111; // 7673 : 255 - 0xff
      13'h1DFA: dout <= 8'b00000000; // 7674 :   0 - 0x0
      13'h1DFB: dout <= 8'b11111111; // 7675 : 255 - 0xff
      13'h1DFC: dout <= 8'b00000000; // 7676 :   0 - 0x0
      13'h1DFD: dout <= 8'b00000000; // 7677 :   0 - 0x0
      13'h1DFE: dout <= 8'b00000000; // 7678 :   0 - 0x0
      13'h1DFF: dout <= 8'b00000000; // 7679 :   0 - 0x0
      13'h1E00: dout <= 8'b00110000; // 7680 :  48 - 0x30 -- Background 0xe0
      13'h1E01: dout <= 8'b11110000; // 7681 : 240 - 0xf0
      13'h1E02: dout <= 8'b00000000; // 7682 :   0 - 0x0
      13'h1E03: dout <= 8'b00000000; // 7683 :   0 - 0x0
      13'h1E04: dout <= 8'b00000000; // 7684 :   0 - 0x0
      13'h1E05: dout <= 8'b11111111; // 7685 : 255 - 0xff
      13'h1E06: dout <= 8'b11111111; // 7686 : 255 - 0xff
      13'h1E07: dout <= 8'b11111111; // 7687 : 255 - 0xff
      13'h1E08: dout <= 8'b00110100; // 7688 :  52 - 0x34
      13'h1E09: dout <= 8'b11110110; // 7689 : 246 - 0xf6
      13'h1E0A: dout <= 8'b00000010; // 7690 :   2 - 0x2
      13'h1E0B: dout <= 8'b11111111; // 7691 : 255 - 0xff
      13'h1E0C: dout <= 8'b00000000; // 7692 :   0 - 0x0
      13'h1E0D: dout <= 8'b00000000; // 7693 :   0 - 0x0
      13'h1E0E: dout <= 8'b00000000; // 7694 :   0 - 0x0
      13'h1E0F: dout <= 8'b00000000; // 7695 :   0 - 0x0
      13'h1E10: dout <= 8'b11111111; // 7696 : 255 - 0xff -- Background 0xe1
      13'h1E11: dout <= 8'b11111111; // 7697 : 255 - 0xff
      13'h1E12: dout <= 8'b00000000; // 7698 :   0 - 0x0
      13'h1E13: dout <= 8'b00000000; // 7699 :   0 - 0x0
      13'h1E14: dout <= 8'b00000000; // 7700 :   0 - 0x0
      13'h1E15: dout <= 8'b11111111; // 7701 : 255 - 0xff
      13'h1E16: dout <= 8'b11111111; // 7702 : 255 - 0xff
      13'h1E17: dout <= 8'b11111111; // 7703 : 255 - 0xff
      13'h1E18: dout <= 8'b11111111; // 7704 : 255 - 0xff
      13'h1E19: dout <= 8'b11111111; // 7705 : 255 - 0xff
      13'h1E1A: dout <= 8'b00000000; // 7706 :   0 - 0x0
      13'h1E1B: dout <= 8'b01111111; // 7707 : 127 - 0x7f
      13'h1E1C: dout <= 8'b00000000; // 7708 :   0 - 0x0
      13'h1E1D: dout <= 8'b00000000; // 7709 :   0 - 0x0
      13'h1E1E: dout <= 8'b00000000; // 7710 :   0 - 0x0
      13'h1E1F: dout <= 8'b00000000; // 7711 :   0 - 0x0
      13'h1E20: dout <= 8'b11100001; // 7712 : 225 - 0xe1 -- Background 0xe2
      13'h1E21: dout <= 8'b11111111; // 7713 : 255 - 0xff
      13'h1E22: dout <= 8'b00000000; // 7714 :   0 - 0x0
      13'h1E23: dout <= 8'b00000000; // 7715 :   0 - 0x0
      13'h1E24: dout <= 8'b00000000; // 7716 :   0 - 0x0
      13'h1E25: dout <= 8'b11111111; // 7717 : 255 - 0xff
      13'h1E26: dout <= 8'b11111111; // 7718 : 255 - 0xff
      13'h1E27: dout <= 8'b11111111; // 7719 : 255 - 0xff
      13'h1E28: dout <= 8'b11100001; // 7720 : 225 - 0xe1
      13'h1E29: dout <= 8'b11111111; // 7721 : 255 - 0xff
      13'h1E2A: dout <= 8'b00000000; // 7722 :   0 - 0x0
      13'h1E2B: dout <= 8'b11111111; // 7723 : 255 - 0xff
      13'h1E2C: dout <= 8'b00000000; // 7724 :   0 - 0x0
      13'h1E2D: dout <= 8'b00000000; // 7725 :   0 - 0x0
      13'h1E2E: dout <= 8'b00000000; // 7726 :   0 - 0x0
      13'h1E2F: dout <= 8'b00000000; // 7727 :   0 - 0x0
      13'h1E30: dout <= 8'b00011111; // 7728 :  31 - 0x1f -- Background 0xe3
      13'h1E31: dout <= 8'b00011111; // 7729 :  31 - 0x1f
      13'h1E32: dout <= 8'b00011111; // 7730 :  31 - 0x1f
      13'h1E33: dout <= 8'b00011111; // 7731 :  31 - 0x1f
      13'h1E34: dout <= 8'b00011111; // 7732 :  31 - 0x1f
      13'h1E35: dout <= 8'b11111111; // 7733 : 255 - 0xff
      13'h1E36: dout <= 8'b11111111; // 7734 : 255 - 0xff
      13'h1E37: dout <= 8'b11111111; // 7735 : 255 - 0xff
      13'h1E38: dout <= 8'b01000000; // 7736 :  64 - 0x40
      13'h1E39: dout <= 8'b01000000; // 7737 :  64 - 0x40
      13'h1E3A: dout <= 8'b01000000; // 7738 :  64 - 0x40
      13'h1E3B: dout <= 8'b11000000; // 7739 : 192 - 0xc0
      13'h1E3C: dout <= 8'b00000000; // 7740 :   0 - 0x0
      13'h1E3D: dout <= 8'b00000000; // 7741 :   0 - 0x0
      13'h1E3E: dout <= 8'b00000000; // 7742 :   0 - 0x0
      13'h1E3F: dout <= 8'b00000000; // 7743 :   0 - 0x0
      13'h1E40: dout <= 8'b00000000; // 7744 :   0 - 0x0 -- Background 0xe4
      13'h1E41: dout <= 8'b00011111; // 7745 :  31 - 0x1f
      13'h1E42: dout <= 8'b00111111; // 7746 :  63 - 0x3f
      13'h1E43: dout <= 8'b01111000; // 7747 : 120 - 0x78
      13'h1E44: dout <= 8'b01110111; // 7748 : 119 - 0x77
      13'h1E45: dout <= 8'b01101111; // 7749 : 111 - 0x6f
      13'h1E46: dout <= 8'b01101111; // 7750 : 111 - 0x6f
      13'h1E47: dout <= 8'b01101111; // 7751 : 111 - 0x6f
      13'h1E48: dout <= 8'b00000000; // 7752 :   0 - 0x0
      13'h1E49: dout <= 8'b00000000; // 7753 :   0 - 0x0
      13'h1E4A: dout <= 8'b00000000; // 7754 :   0 - 0x0
      13'h1E4B: dout <= 8'b00000000; // 7755 :   0 - 0x0
      13'h1E4C: dout <= 8'b00000111; // 7756 :   7 - 0x7
      13'h1E4D: dout <= 8'b00001111; // 7757 :  15 - 0xf
      13'h1E4E: dout <= 8'b00001111; // 7758 :  15 - 0xf
      13'h1E4F: dout <= 8'b00001111; // 7759 :  15 - 0xf
      13'h1E50: dout <= 8'b00000000; // 7760 :   0 - 0x0 -- Background 0xe5
      13'h1E51: dout <= 8'b11111000; // 7761 : 248 - 0xf8
      13'h1E52: dout <= 8'b11111100; // 7762 : 252 - 0xfc
      13'h1E53: dout <= 8'b00011110; // 7763 :  30 - 0x1e
      13'h1E54: dout <= 8'b11101110; // 7764 : 238 - 0xee
      13'h1E55: dout <= 8'b11110110; // 7765 : 246 - 0xf6
      13'h1E56: dout <= 8'b11110110; // 7766 : 246 - 0xf6
      13'h1E57: dout <= 8'b11110110; // 7767 : 246 - 0xf6
      13'h1E58: dout <= 8'b00000000; // 7768 :   0 - 0x0
      13'h1E59: dout <= 8'b00000000; // 7769 :   0 - 0x0
      13'h1E5A: dout <= 8'b00000000; // 7770 :   0 - 0x0
      13'h1E5B: dout <= 8'b00000000; // 7771 :   0 - 0x0
      13'h1E5C: dout <= 8'b11100000; // 7772 : 224 - 0xe0
      13'h1E5D: dout <= 8'b11110000; // 7773 : 240 - 0xf0
      13'h1E5E: dout <= 8'b11110000; // 7774 : 240 - 0xf0
      13'h1E5F: dout <= 8'b11110000; // 7775 : 240 - 0xf0
      13'h1E60: dout <= 8'b11110110; // 7776 : 246 - 0xf6 -- Background 0xe6
      13'h1E61: dout <= 8'b11110110; // 7777 : 246 - 0xf6
      13'h1E62: dout <= 8'b11110110; // 7778 : 246 - 0xf6
      13'h1E63: dout <= 8'b11101110; // 7779 : 238 - 0xee
      13'h1E64: dout <= 8'b00011110; // 7780 :  30 - 0x1e
      13'h1E65: dout <= 8'b11111100; // 7781 : 252 - 0xfc
      13'h1E66: dout <= 8'b11111000; // 7782 : 248 - 0xf8
      13'h1E67: dout <= 8'b00000000; // 7783 :   0 - 0x0
      13'h1E68: dout <= 8'b11110000; // 7784 : 240 - 0xf0
      13'h1E69: dout <= 8'b11110000; // 7785 : 240 - 0xf0
      13'h1E6A: dout <= 8'b11110000; // 7786 : 240 - 0xf0
      13'h1E6B: dout <= 8'b11100000; // 7787 : 224 - 0xe0
      13'h1E6C: dout <= 8'b00000000; // 7788 :   0 - 0x0
      13'h1E6D: dout <= 8'b00000000; // 7789 :   0 - 0x0
      13'h1E6E: dout <= 8'b00000000; // 7790 :   0 - 0x0
      13'h1E6F: dout <= 8'b00000000; // 7791 :   0 - 0x0
      13'h1E70: dout <= 8'b01101111; // 7792 : 111 - 0x6f -- Background 0xe7
      13'h1E71: dout <= 8'b01101111; // 7793 : 111 - 0x6f
      13'h1E72: dout <= 8'b01101111; // 7794 : 111 - 0x6f
      13'h1E73: dout <= 8'b01110111; // 7795 : 119 - 0x77
      13'h1E74: dout <= 8'b01111000; // 7796 : 120 - 0x78
      13'h1E75: dout <= 8'b00111111; // 7797 :  63 - 0x3f
      13'h1E76: dout <= 8'b00011111; // 7798 :  31 - 0x1f
      13'h1E77: dout <= 8'b00000000; // 7799 :   0 - 0x0
      13'h1E78: dout <= 8'b00001111; // 7800 :  15 - 0xf
      13'h1E79: dout <= 8'b00001111; // 7801 :  15 - 0xf
      13'h1E7A: dout <= 8'b00001111; // 7802 :  15 - 0xf
      13'h1E7B: dout <= 8'b00000111; // 7803 :   7 - 0x7
      13'h1E7C: dout <= 8'b00000000; // 7804 :   0 - 0x0
      13'h1E7D: dout <= 8'b00000000; // 7805 :   0 - 0x0
      13'h1E7E: dout <= 8'b00000000; // 7806 :   0 - 0x0
      13'h1E7F: dout <= 8'b00000000; // 7807 :   0 - 0x0
      13'h1E80: dout <= 8'b00000000; // 7808 :   0 - 0x0 -- Background 0xe8
      13'h1E81: dout <= 8'b11111111; // 7809 : 255 - 0xff
      13'h1E82: dout <= 8'b11111111; // 7810 : 255 - 0xff
      13'h1E83: dout <= 8'b00000000; // 7811 :   0 - 0x0
      13'h1E84: dout <= 8'b11111111; // 7812 : 255 - 0xff
      13'h1E85: dout <= 8'b11111111; // 7813 : 255 - 0xff
      13'h1E86: dout <= 8'b11111111; // 7814 : 255 - 0xff
      13'h1E87: dout <= 8'b11111111; // 7815 : 255 - 0xff
      13'h1E88: dout <= 8'b00000000; // 7816 :   0 - 0x0
      13'h1E89: dout <= 8'b00000000; // 7817 :   0 - 0x0
      13'h1E8A: dout <= 8'b00000000; // 7818 :   0 - 0x0
      13'h1E8B: dout <= 8'b00000000; // 7819 :   0 - 0x0
      13'h1E8C: dout <= 8'b11111111; // 7820 : 255 - 0xff
      13'h1E8D: dout <= 8'b11111111; // 7821 : 255 - 0xff
      13'h1E8E: dout <= 8'b11111111; // 7822 : 255 - 0xff
      13'h1E8F: dout <= 8'b11111111; // 7823 : 255 - 0xff
      13'h1E90: dout <= 8'b11110110; // 7824 : 246 - 0xf6 -- Background 0xe9
      13'h1E91: dout <= 8'b11110110; // 7825 : 246 - 0xf6
      13'h1E92: dout <= 8'b11110110; // 7826 : 246 - 0xf6
      13'h1E93: dout <= 8'b11110110; // 7827 : 246 - 0xf6
      13'h1E94: dout <= 8'b11110110; // 7828 : 246 - 0xf6
      13'h1E95: dout <= 8'b11110110; // 7829 : 246 - 0xf6
      13'h1E96: dout <= 8'b11110110; // 7830 : 246 - 0xf6
      13'h1E97: dout <= 8'b11110110; // 7831 : 246 - 0xf6
      13'h1E98: dout <= 8'b11110000; // 7832 : 240 - 0xf0
      13'h1E99: dout <= 8'b11110000; // 7833 : 240 - 0xf0
      13'h1E9A: dout <= 8'b11110000; // 7834 : 240 - 0xf0
      13'h1E9B: dout <= 8'b11110000; // 7835 : 240 - 0xf0
      13'h1E9C: dout <= 8'b11110000; // 7836 : 240 - 0xf0
      13'h1E9D: dout <= 8'b11110000; // 7837 : 240 - 0xf0
      13'h1E9E: dout <= 8'b11110000; // 7838 : 240 - 0xf0
      13'h1E9F: dout <= 8'b11110000; // 7839 : 240 - 0xf0
      13'h1EA0: dout <= 8'b11111111; // 7840 : 255 - 0xff -- Background 0xea
      13'h1EA1: dout <= 8'b11111111; // 7841 : 255 - 0xff
      13'h1EA2: dout <= 8'b11111111; // 7842 : 255 - 0xff
      13'h1EA3: dout <= 8'b11111111; // 7843 : 255 - 0xff
      13'h1EA4: dout <= 8'b00000000; // 7844 :   0 - 0x0
      13'h1EA5: dout <= 8'b11111111; // 7845 : 255 - 0xff
      13'h1EA6: dout <= 8'b11111111; // 7846 : 255 - 0xff
      13'h1EA7: dout <= 8'b00000000; // 7847 :   0 - 0x0
      13'h1EA8: dout <= 8'b11111111; // 7848 : 255 - 0xff
      13'h1EA9: dout <= 8'b11111111; // 7849 : 255 - 0xff
      13'h1EAA: dout <= 8'b11111111; // 7850 : 255 - 0xff
      13'h1EAB: dout <= 8'b11111111; // 7851 : 255 - 0xff
      13'h1EAC: dout <= 8'b00000000; // 7852 :   0 - 0x0
      13'h1EAD: dout <= 8'b00000000; // 7853 :   0 - 0x0
      13'h1EAE: dout <= 8'b00000000; // 7854 :   0 - 0x0
      13'h1EAF: dout <= 8'b00000000; // 7855 :   0 - 0x0
      13'h1EB0: dout <= 8'b01101111; // 7856 : 111 - 0x6f -- Background 0xeb
      13'h1EB1: dout <= 8'b01101111; // 7857 : 111 - 0x6f
      13'h1EB2: dout <= 8'b01101111; // 7858 : 111 - 0x6f
      13'h1EB3: dout <= 8'b01101111; // 7859 : 111 - 0x6f
      13'h1EB4: dout <= 8'b01101111; // 7860 : 111 - 0x6f
      13'h1EB5: dout <= 8'b01101111; // 7861 : 111 - 0x6f
      13'h1EB6: dout <= 8'b01101111; // 7862 : 111 - 0x6f
      13'h1EB7: dout <= 8'b01101111; // 7863 : 111 - 0x6f
      13'h1EB8: dout <= 8'b00001111; // 7864 :  15 - 0xf
      13'h1EB9: dout <= 8'b00001111; // 7865 :  15 - 0xf
      13'h1EBA: dout <= 8'b00001111; // 7866 :  15 - 0xf
      13'h1EBB: dout <= 8'b00001111; // 7867 :  15 - 0xf
      13'h1EBC: dout <= 8'b00001111; // 7868 :  15 - 0xf
      13'h1EBD: dout <= 8'b00001111; // 7869 :  15 - 0xf
      13'h1EBE: dout <= 8'b00001111; // 7870 :  15 - 0xf
      13'h1EBF: dout <= 8'b00001111; // 7871 :  15 - 0xf
      13'h1EC0: dout <= 8'b00000000; // 7872 :   0 - 0x0 -- Background 0xec
      13'h1EC1: dout <= 8'b00000000; // 7873 :   0 - 0x0
      13'h1EC2: dout <= 8'b00000000; // 7874 :   0 - 0x0
      13'h1EC3: dout <= 8'b00000000; // 7875 :   0 - 0x0
      13'h1EC4: dout <= 8'b00000000; // 7876 :   0 - 0x0
      13'h1EC5: dout <= 8'b00000000; // 7877 :   0 - 0x0
      13'h1EC6: dout <= 8'b00000000; // 7878 :   0 - 0x0
      13'h1EC7: dout <= 8'b00000000; // 7879 :   0 - 0x0
      13'h1EC8: dout <= 8'b00000000; // 7880 :   0 - 0x0
      13'h1EC9: dout <= 8'b00000000; // 7881 :   0 - 0x0
      13'h1ECA: dout <= 8'b00000000; // 7882 :   0 - 0x0
      13'h1ECB: dout <= 8'b00000000; // 7883 :   0 - 0x0
      13'h1ECC: dout <= 8'b00000000; // 7884 :   0 - 0x0
      13'h1ECD: dout <= 8'b00000000; // 7885 :   0 - 0x0
      13'h1ECE: dout <= 8'b00000000; // 7886 :   0 - 0x0
      13'h1ECF: dout <= 8'b00000000; // 7887 :   0 - 0x0
      13'h1ED0: dout <= 8'b00000000; // 7888 :   0 - 0x0 -- Background 0xed
      13'h1ED1: dout <= 8'b00000000; // 7889 :   0 - 0x0
      13'h1ED2: dout <= 8'b00000000; // 7890 :   0 - 0x0
      13'h1ED3: dout <= 8'b00000000; // 7891 :   0 - 0x0
      13'h1ED4: dout <= 8'b00000000; // 7892 :   0 - 0x0
      13'h1ED5: dout <= 8'b00000000; // 7893 :   0 - 0x0
      13'h1ED6: dout <= 8'b00000000; // 7894 :   0 - 0x0
      13'h1ED7: dout <= 8'b00000000; // 7895 :   0 - 0x0
      13'h1ED8: dout <= 8'b00000000; // 7896 :   0 - 0x0
      13'h1ED9: dout <= 8'b00000000; // 7897 :   0 - 0x0
      13'h1EDA: dout <= 8'b00000000; // 7898 :   0 - 0x0
      13'h1EDB: dout <= 8'b00000000; // 7899 :   0 - 0x0
      13'h1EDC: dout <= 8'b00000000; // 7900 :   0 - 0x0
      13'h1EDD: dout <= 8'b00000000; // 7901 :   0 - 0x0
      13'h1EDE: dout <= 8'b00000000; // 7902 :   0 - 0x0
      13'h1EDF: dout <= 8'b00000000; // 7903 :   0 - 0x0
      13'h1EE0: dout <= 8'b00000000; // 7904 :   0 - 0x0 -- Background 0xee
      13'h1EE1: dout <= 8'b00000000; // 7905 :   0 - 0x0
      13'h1EE2: dout <= 8'b00000000; // 7906 :   0 - 0x0
      13'h1EE3: dout <= 8'b00000000; // 7907 :   0 - 0x0
      13'h1EE4: dout <= 8'b00000000; // 7908 :   0 - 0x0
      13'h1EE5: dout <= 8'b00000000; // 7909 :   0 - 0x0
      13'h1EE6: dout <= 8'b00000000; // 7910 :   0 - 0x0
      13'h1EE7: dout <= 8'b00000000; // 7911 :   0 - 0x0
      13'h1EE8: dout <= 8'b00000000; // 7912 :   0 - 0x0
      13'h1EE9: dout <= 8'b00000000; // 7913 :   0 - 0x0
      13'h1EEA: dout <= 8'b00000000; // 7914 :   0 - 0x0
      13'h1EEB: dout <= 8'b00000000; // 7915 :   0 - 0x0
      13'h1EEC: dout <= 8'b00000000; // 7916 :   0 - 0x0
      13'h1EED: dout <= 8'b00000000; // 7917 :   0 - 0x0
      13'h1EEE: dout <= 8'b00000000; // 7918 :   0 - 0x0
      13'h1EEF: dout <= 8'b00000000; // 7919 :   0 - 0x0
      13'h1EF0: dout <= 8'b00000000; // 7920 :   0 - 0x0 -- Background 0xef
      13'h1EF1: dout <= 8'b00000000; // 7921 :   0 - 0x0
      13'h1EF2: dout <= 8'b00000000; // 7922 :   0 - 0x0
      13'h1EF3: dout <= 8'b00000000; // 7923 :   0 - 0x0
      13'h1EF4: dout <= 8'b00000000; // 7924 :   0 - 0x0
      13'h1EF5: dout <= 8'b00000000; // 7925 :   0 - 0x0
      13'h1EF6: dout <= 8'b00000000; // 7926 :   0 - 0x0
      13'h1EF7: dout <= 8'b00000000; // 7927 :   0 - 0x0
      13'h1EF8: dout <= 8'b00000000; // 7928 :   0 - 0x0
      13'h1EF9: dout <= 8'b00000000; // 7929 :   0 - 0x0
      13'h1EFA: dout <= 8'b00000000; // 7930 :   0 - 0x0
      13'h1EFB: dout <= 8'b00000000; // 7931 :   0 - 0x0
      13'h1EFC: dout <= 8'b00000000; // 7932 :   0 - 0x0
      13'h1EFD: dout <= 8'b00000000; // 7933 :   0 - 0x0
      13'h1EFE: dout <= 8'b00000000; // 7934 :   0 - 0x0
      13'h1EFF: dout <= 8'b00000000; // 7935 :   0 - 0x0
      13'h1F00: dout <= 8'b11111111; // 7936 : 255 - 0xff -- Background 0xf0
      13'h1F01: dout <= 8'b11111111; // 7937 : 255 - 0xff
      13'h1F02: dout <= 8'b11111111; // 7938 : 255 - 0xff
      13'h1F03: dout <= 8'b11111111; // 7939 : 255 - 0xff
      13'h1F04: dout <= 8'b11111111; // 7940 : 255 - 0xff
      13'h1F05: dout <= 8'b11111111; // 7941 : 255 - 0xff
      13'h1F06: dout <= 8'b11111111; // 7942 : 255 - 0xff
      13'h1F07: dout <= 8'b11111111; // 7943 : 255 - 0xff
      13'h1F08: dout <= 8'b11111111; // 7944 : 255 - 0xff
      13'h1F09: dout <= 8'b11111111; // 7945 : 255 - 0xff
      13'h1F0A: dout <= 8'b11111111; // 7946 : 255 - 0xff
      13'h1F0B: dout <= 8'b11111111; // 7947 : 255 - 0xff
      13'h1F0C: dout <= 8'b11111111; // 7948 : 255 - 0xff
      13'h1F0D: dout <= 8'b11111111; // 7949 : 255 - 0xff
      13'h1F0E: dout <= 8'b11111111; // 7950 : 255 - 0xff
      13'h1F0F: dout <= 8'b11111111; // 7951 : 255 - 0xff
      13'h1F10: dout <= 8'b11111111; // 7952 : 255 - 0xff -- Background 0xf1
      13'h1F11: dout <= 8'b11111111; // 7953 : 255 - 0xff
      13'h1F12: dout <= 8'b11111111; // 7954 : 255 - 0xff
      13'h1F13: dout <= 8'b11111111; // 7955 : 255 - 0xff
      13'h1F14: dout <= 8'b11111111; // 7956 : 255 - 0xff
      13'h1F15: dout <= 8'b11111111; // 7957 : 255 - 0xff
      13'h1F16: dout <= 8'b11111111; // 7958 : 255 - 0xff
      13'h1F17: dout <= 8'b11111111; // 7959 : 255 - 0xff
      13'h1F18: dout <= 8'b11111111; // 7960 : 255 - 0xff
      13'h1F19: dout <= 8'b11111111; // 7961 : 255 - 0xff
      13'h1F1A: dout <= 8'b11111111; // 7962 : 255 - 0xff
      13'h1F1B: dout <= 8'b11111111; // 7963 : 255 - 0xff
      13'h1F1C: dout <= 8'b11111111; // 7964 : 255 - 0xff
      13'h1F1D: dout <= 8'b11111111; // 7965 : 255 - 0xff
      13'h1F1E: dout <= 8'b11111111; // 7966 : 255 - 0xff
      13'h1F1F: dout <= 8'b11111111; // 7967 : 255 - 0xff
      13'h1F20: dout <= 8'b11111111; // 7968 : 255 - 0xff -- Background 0xf2
      13'h1F21: dout <= 8'b11111111; // 7969 : 255 - 0xff
      13'h1F22: dout <= 8'b11111111; // 7970 : 255 - 0xff
      13'h1F23: dout <= 8'b11111111; // 7971 : 255 - 0xff
      13'h1F24: dout <= 8'b11111111; // 7972 : 255 - 0xff
      13'h1F25: dout <= 8'b11111111; // 7973 : 255 - 0xff
      13'h1F26: dout <= 8'b11111111; // 7974 : 255 - 0xff
      13'h1F27: dout <= 8'b11111111; // 7975 : 255 - 0xff
      13'h1F28: dout <= 8'b11111111; // 7976 : 255 - 0xff
      13'h1F29: dout <= 8'b11111111; // 7977 : 255 - 0xff
      13'h1F2A: dout <= 8'b11111111; // 7978 : 255 - 0xff
      13'h1F2B: dout <= 8'b11111111; // 7979 : 255 - 0xff
      13'h1F2C: dout <= 8'b11111111; // 7980 : 255 - 0xff
      13'h1F2D: dout <= 8'b11111111; // 7981 : 255 - 0xff
      13'h1F2E: dout <= 8'b11111111; // 7982 : 255 - 0xff
      13'h1F2F: dout <= 8'b11111111; // 7983 : 255 - 0xff
      13'h1F30: dout <= 8'b11111111; // 7984 : 255 - 0xff -- Background 0xf3
      13'h1F31: dout <= 8'b11111111; // 7985 : 255 - 0xff
      13'h1F32: dout <= 8'b11111111; // 7986 : 255 - 0xff
      13'h1F33: dout <= 8'b11111111; // 7987 : 255 - 0xff
      13'h1F34: dout <= 8'b11111111; // 7988 : 255 - 0xff
      13'h1F35: dout <= 8'b11111111; // 7989 : 255 - 0xff
      13'h1F36: dout <= 8'b11111111; // 7990 : 255 - 0xff
      13'h1F37: dout <= 8'b11111111; // 7991 : 255 - 0xff
      13'h1F38: dout <= 8'b11111111; // 7992 : 255 - 0xff
      13'h1F39: dout <= 8'b11111111; // 7993 : 255 - 0xff
      13'h1F3A: dout <= 8'b11111111; // 7994 : 255 - 0xff
      13'h1F3B: dout <= 8'b11111111; // 7995 : 255 - 0xff
      13'h1F3C: dout <= 8'b11111111; // 7996 : 255 - 0xff
      13'h1F3D: dout <= 8'b11111111; // 7997 : 255 - 0xff
      13'h1F3E: dout <= 8'b11111111; // 7998 : 255 - 0xff
      13'h1F3F: dout <= 8'b11111111; // 7999 : 255 - 0xff
      13'h1F40: dout <= 8'b11111111; // 8000 : 255 - 0xff -- Background 0xf4
      13'h1F41: dout <= 8'b11111111; // 8001 : 255 - 0xff
      13'h1F42: dout <= 8'b11111111; // 8002 : 255 - 0xff
      13'h1F43: dout <= 8'b11111111; // 8003 : 255 - 0xff
      13'h1F44: dout <= 8'b11111111; // 8004 : 255 - 0xff
      13'h1F45: dout <= 8'b11111111; // 8005 : 255 - 0xff
      13'h1F46: dout <= 8'b11111111; // 8006 : 255 - 0xff
      13'h1F47: dout <= 8'b11111111; // 8007 : 255 - 0xff
      13'h1F48: dout <= 8'b11111111; // 8008 : 255 - 0xff
      13'h1F49: dout <= 8'b11111111; // 8009 : 255 - 0xff
      13'h1F4A: dout <= 8'b11111111; // 8010 : 255 - 0xff
      13'h1F4B: dout <= 8'b11111111; // 8011 : 255 - 0xff
      13'h1F4C: dout <= 8'b11111111; // 8012 : 255 - 0xff
      13'h1F4D: dout <= 8'b11111111; // 8013 : 255 - 0xff
      13'h1F4E: dout <= 8'b11111111; // 8014 : 255 - 0xff
      13'h1F4F: dout <= 8'b11111111; // 8015 : 255 - 0xff
      13'h1F50: dout <= 8'b11111111; // 8016 : 255 - 0xff -- Background 0xf5
      13'h1F51: dout <= 8'b11111111; // 8017 : 255 - 0xff
      13'h1F52: dout <= 8'b11111111; // 8018 : 255 - 0xff
      13'h1F53: dout <= 8'b11111111; // 8019 : 255 - 0xff
      13'h1F54: dout <= 8'b11111111; // 8020 : 255 - 0xff
      13'h1F55: dout <= 8'b11111111; // 8021 : 255 - 0xff
      13'h1F56: dout <= 8'b11111111; // 8022 : 255 - 0xff
      13'h1F57: dout <= 8'b11111111; // 8023 : 255 - 0xff
      13'h1F58: dout <= 8'b11111111; // 8024 : 255 - 0xff
      13'h1F59: dout <= 8'b11111111; // 8025 : 255 - 0xff
      13'h1F5A: dout <= 8'b11111111; // 8026 : 255 - 0xff
      13'h1F5B: dout <= 8'b11111111; // 8027 : 255 - 0xff
      13'h1F5C: dout <= 8'b11111111; // 8028 : 255 - 0xff
      13'h1F5D: dout <= 8'b11111111; // 8029 : 255 - 0xff
      13'h1F5E: dout <= 8'b11111111; // 8030 : 255 - 0xff
      13'h1F5F: dout <= 8'b11111111; // 8031 : 255 - 0xff
      13'h1F60: dout <= 8'b11111111; // 8032 : 255 - 0xff -- Background 0xf6
      13'h1F61: dout <= 8'b11111111; // 8033 : 255 - 0xff
      13'h1F62: dout <= 8'b11111111; // 8034 : 255 - 0xff
      13'h1F63: dout <= 8'b11111111; // 8035 : 255 - 0xff
      13'h1F64: dout <= 8'b11111111; // 8036 : 255 - 0xff
      13'h1F65: dout <= 8'b11111111; // 8037 : 255 - 0xff
      13'h1F66: dout <= 8'b11111111; // 8038 : 255 - 0xff
      13'h1F67: dout <= 8'b11111111; // 8039 : 255 - 0xff
      13'h1F68: dout <= 8'b11111111; // 8040 : 255 - 0xff
      13'h1F69: dout <= 8'b11111111; // 8041 : 255 - 0xff
      13'h1F6A: dout <= 8'b11111111; // 8042 : 255 - 0xff
      13'h1F6B: dout <= 8'b11111111; // 8043 : 255 - 0xff
      13'h1F6C: dout <= 8'b11111111; // 8044 : 255 - 0xff
      13'h1F6D: dout <= 8'b11111111; // 8045 : 255 - 0xff
      13'h1F6E: dout <= 8'b11111111; // 8046 : 255 - 0xff
      13'h1F6F: dout <= 8'b11111111; // 8047 : 255 - 0xff
      13'h1F70: dout <= 8'b11111111; // 8048 : 255 - 0xff -- Background 0xf7
      13'h1F71: dout <= 8'b11111111; // 8049 : 255 - 0xff
      13'h1F72: dout <= 8'b11111111; // 8050 : 255 - 0xff
      13'h1F73: dout <= 8'b11111111; // 8051 : 255 - 0xff
      13'h1F74: dout <= 8'b11111111; // 8052 : 255 - 0xff
      13'h1F75: dout <= 8'b11111111; // 8053 : 255 - 0xff
      13'h1F76: dout <= 8'b11111111; // 8054 : 255 - 0xff
      13'h1F77: dout <= 8'b11111111; // 8055 : 255 - 0xff
      13'h1F78: dout <= 8'b11111111; // 8056 : 255 - 0xff
      13'h1F79: dout <= 8'b11111111; // 8057 : 255 - 0xff
      13'h1F7A: dout <= 8'b11111111; // 8058 : 255 - 0xff
      13'h1F7B: dout <= 8'b11111111; // 8059 : 255 - 0xff
      13'h1F7C: dout <= 8'b11111111; // 8060 : 255 - 0xff
      13'h1F7D: dout <= 8'b11111111; // 8061 : 255 - 0xff
      13'h1F7E: dout <= 8'b11111111; // 8062 : 255 - 0xff
      13'h1F7F: dout <= 8'b11111111; // 8063 : 255 - 0xff
      13'h1F80: dout <= 8'b11111111; // 8064 : 255 - 0xff -- Background 0xf8
      13'h1F81: dout <= 8'b11111111; // 8065 : 255 - 0xff
      13'h1F82: dout <= 8'b11111111; // 8066 : 255 - 0xff
      13'h1F83: dout <= 8'b11111111; // 8067 : 255 - 0xff
      13'h1F84: dout <= 8'b11111111; // 8068 : 255 - 0xff
      13'h1F85: dout <= 8'b11111111; // 8069 : 255 - 0xff
      13'h1F86: dout <= 8'b11111111; // 8070 : 255 - 0xff
      13'h1F87: dout <= 8'b11111111; // 8071 : 255 - 0xff
      13'h1F88: dout <= 8'b11111111; // 8072 : 255 - 0xff
      13'h1F89: dout <= 8'b11111111; // 8073 : 255 - 0xff
      13'h1F8A: dout <= 8'b11111111; // 8074 : 255 - 0xff
      13'h1F8B: dout <= 8'b11111111; // 8075 : 255 - 0xff
      13'h1F8C: dout <= 8'b11111111; // 8076 : 255 - 0xff
      13'h1F8D: dout <= 8'b11111111; // 8077 : 255 - 0xff
      13'h1F8E: dout <= 8'b11111111; // 8078 : 255 - 0xff
      13'h1F8F: dout <= 8'b11111111; // 8079 : 255 - 0xff
      13'h1F90: dout <= 8'b11111111; // 8080 : 255 - 0xff -- Background 0xf9
      13'h1F91: dout <= 8'b11111111; // 8081 : 255 - 0xff
      13'h1F92: dout <= 8'b11111111; // 8082 : 255 - 0xff
      13'h1F93: dout <= 8'b11111111; // 8083 : 255 - 0xff
      13'h1F94: dout <= 8'b11111111; // 8084 : 255 - 0xff
      13'h1F95: dout <= 8'b11111111; // 8085 : 255 - 0xff
      13'h1F96: dout <= 8'b11111111; // 8086 : 255 - 0xff
      13'h1F97: dout <= 8'b11111111; // 8087 : 255 - 0xff
      13'h1F98: dout <= 8'b11111111; // 8088 : 255 - 0xff
      13'h1F99: dout <= 8'b11111111; // 8089 : 255 - 0xff
      13'h1F9A: dout <= 8'b11111111; // 8090 : 255 - 0xff
      13'h1F9B: dout <= 8'b11111111; // 8091 : 255 - 0xff
      13'h1F9C: dout <= 8'b11111111; // 8092 : 255 - 0xff
      13'h1F9D: dout <= 8'b11111111; // 8093 : 255 - 0xff
      13'h1F9E: dout <= 8'b11111111; // 8094 : 255 - 0xff
      13'h1F9F: dout <= 8'b11111111; // 8095 : 255 - 0xff
      13'h1FA0: dout <= 8'b11111111; // 8096 : 255 - 0xff -- Background 0xfa
      13'h1FA1: dout <= 8'b11111111; // 8097 : 255 - 0xff
      13'h1FA2: dout <= 8'b11111111; // 8098 : 255 - 0xff
      13'h1FA3: dout <= 8'b11111111; // 8099 : 255 - 0xff
      13'h1FA4: dout <= 8'b11111111; // 8100 : 255 - 0xff
      13'h1FA5: dout <= 8'b11111111; // 8101 : 255 - 0xff
      13'h1FA6: dout <= 8'b11111111; // 8102 : 255 - 0xff
      13'h1FA7: dout <= 8'b11111111; // 8103 : 255 - 0xff
      13'h1FA8: dout <= 8'b11111111; // 8104 : 255 - 0xff
      13'h1FA9: dout <= 8'b11111111; // 8105 : 255 - 0xff
      13'h1FAA: dout <= 8'b11111111; // 8106 : 255 - 0xff
      13'h1FAB: dout <= 8'b11111111; // 8107 : 255 - 0xff
      13'h1FAC: dout <= 8'b11111111; // 8108 : 255 - 0xff
      13'h1FAD: dout <= 8'b11111111; // 8109 : 255 - 0xff
      13'h1FAE: dout <= 8'b11111111; // 8110 : 255 - 0xff
      13'h1FAF: dout <= 8'b11111111; // 8111 : 255 - 0xff
      13'h1FB0: dout <= 8'b11111111; // 8112 : 255 - 0xff -- Background 0xfb
      13'h1FB1: dout <= 8'b11111111; // 8113 : 255 - 0xff
      13'h1FB2: dout <= 8'b11111111; // 8114 : 255 - 0xff
      13'h1FB3: dout <= 8'b11111111; // 8115 : 255 - 0xff
      13'h1FB4: dout <= 8'b11111111; // 8116 : 255 - 0xff
      13'h1FB5: dout <= 8'b11111111; // 8117 : 255 - 0xff
      13'h1FB6: dout <= 8'b11111111; // 8118 : 255 - 0xff
      13'h1FB7: dout <= 8'b11111111; // 8119 : 255 - 0xff
      13'h1FB8: dout <= 8'b11111111; // 8120 : 255 - 0xff
      13'h1FB9: dout <= 8'b11111111; // 8121 : 255 - 0xff
      13'h1FBA: dout <= 8'b11111111; // 8122 : 255 - 0xff
      13'h1FBB: dout <= 8'b11111111; // 8123 : 255 - 0xff
      13'h1FBC: dout <= 8'b11111111; // 8124 : 255 - 0xff
      13'h1FBD: dout <= 8'b11111111; // 8125 : 255 - 0xff
      13'h1FBE: dout <= 8'b11111111; // 8126 : 255 - 0xff
      13'h1FBF: dout <= 8'b11111111; // 8127 : 255 - 0xff
      13'h1FC0: dout <= 8'b11111111; // 8128 : 255 - 0xff -- Background 0xfc
      13'h1FC1: dout <= 8'b11111111; // 8129 : 255 - 0xff
      13'h1FC2: dout <= 8'b11111111; // 8130 : 255 - 0xff
      13'h1FC3: dout <= 8'b11111111; // 8131 : 255 - 0xff
      13'h1FC4: dout <= 8'b11111111; // 8132 : 255 - 0xff
      13'h1FC5: dout <= 8'b11111111; // 8133 : 255 - 0xff
      13'h1FC6: dout <= 8'b11111111; // 8134 : 255 - 0xff
      13'h1FC7: dout <= 8'b11111111; // 8135 : 255 - 0xff
      13'h1FC8: dout <= 8'b11111111; // 8136 : 255 - 0xff
      13'h1FC9: dout <= 8'b11111111; // 8137 : 255 - 0xff
      13'h1FCA: dout <= 8'b11111111; // 8138 : 255 - 0xff
      13'h1FCB: dout <= 8'b11111111; // 8139 : 255 - 0xff
      13'h1FCC: dout <= 8'b11111111; // 8140 : 255 - 0xff
      13'h1FCD: dout <= 8'b11111111; // 8141 : 255 - 0xff
      13'h1FCE: dout <= 8'b11111111; // 8142 : 255 - 0xff
      13'h1FCF: dout <= 8'b11111111; // 8143 : 255 - 0xff
      13'h1FD0: dout <= 8'b11111111; // 8144 : 255 - 0xff -- Background 0xfd
      13'h1FD1: dout <= 8'b11111111; // 8145 : 255 - 0xff
      13'h1FD2: dout <= 8'b11111111; // 8146 : 255 - 0xff
      13'h1FD3: dout <= 8'b11111111; // 8147 : 255 - 0xff
      13'h1FD4: dout <= 8'b11111111; // 8148 : 255 - 0xff
      13'h1FD5: dout <= 8'b11111111; // 8149 : 255 - 0xff
      13'h1FD6: dout <= 8'b11111111; // 8150 : 255 - 0xff
      13'h1FD7: dout <= 8'b11111111; // 8151 : 255 - 0xff
      13'h1FD8: dout <= 8'b11111111; // 8152 : 255 - 0xff
      13'h1FD9: dout <= 8'b11111111; // 8153 : 255 - 0xff
      13'h1FDA: dout <= 8'b11111111; // 8154 : 255 - 0xff
      13'h1FDB: dout <= 8'b11111111; // 8155 : 255 - 0xff
      13'h1FDC: dout <= 8'b11111111; // 8156 : 255 - 0xff
      13'h1FDD: dout <= 8'b11111111; // 8157 : 255 - 0xff
      13'h1FDE: dout <= 8'b11111111; // 8158 : 255 - 0xff
      13'h1FDF: dout <= 8'b11111111; // 8159 : 255 - 0xff
      13'h1FE0: dout <= 8'b11111111; // 8160 : 255 - 0xff -- Background 0xfe
      13'h1FE1: dout <= 8'b11111111; // 8161 : 255 - 0xff
      13'h1FE2: dout <= 8'b11111111; // 8162 : 255 - 0xff
      13'h1FE3: dout <= 8'b11111111; // 8163 : 255 - 0xff
      13'h1FE4: dout <= 8'b11111111; // 8164 : 255 - 0xff
      13'h1FE5: dout <= 8'b11111111; // 8165 : 255 - 0xff
      13'h1FE6: dout <= 8'b11111111; // 8166 : 255 - 0xff
      13'h1FE7: dout <= 8'b11111111; // 8167 : 255 - 0xff
      13'h1FE8: dout <= 8'b11111111; // 8168 : 255 - 0xff
      13'h1FE9: dout <= 8'b11111111; // 8169 : 255 - 0xff
      13'h1FEA: dout <= 8'b11111111; // 8170 : 255 - 0xff
      13'h1FEB: dout <= 8'b11111111; // 8171 : 255 - 0xff
      13'h1FEC: dout <= 8'b11111111; // 8172 : 255 - 0xff
      13'h1FED: dout <= 8'b11111111; // 8173 : 255 - 0xff
      13'h1FEE: dout <= 8'b11111111; // 8174 : 255 - 0xff
      13'h1FEF: dout <= 8'b11111111; // 8175 : 255 - 0xff
      13'h1FF0: dout <= 8'b11111111; // 8176 : 255 - 0xff -- Background 0xff
      13'h1FF1: dout <= 8'b11111111; // 8177 : 255 - 0xff
      13'h1FF2: dout <= 8'b11111111; // 8178 : 255 - 0xff
      13'h1FF3: dout <= 8'b11111111; // 8179 : 255 - 0xff
      13'h1FF4: dout <= 8'b11111111; // 8180 : 255 - 0xff
      13'h1FF5: dout <= 8'b11111111; // 8181 : 255 - 0xff
      13'h1FF6: dout <= 8'b11111111; // 8182 : 255 - 0xff
      13'h1FF7: dout <= 8'b11111111; // 8183 : 255 - 0xff
      13'h1FF8: dout <= 8'b11111111; // 8184 : 255 - 0xff
      13'h1FF9: dout <= 8'b11111111; // 8185 : 255 - 0xff
      13'h1FFA: dout <= 8'b11111111; // 8186 : 255 - 0xff
      13'h1FFB: dout <= 8'b11111111; // 8187 : 255 - 0xff
      13'h1FFC: dout <= 8'b11111111; // 8188 : 255 - 0xff
      13'h1FFD: dout <= 8'b11111111; // 8189 : 255 - 0xff
      13'h1FFE: dout <= 8'b11111111; // 8190 : 255 - 0xff
      13'h1FFF: dout <= 8'b11111111; // 8191 : 255 - 0xff
    endcase
  end

endmodule
