--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE WITH ONLY ONE COLOR PLANE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: sprilo_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_SPRILO_color0 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_SPRILO_color0;

architecture BEHAVIORAL of ROM_PTABLE_SPRILO_color0 is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
    "00000000", --    0 -  0x0  :    0 - 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000000", --   16 - 0x10  :    0 - 0x0
    "00000000", --   17 - 0x11  :    0 - 0x0
    "00000000", --   18 - 0x12  :    0 - 0x0
    "00000000", --   19 - 0x13  :    0 - 0x0
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00000000", --   21 - 0x15  :    0 - 0x0
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0
    "00000000", --   33 - 0x21  :    0 - 0x0
    "00000000", --   34 - 0x22  :    0 - 0x0
    "00000000", --   35 - 0x23  :    0 - 0x0
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00000000", --   51 - 0x33  :    0 - 0x0
    "00000000", --   52 - 0x34  :    0 - 0x0
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000000", --   54 - 0x36  :    0 - 0x0
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0
    "01111110", --   65 - 0x41  :  126 - 0x7e
    "01111110", --   66 - 0x42  :  126 - 0x7e
    "00111100", --   67 - 0x43  :   60 - 0x3c
    "00111100", --   68 - 0x44  :   60 - 0x3c
    "01111110", --   69 - 0x45  :  126 - 0x7e
    "01011010", --   70 - 0x46  :   90 - 0x5a
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0
    "01100110", --   73 - 0x49  :  102 - 0x66
    "01111100", --   74 - 0x4a  :  124 - 0x7c
    "01111110", --   75 - 0x4b  :  126 - 0x7e
    "01111110", --   76 - 0x4c  :  126 - 0x7e
    "01111100", --   77 - 0x4d  :  124 - 0x7c
    "01100110", --   78 - 0x4e  :  102 - 0x66
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00010000", --   80 - 0x50  :   16 - 0x10
    "00011000", --   81 - 0x51  :   24 - 0x18
    "00111000", --   82 - 0x52  :   56 - 0x38
    "11111110", --   83 - 0x53  :  254 - 0xfe
    "01111101", --   84 - 0x54  :  125 - 0x7d
    "00011100", --   85 - 0x55  :   28 - 0x1c
    "00010000", --   86 - 0x56  :   16 - 0x10
    "00001000", --   87 - 0x57  :    8 - 0x8
    "00000000", --   88 - 0x58  :    0 - 0x0
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "00000000", --  144 - 0x90  :    0 - 0x0
    "00000000", --  145 - 0x91  :    0 - 0x0
    "00000000", --  146 - 0x92  :    0 - 0x0
    "00000000", --  147 - 0x93  :    0 - 0x0
    "00000000", --  148 - 0x94  :    0 - 0x0
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "00000000", --  164 - 0xa4  :    0 - 0x0
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "00000000", --  194 - 0xc2  :    0 - 0x0
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00000000", --  196 - 0xc4  :    0 - 0x0
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00000000", --  208 - 0xd0  :    0 - 0x0
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00000000", --  211 - 0xd3  :    0 - 0x0
    "00000000", --  212 - 0xd4  :    0 - 0x0
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00000000", --  228 - 0xe4  :    0 - 0x0
    "00000000", --  229 - 0xe5  :    0 - 0x0
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0
    "00000000", --  241 - 0xf1  :    0 - 0x0
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "00000000", --  243 - 0xf3  :    0 - 0x0
    "00000000", --  244 - 0xf4  :    0 - 0x0
    "00000000", --  245 - 0xf5  :    0 - 0x0
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00000000", --  272 - 0x110  :    0 - 0x0
    "00000000", --  273 - 0x111  :    0 - 0x0
    "00000000", --  274 - 0x112  :    0 - 0x0
    "00000000", --  275 - 0x113  :    0 - 0x0
    "00000000", --  276 - 0x114  :    0 - 0x0
    "00000000", --  277 - 0x115  :    0 - 0x0
    "00000000", --  278 - 0x116  :    0 - 0x0
    "00000000", --  279 - 0x117  :    0 - 0x0
    "00000000", --  280 - 0x118  :    0 - 0x0
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00000000", --  283 - 0x11b  :    0 - 0x0
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000000", --  298 - 0x12a  :    0 - 0x0
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0
    "00000000", --  305 - 0x131  :    0 - 0x0
    "00000000", --  306 - 0x132  :    0 - 0x0
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "00000000", --  309 - 0x135  :    0 - 0x0
    "00000000", --  310 - 0x136  :    0 - 0x0
    "00000000", --  311 - 0x137  :    0 - 0x0
    "00000000", --  312 - 0x138  :    0 - 0x0
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "00000000", --  324 - 0x144  :    0 - 0x0
    "00000000", --  325 - 0x145  :    0 - 0x0
    "00000000", --  326 - 0x146  :    0 - 0x0
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00000000", --  328 - 0x148  :    0 - 0x0
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000000", --  330 - 0x14a  :    0 - 0x0
    "00000000", --  331 - 0x14b  :    0 - 0x0
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00000000", --  336 - 0x150  :    0 - 0x0
    "00000000", --  337 - 0x151  :    0 - 0x0
    "00000000", --  338 - 0x152  :    0 - 0x0
    "00000000", --  339 - 0x153  :    0 - 0x0
    "00000000", --  340 - 0x154  :    0 - 0x0
    "00000000", --  341 - 0x155  :    0 - 0x0
    "00000000", --  342 - 0x156  :    0 - 0x0
    "00000000", --  343 - 0x157  :    0 - 0x0
    "00000000", --  344 - 0x158  :    0 - 0x0
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000000", --  376 - 0x178  :    0 - 0x0
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00000000", --  379 - 0x17b  :    0 - 0x0
    "00000000", --  380 - 0x17c  :    0 - 0x0
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000000", --  384 - 0x180  :    0 - 0x0
    "00000000", --  385 - 0x181  :    0 - 0x0
    "00000000", --  386 - 0x182  :    0 - 0x0
    "00000000", --  387 - 0x183  :    0 - 0x0
    "00000000", --  388 - 0x184  :    0 - 0x0
    "00000000", --  389 - 0x185  :    0 - 0x0
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00000000", --  400 - 0x190  :    0 - 0x0
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000000", --  403 - 0x193  :    0 - 0x0
    "00000000", --  404 - 0x194  :    0 - 0x0
    "00000000", --  405 - 0x195  :    0 - 0x0
    "00000000", --  406 - 0x196  :    0 - 0x0
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00000000", --  408 - 0x198  :    0 - 0x0
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "00000000", --  411 - 0x19b  :    0 - 0x0
    "00000000", --  412 - 0x19c  :    0 - 0x0
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00000000", --  416 - 0x1a0  :    0 - 0x0
    "00000000", --  417 - 0x1a1  :    0 - 0x0
    "00000000", --  418 - 0x1a2  :    0 - 0x0
    "00000000", --  419 - 0x1a3  :    0 - 0x0
    "00000000", --  420 - 0x1a4  :    0 - 0x0
    "00000000", --  421 - 0x1a5  :    0 - 0x0
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "00000000", --  424 - 0x1a8  :    0 - 0x0
    "00000000", --  425 - 0x1a9  :    0 - 0x0
    "00000000", --  426 - 0x1aa  :    0 - 0x0
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00000000", --  434 - 0x1b2  :    0 - 0x0
    "00000000", --  435 - 0x1b3  :    0 - 0x0
    "00000000", --  436 - 0x1b4  :    0 - 0x0
    "00000000", --  437 - 0x1b5  :    0 - 0x0
    "00000000", --  438 - 0x1b6  :    0 - 0x0
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "00000000", --  440 - 0x1b8  :    0 - 0x0
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "00000000", --  453 - 0x1c5  :    0 - 0x0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "00000000", --  467 - 0x1d3  :    0 - 0x0
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "00000000", --  469 - 0x1d5  :    0 - 0x0
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "00000000", --  485 - 0x1e5  :    0 - 0x0
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00000000", --  500 - 0x1f4  :    0 - 0x0
    "00000000", --  501 - 0x1f5  :    0 - 0x0
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "00000000", --  504 - 0x1f8  :    0 - 0x0
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00000000", --  528 - 0x210  :    0 - 0x0
    "00000000", --  529 - 0x211  :    0 - 0x0
    "00000000", --  530 - 0x212  :    0 - 0x0
    "00000000", --  531 - 0x213  :    0 - 0x0
    "00000000", --  532 - 0x214  :    0 - 0x0
    "00000000", --  533 - 0x215  :    0 - 0x0
    "00000000", --  534 - 0x216  :    0 - 0x0
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00000000", --  536 - 0x218  :    0 - 0x0
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000000", --  544 - 0x220  :    0 - 0x0
    "00000000", --  545 - 0x221  :    0 - 0x0
    "00000000", --  546 - 0x222  :    0 - 0x0
    "00000000", --  547 - 0x223  :    0 - 0x0
    "00000000", --  548 - 0x224  :    0 - 0x0
    "00000000", --  549 - 0x225  :    0 - 0x0
    "00000000", --  550 - 0x226  :    0 - 0x0
    "00000000", --  551 - 0x227  :    0 - 0x0
    "00000000", --  552 - 0x228  :    0 - 0x0
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000000", --  560 - 0x230  :    0 - 0x0
    "00000000", --  561 - 0x231  :    0 - 0x0
    "00000000", --  562 - 0x232  :    0 - 0x0
    "00000000", --  563 - 0x233  :    0 - 0x0
    "00000000", --  564 - 0x234  :    0 - 0x0
    "00000000", --  565 - 0x235  :    0 - 0x0
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00000000", --  568 - 0x238  :    0 - 0x0
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00000000", --  584 - 0x248  :    0 - 0x0
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000000", --  592 - 0x250  :    0 - 0x0
    "00000000", --  593 - 0x251  :    0 - 0x0
    "00000000", --  594 - 0x252  :    0 - 0x0
    "00000000", --  595 - 0x253  :    0 - 0x0
    "00000000", --  596 - 0x254  :    0 - 0x0
    "00000000", --  597 - 0x255  :    0 - 0x0
    "00000000", --  598 - 0x256  :    0 - 0x0
    "00000000", --  599 - 0x257  :    0 - 0x0
    "00000000", --  600 - 0x258  :    0 - 0x0
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0
    "00000000", --  609 - 0x261  :    0 - 0x0
    "00000000", --  610 - 0x262  :    0 - 0x0
    "00000000", --  611 - 0x263  :    0 - 0x0
    "00000000", --  612 - 0x264  :    0 - 0x0
    "00000000", --  613 - 0x265  :    0 - 0x0
    "00000000", --  614 - 0x266  :    0 - 0x0
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0
    "00000000", --  625 - 0x271  :    0 - 0x0
    "00000000", --  626 - 0x272  :    0 - 0x0
    "00000000", --  627 - 0x273  :    0 - 0x0
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000000", --  629 - 0x275  :    0 - 0x0
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0
    "00000000", --  633 - 0x279  :    0 - 0x0
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "00000000", --  635 - 0x27b  :    0 - 0x0
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0
    "00000000", --  657 - 0x291  :    0 - 0x0
    "00000000", --  658 - 0x292  :    0 - 0x0
    "00000000", --  659 - 0x293  :    0 - 0x0
    "00000000", --  660 - 0x294  :    0 - 0x0
    "00000000", --  661 - 0x295  :    0 - 0x0
    "00000000", --  662 - 0x296  :    0 - 0x0
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00000000", --  672 - 0x2a0  :    0 - 0x0
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "00000000", --  674 - 0x2a2  :    0 - 0x0
    "00000000", --  675 - 0x2a3  :    0 - 0x0
    "00000000", --  676 - 0x2a4  :    0 - 0x0
    "00000000", --  677 - 0x2a5  :    0 - 0x0
    "00000000", --  678 - 0x2a6  :    0 - 0x0
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "00000000", --  680 - 0x2a8  :    0 - 0x0
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "00000000", --  686 - 0x2ae  :    0 - 0x0
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "00000000", --  688 - 0x2b0  :    0 - 0x0
    "00000000", --  689 - 0x2b1  :    0 - 0x0
    "00000000", --  690 - 0x2b2  :    0 - 0x0
    "00000000", --  691 - 0x2b3  :    0 - 0x0
    "00000000", --  692 - 0x2b4  :    0 - 0x0
    "00000000", --  693 - 0x2b5  :    0 - 0x0
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "00000000", --  696 - 0x2b8  :    0 - 0x0
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000000", --  704 - 0x2c0  :    0 - 0x0
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "00000000", --  707 - 0x2c3  :    0 - 0x0
    "00000000", --  708 - 0x2c4  :    0 - 0x0
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000000", --  752 - 0x2f0  :    0 - 0x0
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00000000", --  754 - 0x2f2  :    0 - 0x0
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "00000000", --  756 - 0x2f4  :    0 - 0x0
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "00000000", --  764 - 0x2fc  :    0 - 0x0
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00000000", --  770 - 0x302  :    0 - 0x0
    "00000000", --  771 - 0x303  :    0 - 0x0
    "00000000", --  772 - 0x304  :    0 - 0x0
    "00000000", --  773 - 0x305  :    0 - 0x0
    "00000000", --  774 - 0x306  :    0 - 0x0
    "00000000", --  775 - 0x307  :    0 - 0x0
    "00000000", --  776 - 0x308  :    0 - 0x0
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000000", --  779 - 0x30b  :    0 - 0x0
    "00000000", --  780 - 0x30c  :    0 - 0x0
    "00000000", --  781 - 0x30d  :    0 - 0x0
    "00000000", --  782 - 0x30e  :    0 - 0x0
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00000000", --  784 - 0x310  :    0 - 0x0
    "00000000", --  785 - 0x311  :    0 - 0x0
    "00000000", --  786 - 0x312  :    0 - 0x0
    "00000000", --  787 - 0x313  :    0 - 0x0
    "00000000", --  788 - 0x314  :    0 - 0x0
    "00000000", --  789 - 0x315  :    0 - 0x0
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "00000000", --  804 - 0x324  :    0 - 0x0
    "00000000", --  805 - 0x325  :    0 - 0x0
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "00000000", --  813 - 0x32d  :    0 - 0x0
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00000000", --  816 - 0x330  :    0 - 0x0
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000000", --  818 - 0x332  :    0 - 0x0
    "00000000", --  819 - 0x333  :    0 - 0x0
    "00000000", --  820 - 0x334  :    0 - 0x0
    "00000000", --  821 - 0x335  :    0 - 0x0
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000000", --  824 - 0x338  :    0 - 0x0
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "00000000", --  868 - 0x364  :    0 - 0x0
    "00000000", --  869 - 0x365  :    0 - 0x0
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00000000", --  888 - 0x378  :    0 - 0x0
    "00000000", --  889 - 0x379  :    0 - 0x0
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000000", -- 1024 - 0x400  :    0 - 0x0
    "00000000", -- 1025 - 0x401  :    0 - 0x0
    "00000000", -- 1026 - 0x402  :    0 - 0x0
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00000000", -- 1029 - 0x405  :    0 - 0x0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00000000", -- 1032 - 0x408  :    0 - 0x0
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "00000000", -- 1045 - 0x415  :    0 - 0x0
    "00000000", -- 1046 - 0x416  :    0 - 0x0
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0
    "00000000", -- 1057 - 0x421  :    0 - 0x0
    "00000000", -- 1058 - 0x422  :    0 - 0x0
    "00000000", -- 1059 - 0x423  :    0 - 0x0
    "00000000", -- 1060 - 0x424  :    0 - 0x0
    "00000000", -- 1061 - 0x425  :    0 - 0x0
    "00000000", -- 1062 - 0x426  :    0 - 0x0
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0
    "00000000", -- 1089 - 0x441  :    0 - 0x0
    "00000000", -- 1090 - 0x442  :    0 - 0x0
    "00000000", -- 1091 - 0x443  :    0 - 0x0
    "00000000", -- 1092 - 0x444  :    0 - 0x0
    "00000000", -- 1093 - 0x445  :    0 - 0x0
    "00000000", -- 1094 - 0x446  :    0 - 0x0
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00000000", -- 1096 - 0x448  :    0 - 0x0
    "00000000", -- 1097 - 0x449  :    0 - 0x0
    "00000000", -- 1098 - 0x44a  :    0 - 0x0
    "00000000", -- 1099 - 0x44b  :    0 - 0x0
    "00000000", -- 1100 - 0x44c  :    0 - 0x0
    "00000000", -- 1101 - 0x44d  :    0 - 0x0
    "00000000", -- 1102 - 0x44e  :    0 - 0x0
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0
    "00000000", -- 1105 - 0x451  :    0 - 0x0
    "00000000", -- 1106 - 0x452  :    0 - 0x0
    "00000000", -- 1107 - 0x453  :    0 - 0x0
    "00000000", -- 1108 - 0x454  :    0 - 0x0
    "00000000", -- 1109 - 0x455  :    0 - 0x0
    "00000000", -- 1110 - 0x456  :    0 - 0x0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00000000", -- 1112 - 0x458  :    0 - 0x0
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "00000000", -- 1114 - 0x45a  :    0 - 0x0
    "00000000", -- 1115 - 0x45b  :    0 - 0x0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00000000", -- 1117 - 0x45d  :    0 - 0x0
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000000", -- 1120 - 0x460  :    0 - 0x0
    "00000000", -- 1121 - 0x461  :    0 - 0x0
    "00000000", -- 1122 - 0x462  :    0 - 0x0
    "00000000", -- 1123 - 0x463  :    0 - 0x0
    "00000000", -- 1124 - 0x464  :    0 - 0x0
    "00000000", -- 1125 - 0x465  :    0 - 0x0
    "00000000", -- 1126 - 0x466  :    0 - 0x0
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000000", -- 1128 - 0x468  :    0 - 0x0
    "00000000", -- 1129 - 0x469  :    0 - 0x0
    "00000000", -- 1130 - 0x46a  :    0 - 0x0
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0
    "00000000", -- 1137 - 0x471  :    0 - 0x0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "00000000", -- 1140 - 0x474  :    0 - 0x0
    "00000000", -- 1141 - 0x475  :    0 - 0x0
    "00000000", -- 1142 - 0x476  :    0 - 0x0
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000000", -- 1144 - 0x478  :    0 - 0x0
    "00000000", -- 1145 - 0x479  :    0 - 0x0
    "00000000", -- 1146 - 0x47a  :    0 - 0x0
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00000000", -- 1156 - 0x484  :    0 - 0x0
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "00000000", -- 1158 - 0x486  :    0 - 0x0
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0
    "00000000", -- 1169 - 0x491  :    0 - 0x0
    "00000000", -- 1170 - 0x492  :    0 - 0x0
    "00000000", -- 1171 - 0x493  :    0 - 0x0
    "00000000", -- 1172 - 0x494  :    0 - 0x0
    "00000000", -- 1173 - 0x495  :    0 - 0x0
    "00000000", -- 1174 - 0x496  :    0 - 0x0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "00000000", -- 1176 - 0x498  :    0 - 0x0
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000000", -- 1186 - 0x4a2  :    0 - 0x0
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00000000", -- 1188 - 0x4a4  :    0 - 0x0
    "00000000", -- 1189 - 0x4a5  :    0 - 0x0
    "00000000", -- 1190 - 0x4a6  :    0 - 0x0
    "00000000", -- 1191 - 0x4a7  :    0 - 0x0
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00000000", -- 1194 - 0x4aa  :    0 - 0x0
    "00000000", -- 1195 - 0x4ab  :    0 - 0x0
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0
    "00000000", -- 1201 - 0x4b1  :    0 - 0x0
    "00000000", -- 1202 - 0x4b2  :    0 - 0x0
    "00000000", -- 1203 - 0x4b3  :    0 - 0x0
    "00000000", -- 1204 - 0x4b4  :    0 - 0x0
    "00000000", -- 1205 - 0x4b5  :    0 - 0x0
    "00000000", -- 1206 - 0x4b6  :    0 - 0x0
    "00000000", -- 1207 - 0x4b7  :    0 - 0x0
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0
    "00000000", -- 1217 - 0x4c1  :    0 - 0x0
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000000", -- 1219 - 0x4c3  :    0 - 0x0
    "00000000", -- 1220 - 0x4c4  :    0 - 0x0
    "00000000", -- 1221 - 0x4c5  :    0 - 0x0
    "00000000", -- 1222 - 0x4c6  :    0 - 0x0
    "00000000", -- 1223 - 0x4c7  :    0 - 0x0
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "00000000", -- 1228 - 0x4cc  :    0 - 0x0
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00000000", -- 1235 - 0x4d3  :    0 - 0x0
    "00000000", -- 1236 - 0x4d4  :    0 - 0x0
    "00000000", -- 1237 - 0x4d5  :    0 - 0x0
    "00000000", -- 1238 - 0x4d6  :    0 - 0x0
    "00000000", -- 1239 - 0x4d7  :    0 - 0x0
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0
    "00000000", -- 1249 - 0x4e1  :    0 - 0x0
    "00000000", -- 1250 - 0x4e2  :    0 - 0x0
    "00000000", -- 1251 - 0x4e3  :    0 - 0x0
    "00000000", -- 1252 - 0x4e4  :    0 - 0x0
    "00000000", -- 1253 - 0x4e5  :    0 - 0x0
    "00000000", -- 1254 - 0x4e6  :    0 - 0x0
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0
    "00000000", -- 1257 - 0x4e9  :    0 - 0x0
    "00000000", -- 1258 - 0x4ea  :    0 - 0x0
    "00000000", -- 1259 - 0x4eb  :    0 - 0x0
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00000000", -- 1261 - 0x4ed  :    0 - 0x0
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0
    "00000000", -- 1265 - 0x4f1  :    0 - 0x0
    "00000000", -- 1266 - 0x4f2  :    0 - 0x0
    "00000000", -- 1267 - 0x4f3  :    0 - 0x0
    "00000000", -- 1268 - 0x4f4  :    0 - 0x0
    "00000000", -- 1269 - 0x4f5  :    0 - 0x0
    "00000000", -- 1270 - 0x4f6  :    0 - 0x0
    "00000000", -- 1271 - 0x4f7  :    0 - 0x0
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0
    "00000000", -- 1281 - 0x501  :    0 - 0x0
    "00000000", -- 1282 - 0x502  :    0 - 0x0
    "00000000", -- 1283 - 0x503  :    0 - 0x0
    "00000000", -- 1284 - 0x504  :    0 - 0x0
    "00000000", -- 1285 - 0x505  :    0 - 0x0
    "00000000", -- 1286 - 0x506  :    0 - 0x0
    "00000000", -- 1287 - 0x507  :    0 - 0x0
    "00000000", -- 1288 - 0x508  :    0 - 0x0
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00000000", -- 1290 - 0x50a  :    0 - 0x0
    "00000000", -- 1291 - 0x50b  :    0 - 0x0
    "00000000", -- 1292 - 0x50c  :    0 - 0x0
    "00000000", -- 1293 - 0x50d  :    0 - 0x0
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00000000", -- 1296 - 0x510  :    0 - 0x0
    "00000000", -- 1297 - 0x511  :    0 - 0x0
    "00000000", -- 1298 - 0x512  :    0 - 0x0
    "00000000", -- 1299 - 0x513  :    0 - 0x0
    "00000000", -- 1300 - 0x514  :    0 - 0x0
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "00000000", -- 1302 - 0x516  :    0 - 0x0
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "00000000", -- 1304 - 0x518  :    0 - 0x0
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "00000000", -- 1306 - 0x51a  :    0 - 0x0
    "00000000", -- 1307 - 0x51b  :    0 - 0x0
    "00000000", -- 1308 - 0x51c  :    0 - 0x0
    "00000000", -- 1309 - 0x51d  :    0 - 0x0
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00000000", -- 1312 - 0x520  :    0 - 0x0
    "00000000", -- 1313 - 0x521  :    0 - 0x0
    "00000000", -- 1314 - 0x522  :    0 - 0x0
    "00000000", -- 1315 - 0x523  :    0 - 0x0
    "00000000", -- 1316 - 0x524  :    0 - 0x0
    "00000000", -- 1317 - 0x525  :    0 - 0x0
    "00000000", -- 1318 - 0x526  :    0 - 0x0
    "00000000", -- 1319 - 0x527  :    0 - 0x0
    "00000000", -- 1320 - 0x528  :    0 - 0x0
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "00000000", -- 1324 - 0x52c  :    0 - 0x0
    "00000000", -- 1325 - 0x52d  :    0 - 0x0
    "00000000", -- 1326 - 0x52e  :    0 - 0x0
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00000000", -- 1328 - 0x530  :    0 - 0x0
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "00000000", -- 1331 - 0x533  :    0 - 0x0
    "00000000", -- 1332 - 0x534  :    0 - 0x0
    "00000000", -- 1333 - 0x535  :    0 - 0x0
    "00000000", -- 1334 - 0x536  :    0 - 0x0
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "00000000", -- 1336 - 0x538  :    0 - 0x0
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "00000000", -- 1338 - 0x53a  :    0 - 0x0
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00000000", -- 1344 - 0x540  :    0 - 0x0
    "00000000", -- 1345 - 0x541  :    0 - 0x0
    "00000000", -- 1346 - 0x542  :    0 - 0x0
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00000000", -- 1349 - 0x545  :    0 - 0x0
    "00000000", -- 1350 - 0x546  :    0 - 0x0
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "00000000", -- 1352 - 0x548  :    0 - 0x0
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "00000000", -- 1354 - 0x54a  :    0 - 0x0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "00000000", -- 1357 - 0x54d  :    0 - 0x0
    "00000000", -- 1358 - 0x54e  :    0 - 0x0
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "00000000", -- 1380 - 0x564  :    0 - 0x0
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "00000000", -- 1386 - 0x56a  :    0 - 0x0
    "00000000", -- 1387 - 0x56b  :    0 - 0x0
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000000", -- 1396 - 0x574  :    0 - 0x0
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "00000000", -- 1408 - 0x580  :    0 - 0x0
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "00000000", -- 1410 - 0x582  :    0 - 0x0
    "00000000", -- 1411 - 0x583  :    0 - 0x0
    "00000000", -- 1412 - 0x584  :    0 - 0x0
    "00000000", -- 1413 - 0x585  :    0 - 0x0
    "00000000", -- 1414 - 0x586  :    0 - 0x0
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00000000", -- 1416 - 0x588  :    0 - 0x0
    "00000000", -- 1417 - 0x589  :    0 - 0x0
    "00000000", -- 1418 - 0x58a  :    0 - 0x0
    "00000000", -- 1419 - 0x58b  :    0 - 0x0
    "00000000", -- 1420 - 0x58c  :    0 - 0x0
    "00000000", -- 1421 - 0x58d  :    0 - 0x0
    "00000000", -- 1422 - 0x58e  :    0 - 0x0
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "00000000", -- 1424 - 0x590  :    0 - 0x0
    "00000000", -- 1425 - 0x591  :    0 - 0x0
    "00000000", -- 1426 - 0x592  :    0 - 0x0
    "00000000", -- 1427 - 0x593  :    0 - 0x0
    "00000000", -- 1428 - 0x594  :    0 - 0x0
    "00000000", -- 1429 - 0x595  :    0 - 0x0
    "00000000", -- 1430 - 0x596  :    0 - 0x0
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00000000", -- 1432 - 0x598  :    0 - 0x0
    "00000000", -- 1433 - 0x599  :    0 - 0x0
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00000000", -- 1435 - 0x59b  :    0 - 0x0
    "00000000", -- 1436 - 0x59c  :    0 - 0x0
    "00000000", -- 1437 - 0x59d  :    0 - 0x0
    "00000000", -- 1438 - 0x59e  :    0 - 0x0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "00000000", -- 1442 - 0x5a2  :    0 - 0x0
    "00000000", -- 1443 - 0x5a3  :    0 - 0x0
    "00000000", -- 1444 - 0x5a4  :    0 - 0x0
    "00000000", -- 1445 - 0x5a5  :    0 - 0x0
    "00000000", -- 1446 - 0x5a6  :    0 - 0x0
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "00000000", -- 1450 - 0x5aa  :    0 - 0x0
    "00000000", -- 1451 - 0x5ab  :    0 - 0x0
    "00000000", -- 1452 - 0x5ac  :    0 - 0x0
    "00000000", -- 1453 - 0x5ad  :    0 - 0x0
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00000000", -- 1461 - 0x5b5  :    0 - 0x0
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "00000000", -- 1466 - 0x5ba  :    0 - 0x0
    "00000000", -- 1467 - 0x5bb  :    0 - 0x0
    "00000000", -- 1468 - 0x5bc  :    0 - 0x0
    "00000000", -- 1469 - 0x5bd  :    0 - 0x0
    "00000000", -- 1470 - 0x5be  :    0 - 0x0
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0
    "00000000", -- 1473 - 0x5c1  :    0 - 0x0
    "00000000", -- 1474 - 0x5c2  :    0 - 0x0
    "00000000", -- 1475 - 0x5c3  :    0 - 0x0
    "00000000", -- 1476 - 0x5c4  :    0 - 0x0
    "00000000", -- 1477 - 0x5c5  :    0 - 0x0
    "00000000", -- 1478 - 0x5c6  :    0 - 0x0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "00000000", -- 1482 - 0x5ca  :    0 - 0x0
    "00000000", -- 1483 - 0x5cb  :    0 - 0x0
    "00000000", -- 1484 - 0x5cc  :    0 - 0x0
    "00000000", -- 1485 - 0x5cd  :    0 - 0x0
    "00000000", -- 1486 - 0x5ce  :    0 - 0x0
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0
    "00000000", -- 1489 - 0x5d1  :    0 - 0x0
    "00000000", -- 1490 - 0x5d2  :    0 - 0x0
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "00000000", -- 1492 - 0x5d4  :    0 - 0x0
    "00000000", -- 1493 - 0x5d5  :    0 - 0x0
    "00000000", -- 1494 - 0x5d6  :    0 - 0x0
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0
    "00000000", -- 1505 - 0x5e1  :    0 - 0x0
    "00000000", -- 1506 - 0x5e2  :    0 - 0x0
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "00000000", -- 1508 - 0x5e4  :    0 - 0x0
    "00000000", -- 1509 - 0x5e5  :    0 - 0x0
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00000000", -- 1514 - 0x5ea  :    0 - 0x0
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "00000000", -- 1516 - 0x5ec  :    0 - 0x0
    "00000000", -- 1517 - 0x5ed  :    0 - 0x0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000000", -- 1542 - 0x606  :    0 - 0x0
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00000000", -- 1544 - 0x608  :    0 - 0x0
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000000", -- 1578 - 0x62a  :    0 - 0x0
    "00000000", -- 1579 - 0x62b  :    0 - 0x0
    "00000000", -- 1580 - 0x62c  :    0 - 0x0
    "00000000", -- 1581 - 0x62d  :    0 - 0x0
    "00000000", -- 1582 - 0x62e  :    0 - 0x0
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "00000000", -- 1584 - 0x630  :    0 - 0x0
    "00000000", -- 1585 - 0x631  :    0 - 0x0
    "00000000", -- 1586 - 0x632  :    0 - 0x0
    "00000000", -- 1587 - 0x633  :    0 - 0x0
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "00000000", -- 1589 - 0x635  :    0 - 0x0
    "00000000", -- 1590 - 0x636  :    0 - 0x0
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00000000", -- 1592 - 0x638  :    0 - 0x0
    "00000000", -- 1593 - 0x639  :    0 - 0x0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "00000000", -- 1596 - 0x63c  :    0 - 0x0
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00000000", -- 1608 - 0x648  :    0 - 0x0
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "00000000", -- 1622 - 0x656  :    0 - 0x0
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00000000", -- 1680 - 0x690  :    0 - 0x0
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00000000", -- 1685 - 0x695  :    0 - 0x0
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00000000", -- 1688 - 0x698  :    0 - 0x0
    "00000000", -- 1689 - 0x699  :    0 - 0x0
    "00000000", -- 1690 - 0x69a  :    0 - 0x0
    "00000000", -- 1691 - 0x69b  :    0 - 0x0
    "00000000", -- 1692 - 0x69c  :    0 - 0x0
    "00000000", -- 1693 - 0x69d  :    0 - 0x0
    "00000000", -- 1694 - 0x69e  :    0 - 0x0
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0
    "00000000", -- 1705 - 0x6a9  :    0 - 0x0
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "00000000", -- 1715 - 0x6b3  :    0 - 0x0
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "00000000", -- 1720 - 0x6b8  :    0 - 0x0
    "00000000", -- 1721 - 0x6b9  :    0 - 0x0
    "00000000", -- 1722 - 0x6ba  :    0 - 0x0
    "00000000", -- 1723 - 0x6bb  :    0 - 0x0
    "00000000", -- 1724 - 0x6bc  :    0 - 0x0
    "00000000", -- 1725 - 0x6bd  :    0 - 0x0
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000000", -- 1734 - 0x6c6  :    0 - 0x0
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "00000000", -- 1738 - 0x6ca  :    0 - 0x0
    "00000000", -- 1739 - 0x6cb  :    0 - 0x0
    "00000000", -- 1740 - 0x6cc  :    0 - 0x0
    "00000000", -- 1741 - 0x6cd  :    0 - 0x0
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0
    "00000000", -- 1753 - 0x6d9  :    0 - 0x0
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "00000000", -- 1755 - 0x6db  :    0 - 0x0
    "00000000", -- 1756 - 0x6dc  :    0 - 0x0
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00000000", -- 1773 - 0x6ed  :    0 - 0x0
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0
    "00000000", -- 1777 - 0x6f1  :    0 - 0x0
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00000000", -- 1779 - 0x6f3  :    0 - 0x0
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "00000000", -- 1781 - 0x6f5  :    0 - 0x0
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "00000000", -- 1784 - 0x6f8  :    0 - 0x0
    "00000000", -- 1785 - 0x6f9  :    0 - 0x0
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "00000000", -- 1787 - 0x6fb  :    0 - 0x0
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "00000000", -- 1789 - 0x6fd  :    0 - 0x0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00000000", -- 1792 - 0x700  :    0 - 0x0
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000000", -- 1816 - 0x718  :    0 - 0x0
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000000", -- 1828 - 0x724  :    0 - 0x0
    "00000000", -- 1829 - 0x725  :    0 - 0x0
    "00000000", -- 1830 - 0x726  :    0 - 0x0
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "00000000", -- 1840 - 0x730  :    0 - 0x0
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "00000000", -- 1845 - 0x735  :    0 - 0x0
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000", -- 2047 - 0x7ff  :    0 - 0x0
    "00111110", -- 2048 - 0x800  :   62 - 0x3e
    "01111111", -- 2049 - 0x801  :  127 - 0x7f
    "01110111", -- 2050 - 0x802  :  119 - 0x77
    "01111111", -- 2051 - 0x803  :  127 - 0x7f
    "01111111", -- 2052 - 0x804  :  127 - 0x7f
    "01110111", -- 2053 - 0x805  :  119 - 0x77
    "01111111", -- 2054 - 0x806  :  127 - 0x7f
    "00111110", -- 2055 - 0x807  :   62 - 0x3e
    "00011100", -- 2056 - 0x808  :   28 - 0x1c
    "00111100", -- 2057 - 0x809  :   60 - 0x3c
    "01111100", -- 2058 - 0x80a  :  124 - 0x7c
    "00011100", -- 2059 - 0x80b  :   28 - 0x1c
    "00011100", -- 2060 - 0x80c  :   28 - 0x1c
    "00011100", -- 2061 - 0x80d  :   28 - 0x1c
    "01111111", -- 2062 - 0x80e  :  127 - 0x7f
    "01111111", -- 2063 - 0x80f  :  127 - 0x7f
    "00111110", -- 2064 - 0x810  :   62 - 0x3e
    "01111111", -- 2065 - 0x811  :  127 - 0x7f
    "00000111", -- 2066 - 0x812  :    7 - 0x7
    "00111111", -- 2067 - 0x813  :   63 - 0x3f
    "01111111", -- 2068 - 0x814  :  127 - 0x7f
    "01110000", -- 2069 - 0x815  :  112 - 0x70
    "01111111", -- 2070 - 0x816  :  127 - 0x7f
    "01111111", -- 2071 - 0x817  :  127 - 0x7f
    "00111110", -- 2072 - 0x818  :   62 - 0x3e
    "01111111", -- 2073 - 0x819  :  127 - 0x7f
    "00000111", -- 2074 - 0x81a  :    7 - 0x7
    "00011111", -- 2075 - 0x81b  :   31 - 0x1f
    "00011111", -- 2076 - 0x81c  :   31 - 0x1f
    "00000111", -- 2077 - 0x81d  :    7 - 0x7
    "01111111", -- 2078 - 0x81e  :  127 - 0x7f
    "00111110", -- 2079 - 0x81f  :   62 - 0x3e
    "00110000", -- 2080 - 0x820  :   48 - 0x30
    "01110000", -- 2081 - 0x821  :  112 - 0x70
    "01110111", -- 2082 - 0x822  :  119 - 0x77
    "01110111", -- 2083 - 0x823  :  119 - 0x77
    "01111111", -- 2084 - 0x824  :  127 - 0x7f
    "01111111", -- 2085 - 0x825  :  127 - 0x7f
    "00000111", -- 2086 - 0x826  :    7 - 0x7
    "00000111", -- 2087 - 0x827  :    7 - 0x7
    "01111111", -- 2088 - 0x828  :  127 - 0x7f
    "01111111", -- 2089 - 0x829  :  127 - 0x7f
    "01110000", -- 2090 - 0x82a  :  112 - 0x70
    "01111110", -- 2091 - 0x82b  :  126 - 0x7e
    "01111111", -- 2092 - 0x82c  :  127 - 0x7f
    "00000111", -- 2093 - 0x82d  :    7 - 0x7
    "01111111", -- 2094 - 0x82e  :  127 - 0x7f
    "00111110", -- 2095 - 0x82f  :   62 - 0x3e
    "00111110", -- 2096 - 0x830  :   62 - 0x3e
    "01111111", -- 2097 - 0x831  :  127 - 0x7f
    "01110000", -- 2098 - 0x832  :  112 - 0x70
    "01111110", -- 2099 - 0x833  :  126 - 0x7e
    "01111111", -- 2100 - 0x834  :  127 - 0x7f
    "01110111", -- 2101 - 0x835  :  119 - 0x77
    "01111111", -- 2102 - 0x836  :  127 - 0x7f
    "00111110", -- 2103 - 0x837  :   62 - 0x3e
    "01111111", -- 2104 - 0x838  :  127 - 0x7f
    "01111111", -- 2105 - 0x839  :  127 - 0x7f
    "00000111", -- 2106 - 0x83a  :    7 - 0x7
    "00001110", -- 2107 - 0x83b  :   14 - 0xe
    "00001110", -- 2108 - 0x83c  :   14 - 0xe
    "00011100", -- 2109 - 0x83d  :   28 - 0x1c
    "00011100", -- 2110 - 0x83e  :   28 - 0x1c
    "00011100", -- 2111 - 0x83f  :   28 - 0x1c
    "00111110", -- 2112 - 0x840  :   62 - 0x3e
    "01111111", -- 2113 - 0x841  :  127 - 0x7f
    "01110111", -- 2114 - 0x842  :  119 - 0x77
    "00111110", -- 2115 - 0x843  :   62 - 0x3e
    "01111111", -- 2116 - 0x844  :  127 - 0x7f
    "01110111", -- 2117 - 0x845  :  119 - 0x77
    "01111111", -- 2118 - 0x846  :  127 - 0x7f
    "00111110", -- 2119 - 0x847  :   62 - 0x3e
    "00111110", -- 2120 - 0x848  :   62 - 0x3e
    "01111111", -- 2121 - 0x849  :  127 - 0x7f
    "01110111", -- 2122 - 0x84a  :  119 - 0x77
    "01111111", -- 2123 - 0x84b  :  127 - 0x7f
    "00111111", -- 2124 - 0x84c  :   63 - 0x3f
    "00000111", -- 2125 - 0x84d  :    7 - 0x7
    "01111111", -- 2126 - 0x84e  :  127 - 0x7f
    "00111110", -- 2127 - 0x84f  :   62 - 0x3e
    "00000000", -- 2128 - 0x850  :    0 - 0x0
    "00000000", -- 2129 - 0x851  :    0 - 0x0
    "00000000", -- 2130 - 0x852  :    0 - 0x0
    "00000000", -- 2131 - 0x853  :    0 - 0x0
    "00000000", -- 2132 - 0x854  :    0 - 0x0
    "00110000", -- 2133 - 0x855  :   48 - 0x30
    "01111000", -- 2134 - 0x856  :  120 - 0x78
    "00110000", -- 2135 - 0x857  :   48 - 0x30
    "01110000", -- 2136 - 0x858  :  112 - 0x70
    "11111000", -- 2137 - 0x859  :  248 - 0xf8
    "11111000", -- 2138 - 0x85a  :  248 - 0xf8
    "11111000", -- 2139 - 0x85b  :  248 - 0xf8
    "01110000", -- 2140 - 0x85c  :  112 - 0x70
    "00000000", -- 2141 - 0x85d  :    0 - 0x0
    "01110000", -- 2142 - 0x85e  :  112 - 0x70
    "01110000", -- 2143 - 0x85f  :  112 - 0x70
    "01111000", -- 2144 - 0x860  :  120 - 0x78
    "11111100", -- 2145 - 0x861  :  252 - 0xfc
    "00011100", -- 2146 - 0x862  :   28 - 0x1c
    "00111000", -- 2147 - 0x863  :   56 - 0x38
    "00110000", -- 2148 - 0x864  :   48 - 0x30
    "00000000", -- 2149 - 0x865  :    0 - 0x0
    "01110000", -- 2150 - 0x866  :  112 - 0x70
    "01110000", -- 2151 - 0x867  :  112 - 0x70
    "00111100", -- 2152 - 0x868  :   60 - 0x3c
    "01111110", -- 2153 - 0x869  :  126 - 0x7e
    "11011011", -- 2154 - 0x86a  :  219 - 0xdb
    "11011111", -- 2155 - 0x86b  :  223 - 0xdf
    "11000011", -- 2156 - 0x86c  :  195 - 0xc3
    "01100110", -- 2157 - 0x86d  :  102 - 0x66
    "00111100", -- 2158 - 0x86e  :   60 - 0x3c
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "00000000", -- 2160 - 0x870  :    0 - 0x0
    "00000000", -- 2161 - 0x871  :    0 - 0x0
    "00000000", -- 2162 - 0x872  :    0 - 0x0
    "00111100", -- 2163 - 0x873  :   60 - 0x3c
    "00111110", -- 2164 - 0x874  :   62 - 0x3e
    "00011110", -- 2165 - 0x875  :   30 - 0x1e
    "00000000", -- 2166 - 0x876  :    0 - 0x0
    "00000000", -- 2167 - 0x877  :    0 - 0x0
    "11111111", -- 2168 - 0x878  :  255 - 0xff
    "11111111", -- 2169 - 0x879  :  255 - 0xff
    "11111111", -- 2170 - 0x87a  :  255 - 0xff
    "11111111", -- 2171 - 0x87b  :  255 - 0xff
    "11111111", -- 2172 - 0x87c  :  255 - 0xff
    "11111111", -- 2173 - 0x87d  :  255 - 0xff
    "11100000", -- 2174 - 0x87e  :  224 - 0xe0
    "11100000", -- 2175 - 0x87f  :  224 - 0xe0
    "00001110", -- 2176 - 0x880  :   14 - 0xe
    "00001110", -- 2177 - 0x881  :   14 - 0xe
    "00011100", -- 2178 - 0x882  :   28 - 0x1c
    "00011100", -- 2179 - 0x883  :   28 - 0x1c
    "00011100", -- 2180 - 0x884  :   28 - 0x1c
    "00011100", -- 2181 - 0x885  :   28 - 0x1c
    "00111000", -- 2182 - 0x886  :   56 - 0x38
    "00111000", -- 2183 - 0x887  :   56 - 0x38
    "00011100", -- 2184 - 0x888  :   28 - 0x1c
    "00111110", -- 2185 - 0x889  :   62 - 0x3e
    "01110111", -- 2186 - 0x88a  :  119 - 0x77
    "01110111", -- 2187 - 0x88b  :  119 - 0x77
    "01111111", -- 2188 - 0x88c  :  127 - 0x7f
    "01111111", -- 2189 - 0x88d  :  127 - 0x7f
    "01110111", -- 2190 - 0x88e  :  119 - 0x77
    "01110111", -- 2191 - 0x88f  :  119 - 0x77
    "01111110", -- 2192 - 0x890  :  126 - 0x7e
    "01110111", -- 2193 - 0x891  :  119 - 0x77
    "01110111", -- 2194 - 0x892  :  119 - 0x77
    "01111110", -- 2195 - 0x893  :  126 - 0x7e
    "01111110", -- 2196 - 0x894  :  126 - 0x7e
    "01110111", -- 2197 - 0x895  :  119 - 0x77
    "01110111", -- 2198 - 0x896  :  119 - 0x77
    "01111110", -- 2199 - 0x897  :  126 - 0x7e
    "00111110", -- 2200 - 0x898  :   62 - 0x3e
    "01111111", -- 2201 - 0x899  :  127 - 0x7f
    "01110111", -- 2202 - 0x89a  :  119 - 0x77
    "01110000", -- 2203 - 0x89b  :  112 - 0x70
    "01110000", -- 2204 - 0x89c  :  112 - 0x70
    "01110111", -- 2205 - 0x89d  :  119 - 0x77
    "01111111", -- 2206 - 0x89e  :  127 - 0x7f
    "00111110", -- 2207 - 0x89f  :   62 - 0x3e
    "01111110", -- 2208 - 0x8a0  :  126 - 0x7e
    "01111111", -- 2209 - 0x8a1  :  127 - 0x7f
    "01110111", -- 2210 - 0x8a2  :  119 - 0x77
    "01110111", -- 2211 - 0x8a3  :  119 - 0x77
    "01110111", -- 2212 - 0x8a4  :  119 - 0x77
    "01110111", -- 2213 - 0x8a5  :  119 - 0x77
    "01111111", -- 2214 - 0x8a6  :  127 - 0x7f
    "01111110", -- 2215 - 0x8a7  :  126 - 0x7e
    "01111111", -- 2216 - 0x8a8  :  127 - 0x7f
    "01111111", -- 2217 - 0x8a9  :  127 - 0x7f
    "01110000", -- 2218 - 0x8aa  :  112 - 0x70
    "01111100", -- 2219 - 0x8ab  :  124 - 0x7c
    "01111100", -- 2220 - 0x8ac  :  124 - 0x7c
    "01110000", -- 2221 - 0x8ad  :  112 - 0x70
    "01111111", -- 2222 - 0x8ae  :  127 - 0x7f
    "01111111", -- 2223 - 0x8af  :  127 - 0x7f
    "01111111", -- 2224 - 0x8b0  :  127 - 0x7f
    "01111111", -- 2225 - 0x8b1  :  127 - 0x7f
    "01110000", -- 2226 - 0x8b2  :  112 - 0x70
    "01111100", -- 2227 - 0x8b3  :  124 - 0x7c
    "01111100", -- 2228 - 0x8b4  :  124 - 0x7c
    "01110000", -- 2229 - 0x8b5  :  112 - 0x70
    "01110000", -- 2230 - 0x8b6  :  112 - 0x70
    "01110000", -- 2231 - 0x8b7  :  112 - 0x70
    "00111110", -- 2232 - 0x8b8  :   62 - 0x3e
    "01111111", -- 2233 - 0x8b9  :  127 - 0x7f
    "01110111", -- 2234 - 0x8ba  :  119 - 0x77
    "01110000", -- 2235 - 0x8bb  :  112 - 0x70
    "01111111", -- 2236 - 0x8bc  :  127 - 0x7f
    "01110111", -- 2237 - 0x8bd  :  119 - 0x77
    "01111111", -- 2238 - 0x8be  :  127 - 0x7f
    "00111110", -- 2239 - 0x8bf  :   62 - 0x3e
    "01110111", -- 2240 - 0x8c0  :  119 - 0x77
    "01110111", -- 2241 - 0x8c1  :  119 - 0x77
    "01110111", -- 2242 - 0x8c2  :  119 - 0x77
    "01111111", -- 2243 - 0x8c3  :  127 - 0x7f
    "01111111", -- 2244 - 0x8c4  :  127 - 0x7f
    "01110111", -- 2245 - 0x8c5  :  119 - 0x77
    "01110111", -- 2246 - 0x8c6  :  119 - 0x77
    "01110111", -- 2247 - 0x8c7  :  119 - 0x77
    "00111110", -- 2248 - 0x8c8  :   62 - 0x3e
    "00111110", -- 2249 - 0x8c9  :   62 - 0x3e
    "00011100", -- 2250 - 0x8ca  :   28 - 0x1c
    "00011100", -- 2251 - 0x8cb  :   28 - 0x1c
    "00011100", -- 2252 - 0x8cc  :   28 - 0x1c
    "00011100", -- 2253 - 0x8cd  :   28 - 0x1c
    "00111110", -- 2254 - 0x8ce  :   62 - 0x3e
    "00111110", -- 2255 - 0x8cf  :   62 - 0x3e
    "00000111", -- 2256 - 0x8d0  :    7 - 0x7
    "00000111", -- 2257 - 0x8d1  :    7 - 0x7
    "00000111", -- 2258 - 0x8d2  :    7 - 0x7
    "00000111", -- 2259 - 0x8d3  :    7 - 0x7
    "00000111", -- 2260 - 0x8d4  :    7 - 0x7
    "01110111", -- 2261 - 0x8d5  :  119 - 0x77
    "01111111", -- 2262 - 0x8d6  :  127 - 0x7f
    "00111110", -- 2263 - 0x8d7  :   62 - 0x3e
    "01110011", -- 2264 - 0x8d8  :  115 - 0x73
    "01110111", -- 2265 - 0x8d9  :  119 - 0x77
    "01111110", -- 2266 - 0x8da  :  126 - 0x7e
    "01111100", -- 2267 - 0x8db  :  124 - 0x7c
    "01111110", -- 2268 - 0x8dc  :  126 - 0x7e
    "01110111", -- 2269 - 0x8dd  :  119 - 0x77
    "01110111", -- 2270 - 0x8de  :  119 - 0x77
    "01110111", -- 2271 - 0x8df  :  119 - 0x77
    "01110000", -- 2272 - 0x8e0  :  112 - 0x70
    "01110000", -- 2273 - 0x8e1  :  112 - 0x70
    "01110000", -- 2274 - 0x8e2  :  112 - 0x70
    "01110000", -- 2275 - 0x8e3  :  112 - 0x70
    "01110000", -- 2276 - 0x8e4  :  112 - 0x70
    "01110000", -- 2277 - 0x8e5  :  112 - 0x70
    "01111111", -- 2278 - 0x8e6  :  127 - 0x7f
    "01111111", -- 2279 - 0x8e7  :  127 - 0x7f
    "11100111", -- 2280 - 0x8e8  :  231 - 0xe7
    "11111111", -- 2281 - 0x8e9  :  255 - 0xff
    "11111111", -- 2282 - 0x8ea  :  255 - 0xff
    "11111111", -- 2283 - 0x8eb  :  255 - 0xff
    "11111111", -- 2284 - 0x8ec  :  255 - 0xff
    "11100111", -- 2285 - 0x8ed  :  231 - 0xe7
    "11100111", -- 2286 - 0x8ee  :  231 - 0xe7
    "11100111", -- 2287 - 0x8ef  :  231 - 0xe7
    "01110111", -- 2288 - 0x8f0  :  119 - 0x77
    "01110111", -- 2289 - 0x8f1  :  119 - 0x77
    "01111111", -- 2290 - 0x8f2  :  127 - 0x7f
    "01111111", -- 2291 - 0x8f3  :  127 - 0x7f
    "01111111", -- 2292 - 0x8f4  :  127 - 0x7f
    "01111111", -- 2293 - 0x8f5  :  127 - 0x7f
    "01110111", -- 2294 - 0x8f6  :  119 - 0x77
    "01110111", -- 2295 - 0x8f7  :  119 - 0x77
    "00111100", -- 2296 - 0x8f8  :   60 - 0x3c
    "01111110", -- 2297 - 0x8f9  :  126 - 0x7e
    "11100111", -- 2298 - 0x8fa  :  231 - 0xe7
    "11100111", -- 2299 - 0x8fb  :  231 - 0xe7
    "11100111", -- 2300 - 0x8fc  :  231 - 0xe7
    "11100111", -- 2301 - 0x8fd  :  231 - 0xe7
    "01111110", -- 2302 - 0x8fe  :  126 - 0x7e
    "00111100", -- 2303 - 0x8ff  :   60 - 0x3c
    "01111110", -- 2304 - 0x900  :  126 - 0x7e
    "01111111", -- 2305 - 0x901  :  127 - 0x7f
    "01110111", -- 2306 - 0x902  :  119 - 0x77
    "01110111", -- 2307 - 0x903  :  119 - 0x77
    "01111111", -- 2308 - 0x904  :  127 - 0x7f
    "01111110", -- 2309 - 0x905  :  126 - 0x7e
    "01110000", -- 2310 - 0x906  :  112 - 0x70
    "01110000", -- 2311 - 0x907  :  112 - 0x70
    "00111100", -- 2312 - 0x908  :   60 - 0x3c
    "01111110", -- 2313 - 0x909  :  126 - 0x7e
    "11100111", -- 2314 - 0x90a  :  231 - 0xe7
    "11100111", -- 2315 - 0x90b  :  231 - 0xe7
    "11100111", -- 2316 - 0x90c  :  231 - 0xe7
    "11101110", -- 2317 - 0x90d  :  238 - 0xee
    "01111111", -- 2318 - 0x90e  :  127 - 0x7f
    "00111111", -- 2319 - 0x90f  :   63 - 0x3f
    "01111110", -- 2320 - 0x910  :  126 - 0x7e
    "01111111", -- 2321 - 0x911  :  127 - 0x7f
    "01110111", -- 2322 - 0x912  :  119 - 0x77
    "01110111", -- 2323 - 0x913  :  119 - 0x77
    "01111111", -- 2324 - 0x914  :  127 - 0x7f
    "01111110", -- 2325 - 0x915  :  126 - 0x7e
    "01110111", -- 2326 - 0x916  :  119 - 0x77
    "01110111", -- 2327 - 0x917  :  119 - 0x77
    "00111110", -- 2328 - 0x918  :   62 - 0x3e
    "01111111", -- 2329 - 0x919  :  127 - 0x7f
    "01110000", -- 2330 - 0x91a  :  112 - 0x70
    "01111110", -- 2331 - 0x91b  :  126 - 0x7e
    "00111111", -- 2332 - 0x91c  :   63 - 0x3f
    "00000111", -- 2333 - 0x91d  :    7 - 0x7
    "01111111", -- 2334 - 0x91e  :  127 - 0x7f
    "00111110", -- 2335 - 0x91f  :   62 - 0x3e
    "01111111", -- 2336 - 0x920  :  127 - 0x7f
    "01111111", -- 2337 - 0x921  :  127 - 0x7f
    "00011100", -- 2338 - 0x922  :   28 - 0x1c
    "00011100", -- 2339 - 0x923  :   28 - 0x1c
    "00011100", -- 2340 - 0x924  :   28 - 0x1c
    "00011100", -- 2341 - 0x925  :   28 - 0x1c
    "00011100", -- 2342 - 0x926  :   28 - 0x1c
    "00011100", -- 2343 - 0x927  :   28 - 0x1c
    "01110111", -- 2344 - 0x928  :  119 - 0x77
    "01110111", -- 2345 - 0x929  :  119 - 0x77
    "01110111", -- 2346 - 0x92a  :  119 - 0x77
    "01110111", -- 2347 - 0x92b  :  119 - 0x77
    "01110111", -- 2348 - 0x92c  :  119 - 0x77
    "01110111", -- 2349 - 0x92d  :  119 - 0x77
    "01111111", -- 2350 - 0x92e  :  127 - 0x7f
    "00111110", -- 2351 - 0x92f  :   62 - 0x3e
    "01110111", -- 2352 - 0x930  :  119 - 0x77
    "01110111", -- 2353 - 0x931  :  119 - 0x77
    "01110111", -- 2354 - 0x932  :  119 - 0x77
    "01110111", -- 2355 - 0x933  :  119 - 0x77
    "01110111", -- 2356 - 0x934  :  119 - 0x77
    "01110111", -- 2357 - 0x935  :  119 - 0x77
    "00111110", -- 2358 - 0x936  :   62 - 0x3e
    "00011100", -- 2359 - 0x937  :   28 - 0x1c
    "11100111", -- 2360 - 0x938  :  231 - 0xe7
    "11100111", -- 2361 - 0x939  :  231 - 0xe7
    "11100111", -- 2362 - 0x93a  :  231 - 0xe7
    "11100111", -- 2363 - 0x93b  :  231 - 0xe7
    "11110111", -- 2364 - 0x93c  :  247 - 0xf7
    "11111111", -- 2365 - 0x93d  :  255 - 0xff
    "11111111", -- 2366 - 0x93e  :  255 - 0xff
    "01111110", -- 2367 - 0x93f  :  126 - 0x7e
    "01110111", -- 2368 - 0x940  :  119 - 0x77
    "01110111", -- 2369 - 0x941  :  119 - 0x77
    "01110111", -- 2370 - 0x942  :  119 - 0x77
    "00111110", -- 2371 - 0x943  :   62 - 0x3e
    "00111110", -- 2372 - 0x944  :   62 - 0x3e
    "01110111", -- 2373 - 0x945  :  119 - 0x77
    "01110111", -- 2374 - 0x946  :  119 - 0x77
    "01110111", -- 2375 - 0x947  :  119 - 0x77
    "01110111", -- 2376 - 0x948  :  119 - 0x77
    "01110111", -- 2377 - 0x949  :  119 - 0x77
    "01110111", -- 2378 - 0x94a  :  119 - 0x77
    "01111111", -- 2379 - 0x94b  :  127 - 0x7f
    "00111110", -- 2380 - 0x94c  :   62 - 0x3e
    "00011100", -- 2381 - 0x94d  :   28 - 0x1c
    "00011100", -- 2382 - 0x94e  :   28 - 0x1c
    "00011100", -- 2383 - 0x94f  :   28 - 0x1c
    "01111111", -- 2384 - 0x950  :  127 - 0x7f
    "01111111", -- 2385 - 0x951  :  127 - 0x7f
    "00001110", -- 2386 - 0x952  :   14 - 0xe
    "00011100", -- 2387 - 0x953  :   28 - 0x1c
    "00011100", -- 2388 - 0x954  :   28 - 0x1c
    "00111000", -- 2389 - 0x955  :   56 - 0x38
    "01111111", -- 2390 - 0x956  :  127 - 0x7f
    "01111111", -- 2391 - 0x957  :  127 - 0x7f
    "00111110", -- 2392 - 0x958  :   62 - 0x3e
    "01100011", -- 2393 - 0x959  :   99 - 0x63
    "01101111", -- 2394 - 0x95a  :  111 - 0x6f
    "01111111", -- 2395 - 0x95b  :  127 - 0x7f
    "01111111", -- 2396 - 0x95c  :  127 - 0x7f
    "01111110", -- 2397 - 0x95d  :  126 - 0x7e
    "01100000", -- 2398 - 0x95e  :   96 - 0x60
    "00111111", -- 2399 - 0x95f  :   63 - 0x3f
    "00000000", -- 2400 - 0x960  :    0 - 0x0
    "01110000", -- 2401 - 0x961  :  112 - 0x70
    "01111100", -- 2402 - 0x962  :  124 - 0x7c
    "01111111", -- 2403 - 0x963  :  127 - 0x7f
    "01111111", -- 2404 - 0x964  :  127 - 0x7f
    "01111100", -- 2405 - 0x965  :  124 - 0x7c
    "01110000", -- 2406 - 0x966  :  112 - 0x70
    "00000000", -- 2407 - 0x967  :    0 - 0x0
    "00000000", -- 2408 - 0x968  :    0 - 0x0
    "01110000", -- 2409 - 0x969  :  112 - 0x70
    "01110000", -- 2410 - 0x96a  :  112 - 0x70
    "00000000", -- 2411 - 0x96b  :    0 - 0x0
    "00000000", -- 2412 - 0x96c  :    0 - 0x0
    "01110000", -- 2413 - 0x96d  :  112 - 0x70
    "01110000", -- 2414 - 0x96e  :  112 - 0x70
    "00000000", -- 2415 - 0x96f  :    0 - 0x0
    "00000000", -- 2416 - 0x970  :    0 - 0x0
    "00000000", -- 2417 - 0x971  :    0 - 0x0
    "00000000", -- 2418 - 0x972  :    0 - 0x0
    "00000000", -- 2419 - 0x973  :    0 - 0x0
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "00000000", -- 2424 - 0x978  :    0 - 0x0
    "00000000", -- 2425 - 0x979  :    0 - 0x0
    "00000000", -- 2426 - 0x97a  :    0 - 0x0
    "00000000", -- 2427 - 0x97b  :    0 - 0x0
    "00000000", -- 2428 - 0x97c  :    0 - 0x0
    "00000000", -- 2429 - 0x97d  :    0 - 0x0
    "00000000", -- 2430 - 0x97e  :    0 - 0x0
    "00000000", -- 2431 - 0x97f  :    0 - 0x0
    "00000000", -- 2432 - 0x980  :    0 - 0x0
    "00000000", -- 2433 - 0x981  :    0 - 0x0
    "00000000", -- 2434 - 0x982  :    0 - 0x0
    "00000000", -- 2435 - 0x983  :    0 - 0x0
    "00000000", -- 2436 - 0x984  :    0 - 0x0
    "00000000", -- 2437 - 0x985  :    0 - 0x0
    "00000000", -- 2438 - 0x986  :    0 - 0x0
    "00000000", -- 2439 - 0x987  :    0 - 0x0
    "00000000", -- 2440 - 0x988  :    0 - 0x0
    "00000000", -- 2441 - 0x989  :    0 - 0x0
    "00000000", -- 2442 - 0x98a  :    0 - 0x0
    "00000000", -- 2443 - 0x98b  :    0 - 0x0
    "00000000", -- 2444 - 0x98c  :    0 - 0x0
    "00000000", -- 2445 - 0x98d  :    0 - 0x0
    "00000000", -- 2446 - 0x98e  :    0 - 0x0
    "00000000", -- 2447 - 0x98f  :    0 - 0x0
    "00000000", -- 2448 - 0x990  :    0 - 0x0
    "00000000", -- 2449 - 0x991  :    0 - 0x0
    "00000000", -- 2450 - 0x992  :    0 - 0x0
    "00000000", -- 2451 - 0x993  :    0 - 0x0
    "00000000", -- 2452 - 0x994  :    0 - 0x0
    "00000000", -- 2453 - 0x995  :    0 - 0x0
    "00000000", -- 2454 - 0x996  :    0 - 0x0
    "00000000", -- 2455 - 0x997  :    0 - 0x0
    "00000000", -- 2456 - 0x998  :    0 - 0x0
    "00000000", -- 2457 - 0x999  :    0 - 0x0
    "00000000", -- 2458 - 0x99a  :    0 - 0x0
    "00000000", -- 2459 - 0x99b  :    0 - 0x0
    "00000000", -- 2460 - 0x99c  :    0 - 0x0
    "00000000", -- 2461 - 0x99d  :    0 - 0x0
    "00000000", -- 2462 - 0x99e  :    0 - 0x0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "00000000", -- 2464 - 0x9a0  :    0 - 0x0
    "00000000", -- 2465 - 0x9a1  :    0 - 0x0
    "00000000", -- 2466 - 0x9a2  :    0 - 0x0
    "00000000", -- 2467 - 0x9a3  :    0 - 0x0
    "00000000", -- 2468 - 0x9a4  :    0 - 0x0
    "00000000", -- 2469 - 0x9a5  :    0 - 0x0
    "00000000", -- 2470 - 0x9a6  :    0 - 0x0
    "00000000", -- 2471 - 0x9a7  :    0 - 0x0
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "00000000", -- 2474 - 0x9aa  :    0 - 0x0
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00000000", -- 2476 - 0x9ac  :    0 - 0x0
    "00000000", -- 2477 - 0x9ad  :    0 - 0x0
    "00000000", -- 2478 - 0x9ae  :    0 - 0x0
    "00000000", -- 2479 - 0x9af  :    0 - 0x0
    "00000000", -- 2480 - 0x9b0  :    0 - 0x0
    "00000000", -- 2481 - 0x9b1  :    0 - 0x0
    "00000000", -- 2482 - 0x9b2  :    0 - 0x0
    "00000000", -- 2483 - 0x9b3  :    0 - 0x0
    "00000000", -- 2484 - 0x9b4  :    0 - 0x0
    "00000000", -- 2485 - 0x9b5  :    0 - 0x0
    "00000000", -- 2486 - 0x9b6  :    0 - 0x0
    "00000000", -- 2487 - 0x9b7  :    0 - 0x0
    "00000000", -- 2488 - 0x9b8  :    0 - 0x0
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "00000000", -- 2490 - 0x9ba  :    0 - 0x0
    "00000000", -- 2491 - 0x9bb  :    0 - 0x0
    "00000000", -- 2492 - 0x9bc  :    0 - 0x0
    "00000000", -- 2493 - 0x9bd  :    0 - 0x0
    "00000000", -- 2494 - 0x9be  :    0 - 0x0
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000000", -- 2498 - 0x9c2  :    0 - 0x0
    "00000000", -- 2499 - 0x9c3  :    0 - 0x0
    "00000000", -- 2500 - 0x9c4  :    0 - 0x0
    "00000000", -- 2501 - 0x9c5  :    0 - 0x0
    "00000000", -- 2502 - 0x9c6  :    0 - 0x0
    "00000000", -- 2503 - 0x9c7  :    0 - 0x0
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0
    "00000000", -- 2513 - 0x9d1  :    0 - 0x0
    "00000000", -- 2514 - 0x9d2  :    0 - 0x0
    "00000000", -- 2515 - 0x9d3  :    0 - 0x0
    "00000000", -- 2516 - 0x9d4  :    0 - 0x0
    "00000000", -- 2517 - 0x9d5  :    0 - 0x0
    "00000000", -- 2518 - 0x9d6  :    0 - 0x0
    "00000000", -- 2519 - 0x9d7  :    0 - 0x0
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0
    "00000000", -- 2521 - 0x9d9  :    0 - 0x0
    "00000000", -- 2522 - 0x9da  :    0 - 0x0
    "00000000", -- 2523 - 0x9db  :    0 - 0x0
    "00000000", -- 2524 - 0x9dc  :    0 - 0x0
    "00000000", -- 2525 - 0x9dd  :    0 - 0x0
    "00000000", -- 2526 - 0x9de  :    0 - 0x0
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0
    "00000000", -- 2529 - 0x9e1  :    0 - 0x0
    "00000000", -- 2530 - 0x9e2  :    0 - 0x0
    "00000000", -- 2531 - 0x9e3  :    0 - 0x0
    "00000000", -- 2532 - 0x9e4  :    0 - 0x0
    "00000000", -- 2533 - 0x9e5  :    0 - 0x0
    "00000000", -- 2534 - 0x9e6  :    0 - 0x0
    "00000000", -- 2535 - 0x9e7  :    0 - 0x0
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0
    "00000000", -- 2537 - 0x9e9  :    0 - 0x0
    "00000000", -- 2538 - 0x9ea  :    0 - 0x0
    "00000000", -- 2539 - 0x9eb  :    0 - 0x0
    "00000000", -- 2540 - 0x9ec  :    0 - 0x0
    "00000000", -- 2541 - 0x9ed  :    0 - 0x0
    "00000000", -- 2542 - 0x9ee  :    0 - 0x0
    "00000000", -- 2543 - 0x9ef  :    0 - 0x0
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0
    "00000000", -- 2545 - 0x9f1  :    0 - 0x0
    "00000000", -- 2546 - 0x9f2  :    0 - 0x0
    "00000000", -- 2547 - 0x9f3  :    0 - 0x0
    "00000000", -- 2548 - 0x9f4  :    0 - 0x0
    "00000000", -- 2549 - 0x9f5  :    0 - 0x0
    "00000000", -- 2550 - 0x9f6  :    0 - 0x0
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00000000", -- 2560 - 0xa00  :    0 - 0x0
    "00000000", -- 2561 - 0xa01  :    0 - 0x0
    "00000000", -- 2562 - 0xa02  :    0 - 0x0
    "00000000", -- 2563 - 0xa03  :    0 - 0x0
    "00000000", -- 2564 - 0xa04  :    0 - 0x0
    "00000000", -- 2565 - 0xa05  :    0 - 0x0
    "00000000", -- 2566 - 0xa06  :    0 - 0x0
    "00000000", -- 2567 - 0xa07  :    0 - 0x0
    "00000000", -- 2568 - 0xa08  :    0 - 0x0
    "00000000", -- 2569 - 0xa09  :    0 - 0x0
    "00000000", -- 2570 - 0xa0a  :    0 - 0x0
    "00000000", -- 2571 - 0xa0b  :    0 - 0x0
    "00000000", -- 2572 - 0xa0c  :    0 - 0x0
    "00000000", -- 2573 - 0xa0d  :    0 - 0x0
    "00000000", -- 2574 - 0xa0e  :    0 - 0x0
    "00000000", -- 2575 - 0xa0f  :    0 - 0x0
    "00000000", -- 2576 - 0xa10  :    0 - 0x0
    "00000000", -- 2577 - 0xa11  :    0 - 0x0
    "00000000", -- 2578 - 0xa12  :    0 - 0x0
    "00000000", -- 2579 - 0xa13  :    0 - 0x0
    "00000000", -- 2580 - 0xa14  :    0 - 0x0
    "00000000", -- 2581 - 0xa15  :    0 - 0x0
    "00000000", -- 2582 - 0xa16  :    0 - 0x0
    "00000000", -- 2583 - 0xa17  :    0 - 0x0
    "00000000", -- 2584 - 0xa18  :    0 - 0x0
    "00000000", -- 2585 - 0xa19  :    0 - 0x0
    "00000000", -- 2586 - 0xa1a  :    0 - 0x0
    "00000000", -- 2587 - 0xa1b  :    0 - 0x0
    "00000000", -- 2588 - 0xa1c  :    0 - 0x0
    "00000000", -- 2589 - 0xa1d  :    0 - 0x0
    "00000000", -- 2590 - 0xa1e  :    0 - 0x0
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "00000000", -- 2592 - 0xa20  :    0 - 0x0
    "00000000", -- 2593 - 0xa21  :    0 - 0x0
    "00000000", -- 2594 - 0xa22  :    0 - 0x0
    "00000000", -- 2595 - 0xa23  :    0 - 0x0
    "00000000", -- 2596 - 0xa24  :    0 - 0x0
    "00000000", -- 2597 - 0xa25  :    0 - 0x0
    "00000000", -- 2598 - 0xa26  :    0 - 0x0
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00000000", -- 2600 - 0xa28  :    0 - 0x0
    "00000000", -- 2601 - 0xa29  :    0 - 0x0
    "00000000", -- 2602 - 0xa2a  :    0 - 0x0
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "00000000", -- 2608 - 0xa30  :    0 - 0x0
    "00000000", -- 2609 - 0xa31  :    0 - 0x0
    "00000000", -- 2610 - 0xa32  :    0 - 0x0
    "00000000", -- 2611 - 0xa33  :    0 - 0x0
    "00000000", -- 2612 - 0xa34  :    0 - 0x0
    "00000000", -- 2613 - 0xa35  :    0 - 0x0
    "00000000", -- 2614 - 0xa36  :    0 - 0x0
    "00000000", -- 2615 - 0xa37  :    0 - 0x0
    "00000000", -- 2616 - 0xa38  :    0 - 0x0
    "00000000", -- 2617 - 0xa39  :    0 - 0x0
    "00000000", -- 2618 - 0xa3a  :    0 - 0x0
    "00000000", -- 2619 - 0xa3b  :    0 - 0x0
    "00000000", -- 2620 - 0xa3c  :    0 - 0x0
    "00000000", -- 2621 - 0xa3d  :    0 - 0x0
    "00000000", -- 2622 - 0xa3e  :    0 - 0x0
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "00000000", -- 2624 - 0xa40  :    0 - 0x0
    "00000000", -- 2625 - 0xa41  :    0 - 0x0
    "00000000", -- 2626 - 0xa42  :    0 - 0x0
    "00000000", -- 2627 - 0xa43  :    0 - 0x0
    "00000000", -- 2628 - 0xa44  :    0 - 0x0
    "00000000", -- 2629 - 0xa45  :    0 - 0x0
    "00000000", -- 2630 - 0xa46  :    0 - 0x0
    "00000000", -- 2631 - 0xa47  :    0 - 0x0
    "00000000", -- 2632 - 0xa48  :    0 - 0x0
    "00000000", -- 2633 - 0xa49  :    0 - 0x0
    "00000000", -- 2634 - 0xa4a  :    0 - 0x0
    "00000000", -- 2635 - 0xa4b  :    0 - 0x0
    "00000000", -- 2636 - 0xa4c  :    0 - 0x0
    "00000000", -- 2637 - 0xa4d  :    0 - 0x0
    "00000000", -- 2638 - 0xa4e  :    0 - 0x0
    "00000000", -- 2639 - 0xa4f  :    0 - 0x0
    "00000000", -- 2640 - 0xa50  :    0 - 0x0
    "00000000", -- 2641 - 0xa51  :    0 - 0x0
    "00000000", -- 2642 - 0xa52  :    0 - 0x0
    "00000000", -- 2643 - 0xa53  :    0 - 0x0
    "00000000", -- 2644 - 0xa54  :    0 - 0x0
    "00000000", -- 2645 - 0xa55  :    0 - 0x0
    "00000000", -- 2646 - 0xa56  :    0 - 0x0
    "00000000", -- 2647 - 0xa57  :    0 - 0x0
    "00000000", -- 2648 - 0xa58  :    0 - 0x0
    "00000000", -- 2649 - 0xa59  :    0 - 0x0
    "00000000", -- 2650 - 0xa5a  :    0 - 0x0
    "00000000", -- 2651 - 0xa5b  :    0 - 0x0
    "00000000", -- 2652 - 0xa5c  :    0 - 0x0
    "00000000", -- 2653 - 0xa5d  :    0 - 0x0
    "00000000", -- 2654 - 0xa5e  :    0 - 0x0
    "00000000", -- 2655 - 0xa5f  :    0 - 0x0
    "00000000", -- 2656 - 0xa60  :    0 - 0x0
    "00000000", -- 2657 - 0xa61  :    0 - 0x0
    "00000000", -- 2658 - 0xa62  :    0 - 0x0
    "00000000", -- 2659 - 0xa63  :    0 - 0x0
    "00000000", -- 2660 - 0xa64  :    0 - 0x0
    "00000000", -- 2661 - 0xa65  :    0 - 0x0
    "00000000", -- 2662 - 0xa66  :    0 - 0x0
    "00000000", -- 2663 - 0xa67  :    0 - 0x0
    "00000000", -- 2664 - 0xa68  :    0 - 0x0
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "00000000", -- 2666 - 0xa6a  :    0 - 0x0
    "00000000", -- 2667 - 0xa6b  :    0 - 0x0
    "00000000", -- 2668 - 0xa6c  :    0 - 0x0
    "00000000", -- 2669 - 0xa6d  :    0 - 0x0
    "00000000", -- 2670 - 0xa6e  :    0 - 0x0
    "00000000", -- 2671 - 0xa6f  :    0 - 0x0
    "00000000", -- 2672 - 0xa70  :    0 - 0x0
    "00000000", -- 2673 - 0xa71  :    0 - 0x0
    "00000000", -- 2674 - 0xa72  :    0 - 0x0
    "00000000", -- 2675 - 0xa73  :    0 - 0x0
    "00000000", -- 2676 - 0xa74  :    0 - 0x0
    "00000000", -- 2677 - 0xa75  :    0 - 0x0
    "00000000", -- 2678 - 0xa76  :    0 - 0x0
    "00000000", -- 2679 - 0xa77  :    0 - 0x0
    "00000000", -- 2680 - 0xa78  :    0 - 0x0
    "00000000", -- 2681 - 0xa79  :    0 - 0x0
    "00000000", -- 2682 - 0xa7a  :    0 - 0x0
    "00000000", -- 2683 - 0xa7b  :    0 - 0x0
    "00000000", -- 2684 - 0xa7c  :    0 - 0x0
    "00000000", -- 2685 - 0xa7d  :    0 - 0x0
    "00000000", -- 2686 - 0xa7e  :    0 - 0x0
    "00000000", -- 2687 - 0xa7f  :    0 - 0x0
    "00000000", -- 2688 - 0xa80  :    0 - 0x0
    "00000000", -- 2689 - 0xa81  :    0 - 0x0
    "00000000", -- 2690 - 0xa82  :    0 - 0x0
    "00000000", -- 2691 - 0xa83  :    0 - 0x0
    "00000000", -- 2692 - 0xa84  :    0 - 0x0
    "00000000", -- 2693 - 0xa85  :    0 - 0x0
    "00000000", -- 2694 - 0xa86  :    0 - 0x0
    "00000000", -- 2695 - 0xa87  :    0 - 0x0
    "00000000", -- 2696 - 0xa88  :    0 - 0x0
    "00000000", -- 2697 - 0xa89  :    0 - 0x0
    "00000000", -- 2698 - 0xa8a  :    0 - 0x0
    "00000000", -- 2699 - 0xa8b  :    0 - 0x0
    "00000000", -- 2700 - 0xa8c  :    0 - 0x0
    "00000000", -- 2701 - 0xa8d  :    0 - 0x0
    "00000000", -- 2702 - 0xa8e  :    0 - 0x0
    "00000000", -- 2703 - 0xa8f  :    0 - 0x0
    "00000000", -- 2704 - 0xa90  :    0 - 0x0
    "00000000", -- 2705 - 0xa91  :    0 - 0x0
    "00000000", -- 2706 - 0xa92  :    0 - 0x0
    "00000000", -- 2707 - 0xa93  :    0 - 0x0
    "00000000", -- 2708 - 0xa94  :    0 - 0x0
    "00000000", -- 2709 - 0xa95  :    0 - 0x0
    "00000000", -- 2710 - 0xa96  :    0 - 0x0
    "00000000", -- 2711 - 0xa97  :    0 - 0x0
    "00000000", -- 2712 - 0xa98  :    0 - 0x0
    "00000000", -- 2713 - 0xa99  :    0 - 0x0
    "00000000", -- 2714 - 0xa9a  :    0 - 0x0
    "00000000", -- 2715 - 0xa9b  :    0 - 0x0
    "00000000", -- 2716 - 0xa9c  :    0 - 0x0
    "00000000", -- 2717 - 0xa9d  :    0 - 0x0
    "00000000", -- 2718 - 0xa9e  :    0 - 0x0
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "00000000", -- 2720 - 0xaa0  :    0 - 0x0
    "00000000", -- 2721 - 0xaa1  :    0 - 0x0
    "00000000", -- 2722 - 0xaa2  :    0 - 0x0
    "00000000", -- 2723 - 0xaa3  :    0 - 0x0
    "00000000", -- 2724 - 0xaa4  :    0 - 0x0
    "00000000", -- 2725 - 0xaa5  :    0 - 0x0
    "00000000", -- 2726 - 0xaa6  :    0 - 0x0
    "00000000", -- 2727 - 0xaa7  :    0 - 0x0
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "00000000", -- 2730 - 0xaaa  :    0 - 0x0
    "00000000", -- 2731 - 0xaab  :    0 - 0x0
    "00000000", -- 2732 - 0xaac  :    0 - 0x0
    "00000000", -- 2733 - 0xaad  :    0 - 0x0
    "00000000", -- 2734 - 0xaae  :    0 - 0x0
    "00000000", -- 2735 - 0xaaf  :    0 - 0x0
    "00000000", -- 2736 - 0xab0  :    0 - 0x0
    "00000000", -- 2737 - 0xab1  :    0 - 0x0
    "00000000", -- 2738 - 0xab2  :    0 - 0x0
    "00000000", -- 2739 - 0xab3  :    0 - 0x0
    "00000000", -- 2740 - 0xab4  :    0 - 0x0
    "00000000", -- 2741 - 0xab5  :    0 - 0x0
    "00000000", -- 2742 - 0xab6  :    0 - 0x0
    "00000000", -- 2743 - 0xab7  :    0 - 0x0
    "00000000", -- 2744 - 0xab8  :    0 - 0x0
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "00000000", -- 2747 - 0xabb  :    0 - 0x0
    "00000000", -- 2748 - 0xabc  :    0 - 0x0
    "00000000", -- 2749 - 0xabd  :    0 - 0x0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "00000000", -- 2752 - 0xac0  :    0 - 0x0
    "00000000", -- 2753 - 0xac1  :    0 - 0x0
    "00000000", -- 2754 - 0xac2  :    0 - 0x0
    "00000000", -- 2755 - 0xac3  :    0 - 0x0
    "00000000", -- 2756 - 0xac4  :    0 - 0x0
    "00000000", -- 2757 - 0xac5  :    0 - 0x0
    "00000000", -- 2758 - 0xac6  :    0 - 0x0
    "00000000", -- 2759 - 0xac7  :    0 - 0x0
    "00000000", -- 2760 - 0xac8  :    0 - 0x0
    "00000000", -- 2761 - 0xac9  :    0 - 0x0
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000000", -- 2763 - 0xacb  :    0 - 0x0
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "00000000", -- 2768 - 0xad0  :    0 - 0x0
    "00000000", -- 2769 - 0xad1  :    0 - 0x0
    "00000000", -- 2770 - 0xad2  :    0 - 0x0
    "00000000", -- 2771 - 0xad3  :    0 - 0x0
    "00000000", -- 2772 - 0xad4  :    0 - 0x0
    "00000000", -- 2773 - 0xad5  :    0 - 0x0
    "00000000", -- 2774 - 0xad6  :    0 - 0x0
    "00000000", -- 2775 - 0xad7  :    0 - 0x0
    "00000000", -- 2776 - 0xad8  :    0 - 0x0
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "00000000", -- 2778 - 0xada  :    0 - 0x0
    "00000000", -- 2779 - 0xadb  :    0 - 0x0
    "00000000", -- 2780 - 0xadc  :    0 - 0x0
    "00000000", -- 2781 - 0xadd  :    0 - 0x0
    "00000000", -- 2782 - 0xade  :    0 - 0x0
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "00000000", -- 2784 - 0xae0  :    0 - 0x0
    "00000000", -- 2785 - 0xae1  :    0 - 0x0
    "00000000", -- 2786 - 0xae2  :    0 - 0x0
    "00000000", -- 2787 - 0xae3  :    0 - 0x0
    "00000000", -- 2788 - 0xae4  :    0 - 0x0
    "00000000", -- 2789 - 0xae5  :    0 - 0x0
    "00000000", -- 2790 - 0xae6  :    0 - 0x0
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "00000000", -- 2792 - 0xae8  :    0 - 0x0
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000000", -- 2794 - 0xaea  :    0 - 0x0
    "00000000", -- 2795 - 0xaeb  :    0 - 0x0
    "00000000", -- 2796 - 0xaec  :    0 - 0x0
    "00000000", -- 2797 - 0xaed  :    0 - 0x0
    "00000000", -- 2798 - 0xaee  :    0 - 0x0
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "00000000", -- 2800 - 0xaf0  :    0 - 0x0
    "00000000", -- 2801 - 0xaf1  :    0 - 0x0
    "00000000", -- 2802 - 0xaf2  :    0 - 0x0
    "00000000", -- 2803 - 0xaf3  :    0 - 0x0
    "00000000", -- 2804 - 0xaf4  :    0 - 0x0
    "00000000", -- 2805 - 0xaf5  :    0 - 0x0
    "00000000", -- 2806 - 0xaf6  :    0 - 0x0
    "00000000", -- 2807 - 0xaf7  :    0 - 0x0
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0
    "00000000", -- 2809 - 0xaf9  :    0 - 0x0
    "00000000", -- 2810 - 0xafa  :    0 - 0x0
    "00000000", -- 2811 - 0xafb  :    0 - 0x0
    "00000000", -- 2812 - 0xafc  :    0 - 0x0
    "00000000", -- 2813 - 0xafd  :    0 - 0x0
    "00000000", -- 2814 - 0xafe  :    0 - 0x0
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "00000000", -- 2816 - 0xb00  :    0 - 0x0
    "00000000", -- 2817 - 0xb01  :    0 - 0x0
    "00000000", -- 2818 - 0xb02  :    0 - 0x0
    "00000000", -- 2819 - 0xb03  :    0 - 0x0
    "00000000", -- 2820 - 0xb04  :    0 - 0x0
    "00000000", -- 2821 - 0xb05  :    0 - 0x0
    "00000000", -- 2822 - 0xb06  :    0 - 0x0
    "00000000", -- 2823 - 0xb07  :    0 - 0x0
    "00000000", -- 2824 - 0xb08  :    0 - 0x0
    "00000000", -- 2825 - 0xb09  :    0 - 0x0
    "00000000", -- 2826 - 0xb0a  :    0 - 0x0
    "00000000", -- 2827 - 0xb0b  :    0 - 0x0
    "00000000", -- 2828 - 0xb0c  :    0 - 0x0
    "00000000", -- 2829 - 0xb0d  :    0 - 0x0
    "00000000", -- 2830 - 0xb0e  :    0 - 0x0
    "00000000", -- 2831 - 0xb0f  :    0 - 0x0
    "00000000", -- 2832 - 0xb10  :    0 - 0x0
    "00000000", -- 2833 - 0xb11  :    0 - 0x0
    "00000000", -- 2834 - 0xb12  :    0 - 0x0
    "00000000", -- 2835 - 0xb13  :    0 - 0x0
    "00000000", -- 2836 - 0xb14  :    0 - 0x0
    "00000000", -- 2837 - 0xb15  :    0 - 0x0
    "00000000", -- 2838 - 0xb16  :    0 - 0x0
    "00000000", -- 2839 - 0xb17  :    0 - 0x0
    "00000000", -- 2840 - 0xb18  :    0 - 0x0
    "00000000", -- 2841 - 0xb19  :    0 - 0x0
    "00000000", -- 2842 - 0xb1a  :    0 - 0x0
    "00000000", -- 2843 - 0xb1b  :    0 - 0x0
    "00000000", -- 2844 - 0xb1c  :    0 - 0x0
    "00000000", -- 2845 - 0xb1d  :    0 - 0x0
    "00000000", -- 2846 - 0xb1e  :    0 - 0x0
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "00000000", -- 2848 - 0xb20  :    0 - 0x0
    "00000000", -- 2849 - 0xb21  :    0 - 0x0
    "00000000", -- 2850 - 0xb22  :    0 - 0x0
    "00000000", -- 2851 - 0xb23  :    0 - 0x0
    "00000000", -- 2852 - 0xb24  :    0 - 0x0
    "00000000", -- 2853 - 0xb25  :    0 - 0x0
    "00000000", -- 2854 - 0xb26  :    0 - 0x0
    "00000000", -- 2855 - 0xb27  :    0 - 0x0
    "00000000", -- 2856 - 0xb28  :    0 - 0x0
    "00000000", -- 2857 - 0xb29  :    0 - 0x0
    "00000000", -- 2858 - 0xb2a  :    0 - 0x0
    "00000000", -- 2859 - 0xb2b  :    0 - 0x0
    "00000000", -- 2860 - 0xb2c  :    0 - 0x0
    "00000000", -- 2861 - 0xb2d  :    0 - 0x0
    "00000000", -- 2862 - 0xb2e  :    0 - 0x0
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "00000000", -- 2864 - 0xb30  :    0 - 0x0
    "00000000", -- 2865 - 0xb31  :    0 - 0x0
    "00000000", -- 2866 - 0xb32  :    0 - 0x0
    "00000000", -- 2867 - 0xb33  :    0 - 0x0
    "00000000", -- 2868 - 0xb34  :    0 - 0x0
    "00000000", -- 2869 - 0xb35  :    0 - 0x0
    "00000000", -- 2870 - 0xb36  :    0 - 0x0
    "00000000", -- 2871 - 0xb37  :    0 - 0x0
    "00000000", -- 2872 - 0xb38  :    0 - 0x0
    "00000000", -- 2873 - 0xb39  :    0 - 0x0
    "00000000", -- 2874 - 0xb3a  :    0 - 0x0
    "00000000", -- 2875 - 0xb3b  :    0 - 0x0
    "00000000", -- 2876 - 0xb3c  :    0 - 0x0
    "00000000", -- 2877 - 0xb3d  :    0 - 0x0
    "00000000", -- 2878 - 0xb3e  :    0 - 0x0
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "00000000", -- 2880 - 0xb40  :    0 - 0x0
    "00000000", -- 2881 - 0xb41  :    0 - 0x0
    "00000000", -- 2882 - 0xb42  :    0 - 0x0
    "00000000", -- 2883 - 0xb43  :    0 - 0x0
    "00000000", -- 2884 - 0xb44  :    0 - 0x0
    "00000000", -- 2885 - 0xb45  :    0 - 0x0
    "00000000", -- 2886 - 0xb46  :    0 - 0x0
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "00000000", -- 2888 - 0xb48  :    0 - 0x0
    "00000000", -- 2889 - 0xb49  :    0 - 0x0
    "00000000", -- 2890 - 0xb4a  :    0 - 0x0
    "00000000", -- 2891 - 0xb4b  :    0 - 0x0
    "00000000", -- 2892 - 0xb4c  :    0 - 0x0
    "00000000", -- 2893 - 0xb4d  :    0 - 0x0
    "00000000", -- 2894 - 0xb4e  :    0 - 0x0
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "00000000", -- 2896 - 0xb50  :    0 - 0x0
    "00000000", -- 2897 - 0xb51  :    0 - 0x0
    "00000000", -- 2898 - 0xb52  :    0 - 0x0
    "00000000", -- 2899 - 0xb53  :    0 - 0x0
    "00000000", -- 2900 - 0xb54  :    0 - 0x0
    "00000000", -- 2901 - 0xb55  :    0 - 0x0
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "00000000", -- 2904 - 0xb58  :    0 - 0x0
    "00000000", -- 2905 - 0xb59  :    0 - 0x0
    "00000000", -- 2906 - 0xb5a  :    0 - 0x0
    "00000000", -- 2907 - 0xb5b  :    0 - 0x0
    "00000000", -- 2908 - 0xb5c  :    0 - 0x0
    "00000000", -- 2909 - 0xb5d  :    0 - 0x0
    "00000000", -- 2910 - 0xb5e  :    0 - 0x0
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "00000000", -- 2912 - 0xb60  :    0 - 0x0
    "00000000", -- 2913 - 0xb61  :    0 - 0x0
    "00000000", -- 2914 - 0xb62  :    0 - 0x0
    "00000000", -- 2915 - 0xb63  :    0 - 0x0
    "00000000", -- 2916 - 0xb64  :    0 - 0x0
    "00000000", -- 2917 - 0xb65  :    0 - 0x0
    "00000000", -- 2918 - 0xb66  :    0 - 0x0
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "00000000", -- 2920 - 0xb68  :    0 - 0x0
    "00000000", -- 2921 - 0xb69  :    0 - 0x0
    "00000000", -- 2922 - 0xb6a  :    0 - 0x0
    "00000000", -- 2923 - 0xb6b  :    0 - 0x0
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00000000", -- 2928 - 0xb70  :    0 - 0x0
    "00000000", -- 2929 - 0xb71  :    0 - 0x0
    "00000000", -- 2930 - 0xb72  :    0 - 0x0
    "00000000", -- 2931 - 0xb73  :    0 - 0x0
    "00000000", -- 2932 - 0xb74  :    0 - 0x0
    "00000000", -- 2933 - 0xb75  :    0 - 0x0
    "00000000", -- 2934 - 0xb76  :    0 - 0x0
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "00000000", -- 2936 - 0xb78  :    0 - 0x0
    "00000000", -- 2937 - 0xb79  :    0 - 0x0
    "00000000", -- 2938 - 0xb7a  :    0 - 0x0
    "00000000", -- 2939 - 0xb7b  :    0 - 0x0
    "00000000", -- 2940 - 0xb7c  :    0 - 0x0
    "00000000", -- 2941 - 0xb7d  :    0 - 0x0
    "00000000", -- 2942 - 0xb7e  :    0 - 0x0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "00000000", -- 2944 - 0xb80  :    0 - 0x0
    "00000000", -- 2945 - 0xb81  :    0 - 0x0
    "00000000", -- 2946 - 0xb82  :    0 - 0x0
    "00000000", -- 2947 - 0xb83  :    0 - 0x0
    "00000000", -- 2948 - 0xb84  :    0 - 0x0
    "00000000", -- 2949 - 0xb85  :    0 - 0x0
    "00000000", -- 2950 - 0xb86  :    0 - 0x0
    "00000000", -- 2951 - 0xb87  :    0 - 0x0
    "00000000", -- 2952 - 0xb88  :    0 - 0x0
    "00000000", -- 2953 - 0xb89  :    0 - 0x0
    "00000000", -- 2954 - 0xb8a  :    0 - 0x0
    "00000000", -- 2955 - 0xb8b  :    0 - 0x0
    "00000000", -- 2956 - 0xb8c  :    0 - 0x0
    "00000000", -- 2957 - 0xb8d  :    0 - 0x0
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00000000", -- 2960 - 0xb90  :    0 - 0x0
    "00000000", -- 2961 - 0xb91  :    0 - 0x0
    "00000000", -- 2962 - 0xb92  :    0 - 0x0
    "00000000", -- 2963 - 0xb93  :    0 - 0x0
    "00000000", -- 2964 - 0xb94  :    0 - 0x0
    "00000000", -- 2965 - 0xb95  :    0 - 0x0
    "00000000", -- 2966 - 0xb96  :    0 - 0x0
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "00000000", -- 2968 - 0xb98  :    0 - 0x0
    "00000000", -- 2969 - 0xb99  :    0 - 0x0
    "00000000", -- 2970 - 0xb9a  :    0 - 0x0
    "00000000", -- 2971 - 0xb9b  :    0 - 0x0
    "00000000", -- 2972 - 0xb9c  :    0 - 0x0
    "00000000", -- 2973 - 0xb9d  :    0 - 0x0
    "00000000", -- 2974 - 0xb9e  :    0 - 0x0
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "00000000", -- 2976 - 0xba0  :    0 - 0x0
    "00000000", -- 2977 - 0xba1  :    0 - 0x0
    "00000000", -- 2978 - 0xba2  :    0 - 0x0
    "00000000", -- 2979 - 0xba3  :    0 - 0x0
    "00000000", -- 2980 - 0xba4  :    0 - 0x0
    "00000000", -- 2981 - 0xba5  :    0 - 0x0
    "00000000", -- 2982 - 0xba6  :    0 - 0x0
    "00000000", -- 2983 - 0xba7  :    0 - 0x0
    "00000000", -- 2984 - 0xba8  :    0 - 0x0
    "00000000", -- 2985 - 0xba9  :    0 - 0x0
    "00000000", -- 2986 - 0xbaa  :    0 - 0x0
    "00000000", -- 2987 - 0xbab  :    0 - 0x0
    "00000000", -- 2988 - 0xbac  :    0 - 0x0
    "00000000", -- 2989 - 0xbad  :    0 - 0x0
    "00000000", -- 2990 - 0xbae  :    0 - 0x0
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "00000000", -- 2992 - 0xbb0  :    0 - 0x0
    "00000000", -- 2993 - 0xbb1  :    0 - 0x0
    "00000000", -- 2994 - 0xbb2  :    0 - 0x0
    "00000000", -- 2995 - 0xbb3  :    0 - 0x0
    "00000000", -- 2996 - 0xbb4  :    0 - 0x0
    "00000000", -- 2997 - 0xbb5  :    0 - 0x0
    "00000000", -- 2998 - 0xbb6  :    0 - 0x0
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "00000000", -- 3000 - 0xbb8  :    0 - 0x0
    "00000000", -- 3001 - 0xbb9  :    0 - 0x0
    "00000000", -- 3002 - 0xbba  :    0 - 0x0
    "00000000", -- 3003 - 0xbbb  :    0 - 0x0
    "00000000", -- 3004 - 0xbbc  :    0 - 0x0
    "00000000", -- 3005 - 0xbbd  :    0 - 0x0
    "00000000", -- 3006 - 0xbbe  :    0 - 0x0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000000", -- 3011 - 0xbc3  :    0 - 0x0
    "00000000", -- 3012 - 0xbc4  :    0 - 0x0
    "00000000", -- 3013 - 0xbc5  :    0 - 0x0
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000000", -- 3022 - 0xbce  :    0 - 0x0
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0
    "00000000", -- 3025 - 0xbd1  :    0 - 0x0
    "00000000", -- 3026 - 0xbd2  :    0 - 0x0
    "00000000", -- 3027 - 0xbd3  :    0 - 0x0
    "00000000", -- 3028 - 0xbd4  :    0 - 0x0
    "00000000", -- 3029 - 0xbd5  :    0 - 0x0
    "00000000", -- 3030 - 0xbd6  :    0 - 0x0
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0
    "00000000", -- 3033 - 0xbd9  :    0 - 0x0
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00000000", -- 3035 - 0xbdb  :    0 - 0x0
    "00000000", -- 3036 - 0xbdc  :    0 - 0x0
    "00000000", -- 3037 - 0xbdd  :    0 - 0x0
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0
    "00000000", -- 3041 - 0xbe1  :    0 - 0x0
    "00000000", -- 3042 - 0xbe2  :    0 - 0x0
    "00000000", -- 3043 - 0xbe3  :    0 - 0x0
    "00000000", -- 3044 - 0xbe4  :    0 - 0x0
    "00000000", -- 3045 - 0xbe5  :    0 - 0x0
    "00000000", -- 3046 - 0xbe6  :    0 - 0x0
    "00000000", -- 3047 - 0xbe7  :    0 - 0x0
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0
    "00000000", -- 3049 - 0xbe9  :    0 - 0x0
    "00000000", -- 3050 - 0xbea  :    0 - 0x0
    "00000000", -- 3051 - 0xbeb  :    0 - 0x0
    "00000000", -- 3052 - 0xbec  :    0 - 0x0
    "00000000", -- 3053 - 0xbed  :    0 - 0x0
    "00000000", -- 3054 - 0xbee  :    0 - 0x0
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00000000", -- 3058 - 0xbf2  :    0 - 0x0
    "00000000", -- 3059 - 0xbf3  :    0 - 0x0
    "00000000", -- 3060 - 0xbf4  :    0 - 0x0
    "00000000", -- 3061 - 0xbf5  :    0 - 0x0
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0
    "00000000", -- 3065 - 0xbf9  :    0 - 0x0
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00000000", -- 3068 - 0xbfc  :    0 - 0x0
    "00000000", -- 3069 - 0xbfd  :    0 - 0x0
    "00000000", -- 3070 - 0xbfe  :    0 - 0x0
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00000000", -- 3072 - 0xc00  :    0 - 0x0
    "00000000", -- 3073 - 0xc01  :    0 - 0x0
    "00000000", -- 3074 - 0xc02  :    0 - 0x0
    "00000000", -- 3075 - 0xc03  :    0 - 0x0
    "00000000", -- 3076 - 0xc04  :    0 - 0x0
    "00000000", -- 3077 - 0xc05  :    0 - 0x0
    "00000000", -- 3078 - 0xc06  :    0 - 0x0
    "00000000", -- 3079 - 0xc07  :    0 - 0x0
    "00000000", -- 3080 - 0xc08  :    0 - 0x0
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "00000000", -- 3083 - 0xc0b  :    0 - 0x0
    "00000000", -- 3084 - 0xc0c  :    0 - 0x0
    "00000000", -- 3085 - 0xc0d  :    0 - 0x0
    "00000000", -- 3086 - 0xc0e  :    0 - 0x0
    "00000000", -- 3087 - 0xc0f  :    0 - 0x0
    "00000000", -- 3088 - 0xc10  :    0 - 0x0
    "00000000", -- 3089 - 0xc11  :    0 - 0x0
    "00000000", -- 3090 - 0xc12  :    0 - 0x0
    "00000000", -- 3091 - 0xc13  :    0 - 0x0
    "00000000", -- 3092 - 0xc14  :    0 - 0x0
    "00000000", -- 3093 - 0xc15  :    0 - 0x0
    "00000000", -- 3094 - 0xc16  :    0 - 0x0
    "00000000", -- 3095 - 0xc17  :    0 - 0x0
    "00000000", -- 3096 - 0xc18  :    0 - 0x0
    "00000000", -- 3097 - 0xc19  :    0 - 0x0
    "00000000", -- 3098 - 0xc1a  :    0 - 0x0
    "00000000", -- 3099 - 0xc1b  :    0 - 0x0
    "00000000", -- 3100 - 0xc1c  :    0 - 0x0
    "00000000", -- 3101 - 0xc1d  :    0 - 0x0
    "00000000", -- 3102 - 0xc1e  :    0 - 0x0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00000000", -- 3104 - 0xc20  :    0 - 0x0
    "00000000", -- 3105 - 0xc21  :    0 - 0x0
    "00000000", -- 3106 - 0xc22  :    0 - 0x0
    "00000000", -- 3107 - 0xc23  :    0 - 0x0
    "00000000", -- 3108 - 0xc24  :    0 - 0x0
    "00000000", -- 3109 - 0xc25  :    0 - 0x0
    "00000000", -- 3110 - 0xc26  :    0 - 0x0
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "00000000", -- 3115 - 0xc2b  :    0 - 0x0
    "00000000", -- 3116 - 0xc2c  :    0 - 0x0
    "00000000", -- 3117 - 0xc2d  :    0 - 0x0
    "00000000", -- 3118 - 0xc2e  :    0 - 0x0
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "00000000", -- 3120 - 0xc30  :    0 - 0x0
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "00000000", -- 3122 - 0xc32  :    0 - 0x0
    "00000000", -- 3123 - 0xc33  :    0 - 0x0
    "00000000", -- 3124 - 0xc34  :    0 - 0x0
    "00000000", -- 3125 - 0xc35  :    0 - 0x0
    "00000000", -- 3126 - 0xc36  :    0 - 0x0
    "00000000", -- 3127 - 0xc37  :    0 - 0x0
    "00000000", -- 3128 - 0xc38  :    0 - 0x0
    "00000000", -- 3129 - 0xc39  :    0 - 0x0
    "00000000", -- 3130 - 0xc3a  :    0 - 0x0
    "00000000", -- 3131 - 0xc3b  :    0 - 0x0
    "00000000", -- 3132 - 0xc3c  :    0 - 0x0
    "00000000", -- 3133 - 0xc3d  :    0 - 0x0
    "00000000", -- 3134 - 0xc3e  :    0 - 0x0
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00000000", -- 3136 - 0xc40  :    0 - 0x0
    "00000000", -- 3137 - 0xc41  :    0 - 0x0
    "00000000", -- 3138 - 0xc42  :    0 - 0x0
    "00000000", -- 3139 - 0xc43  :    0 - 0x0
    "00000000", -- 3140 - 0xc44  :    0 - 0x0
    "00000000", -- 3141 - 0xc45  :    0 - 0x0
    "00000000", -- 3142 - 0xc46  :    0 - 0x0
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00000000", -- 3144 - 0xc48  :    0 - 0x0
    "00000000", -- 3145 - 0xc49  :    0 - 0x0
    "00000000", -- 3146 - 0xc4a  :    0 - 0x0
    "00000000", -- 3147 - 0xc4b  :    0 - 0x0
    "00000000", -- 3148 - 0xc4c  :    0 - 0x0
    "00000000", -- 3149 - 0xc4d  :    0 - 0x0
    "00000000", -- 3150 - 0xc4e  :    0 - 0x0
    "00000000", -- 3151 - 0xc4f  :    0 - 0x0
    "00000000", -- 3152 - 0xc50  :    0 - 0x0
    "00000000", -- 3153 - 0xc51  :    0 - 0x0
    "00000000", -- 3154 - 0xc52  :    0 - 0x0
    "00000000", -- 3155 - 0xc53  :    0 - 0x0
    "00000000", -- 3156 - 0xc54  :    0 - 0x0
    "00000000", -- 3157 - 0xc55  :    0 - 0x0
    "00000000", -- 3158 - 0xc56  :    0 - 0x0
    "00000000", -- 3159 - 0xc57  :    0 - 0x0
    "00000000", -- 3160 - 0xc58  :    0 - 0x0
    "00000000", -- 3161 - 0xc59  :    0 - 0x0
    "00000000", -- 3162 - 0xc5a  :    0 - 0x0
    "00000000", -- 3163 - 0xc5b  :    0 - 0x0
    "00000000", -- 3164 - 0xc5c  :    0 - 0x0
    "00000000", -- 3165 - 0xc5d  :    0 - 0x0
    "00000000", -- 3166 - 0xc5e  :    0 - 0x0
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "00000000", -- 3168 - 0xc60  :    0 - 0x0
    "00000000", -- 3169 - 0xc61  :    0 - 0x0
    "00000000", -- 3170 - 0xc62  :    0 - 0x0
    "00000000", -- 3171 - 0xc63  :    0 - 0x0
    "00000000", -- 3172 - 0xc64  :    0 - 0x0
    "00000000", -- 3173 - 0xc65  :    0 - 0x0
    "00000000", -- 3174 - 0xc66  :    0 - 0x0
    "00000000", -- 3175 - 0xc67  :    0 - 0x0
    "00000000", -- 3176 - 0xc68  :    0 - 0x0
    "00000000", -- 3177 - 0xc69  :    0 - 0x0
    "00000000", -- 3178 - 0xc6a  :    0 - 0x0
    "00000000", -- 3179 - 0xc6b  :    0 - 0x0
    "00000000", -- 3180 - 0xc6c  :    0 - 0x0
    "00000000", -- 3181 - 0xc6d  :    0 - 0x0
    "00000000", -- 3182 - 0xc6e  :    0 - 0x0
    "00000000", -- 3183 - 0xc6f  :    0 - 0x0
    "00000000", -- 3184 - 0xc70  :    0 - 0x0
    "00000000", -- 3185 - 0xc71  :    0 - 0x0
    "00000000", -- 3186 - 0xc72  :    0 - 0x0
    "00000000", -- 3187 - 0xc73  :    0 - 0x0
    "00000000", -- 3188 - 0xc74  :    0 - 0x0
    "00000000", -- 3189 - 0xc75  :    0 - 0x0
    "00000000", -- 3190 - 0xc76  :    0 - 0x0
    "00000000", -- 3191 - 0xc77  :    0 - 0x0
    "00000000", -- 3192 - 0xc78  :    0 - 0x0
    "00000000", -- 3193 - 0xc79  :    0 - 0x0
    "00000000", -- 3194 - 0xc7a  :    0 - 0x0
    "00000000", -- 3195 - 0xc7b  :    0 - 0x0
    "00000000", -- 3196 - 0xc7c  :    0 - 0x0
    "00000000", -- 3197 - 0xc7d  :    0 - 0x0
    "00000000", -- 3198 - 0xc7e  :    0 - 0x0
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "00000000", -- 3200 - 0xc80  :    0 - 0x0
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000000", -- 3204 - 0xc84  :    0 - 0x0
    "00000000", -- 3205 - 0xc85  :    0 - 0x0
    "00000000", -- 3206 - 0xc86  :    0 - 0x0
    "00000000", -- 3207 - 0xc87  :    0 - 0x0
    "00000000", -- 3208 - 0xc88  :    0 - 0x0
    "00000000", -- 3209 - 0xc89  :    0 - 0x0
    "00000000", -- 3210 - 0xc8a  :    0 - 0x0
    "00000000", -- 3211 - 0xc8b  :    0 - 0x0
    "00000000", -- 3212 - 0xc8c  :    0 - 0x0
    "00000000", -- 3213 - 0xc8d  :    0 - 0x0
    "00000000", -- 3214 - 0xc8e  :    0 - 0x0
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00000000", -- 3216 - 0xc90  :    0 - 0x0
    "00000000", -- 3217 - 0xc91  :    0 - 0x0
    "00000000", -- 3218 - 0xc92  :    0 - 0x0
    "00000000", -- 3219 - 0xc93  :    0 - 0x0
    "00000000", -- 3220 - 0xc94  :    0 - 0x0
    "00000000", -- 3221 - 0xc95  :    0 - 0x0
    "00000000", -- 3222 - 0xc96  :    0 - 0x0
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "00000000", -- 3224 - 0xc98  :    0 - 0x0
    "00000000", -- 3225 - 0xc99  :    0 - 0x0
    "00000000", -- 3226 - 0xc9a  :    0 - 0x0
    "00000000", -- 3227 - 0xc9b  :    0 - 0x0
    "00000000", -- 3228 - 0xc9c  :    0 - 0x0
    "00000000", -- 3229 - 0xc9d  :    0 - 0x0
    "00000000", -- 3230 - 0xc9e  :    0 - 0x0
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00000000", -- 3232 - 0xca0  :    0 - 0x0
    "00000000", -- 3233 - 0xca1  :    0 - 0x0
    "00000000", -- 3234 - 0xca2  :    0 - 0x0
    "00000000", -- 3235 - 0xca3  :    0 - 0x0
    "00000000", -- 3236 - 0xca4  :    0 - 0x0
    "00000000", -- 3237 - 0xca5  :    0 - 0x0
    "00000000", -- 3238 - 0xca6  :    0 - 0x0
    "00000000", -- 3239 - 0xca7  :    0 - 0x0
    "00000000", -- 3240 - 0xca8  :    0 - 0x0
    "00000000", -- 3241 - 0xca9  :    0 - 0x0
    "00000000", -- 3242 - 0xcaa  :    0 - 0x0
    "00000000", -- 3243 - 0xcab  :    0 - 0x0
    "00000000", -- 3244 - 0xcac  :    0 - 0x0
    "00000000", -- 3245 - 0xcad  :    0 - 0x0
    "00000000", -- 3246 - 0xcae  :    0 - 0x0
    "00000000", -- 3247 - 0xcaf  :    0 - 0x0
    "00000000", -- 3248 - 0xcb0  :    0 - 0x0
    "00000000", -- 3249 - 0xcb1  :    0 - 0x0
    "00000000", -- 3250 - 0xcb2  :    0 - 0x0
    "00000000", -- 3251 - 0xcb3  :    0 - 0x0
    "00000000", -- 3252 - 0xcb4  :    0 - 0x0
    "00000000", -- 3253 - 0xcb5  :    0 - 0x0
    "00000000", -- 3254 - 0xcb6  :    0 - 0x0
    "00000000", -- 3255 - 0xcb7  :    0 - 0x0
    "00000000", -- 3256 - 0xcb8  :    0 - 0x0
    "00000000", -- 3257 - 0xcb9  :    0 - 0x0
    "00000000", -- 3258 - 0xcba  :    0 - 0x0
    "00000000", -- 3259 - 0xcbb  :    0 - 0x0
    "00000000", -- 3260 - 0xcbc  :    0 - 0x0
    "00000000", -- 3261 - 0xcbd  :    0 - 0x0
    "00000000", -- 3262 - 0xcbe  :    0 - 0x0
    "00000000", -- 3263 - 0xcbf  :    0 - 0x0
    "00000000", -- 3264 - 0xcc0  :    0 - 0x0
    "00000000", -- 3265 - 0xcc1  :    0 - 0x0
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "00000000", -- 3267 - 0xcc3  :    0 - 0x0
    "00000000", -- 3268 - 0xcc4  :    0 - 0x0
    "00000000", -- 3269 - 0xcc5  :    0 - 0x0
    "00000000", -- 3270 - 0xcc6  :    0 - 0x0
    "00000000", -- 3271 - 0xcc7  :    0 - 0x0
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000000", -- 3274 - 0xcca  :    0 - 0x0
    "00000000", -- 3275 - 0xccb  :    0 - 0x0
    "00000000", -- 3276 - 0xccc  :    0 - 0x0
    "00000000", -- 3277 - 0xccd  :    0 - 0x0
    "00000000", -- 3278 - 0xcce  :    0 - 0x0
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00000000", -- 3282 - 0xcd2  :    0 - 0x0
    "00000000", -- 3283 - 0xcd3  :    0 - 0x0
    "00000000", -- 3284 - 0xcd4  :    0 - 0x0
    "00000000", -- 3285 - 0xcd5  :    0 - 0x0
    "00000000", -- 3286 - 0xcd6  :    0 - 0x0
    "00000000", -- 3287 - 0xcd7  :    0 - 0x0
    "00000000", -- 3288 - 0xcd8  :    0 - 0x0
    "00000000", -- 3289 - 0xcd9  :    0 - 0x0
    "00000000", -- 3290 - 0xcda  :    0 - 0x0
    "00000000", -- 3291 - 0xcdb  :    0 - 0x0
    "00000000", -- 3292 - 0xcdc  :    0 - 0x0
    "00000000", -- 3293 - 0xcdd  :    0 - 0x0
    "00000000", -- 3294 - 0xcde  :    0 - 0x0
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "00000000", -- 3296 - 0xce0  :    0 - 0x0
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "00000000", -- 3299 - 0xce3  :    0 - 0x0
    "00000000", -- 3300 - 0xce4  :    0 - 0x0
    "00000000", -- 3301 - 0xce5  :    0 - 0x0
    "00000000", -- 3302 - 0xce6  :    0 - 0x0
    "00000000", -- 3303 - 0xce7  :    0 - 0x0
    "00000000", -- 3304 - 0xce8  :    0 - 0x0
    "00000000", -- 3305 - 0xce9  :    0 - 0x0
    "00000000", -- 3306 - 0xcea  :    0 - 0x0
    "00000000", -- 3307 - 0xceb  :    0 - 0x0
    "00000000", -- 3308 - 0xcec  :    0 - 0x0
    "00000000", -- 3309 - 0xced  :    0 - 0x0
    "00000000", -- 3310 - 0xcee  :    0 - 0x0
    "00000000", -- 3311 - 0xcef  :    0 - 0x0
    "00000000", -- 3312 - 0xcf0  :    0 - 0x0
    "00000000", -- 3313 - 0xcf1  :    0 - 0x0
    "00000000", -- 3314 - 0xcf2  :    0 - 0x0
    "00000000", -- 3315 - 0xcf3  :    0 - 0x0
    "00000000", -- 3316 - 0xcf4  :    0 - 0x0
    "00000000", -- 3317 - 0xcf5  :    0 - 0x0
    "00000000", -- 3318 - 0xcf6  :    0 - 0x0
    "00000000", -- 3319 - 0xcf7  :    0 - 0x0
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0
    "00000000", -- 3321 - 0xcf9  :    0 - 0x0
    "00000000", -- 3322 - 0xcfa  :    0 - 0x0
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00000000", -- 3328 - 0xd00  :    0 - 0x0
    "00000000", -- 3329 - 0xd01  :    0 - 0x0
    "00000000", -- 3330 - 0xd02  :    0 - 0x0
    "00000000", -- 3331 - 0xd03  :    0 - 0x0
    "00000000", -- 3332 - 0xd04  :    0 - 0x0
    "00000000", -- 3333 - 0xd05  :    0 - 0x0
    "00000000", -- 3334 - 0xd06  :    0 - 0x0
    "00000000", -- 3335 - 0xd07  :    0 - 0x0
    "00000000", -- 3336 - 0xd08  :    0 - 0x0
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "00000000", -- 3338 - 0xd0a  :    0 - 0x0
    "00000000", -- 3339 - 0xd0b  :    0 - 0x0
    "00000000", -- 3340 - 0xd0c  :    0 - 0x0
    "00000000", -- 3341 - 0xd0d  :    0 - 0x0
    "00000000", -- 3342 - 0xd0e  :    0 - 0x0
    "00000000", -- 3343 - 0xd0f  :    0 - 0x0
    "00000000", -- 3344 - 0xd10  :    0 - 0x0
    "00000000", -- 3345 - 0xd11  :    0 - 0x0
    "00000000", -- 3346 - 0xd12  :    0 - 0x0
    "00000000", -- 3347 - 0xd13  :    0 - 0x0
    "00000000", -- 3348 - 0xd14  :    0 - 0x0
    "00000000", -- 3349 - 0xd15  :    0 - 0x0
    "00000000", -- 3350 - 0xd16  :    0 - 0x0
    "00000000", -- 3351 - 0xd17  :    0 - 0x0
    "00000000", -- 3352 - 0xd18  :    0 - 0x0
    "00000000", -- 3353 - 0xd19  :    0 - 0x0
    "00000000", -- 3354 - 0xd1a  :    0 - 0x0
    "00000000", -- 3355 - 0xd1b  :    0 - 0x0
    "00000000", -- 3356 - 0xd1c  :    0 - 0x0
    "00000000", -- 3357 - 0xd1d  :    0 - 0x0
    "00000000", -- 3358 - 0xd1e  :    0 - 0x0
    "00000000", -- 3359 - 0xd1f  :    0 - 0x0
    "00000000", -- 3360 - 0xd20  :    0 - 0x0
    "00000000", -- 3361 - 0xd21  :    0 - 0x0
    "00000000", -- 3362 - 0xd22  :    0 - 0x0
    "00000000", -- 3363 - 0xd23  :    0 - 0x0
    "00000000", -- 3364 - 0xd24  :    0 - 0x0
    "00000000", -- 3365 - 0xd25  :    0 - 0x0
    "00000000", -- 3366 - 0xd26  :    0 - 0x0
    "00000000", -- 3367 - 0xd27  :    0 - 0x0
    "00000000", -- 3368 - 0xd28  :    0 - 0x0
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "00000000", -- 3370 - 0xd2a  :    0 - 0x0
    "00000000", -- 3371 - 0xd2b  :    0 - 0x0
    "00000000", -- 3372 - 0xd2c  :    0 - 0x0
    "00000000", -- 3373 - 0xd2d  :    0 - 0x0
    "00000000", -- 3374 - 0xd2e  :    0 - 0x0
    "00000000", -- 3375 - 0xd2f  :    0 - 0x0
    "00000000", -- 3376 - 0xd30  :    0 - 0x0
    "00000000", -- 3377 - 0xd31  :    0 - 0x0
    "00000000", -- 3378 - 0xd32  :    0 - 0x0
    "00000000", -- 3379 - 0xd33  :    0 - 0x0
    "00000000", -- 3380 - 0xd34  :    0 - 0x0
    "00000000", -- 3381 - 0xd35  :    0 - 0x0
    "00000000", -- 3382 - 0xd36  :    0 - 0x0
    "00000000", -- 3383 - 0xd37  :    0 - 0x0
    "00000000", -- 3384 - 0xd38  :    0 - 0x0
    "00000000", -- 3385 - 0xd39  :    0 - 0x0
    "00000000", -- 3386 - 0xd3a  :    0 - 0x0
    "00000000", -- 3387 - 0xd3b  :    0 - 0x0
    "00000000", -- 3388 - 0xd3c  :    0 - 0x0
    "00000000", -- 3389 - 0xd3d  :    0 - 0x0
    "00000000", -- 3390 - 0xd3e  :    0 - 0x0
    "00000000", -- 3391 - 0xd3f  :    0 - 0x0
    "00000000", -- 3392 - 0xd40  :    0 - 0x0
    "00000000", -- 3393 - 0xd41  :    0 - 0x0
    "00000000", -- 3394 - 0xd42  :    0 - 0x0
    "00000000", -- 3395 - 0xd43  :    0 - 0x0
    "00000000", -- 3396 - 0xd44  :    0 - 0x0
    "00000000", -- 3397 - 0xd45  :    0 - 0x0
    "00000000", -- 3398 - 0xd46  :    0 - 0x0
    "00000000", -- 3399 - 0xd47  :    0 - 0x0
    "00000000", -- 3400 - 0xd48  :    0 - 0x0
    "00000000", -- 3401 - 0xd49  :    0 - 0x0
    "00000000", -- 3402 - 0xd4a  :    0 - 0x0
    "00000000", -- 3403 - 0xd4b  :    0 - 0x0
    "00000000", -- 3404 - 0xd4c  :    0 - 0x0
    "00000000", -- 3405 - 0xd4d  :    0 - 0x0
    "00000000", -- 3406 - 0xd4e  :    0 - 0x0
    "00000000", -- 3407 - 0xd4f  :    0 - 0x0
    "00000000", -- 3408 - 0xd50  :    0 - 0x0
    "00000000", -- 3409 - 0xd51  :    0 - 0x0
    "00000000", -- 3410 - 0xd52  :    0 - 0x0
    "00000000", -- 3411 - 0xd53  :    0 - 0x0
    "00000000", -- 3412 - 0xd54  :    0 - 0x0
    "00000000", -- 3413 - 0xd55  :    0 - 0x0
    "00000000", -- 3414 - 0xd56  :    0 - 0x0
    "00000000", -- 3415 - 0xd57  :    0 - 0x0
    "00000000", -- 3416 - 0xd58  :    0 - 0x0
    "00000000", -- 3417 - 0xd59  :    0 - 0x0
    "00000000", -- 3418 - 0xd5a  :    0 - 0x0
    "00000000", -- 3419 - 0xd5b  :    0 - 0x0
    "00000000", -- 3420 - 0xd5c  :    0 - 0x0
    "00000000", -- 3421 - 0xd5d  :    0 - 0x0
    "00000000", -- 3422 - 0xd5e  :    0 - 0x0
    "00000000", -- 3423 - 0xd5f  :    0 - 0x0
    "00000000", -- 3424 - 0xd60  :    0 - 0x0
    "00000000", -- 3425 - 0xd61  :    0 - 0x0
    "00000000", -- 3426 - 0xd62  :    0 - 0x0
    "00000000", -- 3427 - 0xd63  :    0 - 0x0
    "00000000", -- 3428 - 0xd64  :    0 - 0x0
    "00000000", -- 3429 - 0xd65  :    0 - 0x0
    "00000000", -- 3430 - 0xd66  :    0 - 0x0
    "00000000", -- 3431 - 0xd67  :    0 - 0x0
    "00000000", -- 3432 - 0xd68  :    0 - 0x0
    "00000000", -- 3433 - 0xd69  :    0 - 0x0
    "00000000", -- 3434 - 0xd6a  :    0 - 0x0
    "00000000", -- 3435 - 0xd6b  :    0 - 0x0
    "00000000", -- 3436 - 0xd6c  :    0 - 0x0
    "00000000", -- 3437 - 0xd6d  :    0 - 0x0
    "00000000", -- 3438 - 0xd6e  :    0 - 0x0
    "00000000", -- 3439 - 0xd6f  :    0 - 0x0
    "00000000", -- 3440 - 0xd70  :    0 - 0x0
    "00000000", -- 3441 - 0xd71  :    0 - 0x0
    "00000000", -- 3442 - 0xd72  :    0 - 0x0
    "00000000", -- 3443 - 0xd73  :    0 - 0x0
    "00000000", -- 3444 - 0xd74  :    0 - 0x0
    "00000000", -- 3445 - 0xd75  :    0 - 0x0
    "00000000", -- 3446 - 0xd76  :    0 - 0x0
    "00000000", -- 3447 - 0xd77  :    0 - 0x0
    "00000000", -- 3448 - 0xd78  :    0 - 0x0
    "00000000", -- 3449 - 0xd79  :    0 - 0x0
    "00000000", -- 3450 - 0xd7a  :    0 - 0x0
    "00000000", -- 3451 - 0xd7b  :    0 - 0x0
    "00000000", -- 3452 - 0xd7c  :    0 - 0x0
    "00000000", -- 3453 - 0xd7d  :    0 - 0x0
    "00000000", -- 3454 - 0xd7e  :    0 - 0x0
    "00000000", -- 3455 - 0xd7f  :    0 - 0x0
    "00000000", -- 3456 - 0xd80  :    0 - 0x0
    "00000000", -- 3457 - 0xd81  :    0 - 0x0
    "00000000", -- 3458 - 0xd82  :    0 - 0x0
    "00000000", -- 3459 - 0xd83  :    0 - 0x0
    "00000000", -- 3460 - 0xd84  :    0 - 0x0
    "00000000", -- 3461 - 0xd85  :    0 - 0x0
    "00000000", -- 3462 - 0xd86  :    0 - 0x0
    "00000000", -- 3463 - 0xd87  :    0 - 0x0
    "00000000", -- 3464 - 0xd88  :    0 - 0x0
    "00000000", -- 3465 - 0xd89  :    0 - 0x0
    "00000000", -- 3466 - 0xd8a  :    0 - 0x0
    "00000000", -- 3467 - 0xd8b  :    0 - 0x0
    "00000000", -- 3468 - 0xd8c  :    0 - 0x0
    "00000000", -- 3469 - 0xd8d  :    0 - 0x0
    "00000000", -- 3470 - 0xd8e  :    0 - 0x0
    "00000000", -- 3471 - 0xd8f  :    0 - 0x0
    "00000000", -- 3472 - 0xd90  :    0 - 0x0
    "00000000", -- 3473 - 0xd91  :    0 - 0x0
    "00000000", -- 3474 - 0xd92  :    0 - 0x0
    "00000000", -- 3475 - 0xd93  :    0 - 0x0
    "00000000", -- 3476 - 0xd94  :    0 - 0x0
    "00000000", -- 3477 - 0xd95  :    0 - 0x0
    "00000000", -- 3478 - 0xd96  :    0 - 0x0
    "00000000", -- 3479 - 0xd97  :    0 - 0x0
    "00000000", -- 3480 - 0xd98  :    0 - 0x0
    "00000000", -- 3481 - 0xd99  :    0 - 0x0
    "00000000", -- 3482 - 0xd9a  :    0 - 0x0
    "00000000", -- 3483 - 0xd9b  :    0 - 0x0
    "00000000", -- 3484 - 0xd9c  :    0 - 0x0
    "00000000", -- 3485 - 0xd9d  :    0 - 0x0
    "00000000", -- 3486 - 0xd9e  :    0 - 0x0
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "00000000", -- 3488 - 0xda0  :    0 - 0x0
    "00000000", -- 3489 - 0xda1  :    0 - 0x0
    "00000000", -- 3490 - 0xda2  :    0 - 0x0
    "00000000", -- 3491 - 0xda3  :    0 - 0x0
    "00000000", -- 3492 - 0xda4  :    0 - 0x0
    "00000000", -- 3493 - 0xda5  :    0 - 0x0
    "00000000", -- 3494 - 0xda6  :    0 - 0x0
    "00000000", -- 3495 - 0xda7  :    0 - 0x0
    "00000000", -- 3496 - 0xda8  :    0 - 0x0
    "00000000", -- 3497 - 0xda9  :    0 - 0x0
    "00000000", -- 3498 - 0xdaa  :    0 - 0x0
    "00000000", -- 3499 - 0xdab  :    0 - 0x0
    "00000000", -- 3500 - 0xdac  :    0 - 0x0
    "00000000", -- 3501 - 0xdad  :    0 - 0x0
    "00000000", -- 3502 - 0xdae  :    0 - 0x0
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00000000", -- 3504 - 0xdb0  :    0 - 0x0
    "00000000", -- 3505 - 0xdb1  :    0 - 0x0
    "00000000", -- 3506 - 0xdb2  :    0 - 0x0
    "00000000", -- 3507 - 0xdb3  :    0 - 0x0
    "00000000", -- 3508 - 0xdb4  :    0 - 0x0
    "00000000", -- 3509 - 0xdb5  :    0 - 0x0
    "00000000", -- 3510 - 0xdb6  :    0 - 0x0
    "00000000", -- 3511 - 0xdb7  :    0 - 0x0
    "00000000", -- 3512 - 0xdb8  :    0 - 0x0
    "00000000", -- 3513 - 0xdb9  :    0 - 0x0
    "00000000", -- 3514 - 0xdba  :    0 - 0x0
    "00000000", -- 3515 - 0xdbb  :    0 - 0x0
    "00000000", -- 3516 - 0xdbc  :    0 - 0x0
    "00000000", -- 3517 - 0xdbd  :    0 - 0x0
    "00000000", -- 3518 - 0xdbe  :    0 - 0x0
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0
    "00000000", -- 3521 - 0xdc1  :    0 - 0x0
    "00000000", -- 3522 - 0xdc2  :    0 - 0x0
    "00000000", -- 3523 - 0xdc3  :    0 - 0x0
    "00000000", -- 3524 - 0xdc4  :    0 - 0x0
    "00000000", -- 3525 - 0xdc5  :    0 - 0x0
    "00000000", -- 3526 - 0xdc6  :    0 - 0x0
    "00000000", -- 3527 - 0xdc7  :    0 - 0x0
    "00000000", -- 3528 - 0xdc8  :    0 - 0x0
    "00000000", -- 3529 - 0xdc9  :    0 - 0x0
    "00000000", -- 3530 - 0xdca  :    0 - 0x0
    "00000000", -- 3531 - 0xdcb  :    0 - 0x0
    "00000000", -- 3532 - 0xdcc  :    0 - 0x0
    "00000000", -- 3533 - 0xdcd  :    0 - 0x0
    "00000000", -- 3534 - 0xdce  :    0 - 0x0
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "00000000", -- 3536 - 0xdd0  :    0 - 0x0
    "00000000", -- 3537 - 0xdd1  :    0 - 0x0
    "00000000", -- 3538 - 0xdd2  :    0 - 0x0
    "00000000", -- 3539 - 0xdd3  :    0 - 0x0
    "00000000", -- 3540 - 0xdd4  :    0 - 0x0
    "00000000", -- 3541 - 0xdd5  :    0 - 0x0
    "00000000", -- 3542 - 0xdd6  :    0 - 0x0
    "00000000", -- 3543 - 0xdd7  :    0 - 0x0
    "00000000", -- 3544 - 0xdd8  :    0 - 0x0
    "00000000", -- 3545 - 0xdd9  :    0 - 0x0
    "00000000", -- 3546 - 0xdda  :    0 - 0x0
    "00000000", -- 3547 - 0xddb  :    0 - 0x0
    "00000000", -- 3548 - 0xddc  :    0 - 0x0
    "00000000", -- 3549 - 0xddd  :    0 - 0x0
    "00000000", -- 3550 - 0xdde  :    0 - 0x0
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "00000000", -- 3552 - 0xde0  :    0 - 0x0
    "00000000", -- 3553 - 0xde1  :    0 - 0x0
    "00000000", -- 3554 - 0xde2  :    0 - 0x0
    "00000000", -- 3555 - 0xde3  :    0 - 0x0
    "00000000", -- 3556 - 0xde4  :    0 - 0x0
    "00000000", -- 3557 - 0xde5  :    0 - 0x0
    "00000000", -- 3558 - 0xde6  :    0 - 0x0
    "00000000", -- 3559 - 0xde7  :    0 - 0x0
    "00000000", -- 3560 - 0xde8  :    0 - 0x0
    "00000000", -- 3561 - 0xde9  :    0 - 0x0
    "00000000", -- 3562 - 0xdea  :    0 - 0x0
    "00000000", -- 3563 - 0xdeb  :    0 - 0x0
    "00000000", -- 3564 - 0xdec  :    0 - 0x0
    "00000000", -- 3565 - 0xded  :    0 - 0x0
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "00000000", -- 3568 - 0xdf0  :    0 - 0x0
    "00000000", -- 3569 - 0xdf1  :    0 - 0x0
    "00000000", -- 3570 - 0xdf2  :    0 - 0x0
    "00000000", -- 3571 - 0xdf3  :    0 - 0x0
    "00000000", -- 3572 - 0xdf4  :    0 - 0x0
    "00000000", -- 3573 - 0xdf5  :    0 - 0x0
    "00000000", -- 3574 - 0xdf6  :    0 - 0x0
    "00000000", -- 3575 - 0xdf7  :    0 - 0x0
    "00000000", -- 3576 - 0xdf8  :    0 - 0x0
    "00000000", -- 3577 - 0xdf9  :    0 - 0x0
    "00000000", -- 3578 - 0xdfa  :    0 - 0x0
    "00000000", -- 3579 - 0xdfb  :    0 - 0x0
    "00000000", -- 3580 - 0xdfc  :    0 - 0x0
    "00000000", -- 3581 - 0xdfd  :    0 - 0x0
    "00000000", -- 3582 - 0xdfe  :    0 - 0x0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "00000000", -- 3584 - 0xe00  :    0 - 0x0
    "00000000", -- 3585 - 0xe01  :    0 - 0x0
    "00000000", -- 3586 - 0xe02  :    0 - 0x0
    "00000000", -- 3587 - 0xe03  :    0 - 0x0
    "00000000", -- 3588 - 0xe04  :    0 - 0x0
    "00000000", -- 3589 - 0xe05  :    0 - 0x0
    "00000000", -- 3590 - 0xe06  :    0 - 0x0
    "00000000", -- 3591 - 0xe07  :    0 - 0x0
    "00000000", -- 3592 - 0xe08  :    0 - 0x0
    "00000000", -- 3593 - 0xe09  :    0 - 0x0
    "00000000", -- 3594 - 0xe0a  :    0 - 0x0
    "00000000", -- 3595 - 0xe0b  :    0 - 0x0
    "00000000", -- 3596 - 0xe0c  :    0 - 0x0
    "00000000", -- 3597 - 0xe0d  :    0 - 0x0
    "00000000", -- 3598 - 0xe0e  :    0 - 0x0
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "00000000", -- 3600 - 0xe10  :    0 - 0x0
    "00000000", -- 3601 - 0xe11  :    0 - 0x0
    "00000000", -- 3602 - 0xe12  :    0 - 0x0
    "00000000", -- 3603 - 0xe13  :    0 - 0x0
    "00000000", -- 3604 - 0xe14  :    0 - 0x0
    "00000000", -- 3605 - 0xe15  :    0 - 0x0
    "00000000", -- 3606 - 0xe16  :    0 - 0x0
    "00000000", -- 3607 - 0xe17  :    0 - 0x0
    "00000000", -- 3608 - 0xe18  :    0 - 0x0
    "00000000", -- 3609 - 0xe19  :    0 - 0x0
    "00000000", -- 3610 - 0xe1a  :    0 - 0x0
    "00000000", -- 3611 - 0xe1b  :    0 - 0x0
    "00000000", -- 3612 - 0xe1c  :    0 - 0x0
    "00000000", -- 3613 - 0xe1d  :    0 - 0x0
    "00000000", -- 3614 - 0xe1e  :    0 - 0x0
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "00000000", -- 3616 - 0xe20  :    0 - 0x0
    "00000000", -- 3617 - 0xe21  :    0 - 0x0
    "00000000", -- 3618 - 0xe22  :    0 - 0x0
    "00000000", -- 3619 - 0xe23  :    0 - 0x0
    "00000000", -- 3620 - 0xe24  :    0 - 0x0
    "00000000", -- 3621 - 0xe25  :    0 - 0x0
    "00000000", -- 3622 - 0xe26  :    0 - 0x0
    "00000000", -- 3623 - 0xe27  :    0 - 0x0
    "00000000", -- 3624 - 0xe28  :    0 - 0x0
    "00000000", -- 3625 - 0xe29  :    0 - 0x0
    "00000000", -- 3626 - 0xe2a  :    0 - 0x0
    "00000000", -- 3627 - 0xe2b  :    0 - 0x0
    "00000000", -- 3628 - 0xe2c  :    0 - 0x0
    "00000000", -- 3629 - 0xe2d  :    0 - 0x0
    "00000000", -- 3630 - 0xe2e  :    0 - 0x0
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "00000000", -- 3632 - 0xe30  :    0 - 0x0
    "00000000", -- 3633 - 0xe31  :    0 - 0x0
    "00000000", -- 3634 - 0xe32  :    0 - 0x0
    "00000000", -- 3635 - 0xe33  :    0 - 0x0
    "00000000", -- 3636 - 0xe34  :    0 - 0x0
    "00000000", -- 3637 - 0xe35  :    0 - 0x0
    "00000000", -- 3638 - 0xe36  :    0 - 0x0
    "00000000", -- 3639 - 0xe37  :    0 - 0x0
    "00000000", -- 3640 - 0xe38  :    0 - 0x0
    "00000000", -- 3641 - 0xe39  :    0 - 0x0
    "00000000", -- 3642 - 0xe3a  :    0 - 0x0
    "00000000", -- 3643 - 0xe3b  :    0 - 0x0
    "00000000", -- 3644 - 0xe3c  :    0 - 0x0
    "00000000", -- 3645 - 0xe3d  :    0 - 0x0
    "00000000", -- 3646 - 0xe3e  :    0 - 0x0
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "00000000", -- 3648 - 0xe40  :    0 - 0x0
    "00000000", -- 3649 - 0xe41  :    0 - 0x0
    "00000000", -- 3650 - 0xe42  :    0 - 0x0
    "00000000", -- 3651 - 0xe43  :    0 - 0x0
    "00000000", -- 3652 - 0xe44  :    0 - 0x0
    "00000000", -- 3653 - 0xe45  :    0 - 0x0
    "00000000", -- 3654 - 0xe46  :    0 - 0x0
    "00000000", -- 3655 - 0xe47  :    0 - 0x0
    "00000000", -- 3656 - 0xe48  :    0 - 0x0
    "00000000", -- 3657 - 0xe49  :    0 - 0x0
    "00000000", -- 3658 - 0xe4a  :    0 - 0x0
    "00000000", -- 3659 - 0xe4b  :    0 - 0x0
    "00000000", -- 3660 - 0xe4c  :    0 - 0x0
    "00000000", -- 3661 - 0xe4d  :    0 - 0x0
    "00000000", -- 3662 - 0xe4e  :    0 - 0x0
    "00000000", -- 3663 - 0xe4f  :    0 - 0x0
    "00000000", -- 3664 - 0xe50  :    0 - 0x0
    "00000000", -- 3665 - 0xe51  :    0 - 0x0
    "00000000", -- 3666 - 0xe52  :    0 - 0x0
    "00000000", -- 3667 - 0xe53  :    0 - 0x0
    "00000000", -- 3668 - 0xe54  :    0 - 0x0
    "00000000", -- 3669 - 0xe55  :    0 - 0x0
    "00000000", -- 3670 - 0xe56  :    0 - 0x0
    "00000000", -- 3671 - 0xe57  :    0 - 0x0
    "00000000", -- 3672 - 0xe58  :    0 - 0x0
    "00000000", -- 3673 - 0xe59  :    0 - 0x0
    "00000000", -- 3674 - 0xe5a  :    0 - 0x0
    "00000000", -- 3675 - 0xe5b  :    0 - 0x0
    "00000000", -- 3676 - 0xe5c  :    0 - 0x0
    "00000000", -- 3677 - 0xe5d  :    0 - 0x0
    "00000000", -- 3678 - 0xe5e  :    0 - 0x0
    "00000000", -- 3679 - 0xe5f  :    0 - 0x0
    "00000000", -- 3680 - 0xe60  :    0 - 0x0
    "00000000", -- 3681 - 0xe61  :    0 - 0x0
    "00000000", -- 3682 - 0xe62  :    0 - 0x0
    "00000000", -- 3683 - 0xe63  :    0 - 0x0
    "00000000", -- 3684 - 0xe64  :    0 - 0x0
    "00000000", -- 3685 - 0xe65  :    0 - 0x0
    "00000000", -- 3686 - 0xe66  :    0 - 0x0
    "00000000", -- 3687 - 0xe67  :    0 - 0x0
    "00111111", -- 3688 - 0xe68  :   63 - 0x3f
    "01111111", -- 3689 - 0xe69  :  127 - 0x7f
    "11111111", -- 3690 - 0xe6a  :  255 - 0xff
    "11110000", -- 3691 - 0xe6b  :  240 - 0xf0
    "11100000", -- 3692 - 0xe6c  :  224 - 0xe0
    "11100011", -- 3693 - 0xe6d  :  227 - 0xe3
    "11100111", -- 3694 - 0xe6e  :  231 - 0xe7
    "11100111", -- 3695 - 0xe6f  :  231 - 0xe7
    "11111100", -- 3696 - 0xe70  :  252 - 0xfc
    "11111110", -- 3697 - 0xe71  :  254 - 0xfe
    "11111111", -- 3698 - 0xe72  :  255 - 0xff
    "00001111", -- 3699 - 0xe73  :   15 - 0xf
    "00000111", -- 3700 - 0xe74  :    7 - 0x7
    "11000111", -- 3701 - 0xe75  :  199 - 0xc7
    "11100111", -- 3702 - 0xe76  :  231 - 0xe7
    "11100111", -- 3703 - 0xe77  :  231 - 0xe7
    "00000000", -- 3704 - 0xe78  :    0 - 0x0
    "00000000", -- 3705 - 0xe79  :    0 - 0x0
    "00000000", -- 3706 - 0xe7a  :    0 - 0x0
    "00000000", -- 3707 - 0xe7b  :    0 - 0x0
    "00000000", -- 3708 - 0xe7c  :    0 - 0x0
    "00000000", -- 3709 - 0xe7d  :    0 - 0x0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "00000000", -- 3712 - 0xe80  :    0 - 0x0
    "00000000", -- 3713 - 0xe81  :    0 - 0x0
    "00000000", -- 3714 - 0xe82  :    0 - 0x0
    "00000000", -- 3715 - 0xe83  :    0 - 0x0
    "00000000", -- 3716 - 0xe84  :    0 - 0x0
    "00000000", -- 3717 - 0xe85  :    0 - 0x0
    "00000000", -- 3718 - 0xe86  :    0 - 0x0
    "00000000", -- 3719 - 0xe87  :    0 - 0x0
    "00000000", -- 3720 - 0xe88  :    0 - 0x0
    "00000000", -- 3721 - 0xe89  :    0 - 0x0
    "00000000", -- 3722 - 0xe8a  :    0 - 0x0
    "00000000", -- 3723 - 0xe8b  :    0 - 0x0
    "00000000", -- 3724 - 0xe8c  :    0 - 0x0
    "00000000", -- 3725 - 0xe8d  :    0 - 0x0
    "00000000", -- 3726 - 0xe8e  :    0 - 0x0
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "00000000", -- 3728 - 0xe90  :    0 - 0x0
    "00000000", -- 3729 - 0xe91  :    0 - 0x0
    "00000000", -- 3730 - 0xe92  :    0 - 0x0
    "00000000", -- 3731 - 0xe93  :    0 - 0x0
    "00000000", -- 3732 - 0xe94  :    0 - 0x0
    "00000000", -- 3733 - 0xe95  :    0 - 0x0
    "00000000", -- 3734 - 0xe96  :    0 - 0x0
    "00000000", -- 3735 - 0xe97  :    0 - 0x0
    "00000000", -- 3736 - 0xe98  :    0 - 0x0
    "00000000", -- 3737 - 0xe99  :    0 - 0x0
    "00000000", -- 3738 - 0xe9a  :    0 - 0x0
    "00000000", -- 3739 - 0xe9b  :    0 - 0x0
    "00000000", -- 3740 - 0xe9c  :    0 - 0x0
    "00000000", -- 3741 - 0xe9d  :    0 - 0x0
    "00000000", -- 3742 - 0xe9e  :    0 - 0x0
    "00000000", -- 3743 - 0xe9f  :    0 - 0x0
    "00000000", -- 3744 - 0xea0  :    0 - 0x0
    "00000000", -- 3745 - 0xea1  :    0 - 0x0
    "00000000", -- 3746 - 0xea2  :    0 - 0x0
    "00000000", -- 3747 - 0xea3  :    0 - 0x0
    "00000000", -- 3748 - 0xea4  :    0 - 0x0
    "00000000", -- 3749 - 0xea5  :    0 - 0x0
    "00000000", -- 3750 - 0xea6  :    0 - 0x0
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "00000000", -- 3752 - 0xea8  :    0 - 0x0
    "00000000", -- 3753 - 0xea9  :    0 - 0x0
    "00000000", -- 3754 - 0xeaa  :    0 - 0x0
    "00000000", -- 3755 - 0xeab  :    0 - 0x0
    "00000000", -- 3756 - 0xeac  :    0 - 0x0
    "00000000", -- 3757 - 0xead  :    0 - 0x0
    "00000000", -- 3758 - 0xeae  :    0 - 0x0
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0
    "00000000", -- 3761 - 0xeb1  :    0 - 0x0
    "00000000", -- 3762 - 0xeb2  :    0 - 0x0
    "00000000", -- 3763 - 0xeb3  :    0 - 0x0
    "00000000", -- 3764 - 0xeb4  :    0 - 0x0
    "00000000", -- 3765 - 0xeb5  :    0 - 0x0
    "00000000", -- 3766 - 0xeb6  :    0 - 0x0
    "00000000", -- 3767 - 0xeb7  :    0 - 0x0
    "00000000", -- 3768 - 0xeb8  :    0 - 0x0
    "00000000", -- 3769 - 0xeb9  :    0 - 0x0
    "00000000", -- 3770 - 0xeba  :    0 - 0x0
    "00000000", -- 3771 - 0xebb  :    0 - 0x0
    "00000000", -- 3772 - 0xebc  :    0 - 0x0
    "00000000", -- 3773 - 0xebd  :    0 - 0x0
    "00000000", -- 3774 - 0xebe  :    0 - 0x0
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "00000000", -- 3776 - 0xec0  :    0 - 0x0
    "00000000", -- 3777 - 0xec1  :    0 - 0x0
    "00000000", -- 3778 - 0xec2  :    0 - 0x0
    "00000000", -- 3779 - 0xec3  :    0 - 0x0
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00000000", -- 3781 - 0xec5  :    0 - 0x0
    "00000000", -- 3782 - 0xec6  :    0 - 0x0
    "00000000", -- 3783 - 0xec7  :    0 - 0x0
    "00000000", -- 3784 - 0xec8  :    0 - 0x0
    "00000000", -- 3785 - 0xec9  :    0 - 0x0
    "00000000", -- 3786 - 0xeca  :    0 - 0x0
    "00000000", -- 3787 - 0xecb  :    0 - 0x0
    "00000000", -- 3788 - 0xecc  :    0 - 0x0
    "00000000", -- 3789 - 0xecd  :    0 - 0x0
    "00000000", -- 3790 - 0xece  :    0 - 0x0
    "00000000", -- 3791 - 0xecf  :    0 - 0x0
    "00000000", -- 3792 - 0xed0  :    0 - 0x0
    "00000000", -- 3793 - 0xed1  :    0 - 0x0
    "00000000", -- 3794 - 0xed2  :    0 - 0x0
    "00000000", -- 3795 - 0xed3  :    0 - 0x0
    "00000000", -- 3796 - 0xed4  :    0 - 0x0
    "00000000", -- 3797 - 0xed5  :    0 - 0x0
    "00000000", -- 3798 - 0xed6  :    0 - 0x0
    "00000000", -- 3799 - 0xed7  :    0 - 0x0
    "00000000", -- 3800 - 0xed8  :    0 - 0x0
    "00000000", -- 3801 - 0xed9  :    0 - 0x0
    "00000000", -- 3802 - 0xeda  :    0 - 0x0
    "00000000", -- 3803 - 0xedb  :    0 - 0x0
    "00000000", -- 3804 - 0xedc  :    0 - 0x0
    "00000000", -- 3805 - 0xedd  :    0 - 0x0
    "00000000", -- 3806 - 0xede  :    0 - 0x0
    "00000000", -- 3807 - 0xedf  :    0 - 0x0
    "00000000", -- 3808 - 0xee0  :    0 - 0x0
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000000", -- 3811 - 0xee3  :    0 - 0x0
    "00000000", -- 3812 - 0xee4  :    0 - 0x0
    "00000000", -- 3813 - 0xee5  :    0 - 0x0
    "00000000", -- 3814 - 0xee6  :    0 - 0x0
    "00000000", -- 3815 - 0xee7  :    0 - 0x0
    "11100111", -- 3816 - 0xee8  :  231 - 0xe7
    "11100111", -- 3817 - 0xee9  :  231 - 0xe7
    "11100011", -- 3818 - 0xeea  :  227 - 0xe3
    "11100000", -- 3819 - 0xeeb  :  224 - 0xe0
    "11110000", -- 3820 - 0xeec  :  240 - 0xf0
    "11111111", -- 3821 - 0xeed  :  255 - 0xff
    "01111111", -- 3822 - 0xeee  :  127 - 0x7f
    "00111111", -- 3823 - 0xeef  :   63 - 0x3f
    "11100111", -- 3824 - 0xef0  :  231 - 0xe7
    "11100111", -- 3825 - 0xef1  :  231 - 0xe7
    "11000111", -- 3826 - 0xef2  :  199 - 0xc7
    "00000111", -- 3827 - 0xef3  :    7 - 0x7
    "00001111", -- 3828 - 0xef4  :   15 - 0xf
    "11111111", -- 3829 - 0xef5  :  255 - 0xff
    "11111110", -- 3830 - 0xef6  :  254 - 0xfe
    "11111100", -- 3831 - 0xef7  :  252 - 0xfc
    "00000000", -- 3832 - 0xef8  :    0 - 0x0
    "00000000", -- 3833 - 0xef9  :    0 - 0x0
    "00000000", -- 3834 - 0xefa  :    0 - 0x0
    "00000000", -- 3835 - 0xefb  :    0 - 0x0
    "00000000", -- 3836 - 0xefc  :    0 - 0x0
    "00000000", -- 3837 - 0xefd  :    0 - 0x0
    "00000000", -- 3838 - 0xefe  :    0 - 0x0
    "00000000", -- 3839 - 0xeff  :    0 - 0x0
    "00000000", -- 3840 - 0xf00  :    0 - 0x0
    "00000000", -- 3841 - 0xf01  :    0 - 0x0
    "00000000", -- 3842 - 0xf02  :    0 - 0x0
    "00000000", -- 3843 - 0xf03  :    0 - 0x0
    "00000000", -- 3844 - 0xf04  :    0 - 0x0
    "00000000", -- 3845 - 0xf05  :    0 - 0x0
    "00000000", -- 3846 - 0xf06  :    0 - 0x0
    "00000000", -- 3847 - 0xf07  :    0 - 0x0
    "00000000", -- 3848 - 0xf08  :    0 - 0x0
    "00000000", -- 3849 - 0xf09  :    0 - 0x0
    "00000000", -- 3850 - 0xf0a  :    0 - 0x0
    "00000000", -- 3851 - 0xf0b  :    0 - 0x0
    "00000000", -- 3852 - 0xf0c  :    0 - 0x0
    "00000000", -- 3853 - 0xf0d  :    0 - 0x0
    "00000000", -- 3854 - 0xf0e  :    0 - 0x0
    "00000000", -- 3855 - 0xf0f  :    0 - 0x0
    "00000000", -- 3856 - 0xf10  :    0 - 0x0
    "00000000", -- 3857 - 0xf11  :    0 - 0x0
    "00000000", -- 3858 - 0xf12  :    0 - 0x0
    "00000000", -- 3859 - 0xf13  :    0 - 0x0
    "00000000", -- 3860 - 0xf14  :    0 - 0x0
    "00000000", -- 3861 - 0xf15  :    0 - 0x0
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "00000000", -- 3864 - 0xf18  :    0 - 0x0
    "00000000", -- 3865 - 0xf19  :    0 - 0x0
    "00000000", -- 3866 - 0xf1a  :    0 - 0x0
    "00000000", -- 3867 - 0xf1b  :    0 - 0x0
    "00000000", -- 3868 - 0xf1c  :    0 - 0x0
    "00000000", -- 3869 - 0xf1d  :    0 - 0x0
    "00000000", -- 3870 - 0xf1e  :    0 - 0x0
    "00000000", -- 3871 - 0xf1f  :    0 - 0x0
    "00000000", -- 3872 - 0xf20  :    0 - 0x0
    "00000000", -- 3873 - 0xf21  :    0 - 0x0
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000000", -- 3876 - 0xf24  :    0 - 0x0
    "00000000", -- 3877 - 0xf25  :    0 - 0x0
    "00000000", -- 3878 - 0xf26  :    0 - 0x0
    "00000000", -- 3879 - 0xf27  :    0 - 0x0
    "01111111", -- 3880 - 0xf28  :  127 - 0x7f
    "11111111", -- 3881 - 0xf29  :  255 - 0xff
    "11111111", -- 3882 - 0xf2a  :  255 - 0xff
    "11100000", -- 3883 - 0xf2b  :  224 - 0xe0
    "11100000", -- 3884 - 0xf2c  :  224 - 0xe0
    "11100000", -- 3885 - 0xf2d  :  224 - 0xe0
    "11100000", -- 3886 - 0xf2e  :  224 - 0xe0
    "11100001", -- 3887 - 0xf2f  :  225 - 0xe1
    "11111110", -- 3888 - 0xf30  :  254 - 0xfe
    "11111111", -- 3889 - 0xf31  :  255 - 0xff
    "11111111", -- 3890 - 0xf32  :  255 - 0xff
    "00000111", -- 3891 - 0xf33  :    7 - 0x7
    "00000111", -- 3892 - 0xf34  :    7 - 0x7
    "00000111", -- 3893 - 0xf35  :    7 - 0x7
    "00000111", -- 3894 - 0xf36  :    7 - 0x7
    "10000111", -- 3895 - 0xf37  :  135 - 0x87
    "00011111", -- 3896 - 0xf38  :   31 - 0x1f
    "00100000", -- 3897 - 0xf39  :   32 - 0x20
    "01000000", -- 3898 - 0xf3a  :   64 - 0x40
    "10000000", -- 3899 - 0xf3b  :  128 - 0x80
    "10000000", -- 3900 - 0xf3c  :  128 - 0x80
    "10000011", -- 3901 - 0xf3d  :  131 - 0x83
    "10000111", -- 3902 - 0xf3e  :  135 - 0x87
    "10000111", -- 3903 - 0xf3f  :  135 - 0x87
    "11111000", -- 3904 - 0xf40  :  248 - 0xf8
    "00000100", -- 3905 - 0xf41  :    4 - 0x4
    "00000010", -- 3906 - 0xf42  :    2 - 0x2
    "00000001", -- 3907 - 0xf43  :    1 - 0x1
    "00000001", -- 3908 - 0xf44  :    1 - 0x1
    "11000001", -- 3909 - 0xf45  :  193 - 0xc1
    "11100001", -- 3910 - 0xf46  :  225 - 0xe1
    "11100001", -- 3911 - 0xf47  :  225 - 0xe1
    "00000000", -- 3912 - 0xf48  :    0 - 0x0
    "00000000", -- 3913 - 0xf49  :    0 - 0x0
    "00001000", -- 3914 - 0xf4a  :    8 - 0x8
    "00010100", -- 3915 - 0xf4b  :   20 - 0x14
    "00000000", -- 3916 - 0xf4c  :    0 - 0x0
    "00000000", -- 3917 - 0xf4d  :    0 - 0x0
    "01000000", -- 3918 - 0xf4e  :   64 - 0x40
    "10100000", -- 3919 - 0xf4f  :  160 - 0xa0
    "01000000", -- 3920 - 0xf50  :   64 - 0x40
    "10100010", -- 3921 - 0xf51  :  162 - 0xa2
    "00000101", -- 3922 - 0xf52  :    5 - 0x5
    "00000000", -- 3923 - 0xf53  :    0 - 0x0
    "00000000", -- 3924 - 0xf54  :    0 - 0x0
    "00010000", -- 3925 - 0xf55  :   16 - 0x10
    "00101000", -- 3926 - 0xf56  :   40 - 0x28
    "00000000", -- 3927 - 0xf57  :    0 - 0x0
    "11111111", -- 3928 - 0xf58  :  255 - 0xff
    "11111111", -- 3929 - 0xf59  :  255 - 0xff
    "11111111", -- 3930 - 0xf5a  :  255 - 0xff
    "00000000", -- 3931 - 0xf5b  :    0 - 0x0
    "00000000", -- 3932 - 0xf5c  :    0 - 0x0
    "00000000", -- 3933 - 0xf5d  :    0 - 0x0
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "11111111", -- 3935 - 0xf5f  :  255 - 0xff
    "11100001", -- 3936 - 0xf60  :  225 - 0xe1
    "11100001", -- 3937 - 0xf61  :  225 - 0xe1
    "11100001", -- 3938 - 0xf62  :  225 - 0xe1
    "11100001", -- 3939 - 0xf63  :  225 - 0xe1
    "11100001", -- 3940 - 0xf64  :  225 - 0xe1
    "11100001", -- 3941 - 0xf65  :  225 - 0xe1
    "11100001", -- 3942 - 0xf66  :  225 - 0xe1
    "11100001", -- 3943 - 0xf67  :  225 - 0xe1
    "11111111", -- 3944 - 0xf68  :  255 - 0xff
    "11111111", -- 3945 - 0xf69  :  255 - 0xff
    "11111111", -- 3946 - 0xf6a  :  255 - 0xff
    "00000000", -- 3947 - 0xf6b  :    0 - 0x0
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "11111111", -- 3949 - 0xf6d  :  255 - 0xff
    "11111111", -- 3950 - 0xf6e  :  255 - 0xff
    "11111111", -- 3951 - 0xf6f  :  255 - 0xff
    "11100111", -- 3952 - 0xf70  :  231 - 0xe7
    "11100111", -- 3953 - 0xf71  :  231 - 0xe7
    "11100111", -- 3954 - 0xf72  :  231 - 0xe7
    "11100111", -- 3955 - 0xf73  :  231 - 0xe7
    "11100111", -- 3956 - 0xf74  :  231 - 0xe7
    "11100111", -- 3957 - 0xf75  :  231 - 0xe7
    "11100111", -- 3958 - 0xf76  :  231 - 0xe7
    "11100111", -- 3959 - 0xf77  :  231 - 0xe7
    "11111111", -- 3960 - 0xf78  :  255 - 0xff
    "11111111", -- 3961 - 0xf79  :  255 - 0xff
    "11111111", -- 3962 - 0xf7a  :  255 - 0xff
    "11111111", -- 3963 - 0xf7b  :  255 - 0xff
    "11111111", -- 3964 - 0xf7c  :  255 - 0xff
    "11111111", -- 3965 - 0xf7d  :  255 - 0xff
    "11111111", -- 3966 - 0xf7e  :  255 - 0xff
    "11111111", -- 3967 - 0xf7f  :  255 - 0xff
    "00000000", -- 3968 - 0xf80  :    0 - 0x0
    "00000000", -- 3969 - 0xf81  :    0 - 0x0
    "00000000", -- 3970 - 0xf82  :    0 - 0x0
    "00000000", -- 3971 - 0xf83  :    0 - 0x0
    "00000000", -- 3972 - 0xf84  :    0 - 0x0
    "00000000", -- 3973 - 0xf85  :    0 - 0x0
    "00000000", -- 3974 - 0xf86  :    0 - 0x0
    "00000000", -- 3975 - 0xf87  :    0 - 0x0
    "00000000", -- 3976 - 0xf88  :    0 - 0x0
    "00000000", -- 3977 - 0xf89  :    0 - 0x0
    "00000000", -- 3978 - 0xf8a  :    0 - 0x0
    "00000000", -- 3979 - 0xf8b  :    0 - 0x0
    "00000000", -- 3980 - 0xf8c  :    0 - 0x0
    "00000000", -- 3981 - 0xf8d  :    0 - 0x0
    "00000000", -- 3982 - 0xf8e  :    0 - 0x0
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "00000000", -- 3984 - 0xf90  :    0 - 0x0
    "00000000", -- 3985 - 0xf91  :    0 - 0x0
    "00000000", -- 3986 - 0xf92  :    0 - 0x0
    "00000000", -- 3987 - 0xf93  :    0 - 0x0
    "00000000", -- 3988 - 0xf94  :    0 - 0x0
    "00000000", -- 3989 - 0xf95  :    0 - 0x0
    "00000000", -- 3990 - 0xf96  :    0 - 0x0
    "00000000", -- 3991 - 0xf97  :    0 - 0x0
    "00000000", -- 3992 - 0xf98  :    0 - 0x0
    "00000000", -- 3993 - 0xf99  :    0 - 0x0
    "00000000", -- 3994 - 0xf9a  :    0 - 0x0
    "00000000", -- 3995 - 0xf9b  :    0 - 0x0
    "00000000", -- 3996 - 0xf9c  :    0 - 0x0
    "00000000", -- 3997 - 0xf9d  :    0 - 0x0
    "00000000", -- 3998 - 0xf9e  :    0 - 0x0
    "00000000", -- 3999 - 0xf9f  :    0 - 0x0
    "11100111", -- 4000 - 0xfa0  :  231 - 0xe7
    "10011001", -- 4001 - 0xfa1  :  153 - 0x99
    "10000001", -- 4002 - 0xfa2  :  129 - 0x81
    "11000011", -- 4003 - 0xfa3  :  195 - 0xc3
    "11111111", -- 4004 - 0xfa4  :  255 - 0xff
    "10111101", -- 4005 - 0xfa5  :  189 - 0xbd
    "10000001", -- 4006 - 0xfa6  :  129 - 0x81
    "11000011", -- 4007 - 0xfa7  :  195 - 0xc3
    "11100001", -- 4008 - 0xfa8  :  225 - 0xe1
    "11100000", -- 4009 - 0xfa9  :  224 - 0xe0
    "11100000", -- 4010 - 0xfaa  :  224 - 0xe0
    "11100000", -- 4011 - 0xfab  :  224 - 0xe0
    "11100000", -- 4012 - 0xfac  :  224 - 0xe0
    "11111111", -- 4013 - 0xfad  :  255 - 0xff
    "11111111", -- 4014 - 0xfae  :  255 - 0xff
    "01111111", -- 4015 - 0xfaf  :  127 - 0x7f
    "10000111", -- 4016 - 0xfb0  :  135 - 0x87
    "00000111", -- 4017 - 0xfb1  :    7 - 0x7
    "00000111", -- 4018 - 0xfb2  :    7 - 0x7
    "00000111", -- 4019 - 0xfb3  :    7 - 0x7
    "00000111", -- 4020 - 0xfb4  :    7 - 0x7
    "11111111", -- 4021 - 0xfb5  :  255 - 0xff
    "11111111", -- 4022 - 0xfb6  :  255 - 0xff
    "11111110", -- 4023 - 0xfb7  :  254 - 0xfe
    "10000111", -- 4024 - 0xfb8  :  135 - 0x87
    "10000111", -- 4025 - 0xfb9  :  135 - 0x87
    "10000011", -- 4026 - 0xfba  :  131 - 0x83
    "10000000", -- 4027 - 0xfbb  :  128 - 0x80
    "10000000", -- 4028 - 0xfbc  :  128 - 0x80
    "01000000", -- 4029 - 0xfbd  :   64 - 0x40
    "00100000", -- 4030 - 0xfbe  :   32 - 0x20
    "00011111", -- 4031 - 0xfbf  :   31 - 0x1f
    "11100001", -- 4032 - 0xfc0  :  225 - 0xe1
    "11100001", -- 4033 - 0xfc1  :  225 - 0xe1
    "11000001", -- 4034 - 0xfc2  :  193 - 0xc1
    "00000001", -- 4035 - 0xfc3  :    1 - 0x1
    "00000001", -- 4036 - 0xfc4  :    1 - 0x1
    "00000010", -- 4037 - 0xfc5  :    2 - 0x2
    "00000100", -- 4038 - 0xfc6  :    4 - 0x4
    "11111000", -- 4039 - 0xfc7  :  248 - 0xf8
    "00000000", -- 4040 - 0xfc8  :    0 - 0x0
    "00000010", -- 4041 - 0xfc9  :    2 - 0x2
    "00000101", -- 4042 - 0xfca  :    5 - 0x5
    "00000000", -- 4043 - 0xfcb  :    0 - 0x0
    "00100000", -- 4044 - 0xfcc  :   32 - 0x20
    "01010000", -- 4045 - 0xfcd  :   80 - 0x50
    "00000000", -- 4046 - 0xfce  :    0 - 0x0
    "00000000", -- 4047 - 0xfcf  :    0 - 0x0
    "00000000", -- 4048 - 0xfd0  :    0 - 0x0
    "00000000", -- 4049 - 0xfd1  :    0 - 0x0
    "00000000", -- 4050 - 0xfd2  :    0 - 0x0
    "00000000", -- 4051 - 0xfd3  :    0 - 0x0
    "00000000", -- 4052 - 0xfd4  :    0 - 0x0
    "00000000", -- 4053 - 0xfd5  :    0 - 0x0
    "00000000", -- 4054 - 0xfd6  :    0 - 0x0
    "00000000", -- 4055 - 0xfd7  :    0 - 0x0
    "11111111", -- 4056 - 0xfd8  :  255 - 0xff
    "00000000", -- 4057 - 0xfd9  :    0 - 0x0
    "00000000", -- 4058 - 0xfda  :    0 - 0x0
    "00000000", -- 4059 - 0xfdb  :    0 - 0x0
    "00000000", -- 4060 - 0xfdc  :    0 - 0x0
    "11111111", -- 4061 - 0xfdd  :  255 - 0xff
    "11111111", -- 4062 - 0xfde  :  255 - 0xff
    "11111111", -- 4063 - 0xfdf  :  255 - 0xff
    "10000111", -- 4064 - 0xfe0  :  135 - 0x87
    "10000111", -- 4065 - 0xfe1  :  135 - 0x87
    "10000111", -- 4066 - 0xfe2  :  135 - 0x87
    "10000111", -- 4067 - 0xfe3  :  135 - 0x87
    "10000111", -- 4068 - 0xfe4  :  135 - 0x87
    "10000111", -- 4069 - 0xfe5  :  135 - 0x87
    "10000111", -- 4070 - 0xfe6  :  135 - 0x87
    "10000111", -- 4071 - 0xfe7  :  135 - 0x87
    "11111111", -- 4072 - 0xfe8  :  255 - 0xff
    "11111111", -- 4073 - 0xfe9  :  255 - 0xff
    "11111111", -- 4074 - 0xfea  :  255 - 0xff
    "11000011", -- 4075 - 0xfeb  :  195 - 0xc3
    "11000011", -- 4076 - 0xfec  :  195 - 0xc3
    "11111111", -- 4077 - 0xfed  :  255 - 0xff
    "11111111", -- 4078 - 0xfee  :  255 - 0xff
    "11111111", -- 4079 - 0xfef  :  255 - 0xff
    "11111111", -- 4080 - 0xff0  :  255 - 0xff
    "11111111", -- 4081 - 0xff1  :  255 - 0xff
    "11100111", -- 4082 - 0xff2  :  231 - 0xe7
    "11100111", -- 4083 - 0xff3  :  231 - 0xe7
    "11100111", -- 4084 - 0xff4  :  231 - 0xe7
    "11100111", -- 4085 - 0xff5  :  231 - 0xe7
    "11111111", -- 4086 - 0xff6  :  255 - 0xff
    "11111111", -- 4087 - 0xff7  :  255 - 0xff
    "11111111", -- 4088 - 0xff8  :  255 - 0xff
    "11111111", -- 4089 - 0xff9  :  255 - 0xff
    "11111111", -- 4090 - 0xffa  :  255 - 0xff
    "11111111", -- 4091 - 0xffb  :  255 - 0xff
    "11111111", -- 4092 - 0xffc  :  255 - 0xff
    "11111111", -- 4093 - 0xffd  :  255 - 0xff
    "11111111", -- 4094 - 0xffe  :  255 - 0xff
    "11111111"  -- 4095 - 0xfff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
