//-   Sprites Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: lawnmower_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_LAWN_SPR
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table both color planes
      12'h0: dout <= 8'b11111111; //    0 : 255 - 0xff -- Sprite 0x0
      12'h1: dout <= 8'b11111111; //    1 : 255 - 0xff
      12'h2: dout <= 8'b11111111; //    2 : 255 - 0xff
      12'h3: dout <= 8'b11111111; //    3 : 255 - 0xff
      12'h4: dout <= 8'b11111111; //    4 : 255 - 0xff
      12'h5: dout <= 8'b11111111; //    5 : 255 - 0xff
      12'h6: dout <= 8'b11111111; //    6 : 255 - 0xff
      12'h7: dout <= 8'b11111111; //    7 : 255 - 0xff
      12'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- plane 1
      12'h9: dout <= 8'b00000000; //    9 :   0 - 0x0
      12'hA: dout <= 8'b00000000; //   10 :   0 - 0x0
      12'hB: dout <= 8'b00000000; //   11 :   0 - 0x0
      12'hC: dout <= 8'b00000000; //   12 :   0 - 0x0
      12'hD: dout <= 8'b00000000; //   13 :   0 - 0x0
      12'hE: dout <= 8'b00000000; //   14 :   0 - 0x0
      12'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      12'h10: dout <= 8'b11111111; //   16 : 255 - 0xff -- Sprite 0x1
      12'h11: dout <= 8'b11111111; //   17 : 255 - 0xff
      12'h12: dout <= 8'b11111111; //   18 : 255 - 0xff
      12'h13: dout <= 8'b11111111; //   19 : 255 - 0xff
      12'h14: dout <= 8'b11111111; //   20 : 255 - 0xff
      12'h15: dout <= 8'b11111111; //   21 : 255 - 0xff
      12'h16: dout <= 8'b11111100; //   22 : 252 - 0xfc
      12'h17: dout <= 8'b11111100; //   23 : 252 - 0xfc
      12'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- plane 1
      12'h19: dout <= 8'b00000000; //   25 :   0 - 0x0
      12'h1A: dout <= 8'b00000000; //   26 :   0 - 0x0
      12'h1B: dout <= 8'b00000000; //   27 :   0 - 0x0
      12'h1C: dout <= 8'b00000000; //   28 :   0 - 0x0
      12'h1D: dout <= 8'b00000111; //   29 :   7 - 0x7
      12'h1E: dout <= 8'b00000111; //   30 :   7 - 0x7
      12'h1F: dout <= 8'b00000110; //   31 :   6 - 0x6
      12'h20: dout <= 8'b11111111; //   32 : 255 - 0xff -- Sprite 0x2
      12'h21: dout <= 8'b11111111; //   33 : 255 - 0xff
      12'h22: dout <= 8'b11111111; //   34 : 255 - 0xff
      12'h23: dout <= 8'b11111111; //   35 : 255 - 0xff
      12'h24: dout <= 8'b11111111; //   36 : 255 - 0xff
      12'h25: dout <= 8'b11111111; //   37 : 255 - 0xff
      12'h26: dout <= 8'b00000000; //   38 :   0 - 0x0
      12'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout <= 8'b00000000; //   40 :   0 - 0x0 -- plane 1
      12'h29: dout <= 8'b00000000; //   41 :   0 - 0x0
      12'h2A: dout <= 8'b00000000; //   42 :   0 - 0x0
      12'h2B: dout <= 8'b00000000; //   43 :   0 - 0x0
      12'h2C: dout <= 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout <= 8'b11111111; //   45 : 255 - 0xff
      12'h2E: dout <= 8'b11111111; //   46 : 255 - 0xff
      12'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout <= 8'b11111111; //   48 : 255 - 0xff -- Sprite 0x3
      12'h31: dout <= 8'b11111111; //   49 : 255 - 0xff
      12'h32: dout <= 8'b11111111; //   50 : 255 - 0xff
      12'h33: dout <= 8'b11111111; //   51 : 255 - 0xff
      12'h34: dout <= 8'b11111111; //   52 : 255 - 0xff
      12'h35: dout <= 8'b11111111; //   53 : 255 - 0xff
      12'h36: dout <= 8'b00011111; //   54 :  31 - 0x1f
      12'h37: dout <= 8'b01000111; //   55 :  71 - 0x47
      12'h38: dout <= 8'b00000000; //   56 :   0 - 0x0 -- plane 1
      12'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      12'h3A: dout <= 8'b00000000; //   58 :   0 - 0x0
      12'h3B: dout <= 8'b00000000; //   59 :   0 - 0x0
      12'h3C: dout <= 8'b00000000; //   60 :   0 - 0x0
      12'h3D: dout <= 8'b11100000; //   61 : 224 - 0xe0
      12'h3E: dout <= 8'b11100000; //   62 : 224 - 0xe0
      12'h3F: dout <= 8'b01100000; //   63 :  96 - 0x60
      12'h40: dout <= 8'b11111111; //   64 : 255 - 0xff -- Sprite 0x4
      12'h41: dout <= 8'b11111111; //   65 : 255 - 0xff
      12'h42: dout <= 8'b11111111; //   66 : 255 - 0xff
      12'h43: dout <= 8'b11111111; //   67 : 255 - 0xff
      12'h44: dout <= 8'b11111111; //   68 : 255 - 0xff
      12'h45: dout <= 8'b11111111; //   69 : 255 - 0xff
      12'h46: dout <= 8'b11100000; //   70 : 224 - 0xe0
      12'h47: dout <= 8'b10000000; //   71 : 128 - 0x80
      12'h48: dout <= 8'b00000000; //   72 :   0 - 0x0 -- plane 1
      12'h49: dout <= 8'b00000000; //   73 :   0 - 0x0
      12'h4A: dout <= 8'b00000000; //   74 :   0 - 0x0
      12'h4B: dout <= 8'b00000000; //   75 :   0 - 0x0
      12'h4C: dout <= 8'b00000000; //   76 :   0 - 0x0
      12'h4D: dout <= 8'b00011111; //   77 :  31 - 0x1f
      12'h4E: dout <= 8'b01111111; //   78 : 127 - 0x7f
      12'h4F: dout <= 8'b11110000; //   79 : 240 - 0xf0
      12'h50: dout <= 8'b11111111; //   80 : 255 - 0xff -- Sprite 0x5
      12'h51: dout <= 8'b11111111; //   81 : 255 - 0xff
      12'h52: dout <= 8'b11111111; //   82 : 255 - 0xff
      12'h53: dout <= 8'b11111111; //   83 : 255 - 0xff
      12'h54: dout <= 8'b11111111; //   84 : 255 - 0xff
      12'h55: dout <= 8'b11110111; //   85 : 247 - 0xf7
      12'h56: dout <= 8'b00000001; //   86 :   1 - 0x1
      12'h57: dout <= 8'b00000100; //   87 :   4 - 0x4
      12'h58: dout <= 8'b00000000; //   88 :   0 - 0x0 -- plane 1
      12'h59: dout <= 8'b00000000; //   89 :   0 - 0x0
      12'h5A: dout <= 8'b00000000; //   90 :   0 - 0x0
      12'h5B: dout <= 8'b00000000; //   91 :   0 - 0x0
      12'h5C: dout <= 8'b00000000; //   92 :   0 - 0x0
      12'h5D: dout <= 8'b11111000; //   93 : 248 - 0xf8
      12'h5E: dout <= 8'b11111110; //   94 : 254 - 0xfe
      12'h5F: dout <= 8'b00001111; //   95 :  15 - 0xf
      12'h60: dout <= 8'b11111111; //   96 : 255 - 0xff -- Sprite 0x6
      12'h61: dout <= 8'b11111111; //   97 : 255 - 0xff
      12'h62: dout <= 8'b11111111; //   98 : 255 - 0xff
      12'h63: dout <= 8'b11111111; //   99 : 255 - 0xff
      12'h64: dout <= 8'b11111111; //  100 : 255 - 0xff
      12'h65: dout <= 8'b11011111; //  101 : 223 - 0xdf
      12'h66: dout <= 8'b00011100; //  102 :  28 - 0x1c
      12'h67: dout <= 8'b01000100; //  103 :  68 - 0x44
      12'h68: dout <= 8'b00000000; //  104 :   0 - 0x0 -- plane 1
      12'h69: dout <= 8'b00000000; //  105 :   0 - 0x0
      12'h6A: dout <= 8'b00000000; //  106 :   0 - 0x0
      12'h6B: dout <= 8'b00000000; //  107 :   0 - 0x0
      12'h6C: dout <= 8'b00000000; //  108 :   0 - 0x0
      12'h6D: dout <= 8'b11100111; //  109 : 231 - 0xe7
      12'h6E: dout <= 8'b11100111; //  110 : 231 - 0xe7
      12'h6F: dout <= 8'b01100110; //  111 : 102 - 0x66
      12'h70: dout <= 8'b11111111; //  112 : 255 - 0xff -- Sprite 0x7
      12'h71: dout <= 8'b11111111; //  113 : 255 - 0xff
      12'h72: dout <= 8'b11111111; //  114 : 255 - 0xff
      12'h73: dout <= 8'b11111111; //  115 : 255 - 0xff
      12'h74: dout <= 8'b11111111; //  116 : 255 - 0xff
      12'h75: dout <= 8'b10111111; //  117 : 191 - 0xbf
      12'h76: dout <= 8'b00111100; //  118 :  60 - 0x3c
      12'h77: dout <= 8'b01001100; //  119 :  76 - 0x4c
      12'h78: dout <= 8'b00000000; //  120 :   0 - 0x0 -- plane 1
      12'h79: dout <= 8'b00000000; //  121 :   0 - 0x0
      12'h7A: dout <= 8'b00000000; //  122 :   0 - 0x0
      12'h7B: dout <= 8'b00000000; //  123 :   0 - 0x0
      12'h7C: dout <= 8'b00000000; //  124 :   0 - 0x0
      12'h7D: dout <= 8'b11000111; //  125 : 199 - 0xc7
      12'h7E: dout <= 8'b11000111; //  126 : 199 - 0xc7
      12'h7F: dout <= 8'b01100110; //  127 : 102 - 0x66
      12'h80: dout <= 8'b11111100; //  128 : 252 - 0xfc -- Sprite 0x8
      12'h81: dout <= 8'b11111100; //  129 : 252 - 0xfc
      12'h82: dout <= 8'b11111100; //  130 : 252 - 0xfc
      12'h83: dout <= 8'b11111100; //  131 : 252 - 0xfc
      12'h84: dout <= 8'b11111100; //  132 : 252 - 0xfc
      12'h85: dout <= 8'b11111100; //  133 : 252 - 0xfc
      12'h86: dout <= 8'b11111100; //  134 : 252 - 0xfc
      12'h87: dout <= 8'b11111100; //  135 : 252 - 0xfc
      12'h88: dout <= 8'b00000110; //  136 :   6 - 0x6 -- plane 1
      12'h89: dout <= 8'b00000110; //  137 :   6 - 0x6
      12'h8A: dout <= 8'b00000110; //  138 :   6 - 0x6
      12'h8B: dout <= 8'b00000110; //  139 :   6 - 0x6
      12'h8C: dout <= 8'b00000110; //  140 :   6 - 0x6
      12'h8D: dout <= 8'b00000110; //  141 :   6 - 0x6
      12'h8E: dout <= 8'b00000110; //  142 :   6 - 0x6
      12'h8F: dout <= 8'b00000110; //  143 :   6 - 0x6
      12'h90: dout <= 8'b00010000; //  144 :  16 - 0x10 -- Sprite 0x9
      12'h91: dout <= 8'b00111000; //  145 :  56 - 0x38
      12'h92: dout <= 8'b01111100; //  146 : 124 - 0x7c
      12'h93: dout <= 8'b11111000; //  147 : 248 - 0xf8
      12'h94: dout <= 8'b01110000; //  148 : 112 - 0x70
      12'h95: dout <= 8'b00100010; //  149 :  34 - 0x22
      12'h96: dout <= 8'b00000101; //  150 :   5 - 0x5
      12'h97: dout <= 8'b00000010; //  151 :   2 - 0x2
      12'h98: dout <= 8'b11111111; //  152 : 255 - 0xff -- plane 1
      12'h99: dout <= 8'b11111111; //  153 : 255 - 0xff
      12'h9A: dout <= 8'b11111111; //  154 : 255 - 0xff
      12'h9B: dout <= 8'b11111111; //  155 : 255 - 0xff
      12'h9C: dout <= 8'b11111111; //  156 : 255 - 0xff
      12'h9D: dout <= 8'b11111111; //  157 : 255 - 0xff
      12'h9E: dout <= 8'b11111111; //  158 : 255 - 0xff
      12'h9F: dout <= 8'b11111111; //  159 : 255 - 0xff
      12'hA0: dout <= 8'b01000111; //  160 :  71 - 0x47 -- Sprite 0xa
      12'hA1: dout <= 8'b01000111; //  161 :  71 - 0x47
      12'hA2: dout <= 8'b01000111; //  162 :  71 - 0x47
      12'hA3: dout <= 8'b01000111; //  163 :  71 - 0x47
      12'hA4: dout <= 8'b01000111; //  164 :  71 - 0x47
      12'hA5: dout <= 8'b01000111; //  165 :  71 - 0x47
      12'hA6: dout <= 8'b01000111; //  166 :  71 - 0x47
      12'hA7: dout <= 8'b01000111; //  167 :  71 - 0x47
      12'hA8: dout <= 8'b01100000; //  168 :  96 - 0x60 -- plane 1
      12'hA9: dout <= 8'b01100000; //  169 :  96 - 0x60
      12'hAA: dout <= 8'b01100000; //  170 :  96 - 0x60
      12'hAB: dout <= 8'b01100000; //  171 :  96 - 0x60
      12'hAC: dout <= 8'b01100000; //  172 :  96 - 0x60
      12'hAD: dout <= 8'b01100000; //  173 :  96 - 0x60
      12'hAE: dout <= 8'b01100000; //  174 :  96 - 0x60
      12'hAF: dout <= 8'b01100000; //  175 :  96 - 0x60
      12'hB0: dout <= 8'b11111111; //  176 : 255 - 0xff -- Sprite 0xb
      12'hB1: dout <= 8'b11111110; //  177 : 254 - 0xfe
      12'hB2: dout <= 8'b11111110; //  178 : 254 - 0xfe
      12'hB3: dout <= 8'b11111100; //  179 : 252 - 0xfc
      12'hB4: dout <= 8'b11111100; //  180 : 252 - 0xfc
      12'hB5: dout <= 8'b11111100; //  181 : 252 - 0xfc
      12'hB6: dout <= 8'b11111100; //  182 : 252 - 0xfc
      12'hB7: dout <= 8'b11111100; //  183 : 252 - 0xfc
      12'hB8: dout <= 8'b00000001; //  184 :   1 - 0x1 -- plane 1
      12'hB9: dout <= 8'b00000011; //  185 :   3 - 0x3
      12'hBA: dout <= 8'b00000011; //  186 :   3 - 0x3
      12'hBB: dout <= 8'b00000111; //  187 :   7 - 0x7
      12'hBC: dout <= 8'b00000110; //  188 :   6 - 0x6
      12'hBD: dout <= 8'b00000110; //  189 :   6 - 0x6
      12'hBE: dout <= 8'b00000110; //  190 :   6 - 0x6
      12'hBF: dout <= 8'b00000110; //  191 :   6 - 0x6
      12'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0xc
      12'hC1: dout <= 8'b00001000; //  193 :   8 - 0x8
      12'hC2: dout <= 8'b00011100; //  194 :  28 - 0x1c
      12'hC3: dout <= 8'b00111000; //  195 :  56 - 0x38
      12'hC4: dout <= 8'b01110000; //  196 : 112 - 0x70
      12'hC5: dout <= 8'b00100010; //  197 :  34 - 0x22
      12'hC6: dout <= 8'b00000101; //  198 :   5 - 0x5
      12'hC7: dout <= 8'b00000010; //  199 :   2 - 0x2
      12'hC8: dout <= 8'b11000111; //  200 : 199 - 0xc7 -- plane 1
      12'hC9: dout <= 8'b10011111; //  201 : 159 - 0x9f
      12'hCA: dout <= 8'b00111111; //  202 :  63 - 0x3f
      12'hCB: dout <= 8'b01111111; //  203 : 127 - 0x7f
      12'hCC: dout <= 8'b01111111; //  204 : 127 - 0x7f
      12'hCD: dout <= 8'b11111111; //  205 : 255 - 0xff
      12'hCE: dout <= 8'b11111111; //  206 : 255 - 0xff
      12'hCF: dout <= 8'b11111111; //  207 : 255 - 0xff
      12'hD0: dout <= 8'b00000010; //  208 :   2 - 0x2 -- Sprite 0xd
      12'hD1: dout <= 8'b00110001; //  209 :  49 - 0x31
      12'hD2: dout <= 8'b01111000; //  210 : 120 - 0x78
      12'hD3: dout <= 8'b11111000; //  211 : 248 - 0xf8
      12'hD4: dout <= 8'b01110000; //  212 : 112 - 0x70
      12'hD5: dout <= 8'b00100010; //  213 :  34 - 0x22
      12'hD6: dout <= 8'b00000101; //  214 :   5 - 0x5
      12'hD7: dout <= 8'b00000010; //  215 :   2 - 0x2
      12'hD8: dout <= 8'b11100011; //  216 : 227 - 0xe3 -- plane 1
      12'hD9: dout <= 8'b11111001; //  217 : 249 - 0xf9
      12'hDA: dout <= 8'b11111100; //  218 : 252 - 0xfc
      12'hDB: dout <= 8'b11111110; //  219 : 254 - 0xfe
      12'hDC: dout <= 8'b11111110; //  220 : 254 - 0xfe
      12'hDD: dout <= 8'b11111111; //  221 : 255 - 0xff
      12'hDE: dout <= 8'b11111111; //  222 : 255 - 0xff
      12'hDF: dout <= 8'b11111111; //  223 : 255 - 0xff
      12'hE0: dout <= 8'b01111100; //  224 : 124 - 0x7c -- Sprite 0xe
      12'hE1: dout <= 8'b00111100; //  225 :  60 - 0x3c
      12'hE2: dout <= 8'b10011100; //  226 : 156 - 0x9c
      12'hE3: dout <= 8'b10001100; //  227 : 140 - 0x8c
      12'hE4: dout <= 8'b01001100; //  228 :  76 - 0x4c
      12'hE5: dout <= 8'b01000100; //  229 :  68 - 0x44
      12'hE6: dout <= 8'b01000100; //  230 :  68 - 0x44
      12'hE7: dout <= 8'b01000100; //  231 :  68 - 0x44
      12'hE8: dout <= 8'b10000110; //  232 : 134 - 0x86 -- plane 1
      12'hE9: dout <= 8'b11000110; //  233 : 198 - 0xc6
      12'hEA: dout <= 8'b11000110; //  234 : 198 - 0xc6
      12'hEB: dout <= 8'b11100110; //  235 : 230 - 0xe6
      12'hEC: dout <= 8'b01100110; //  236 : 102 - 0x66
      12'hED: dout <= 8'b01100110; //  237 : 102 - 0x66
      12'hEE: dout <= 8'b01100110; //  238 : 102 - 0x66
      12'hEF: dout <= 8'b01100110; //  239 : 102 - 0x66
      12'hF0: dout <= 8'b01000100; //  240 :  68 - 0x44 -- Sprite 0xf
      12'hF1: dout <= 8'b01000100; //  241 :  68 - 0x44
      12'hF2: dout <= 8'b01000100; //  242 :  68 - 0x44
      12'hF3: dout <= 8'b01000100; //  243 :  68 - 0x44
      12'hF4: dout <= 8'b01000100; //  244 :  68 - 0x44
      12'hF5: dout <= 8'b01000100; //  245 :  68 - 0x44
      12'hF6: dout <= 8'b01000100; //  246 :  68 - 0x44
      12'hF7: dout <= 8'b01000100; //  247 :  68 - 0x44
      12'hF8: dout <= 8'b01100110; //  248 : 102 - 0x66 -- plane 1
      12'hF9: dout <= 8'b01100110; //  249 : 102 - 0x66
      12'hFA: dout <= 8'b01100110; //  250 : 102 - 0x66
      12'hFB: dout <= 8'b01100110; //  251 : 102 - 0x66
      12'hFC: dout <= 8'b01100110; //  252 : 102 - 0x66
      12'hFD: dout <= 8'b01100110; //  253 : 102 - 0x66
      12'hFE: dout <= 8'b01100110; //  254 : 102 - 0x66
      12'hFF: dout <= 8'b01100110; //  255 : 102 - 0x66
      12'h100: dout <= 8'b01001100; //  256 :  76 - 0x4c -- Sprite 0x10
      12'h101: dout <= 8'b00100100; //  257 :  36 - 0x24
      12'h102: dout <= 8'b00100100; //  258 :  36 - 0x24
      12'h103: dout <= 8'b10010100; //  259 : 148 - 0x94
      12'h104: dout <= 8'b00010000; //  260 :  16 - 0x10
      12'h105: dout <= 8'b00001000; //  261 :   8 - 0x8
      12'h106: dout <= 8'b00001000; //  262 :   8 - 0x8
      12'h107: dout <= 8'b00000100; //  263 :   4 - 0x4
      12'h108: dout <= 8'b01100110; //  264 : 102 - 0x66 -- plane 1
      12'h109: dout <= 8'b00110110; //  265 :  54 - 0x36
      12'h10A: dout <= 8'b10110110; //  266 : 182 - 0xb6
      12'h10B: dout <= 8'b10011110; //  267 : 158 - 0x9e
      12'h10C: dout <= 8'b11011110; //  268 : 222 - 0xde
      12'h10D: dout <= 8'b11001110; //  269 : 206 - 0xce
      12'h10E: dout <= 8'b11101110; //  270 : 238 - 0xee
      12'h10F: dout <= 8'b11100110; //  271 : 230 - 0xe6
      12'h110: dout <= 8'b00000000; //  272 :   0 - 0x0 -- Sprite 0x11
      12'h111: dout <= 8'b00111100; //  273 :  60 - 0x3c
      12'h112: dout <= 8'b01000000; //  274 :  64 - 0x40
      12'h113: dout <= 8'b01000100; //  275 :  68 - 0x44
      12'h114: dout <= 8'b01000100; //  276 :  68 - 0x44
      12'h115: dout <= 8'b01000100; //  277 :  68 - 0x44
      12'h116: dout <= 8'b01000100; //  278 :  68 - 0x44
      12'h117: dout <= 8'b01000100; //  279 :  68 - 0x44
      12'h118: dout <= 8'b10000001; //  280 : 129 - 0x81 -- plane 1
      12'h119: dout <= 8'b00111100; //  281 :  60 - 0x3c
      12'h11A: dout <= 8'b01111110; //  282 : 126 - 0x7e
      12'h11B: dout <= 8'b01100110; //  283 : 102 - 0x66
      12'h11C: dout <= 8'b01100110; //  284 : 102 - 0x66
      12'h11D: dout <= 8'b01100110; //  285 : 102 - 0x66
      12'h11E: dout <= 8'b01100110; //  286 : 102 - 0x66
      12'h11F: dout <= 8'b01100110; //  287 : 102 - 0x66
      12'h120: dout <= 8'b00000100; //  288 :   4 - 0x4 -- Sprite 0x12
      12'h121: dout <= 8'b00010010; //  289 :  18 - 0x12
      12'h122: dout <= 8'b00110010; //  290 :  50 - 0x32
      12'h123: dout <= 8'b01111000; //  291 : 120 - 0x78
      12'h124: dout <= 8'b11111000; //  292 : 248 - 0xf8
      12'h125: dout <= 8'b01110000; //  293 : 112 - 0x70
      12'h126: dout <= 8'b00100100; //  294 :  36 - 0x24
      12'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout <= 8'b11110110; //  296 : 246 - 0xf6 -- plane 1
      12'h129: dout <= 8'b11110010; //  297 : 242 - 0xf2
      12'h12A: dout <= 8'b11111010; //  298 : 250 - 0xfa
      12'h12B: dout <= 8'b11111000; //  299 : 248 - 0xf8
      12'h12C: dout <= 8'b11111100; //  300 : 252 - 0xfc
      12'h12D: dout <= 8'b11111100; //  301 : 252 - 0xfc
      12'h12E: dout <= 8'b11111110; //  302 : 254 - 0xfe
      12'h12F: dout <= 8'b11111110; //  303 : 254 - 0xfe
      12'h130: dout <= 8'b01000100; //  304 :  68 - 0x44 -- Sprite 0x13
      12'h131: dout <= 8'b01000100; //  305 :  68 - 0x44
      12'h132: dout <= 8'b01000100; //  306 :  68 - 0x44
      12'h133: dout <= 8'b01000100; //  307 :  68 - 0x44
      12'h134: dout <= 8'b01000100; //  308 :  68 - 0x44
      12'h135: dout <= 8'b01000100; //  309 :  68 - 0x44
      12'h136: dout <= 8'b01000100; //  310 :  68 - 0x44
      12'h137: dout <= 8'b01011100; //  311 :  92 - 0x5c
      12'h138: dout <= 8'b01100110; //  312 : 102 - 0x66 -- plane 1
      12'h139: dout <= 8'b01100110; //  313 : 102 - 0x66
      12'h13A: dout <= 8'b01100110; //  314 : 102 - 0x66
      12'h13B: dout <= 8'b01100110; //  315 : 102 - 0x66
      12'h13C: dout <= 8'b01100110; //  316 : 102 - 0x66
      12'h13D: dout <= 8'b01100110; //  317 : 102 - 0x66
      12'h13E: dout <= 8'b01100110; //  318 : 102 - 0x66
      12'h13F: dout <= 8'b01111110; //  319 : 126 - 0x7e
      12'h140: dout <= 8'b00010000; //  320 :  16 - 0x10 -- Sprite 0x14
      12'h141: dout <= 8'b00111000; //  321 :  56 - 0x38
      12'h142: dout <= 8'b00111100; //  322 :  60 - 0x3c
      12'h143: dout <= 8'b00111000; //  323 :  56 - 0x38
      12'h144: dout <= 8'b00010000; //  324 :  16 - 0x10
      12'h145: dout <= 8'b00000010; //  325 :   2 - 0x2
      12'h146: dout <= 8'b01000101; //  326 :  69 - 0x45
      12'h147: dout <= 8'b01000010; //  327 :  66 - 0x42
      12'h148: dout <= 8'b11111111; //  328 : 255 - 0xff -- plane 1
      12'h149: dout <= 8'b01111111; //  329 : 127 - 0x7f
      12'h14A: dout <= 8'b01111111; //  330 : 127 - 0x7f
      12'h14B: dout <= 8'b00111111; //  331 :  63 - 0x3f
      12'h14C: dout <= 8'b00111111; //  332 :  63 - 0x3f
      12'h14D: dout <= 8'b00011111; //  333 :  31 - 0x1f
      12'h14E: dout <= 8'b01011111; //  334 :  95 - 0x5f
      12'h14F: dout <= 8'b01001111; //  335 :  79 - 0x4f
      12'h150: dout <= 8'b01000100; //  336 :  68 - 0x44 -- Sprite 0x15
      12'h151: dout <= 8'b01000100; //  337 :  68 - 0x44
      12'h152: dout <= 8'b01000100; //  338 :  68 - 0x44
      12'h153: dout <= 8'b01000100; //  339 :  68 - 0x44
      12'h154: dout <= 8'b01000100; //  340 :  68 - 0x44
      12'h155: dout <= 8'b01011100; //  341 :  92 - 0x5c
      12'h156: dout <= 8'b01000000; //  342 :  64 - 0x40
      12'h157: dout <= 8'b00000000; //  343 :   0 - 0x0
      12'h158: dout <= 8'b01100110; //  344 : 102 - 0x66 -- plane 1
      12'h159: dout <= 8'b01100110; //  345 : 102 - 0x66
      12'h15A: dout <= 8'b01100110; //  346 : 102 - 0x66
      12'h15B: dout <= 8'b01100110; //  347 : 102 - 0x66
      12'h15C: dout <= 8'b01100110; //  348 : 102 - 0x66
      12'h15D: dout <= 8'b01111110; //  349 : 126 - 0x7e
      12'h15E: dout <= 8'b01111110; //  350 : 126 - 0x7e
      12'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout <= 8'b01000000; //  352 :  64 - 0x40 -- Sprite 0x16
      12'h161: dout <= 8'b01000000; //  353 :  64 - 0x40
      12'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      12'h163: dout <= 8'b00000000; //  355 :   0 - 0x0
      12'h164: dout <= 8'b00011000; //  356 :  24 - 0x18
      12'h165: dout <= 8'b00111000; //  357 :  56 - 0x38
      12'h166: dout <= 8'b00010000; //  358 :  16 - 0x10
      12'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout <= 8'b01111110; //  360 : 126 - 0x7e -- plane 1
      12'h169: dout <= 8'b01100110; //  361 : 102 - 0x66
      12'h16A: dout <= 8'b01000010; //  362 :  66 - 0x42
      12'h16B: dout <= 8'b00011000; //  363 :  24 - 0x18
      12'h16C: dout <= 8'b00111100; //  364 :  60 - 0x3c
      12'h16D: dout <= 8'b01111110; //  365 : 126 - 0x7e
      12'h16E: dout <= 8'b11111111; //  366 : 255 - 0xff
      12'h16F: dout <= 8'b11111111; //  367 : 255 - 0xff
      12'h170: dout <= 8'b01000000; //  368 :  64 - 0x40 -- Sprite 0x17
      12'h171: dout <= 8'b01000000; //  369 :  64 - 0x40
      12'h172: dout <= 8'b01000000; //  370 :  64 - 0x40
      12'h173: dout <= 8'b01000000; //  371 :  64 - 0x40
      12'h174: dout <= 8'b01010000; //  372 :  80 - 0x50
      12'h175: dout <= 8'b01010000; //  373 :  80 - 0x50
      12'h176: dout <= 8'b01001000; //  374 :  72 - 0x48
      12'h177: dout <= 8'b01001000; //  375 :  72 - 0x48
      12'h178: dout <= 8'b01101111; //  376 : 111 - 0x6f -- plane 1
      12'h179: dout <= 8'b01100111; //  377 : 103 - 0x67
      12'h17A: dout <= 8'b01110111; //  378 : 119 - 0x77
      12'h17B: dout <= 8'b01110011; //  379 : 115 - 0x73
      12'h17C: dout <= 8'b01111011; //  380 : 123 - 0x7b
      12'h17D: dout <= 8'b01111001; //  381 : 121 - 0x79
      12'h17E: dout <= 8'b01101101; //  382 : 109 - 0x6d
      12'h17F: dout <= 8'b01101100; //  383 : 108 - 0x6c
      12'h180: dout <= 8'b01000111; //  384 :  71 - 0x47 -- Sprite 0x18
      12'h181: dout <= 8'b01000111; //  385 :  71 - 0x47
      12'h182: dout <= 8'b01000111; //  386 :  71 - 0x47
      12'h183: dout <= 8'b01000111; //  387 :  71 - 0x47
      12'h184: dout <= 8'b01000111; //  388 :  71 - 0x47
      12'h185: dout <= 8'b01011111; //  389 :  95 - 0x5f
      12'h186: dout <= 8'b00000000; //  390 :   0 - 0x0
      12'h187: dout <= 8'b00000000; //  391 :   0 - 0x0
      12'h188: dout <= 8'b01100000; //  392 :  96 - 0x60 -- plane 1
      12'h189: dout <= 8'b01100000; //  393 :  96 - 0x60
      12'h18A: dout <= 8'b01100000; //  394 :  96 - 0x60
      12'h18B: dout <= 8'b01100000; //  395 :  96 - 0x60
      12'h18C: dout <= 8'b01100000; //  396 :  96 - 0x60
      12'h18D: dout <= 8'b01111111; //  397 : 127 - 0x7f
      12'h18E: dout <= 8'b01111111; //  398 : 127 - 0x7f
      12'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      12'h190: dout <= 8'b11111100; //  400 : 252 - 0xfc -- Sprite 0x19
      12'h191: dout <= 8'b11111100; //  401 : 252 - 0xfc
      12'h192: dout <= 8'b11111100; //  402 : 252 - 0xfc
      12'h193: dout <= 8'b11111100; //  403 : 252 - 0xfc
      12'h194: dout <= 8'b11111100; //  404 : 252 - 0xfc
      12'h195: dout <= 8'b11011100; //  405 : 220 - 0xdc
      12'h196: dout <= 8'b00011100; //  406 :  28 - 0x1c
      12'h197: dout <= 8'b01000100; //  407 :  68 - 0x44
      12'h198: dout <= 8'b00000110; //  408 :   6 - 0x6 -- plane 1
      12'h199: dout <= 8'b00000110; //  409 :   6 - 0x6
      12'h19A: dout <= 8'b00000110; //  410 :   6 - 0x6
      12'h19B: dout <= 8'b00000110; //  411 :   6 - 0x6
      12'h19C: dout <= 8'b00000110; //  412 :   6 - 0x6
      12'h19D: dout <= 8'b11100110; //  413 : 230 - 0xe6
      12'h19E: dout <= 8'b11100110; //  414 : 230 - 0xe6
      12'h19F: dout <= 8'b01100110; //  415 : 102 - 0x66
      12'h1A0: dout <= 8'b00010000; //  416 :  16 - 0x10 -- Sprite 0x1a
      12'h1A1: dout <= 8'b00111000; //  417 :  56 - 0x38
      12'h1A2: dout <= 8'b01111100; //  418 : 124 - 0x7c
      12'h1A3: dout <= 8'b11100000; //  419 : 224 - 0xe0
      12'h1A4: dout <= 8'b01000000; //  420 :  64 - 0x40
      12'h1A5: dout <= 8'b00000000; //  421 :   0 - 0x0
      12'h1A6: dout <= 8'b00010000; //  422 :  16 - 0x10
      12'h1A7: dout <= 8'b00100000; //  423 :  32 - 0x20
      12'h1A8: dout <= 8'b11111111; //  424 : 255 - 0xff -- plane 1
      12'h1A9: dout <= 8'b11111111; //  425 : 255 - 0xff
      12'h1AA: dout <= 8'b11111111; //  426 : 255 - 0xff
      12'h1AB: dout <= 8'b11111111; //  427 : 255 - 0xff
      12'h1AC: dout <= 8'b11100111; //  428 : 231 - 0xe7
      12'h1AD: dout <= 8'b11000011; //  429 : 195 - 0xc3
      12'h1AE: dout <= 8'b10011001; //  430 : 153 - 0x99
      12'h1AF: dout <= 8'b00111100; //  431 :  60 - 0x3c
      12'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x1b
      12'h1B1: dout <= 8'b01111100; //  433 : 124 - 0x7c
      12'h1B2: dout <= 8'b01000000; //  434 :  64 - 0x40
      12'h1B3: dout <= 8'b01000100; //  435 :  68 - 0x44
      12'h1B4: dout <= 8'b01000100; //  436 :  68 - 0x44
      12'h1B5: dout <= 8'b01000100; //  437 :  68 - 0x44
      12'h1B6: dout <= 8'b01000100; //  438 :  68 - 0x44
      12'h1B7: dout <= 8'b01000100; //  439 :  68 - 0x44
      12'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0 -- plane 1
      12'h1B9: dout <= 8'b01111110; //  441 : 126 - 0x7e
      12'h1BA: dout <= 8'b01111110; //  442 : 126 - 0x7e
      12'h1BB: dout <= 8'b01100110; //  443 : 102 - 0x66
      12'h1BC: dout <= 8'b01100110; //  444 : 102 - 0x66
      12'h1BD: dout <= 8'b01100110; //  445 : 102 - 0x66
      12'h1BE: dout <= 8'b01100110; //  446 : 102 - 0x66
      12'h1BF: dout <= 8'b01100110; //  447 : 102 - 0x66
      12'h1C0: dout <= 8'b00010000; //  448 :  16 - 0x10 -- Sprite 0x1c
      12'h1C1: dout <= 8'b00111000; //  449 :  56 - 0x38
      12'h1C2: dout <= 8'b01110001; //  450 : 113 - 0x71
      12'h1C3: dout <= 8'b11100010; //  451 : 226 - 0xe2
      12'h1C4: dout <= 8'b01000100; //  452 :  68 - 0x44
      12'h1C5: dout <= 8'b00001000; //  453 :   8 - 0x8
      12'h1C6: dout <= 8'b00010000; //  454 :  16 - 0x10
      12'h1C7: dout <= 8'b00100000; //  455 :  32 - 0x20
      12'h1C8: dout <= 8'b11111110; //  456 : 254 - 0xfe -- plane 1
      12'h1C9: dout <= 8'b11111100; //  457 : 252 - 0xfc
      12'h1CA: dout <= 8'b11111001; //  458 : 249 - 0xf9
      12'h1CB: dout <= 8'b11110011; //  459 : 243 - 0xf3
      12'h1CC: dout <= 8'b11100111; //  460 : 231 - 0xe7
      12'h1CD: dout <= 8'b11001110; //  461 : 206 - 0xce
      12'h1CE: dout <= 8'b10011100; //  462 : 156 - 0x9c
      12'h1CF: dout <= 8'b00111000; //  463 :  56 - 0x38
      12'h1D0: dout <= 8'b01000000; //  464 :  64 - 0x40 -- Sprite 0x1d
      12'h1D1: dout <= 8'b10000100; //  465 : 132 - 0x84
      12'h1D2: dout <= 8'b00000010; //  466 :   2 - 0x2
      12'h1D3: dout <= 8'b00000111; //  467 :   7 - 0x7
      12'h1D4: dout <= 8'b00001111; //  468 :  15 - 0xf
      12'h1D5: dout <= 8'b00011111; //  469 :  31 - 0x1f
      12'h1D6: dout <= 8'b00111111; //  470 :  63 - 0x3f
      12'h1D7: dout <= 8'b01111111; //  471 : 127 - 0x7f
      12'h1D8: dout <= 8'b01111110; //  472 : 126 - 0x7e -- plane 1
      12'h1D9: dout <= 8'b11100111; //  473 : 231 - 0xe7
      12'h1DA: dout <= 8'b11000011; //  474 : 195 - 0xc3
      12'h1DB: dout <= 8'b10000001; //  475 : 129 - 0x81
      12'h1DC: dout <= 8'b00000000; //  476 :   0 - 0x0
      12'h1DD: dout <= 8'b00000000; //  477 :   0 - 0x0
      12'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b00010000; //  480 :  16 - 0x10 -- Sprite 0x1e
      12'h1E1: dout <= 8'b00011000; //  481 :  24 - 0x18
      12'h1E2: dout <= 8'b00001100; //  482 :  12 - 0xc
      12'h1E3: dout <= 8'b00000110; //  483 :   6 - 0x6
      12'h1E4: dout <= 8'b10000000; //  484 : 128 - 0x80
      12'h1E5: dout <= 8'b11000000; //  485 : 192 - 0xc0
      12'h1E6: dout <= 8'b11100000; //  486 : 224 - 0xe0
      12'h1E7: dout <= 8'b11110000; //  487 : 240 - 0xf0
      12'h1E8: dout <= 8'b01111111; //  488 : 127 - 0x7f -- plane 1
      12'h1E9: dout <= 8'b00111111; //  489 :  63 - 0x3f
      12'h1EA: dout <= 8'b10011111; //  490 : 159 - 0x9f
      12'h1EB: dout <= 8'b11001111; //  491 : 207 - 0xcf
      12'h1EC: dout <= 8'b11100111; //  492 : 231 - 0xe7
      12'h1ED: dout <= 8'b01110011; //  493 : 115 - 0x73
      12'h1EE: dout <= 8'b00111001; //  494 :  57 - 0x39
      12'h1EF: dout <= 8'b00011100; //  495 :  28 - 0x1c
      12'h1F0: dout <= 8'b11111100; //  496 : 252 - 0xfc -- Sprite 0x1f
      12'h1F1: dout <= 8'b11111101; //  497 : 253 - 0xfd
      12'h1F2: dout <= 8'b11111100; //  498 : 252 - 0xfc
      12'h1F3: dout <= 8'b11111110; //  499 : 254 - 0xfe
      12'h1F4: dout <= 8'b11111110; //  500 : 254 - 0xfe
      12'h1F5: dout <= 8'b11111111; //  501 : 255 - 0xff
      12'h1F6: dout <= 8'b11111111; //  502 : 255 - 0xff
      12'h1F7: dout <= 8'b11111111; //  503 : 255 - 0xff
      12'h1F8: dout <= 8'b00000110; //  504 :   6 - 0x6 -- plane 1
      12'h1F9: dout <= 8'b00000111; //  505 :   7 - 0x7
      12'h1FA: dout <= 8'b00000111; //  506 :   7 - 0x7
      12'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      12'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      12'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      12'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout <= 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x20
      12'h201: dout <= 8'b11111111; //  513 : 255 - 0xff
      12'h202: dout <= 8'b00000000; //  514 :   0 - 0x0
      12'h203: dout <= 8'b00000000; //  515 :   0 - 0x0
      12'h204: dout <= 8'b00000000; //  516 :   0 - 0x0
      12'h205: dout <= 8'b11111111; //  517 : 255 - 0xff
      12'h206: dout <= 8'b11111111; //  518 : 255 - 0xff
      12'h207: dout <= 8'b11111111; //  519 : 255 - 0xff
      12'h208: dout <= 8'b00000000; //  520 :   0 - 0x0 -- plane 1
      12'h209: dout <= 8'b11111111; //  521 : 255 - 0xff
      12'h20A: dout <= 8'b11111111; //  522 : 255 - 0xff
      12'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      12'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      12'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      12'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      12'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout <= 8'b01000100; //  528 :  68 - 0x44 -- Sprite 0x21
      12'h211: dout <= 8'b11000101; //  529 : 197 - 0xc5
      12'h212: dout <= 8'b00000000; //  530 :   0 - 0x0
      12'h213: dout <= 8'b00000110; //  531 :   6 - 0x6
      12'h214: dout <= 8'b00000110; //  532 :   6 - 0x6
      12'h215: dout <= 8'b11111111; //  533 : 255 - 0xff
      12'h216: dout <= 8'b11111111; //  534 : 255 - 0xff
      12'h217: dout <= 8'b11111111; //  535 : 255 - 0xff
      12'h218: dout <= 8'b01100110; //  536 : 102 - 0x66 -- plane 1
      12'h219: dout <= 8'b11100111; //  537 : 231 - 0xe7
      12'h21A: dout <= 8'b11100111; //  538 : 231 - 0xe7
      12'h21B: dout <= 8'b00000000; //  539 :   0 - 0x0
      12'h21C: dout <= 8'b00000000; //  540 :   0 - 0x0
      12'h21D: dout <= 8'b00000000; //  541 :   0 - 0x0
      12'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      12'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout <= 8'b01000000; //  544 :  64 - 0x40 -- Sprite 0x22
      12'h221: dout <= 8'b10000001; //  545 : 129 - 0x81
      12'h222: dout <= 8'b00000011; //  546 :   3 - 0x3
      12'h223: dout <= 8'b00000111; //  547 :   7 - 0x7
      12'h224: dout <= 8'b00001111; //  548 :  15 - 0xf
      12'h225: dout <= 8'b11111111; //  549 : 255 - 0xff
      12'h226: dout <= 8'b11111111; //  550 : 255 - 0xff
      12'h227: dout <= 8'b11111111; //  551 : 255 - 0xff
      12'h228: dout <= 8'b01110000; //  552 : 112 - 0x70 -- plane 1
      12'h229: dout <= 8'b11100000; //  553 : 224 - 0xe0
      12'h22A: dout <= 8'b11000000; //  554 : 192 - 0xc0
      12'h22B: dout <= 8'b00000000; //  555 :   0 - 0x0
      12'h22C: dout <= 8'b00000000; //  556 :   0 - 0x0
      12'h22D: dout <= 8'b00000000; //  557 :   0 - 0x0
      12'h22E: dout <= 8'b00000000; //  558 :   0 - 0x0
      12'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout <= 8'b11111000; //  560 : 248 - 0xf8 -- Sprite 0x23
      12'h231: dout <= 8'b11111100; //  561 : 252 - 0xfc
      12'h232: dout <= 8'b11111110; //  562 : 254 - 0xfe
      12'h233: dout <= 8'b11111110; //  563 : 254 - 0xfe
      12'h234: dout <= 8'b11111111; //  564 : 255 - 0xff
      12'h235: dout <= 8'b11111111; //  565 : 255 - 0xff
      12'h236: dout <= 8'b11111111; //  566 : 255 - 0xff
      12'h237: dout <= 8'b11111111; //  567 : 255 - 0xff
      12'h238: dout <= 8'b00001110; //  568 :  14 - 0xe -- plane 1
      12'h239: dout <= 8'b00000111; //  569 :   7 - 0x7
      12'h23A: dout <= 8'b00000011; //  570 :   3 - 0x3
      12'h23B: dout <= 8'b00000000; //  571 :   0 - 0x0
      12'h23C: dout <= 8'b00000000; //  572 :   0 - 0x0
      12'h23D: dout <= 8'b00000000; //  573 :   0 - 0x0
      12'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout <= 8'b01000111; //  576 :  71 - 0x47 -- Sprite 0x24
      12'h241: dout <= 8'b11000111; //  577 : 199 - 0xc7
      12'h242: dout <= 8'b00000111; //  578 :   7 - 0x7
      12'h243: dout <= 8'b00000111; //  579 :   7 - 0x7
      12'h244: dout <= 8'b00000111; //  580 :   7 - 0x7
      12'h245: dout <= 8'b11111111; //  581 : 255 - 0xff
      12'h246: dout <= 8'b11111111; //  582 : 255 - 0xff
      12'h247: dout <= 8'b11111111; //  583 : 255 - 0xff
      12'h248: dout <= 8'b01100000; //  584 :  96 - 0x60 -- plane 1
      12'h249: dout <= 8'b11100000; //  585 : 224 - 0xe0
      12'h24A: dout <= 8'b11100000; //  586 : 224 - 0xe0
      12'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      12'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      12'h24D: dout <= 8'b00000000; //  589 :   0 - 0x0
      12'h24E: dout <= 8'b00000000; //  590 :   0 - 0x0
      12'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout <= 8'b11111111; //  592 : 255 - 0xff -- Sprite 0x25
      12'h251: dout <= 8'b11111111; //  593 : 255 - 0xff
      12'h252: dout <= 8'b11111111; //  594 : 255 - 0xff
      12'h253: dout <= 8'b11111111; //  595 : 255 - 0xff
      12'h254: dout <= 8'b11111111; //  596 : 255 - 0xff
      12'h255: dout <= 8'b11111111; //  597 : 255 - 0xff
      12'h256: dout <= 8'b00011111; //  598 :  31 - 0x1f
      12'h257: dout <= 8'b00001111; //  599 :  15 - 0xf
      12'h258: dout <= 8'b00000000; //  600 :   0 - 0x0 -- plane 1
      12'h259: dout <= 8'b00000000; //  601 :   0 - 0x0
      12'h25A: dout <= 8'b00000000; //  602 :   0 - 0x0
      12'h25B: dout <= 8'b00000000; //  603 :   0 - 0x0
      12'h25C: dout <= 8'b00000000; //  604 :   0 - 0x0
      12'h25D: dout <= 8'b11000000; //  605 : 192 - 0xc0
      12'h25E: dout <= 8'b11100000; //  606 : 224 - 0xe0
      12'h25F: dout <= 8'b01110000; //  607 : 112 - 0x70
      12'h260: dout <= 8'b11111111; //  608 : 255 - 0xff -- Sprite 0x26
      12'h261: dout <= 8'b11111111; //  609 : 255 - 0xff
      12'h262: dout <= 8'b11111111; //  610 : 255 - 0xff
      12'h263: dout <= 8'b11111111; //  611 : 255 - 0xff
      12'h264: dout <= 8'b11111111; //  612 : 255 - 0xff
      12'h265: dout <= 8'b11111111; //  613 : 255 - 0xff
      12'h266: dout <= 8'b11111100; //  614 : 252 - 0xfc
      12'h267: dout <= 8'b11111000; //  615 : 248 - 0xf8
      12'h268: dout <= 8'b00000000; //  616 :   0 - 0x0 -- plane 1
      12'h269: dout <= 8'b00000000; //  617 :   0 - 0x0
      12'h26A: dout <= 8'b00000000; //  618 :   0 - 0x0
      12'h26B: dout <= 8'b00000000; //  619 :   0 - 0x0
      12'h26C: dout <= 8'b00000000; //  620 :   0 - 0x0
      12'h26D: dout <= 8'b00000011; //  621 :   3 - 0x3
      12'h26E: dout <= 8'b00000111; //  622 :   7 - 0x7
      12'h26F: dout <= 8'b00001110; //  623 :  14 - 0xe
      12'h270: dout <= 8'b00100111; //  624 :  39 - 0x27 -- Sprite 0x27
      12'h271: dout <= 8'b00010011; //  625 :  19 - 0x13
      12'h272: dout <= 8'b00001001; //  626 :   9 - 0x9
      12'h273: dout <= 8'b11000100; //  627 : 196 - 0xc4
      12'h274: dout <= 8'b01100010; //  628 :  98 - 0x62
      12'h275: dout <= 8'b00100001; //  629 :  33 - 0x21
      12'h276: dout <= 8'b00000000; //  630 :   0 - 0x0
      12'h277: dout <= 8'b00000000; //  631 :   0 - 0x0
      12'h278: dout <= 8'b00111000; //  632 :  56 - 0x38 -- plane 1
      12'h279: dout <= 8'b10011100; //  633 : 156 - 0x9c
      12'h27A: dout <= 8'b11001110; //  634 : 206 - 0xce
      12'h27B: dout <= 8'b11100111; //  635 : 231 - 0xe7
      12'h27C: dout <= 8'b11110011; //  636 : 243 - 0xf3
      12'h27D: dout <= 8'b11111001; //  637 : 249 - 0xf9
      12'h27E: dout <= 8'b11111100; //  638 : 252 - 0xfc
      12'h27F: dout <= 8'b11111110; //  639 : 254 - 0xfe
      12'h280: dout <= 8'b11111111; //  640 : 255 - 0xff -- Sprite 0x28
      12'h281: dout <= 8'b11111111; //  641 : 255 - 0xff
      12'h282: dout <= 8'b11111111; //  642 : 255 - 0xff
      12'h283: dout <= 8'b11111111; //  643 : 255 - 0xff
      12'h284: dout <= 8'b01111111; //  644 : 127 - 0x7f
      12'h285: dout <= 8'b00111110; //  645 :  62 - 0x3e
      12'h286: dout <= 8'b10011100; //  646 : 156 - 0x9c
      12'h287: dout <= 8'b01001000; //  647 :  72 - 0x48
      12'h288: dout <= 8'b00000000; //  648 :   0 - 0x0 -- plane 1
      12'h289: dout <= 8'b00000000; //  649 :   0 - 0x0
      12'h28A: dout <= 8'b00000000; //  650 :   0 - 0x0
      12'h28B: dout <= 8'b00000000; //  651 :   0 - 0x0
      12'h28C: dout <= 8'b10000001; //  652 : 129 - 0x81
      12'h28D: dout <= 8'b11000011; //  653 : 195 - 0xc3
      12'h28E: dout <= 8'b11100111; //  654 : 231 - 0xe7
      12'h28F: dout <= 8'b01111110; //  655 : 126 - 0x7e
      12'h290: dout <= 8'b11110000; //  656 : 240 - 0xf0 -- Sprite 0x29
      12'h291: dout <= 8'b11100000; //  657 : 224 - 0xe0
      12'h292: dout <= 8'b11000000; //  658 : 192 - 0xc0
      12'h293: dout <= 8'b10000000; //  659 : 128 - 0x80
      12'h294: dout <= 8'b00000000; //  660 :   0 - 0x0
      12'h295: dout <= 8'b00000010; //  661 :   2 - 0x2
      12'h296: dout <= 8'b00000101; //  662 :   5 - 0x5
      12'h297: dout <= 8'b00000010; //  663 :   2 - 0x2
      12'h298: dout <= 8'b00011100; //  664 :  28 - 0x1c -- plane 1
      12'h299: dout <= 8'b00111001; //  665 :  57 - 0x39
      12'h29A: dout <= 8'b01110011; //  666 : 115 - 0x73
      12'h29B: dout <= 8'b11100111; //  667 : 231 - 0xe7
      12'h29C: dout <= 8'b11001111; //  668 : 207 - 0xcf
      12'h29D: dout <= 8'b10011111; //  669 : 159 - 0x9f
      12'h29E: dout <= 8'b00111111; //  670 :  63 - 0x3f
      12'h29F: dout <= 8'b01111111; //  671 : 127 - 0x7f
      12'h2A0: dout <= 8'b01000111; //  672 :  71 - 0x47 -- Sprite 0x2a
      12'h2A1: dout <= 8'b01000110; //  673 :  70 - 0x46
      12'h2A2: dout <= 8'b01000110; //  674 :  70 - 0x46
      12'h2A3: dout <= 8'b01000100; //  675 :  68 - 0x44
      12'h2A4: dout <= 8'b01000100; //  676 :  68 - 0x44
      12'h2A5: dout <= 8'b01000100; //  677 :  68 - 0x44
      12'h2A6: dout <= 8'b01000100; //  678 :  68 - 0x44
      12'h2A7: dout <= 8'b01000100; //  679 :  68 - 0x44
      12'h2A8: dout <= 8'b01100001; //  680 :  97 - 0x61 -- plane 1
      12'h2A9: dout <= 8'b01100011; //  681 :  99 - 0x63
      12'h2AA: dout <= 8'b01100011; //  682 :  99 - 0x63
      12'h2AB: dout <= 8'b01100111; //  683 : 103 - 0x67
      12'h2AC: dout <= 8'b01100110; //  684 : 102 - 0x66
      12'h2AD: dout <= 8'b01100110; //  685 : 102 - 0x66
      12'h2AE: dout <= 8'b01100110; //  686 : 102 - 0x66
      12'h2AF: dout <= 8'b01100110; //  687 : 102 - 0x66
      12'h2B0: dout <= 8'b01111111; //  688 : 127 - 0x7f -- Sprite 0x2b
      12'h2B1: dout <= 8'b00111111; //  689 :  63 - 0x3f
      12'h2B2: dout <= 8'b10011111; //  690 : 159 - 0x9f
      12'h2B3: dout <= 8'b10001111; //  691 : 143 - 0x8f
      12'h2B4: dout <= 8'b01001111; //  692 :  79 - 0x4f
      12'h2B5: dout <= 8'b01000111; //  693 :  71 - 0x47
      12'h2B6: dout <= 8'b01000111; //  694 :  71 - 0x47
      12'h2B7: dout <= 8'b01000111; //  695 :  71 - 0x47
      12'h2B8: dout <= 8'b10000000; //  696 : 128 - 0x80 -- plane 1
      12'h2B9: dout <= 8'b11000000; //  697 : 192 - 0xc0
      12'h2BA: dout <= 8'b11000000; //  698 : 192 - 0xc0
      12'h2BB: dout <= 8'b11100000; //  699 : 224 - 0xe0
      12'h2BC: dout <= 8'b01100000; //  700 :  96 - 0x60
      12'h2BD: dout <= 8'b01100000; //  701 :  96 - 0x60
      12'h2BE: dout <= 8'b01100000; //  702 :  96 - 0x60
      12'h2BF: dout <= 8'b01100000; //  703 :  96 - 0x60
      12'h2C0: dout <= 8'b00100000; //  704 :  32 - 0x20 -- Sprite 0x2c
      12'h2C1: dout <= 8'b00010000; //  705 :  16 - 0x10
      12'h2C2: dout <= 8'b00000000; //  706 :   0 - 0x0
      12'h2C3: dout <= 8'b11000000; //  707 : 192 - 0xc0
      12'h2C4: dout <= 8'b01100000; //  708 :  96 - 0x60
      12'h2C5: dout <= 8'b00100010; //  709 :  34 - 0x22
      12'h2C6: dout <= 8'b00000101; //  710 :   5 - 0x5
      12'h2C7: dout <= 8'b00000010; //  711 :   2 - 0x2
      12'h2C8: dout <= 8'b00111100; //  712 :  60 - 0x3c -- plane 1
      12'h2C9: dout <= 8'b10011001; //  713 : 153 - 0x99
      12'h2CA: dout <= 8'b11000011; //  714 : 195 - 0xc3
      12'h2CB: dout <= 8'b11100111; //  715 : 231 - 0xe7
      12'h2CC: dout <= 8'b11111111; //  716 : 255 - 0xff
      12'h2CD: dout <= 8'b11111111; //  717 : 255 - 0xff
      12'h2CE: dout <= 8'b11111111; //  718 : 255 - 0xff
      12'h2CF: dout <= 8'b11111111; //  719 : 255 - 0xff
      12'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x2d
      12'h2D1: dout <= 8'b01111111; //  721 : 127 - 0x7f
      12'h2D2: dout <= 8'b01000000; //  722 :  64 - 0x40
      12'h2D3: dout <= 8'b01000000; //  723 :  64 - 0x40
      12'h2D4: dout <= 8'b01000000; //  724 :  64 - 0x40
      12'h2D5: dout <= 8'b01000111; //  725 :  71 - 0x47
      12'h2D6: dout <= 8'b01000111; //  726 :  71 - 0x47
      12'h2D7: dout <= 8'b01000111; //  727 :  71 - 0x47
      12'h2D8: dout <= 8'b00000000; //  728 :   0 - 0x0 -- plane 1
      12'h2D9: dout <= 8'b01111111; //  729 : 127 - 0x7f
      12'h2DA: dout <= 8'b01111111; //  730 : 127 - 0x7f
      12'h2DB: dout <= 8'b01100000; //  731 :  96 - 0x60
      12'h2DC: dout <= 8'b01100000; //  732 :  96 - 0x60
      12'h2DD: dout <= 8'b01100000; //  733 :  96 - 0x60
      12'h2DE: dout <= 8'b01100000; //  734 :  96 - 0x60
      12'h2DF: dout <= 8'b01100000; //  735 :  96 - 0x60
      12'h2E0: dout <= 8'b01000100; //  736 :  68 - 0x44 -- Sprite 0x2e
      12'h2E1: dout <= 8'b11000100; //  737 : 196 - 0xc4
      12'h2E2: dout <= 8'b00000100; //  738 :   4 - 0x4
      12'h2E3: dout <= 8'b00000100; //  739 :   4 - 0x4
      12'h2E4: dout <= 8'b00000100; //  740 :   4 - 0x4
      12'h2E5: dout <= 8'b11111100; //  741 : 252 - 0xfc
      12'h2E6: dout <= 8'b11111100; //  742 : 252 - 0xfc
      12'h2E7: dout <= 8'b11111100; //  743 : 252 - 0xfc
      12'h2E8: dout <= 8'b01100110; //  744 : 102 - 0x66 -- plane 1
      12'h2E9: dout <= 8'b11100110; //  745 : 230 - 0xe6
      12'h2EA: dout <= 8'b11100110; //  746 : 230 - 0xe6
      12'h2EB: dout <= 8'b00000110; //  747 :   6 - 0x6
      12'h2EC: dout <= 8'b00000110; //  748 :   6 - 0x6
      12'h2ED: dout <= 8'b00000110; //  749 :   6 - 0x6
      12'h2EE: dout <= 8'b00000110; //  750 :   6 - 0x6
      12'h2EF: dout <= 8'b00000110; //  751 :   6 - 0x6
      12'h2F0: dout <= 8'b00000001; //  752 :   1 - 0x1 -- Sprite 0x2f
      12'h2F1: dout <= 8'b01111100; //  753 : 124 - 0x7c
      12'h2F2: dout <= 8'b01000000; //  754 :  64 - 0x40
      12'h2F3: dout <= 8'b01000100; //  755 :  68 - 0x44
      12'h2F4: dout <= 8'b01000100; //  756 :  68 - 0x44
      12'h2F5: dout <= 8'b01000100; //  757 :  68 - 0x44
      12'h2F6: dout <= 8'b01000100; //  758 :  68 - 0x44
      12'h2F7: dout <= 8'b01000100; //  759 :  68 - 0x44
      12'h2F8: dout <= 8'b00000001; //  760 :   1 - 0x1 -- plane 1
      12'h2F9: dout <= 8'b01111100; //  761 : 124 - 0x7c
      12'h2FA: dout <= 8'b01111110; //  762 : 126 - 0x7e
      12'h2FB: dout <= 8'b01100110; //  763 : 102 - 0x66
      12'h2FC: dout <= 8'b01100110; //  764 : 102 - 0x66
      12'h2FD: dout <= 8'b01100110; //  765 : 102 - 0x66
      12'h2FE: dout <= 8'b01100110; //  766 : 102 - 0x66
      12'h2FF: dout <= 8'b01100110; //  767 : 102 - 0x66
      12'h300: dout <= 8'b00010000; //  768 :  16 - 0x10 -- Sprite 0x30
      12'h301: dout <= 8'b00111000; //  769 :  56 - 0x38
      12'h302: dout <= 8'b00111100; //  770 :  60 - 0x3c
      12'h303: dout <= 8'b00011000; //  771 :  24 - 0x18
      12'h304: dout <= 8'b00000000; //  772 :   0 - 0x0
      12'h305: dout <= 8'b01000010; //  773 :  66 - 0x42
      12'h306: dout <= 8'b01000100; //  774 :  68 - 0x44
      12'h307: dout <= 8'b01001000; //  775 :  72 - 0x48
      12'h308: dout <= 8'b11111111; //  776 : 255 - 0xff -- plane 1
      12'h309: dout <= 8'b11111111; //  777 : 255 - 0xff
      12'h30A: dout <= 8'b01111110; //  778 : 126 - 0x7e
      12'h30B: dout <= 8'b00111100; //  779 :  60 - 0x3c
      12'h30C: dout <= 8'b00011000; //  780 :  24 - 0x18
      12'h30D: dout <= 8'b01000010; //  781 :  66 - 0x42
      12'h30E: dout <= 8'b01100110; //  782 : 102 - 0x66
      12'h30F: dout <= 8'b01111110; //  783 : 126 - 0x7e
      12'h310: dout <= 8'b01000111; //  784 :  71 - 0x47 -- Sprite 0x31
      12'h311: dout <= 8'b01011111; //  785 :  95 - 0x5f
      12'h312: dout <= 8'b00000000; //  786 :   0 - 0x0
      12'h313: dout <= 8'b00000000; //  787 :   0 - 0x0
      12'h314: dout <= 8'b01110000; //  788 : 112 - 0x70
      12'h315: dout <= 8'b00100010; //  789 :  34 - 0x22
      12'h316: dout <= 8'b00000101; //  790 :   5 - 0x5
      12'h317: dout <= 8'b00000010; //  791 :   2 - 0x2
      12'h318: dout <= 8'b01100000; //  792 :  96 - 0x60 -- plane 1
      12'h319: dout <= 8'b01111111; //  793 : 127 - 0x7f
      12'h31A: dout <= 8'b01111111; //  794 : 127 - 0x7f
      12'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      12'h31C: dout <= 8'b11111111; //  796 : 255 - 0xff
      12'h31D: dout <= 8'b11111111; //  797 : 255 - 0xff
      12'h31E: dout <= 8'b11111111; //  798 : 255 - 0xff
      12'h31F: dout <= 8'b11111111; //  799 : 255 - 0xff
      12'h320: dout <= 8'b11111111; //  800 : 255 - 0xff -- Sprite 0x32
      12'h321: dout <= 8'b11111111; //  801 : 255 - 0xff
      12'h322: dout <= 8'b00000000; //  802 :   0 - 0x0
      12'h323: dout <= 8'b00000000; //  803 :   0 - 0x0
      12'h324: dout <= 8'b01110000; //  804 : 112 - 0x70
      12'h325: dout <= 8'b00100010; //  805 :  34 - 0x22
      12'h326: dout <= 8'b00000101; //  806 :   5 - 0x5
      12'h327: dout <= 8'b00000010; //  807 :   2 - 0x2
      12'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- plane 1
      12'h329: dout <= 8'b11111111; //  809 : 255 - 0xff
      12'h32A: dout <= 8'b11111111; //  810 : 255 - 0xff
      12'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      12'h32C: dout <= 8'b11111111; //  812 : 255 - 0xff
      12'h32D: dout <= 8'b11111111; //  813 : 255 - 0xff
      12'h32E: dout <= 8'b11111111; //  814 : 255 - 0xff
      12'h32F: dout <= 8'b11111111; //  815 : 255 - 0xff
      12'h330: dout <= 8'b11111111; //  816 : 255 - 0xff -- Sprite 0x33
      12'h331: dout <= 8'b11011111; //  817 : 223 - 0xdf
      12'h332: dout <= 8'b00011111; //  818 :  31 - 0x1f
      12'h333: dout <= 8'b01000111; //  819 :  71 - 0x47
      12'h334: dout <= 8'b01000111; //  820 :  71 - 0x47
      12'h335: dout <= 8'b01000111; //  821 :  71 - 0x47
      12'h336: dout <= 8'b01000111; //  822 :  71 - 0x47
      12'h337: dout <= 8'b01000111; //  823 :  71 - 0x47
      12'h338: dout <= 8'b00000000; //  824 :   0 - 0x0 -- plane 1
      12'h339: dout <= 8'b11100000; //  825 : 224 - 0xe0
      12'h33A: dout <= 8'b11100000; //  826 : 224 - 0xe0
      12'h33B: dout <= 8'b01100000; //  827 :  96 - 0x60
      12'h33C: dout <= 8'b01100000; //  828 :  96 - 0x60
      12'h33D: dout <= 8'b01100000; //  829 :  96 - 0x60
      12'h33E: dout <= 8'b01100000; //  830 :  96 - 0x60
      12'h33F: dout <= 8'b01100000; //  831 :  96 - 0x60
      12'h340: dout <= 8'b01000100; //  832 :  68 - 0x44 -- Sprite 0x34
      12'h341: dout <= 8'b01000100; //  833 :  68 - 0x44
      12'h342: dout <= 8'b01000100; //  834 :  68 - 0x44
      12'h343: dout <= 8'b01000100; //  835 :  68 - 0x44
      12'h344: dout <= 8'b01000100; //  836 :  68 - 0x44
      12'h345: dout <= 8'b01000100; //  837 :  68 - 0x44
      12'h346: dout <= 8'b01000100; //  838 :  68 - 0x44
      12'h347: dout <= 8'b01000100; //  839 :  68 - 0x44
      12'h348: dout <= 8'b01111110; //  840 : 126 - 0x7e -- plane 1
      12'h349: dout <= 8'b01100110; //  841 : 102 - 0x66
      12'h34A: dout <= 8'b01100110; //  842 : 102 - 0x66
      12'h34B: dout <= 8'b01100110; //  843 : 102 - 0x66
      12'h34C: dout <= 8'b01100110; //  844 : 102 - 0x66
      12'h34D: dout <= 8'b01100110; //  845 : 102 - 0x66
      12'h34E: dout <= 8'b01100110; //  846 : 102 - 0x66
      12'h34F: dout <= 8'b01100110; //  847 : 102 - 0x66
      12'h350: dout <= 8'b00010000; //  848 :  16 - 0x10 -- Sprite 0x35
      12'h351: dout <= 8'b00111000; //  849 :  56 - 0x38
      12'h352: dout <= 8'b01111100; //  850 : 124 - 0x7c
      12'h353: dout <= 8'b11111000; //  851 : 248 - 0xf8
      12'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout <= 8'b01111111; //  853 : 127 - 0x7f
      12'h356: dout <= 8'b01000000; //  854 :  64 - 0x40
      12'h357: dout <= 8'b01000000; //  855 :  64 - 0x40
      12'h358: dout <= 8'b11111111; //  856 : 255 - 0xff -- plane 1
      12'h359: dout <= 8'b11111111; //  857 : 255 - 0xff
      12'h35A: dout <= 8'b11111111; //  858 : 255 - 0xff
      12'h35B: dout <= 8'b11111111; //  859 : 255 - 0xff
      12'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout <= 8'b01111111; //  861 : 127 - 0x7f
      12'h35E: dout <= 8'b01111111; //  862 : 127 - 0x7f
      12'h35F: dout <= 8'b01100000; //  863 :  96 - 0x60
      12'h360: dout <= 8'b00010000; //  864 :  16 - 0x10 -- Sprite 0x36
      12'h361: dout <= 8'b00111000; //  865 :  56 - 0x38
      12'h362: dout <= 8'b01111100; //  866 : 124 - 0x7c
      12'h363: dout <= 8'b11111000; //  867 : 248 - 0xf8
      12'h364: dout <= 8'b00000000; //  868 :   0 - 0x0
      12'h365: dout <= 8'b11111111; //  869 : 255 - 0xff
      12'h366: dout <= 8'b00000000; //  870 :   0 - 0x0
      12'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      12'h368: dout <= 8'b11111111; //  872 : 255 - 0xff -- plane 1
      12'h369: dout <= 8'b11111111; //  873 : 255 - 0xff
      12'h36A: dout <= 8'b11111111; //  874 : 255 - 0xff
      12'h36B: dout <= 8'b11111111; //  875 : 255 - 0xff
      12'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      12'h36D: dout <= 8'b11111111; //  877 : 255 - 0xff
      12'h36E: dout <= 8'b11111111; //  878 : 255 - 0xff
      12'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout <= 8'b01000111; //  880 :  71 - 0x47 -- Sprite 0x37
      12'h371: dout <= 8'b01000111; //  881 :  71 - 0x47
      12'h372: dout <= 8'b01000111; //  882 :  71 - 0x47
      12'h373: dout <= 8'b01000111; //  883 :  71 - 0x47
      12'h374: dout <= 8'b01000111; //  884 :  71 - 0x47
      12'h375: dout <= 8'b11000111; //  885 : 199 - 0xc7
      12'h376: dout <= 8'b00000111; //  886 :   7 - 0x7
      12'h377: dout <= 8'b00000111; //  887 :   7 - 0x7
      12'h378: dout <= 8'b01100000; //  888 :  96 - 0x60 -- plane 1
      12'h379: dout <= 8'b01100000; //  889 :  96 - 0x60
      12'h37A: dout <= 8'b01100000; //  890 :  96 - 0x60
      12'h37B: dout <= 8'b01100000; //  891 :  96 - 0x60
      12'h37C: dout <= 8'b01100000; //  892 :  96 - 0x60
      12'h37D: dout <= 8'b11100000; //  893 : 224 - 0xe0
      12'h37E: dout <= 8'b11100000; //  894 : 224 - 0xe0
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b01000100; //  896 :  68 - 0x44 -- Sprite 0x38
      12'h381: dout <= 8'b01000100; //  897 :  68 - 0x44
      12'h382: dout <= 8'b01000100; //  898 :  68 - 0x44
      12'h383: dout <= 8'b01000100; //  899 :  68 - 0x44
      12'h384: dout <= 8'b01000100; //  900 :  68 - 0x44
      12'h385: dout <= 8'b01011000; //  901 :  88 - 0x58
      12'h386: dout <= 8'b00000000; //  902 :   0 - 0x0
      12'h387: dout <= 8'b00000000; //  903 :   0 - 0x0
      12'h388: dout <= 8'b01100110; //  904 : 102 - 0x66 -- plane 1
      12'h389: dout <= 8'b01100110; //  905 : 102 - 0x66
      12'h38A: dout <= 8'b01100110; //  906 : 102 - 0x66
      12'h38B: dout <= 8'b01100110; //  907 : 102 - 0x66
      12'h38C: dout <= 8'b01100110; //  908 : 102 - 0x66
      12'h38D: dout <= 8'b01111110; //  909 : 126 - 0x7e
      12'h38E: dout <= 8'b01111100; //  910 : 124 - 0x7c
      12'h38F: dout <= 8'b00000001; //  911 :   1 - 0x1
      12'h390: dout <= 8'b00010000; //  912 :  16 - 0x10 -- Sprite 0x39
      12'h391: dout <= 8'b00111000; //  913 :  56 - 0x38
      12'h392: dout <= 8'b01111100; //  914 : 124 - 0x7c
      12'h393: dout <= 8'b11111000; //  915 : 248 - 0xf8
      12'h394: dout <= 8'b01110000; //  916 : 112 - 0x70
      12'h395: dout <= 8'b00100010; //  917 :  34 - 0x22
      12'h396: dout <= 8'b00000100; //  918 :   4 - 0x4
      12'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout <= 8'b11111111; //  920 : 255 - 0xff -- plane 1
      12'h399: dout <= 8'b11111111; //  921 : 255 - 0xff
      12'h39A: dout <= 8'b11111111; //  922 : 255 - 0xff
      12'h39B: dout <= 8'b11111111; //  923 : 255 - 0xff
      12'h39C: dout <= 8'b11111111; //  924 : 255 - 0xff
      12'h39D: dout <= 8'b11111111; //  925 : 255 - 0xff
      12'h39E: dout <= 8'b11111111; //  926 : 255 - 0xff
      12'h39F: dout <= 8'b11111110; //  927 : 254 - 0xfe
      12'h3A0: dout <= 8'b01000100; //  928 :  68 - 0x44 -- Sprite 0x3a
      12'h3A1: dout <= 8'b01000100; //  929 :  68 - 0x44
      12'h3A2: dout <= 8'b01000100; //  930 :  68 - 0x44
      12'h3A3: dout <= 8'b01000100; //  931 :  68 - 0x44
      12'h3A4: dout <= 8'b01000100; //  932 :  68 - 0x44
      12'h3A5: dout <= 8'b01011000; //  933 :  88 - 0x58
      12'h3A6: dout <= 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout <= 8'b01100110; //  936 : 102 - 0x66 -- plane 1
      12'h3A9: dout <= 8'b01100110; //  937 : 102 - 0x66
      12'h3AA: dout <= 8'b01100110; //  938 : 102 - 0x66
      12'h3AB: dout <= 8'b01100110; //  939 : 102 - 0x66
      12'h3AC: dout <= 8'b01100110; //  940 : 102 - 0x66
      12'h3AD: dout <= 8'b01111110; //  941 : 126 - 0x7e
      12'h3AE: dout <= 8'b00111100; //  942 :  60 - 0x3c
      12'h3AF: dout <= 8'b10000001; //  943 : 129 - 0x81
      12'h3B0: dout <= 8'b01000000; //  944 :  64 - 0x40 -- Sprite 0x3b
      12'h3B1: dout <= 8'b01000111; //  945 :  71 - 0x47
      12'h3B2: dout <= 8'b01000111; //  946 :  71 - 0x47
      12'h3B3: dout <= 8'b01000111; //  947 :  71 - 0x47
      12'h3B4: dout <= 8'b01000111; //  948 :  71 - 0x47
      12'h3B5: dout <= 8'b01011111; //  949 :  95 - 0x5f
      12'h3B6: dout <= 8'b00000000; //  950 :   0 - 0x0
      12'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout <= 8'b01100000; //  952 :  96 - 0x60 -- plane 1
      12'h3B9: dout <= 8'b01100000; //  953 :  96 - 0x60
      12'h3BA: dout <= 8'b01100000; //  954 :  96 - 0x60
      12'h3BB: dout <= 8'b01100000; //  955 :  96 - 0x60
      12'h3BC: dout <= 8'b01100000; //  956 :  96 - 0x60
      12'h3BD: dout <= 8'b01111111; //  957 : 127 - 0x7f
      12'h3BE: dout <= 8'b01111111; //  958 : 127 - 0x7f
      12'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x3c
      12'h3C1: dout <= 8'b11111111; //  961 : 255 - 0xff
      12'h3C2: dout <= 8'b11111111; //  962 : 255 - 0xff
      12'h3C3: dout <= 8'b11111111; //  963 : 255 - 0xff
      12'h3C4: dout <= 8'b11111111; //  964 : 255 - 0xff
      12'h3C5: dout <= 8'b11111111; //  965 : 255 - 0xff
      12'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- plane 1
      12'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout <= 8'b11111111; //  973 : 255 - 0xff
      12'h3CE: dout <= 8'b11111111; //  974 : 255 - 0xff
      12'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout <= 8'b00000111; //  976 :   7 - 0x7 -- Sprite 0x3d
      12'h3D1: dout <= 8'b11111111; //  977 : 255 - 0xff
      12'h3D2: dout <= 8'b11111111; //  978 : 255 - 0xff
      12'h3D3: dout <= 8'b11111111; //  979 : 255 - 0xff
      12'h3D4: dout <= 8'b11111111; //  980 : 255 - 0xff
      12'h3D5: dout <= 8'b11111111; //  981 : 255 - 0xff
      12'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0 -- plane 1
      12'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout <= 8'b11111111; //  989 : 255 - 0xff
      12'h3DE: dout <= 8'b11111111; //  990 : 255 - 0xff
      12'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout <= 8'b00010000; //  992 :  16 - 0x10 -- Sprite 0x3e
      12'h3E1: dout <= 8'b00111000; //  993 :  56 - 0x38
      12'h3E2: dout <= 8'b01110001; //  994 : 113 - 0x71
      12'h3E3: dout <= 8'b11100010; //  995 : 226 - 0xe2
      12'h3E4: dout <= 8'b01100010; //  996 :  98 - 0x62
      12'h3E5: dout <= 8'b00100001; //  997 :  33 - 0x21
      12'h3E6: dout <= 8'b00000000; //  998 :   0 - 0x0
      12'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      12'h3E8: dout <= 8'b11111110; // 1000 : 254 - 0xfe -- plane 1
      12'h3E9: dout <= 8'b11111100; // 1001 : 252 - 0xfc
      12'h3EA: dout <= 8'b11111001; // 1002 : 249 - 0xf9
      12'h3EB: dout <= 8'b11110011; // 1003 : 243 - 0xf3
      12'h3EC: dout <= 8'b11110011; // 1004 : 243 - 0xf3
      12'h3ED: dout <= 8'b11111001; // 1005 : 249 - 0xf9
      12'h3EE: dout <= 8'b11111100; // 1006 : 252 - 0xfc
      12'h3EF: dout <= 8'b11111110; // 1007 : 254 - 0xfe
      12'h3F0: dout <= 8'b10000111; // 1008 : 135 - 0x87 -- Sprite 0x3f
      12'h3F1: dout <= 8'b10000111; // 1009 : 135 - 0x87
      12'h3F2: dout <= 8'b00000111; // 1010 :   7 - 0x7
      12'h3F3: dout <= 8'b00001111; // 1011 :  15 - 0xf
      12'h3F4: dout <= 8'b00001111; // 1012 :  15 - 0xf
      12'h3F5: dout <= 8'b00011111; // 1013 :  31 - 0x1f
      12'h3F6: dout <= 8'b10011111; // 1014 : 159 - 0x9f
      12'h3F7: dout <= 8'b10001111; // 1015 : 143 - 0x8f
      12'h3F8: dout <= 8'b11100000; // 1016 : 224 - 0xe0 -- plane 1
      12'h3F9: dout <= 8'b11000000; // 1017 : 192 - 0xc0
      12'h3FA: dout <= 8'b11000000; // 1018 : 192 - 0xc0
      12'h3FB: dout <= 8'b10000000; // 1019 : 128 - 0x80
      12'h3FC: dout <= 8'b10000000; // 1020 : 128 - 0x80
      12'h3FD: dout <= 8'b11000000; // 1021 : 192 - 0xc0
      12'h3FE: dout <= 8'b11000000; // 1022 : 192 - 0xc0
      12'h3FF: dout <= 8'b11100000; // 1023 : 224 - 0xe0
      12'h400: dout <= 8'b01000100; // 1024 :  68 - 0x44 -- Sprite 0x40
      12'h401: dout <= 8'b01000100; // 1025 :  68 - 0x44
      12'h402: dout <= 8'b01000100; // 1026 :  68 - 0x44
      12'h403: dout <= 8'b01000100; // 1027 :  68 - 0x44
      12'h404: dout <= 8'b01000100; // 1028 :  68 - 0x44
      12'h405: dout <= 8'b01000110; // 1029 :  70 - 0x46
      12'h406: dout <= 8'b01000110; // 1030 :  70 - 0x46
      12'h407: dout <= 8'b01000111; // 1031 :  71 - 0x47
      12'h408: dout <= 8'b01100110; // 1032 : 102 - 0x66 -- plane 1
      12'h409: dout <= 8'b01100110; // 1033 : 102 - 0x66
      12'h40A: dout <= 8'b01100110; // 1034 : 102 - 0x66
      12'h40B: dout <= 8'b01100110; // 1035 : 102 - 0x66
      12'h40C: dout <= 8'b01100111; // 1036 : 103 - 0x67
      12'h40D: dout <= 8'b01100011; // 1037 :  99 - 0x63
      12'h40E: dout <= 8'b01100011; // 1038 :  99 - 0x63
      12'h40F: dout <= 8'b01100001; // 1039 :  97 - 0x61
      12'h410: dout <= 8'b00010000; // 1040 :  16 - 0x10 -- Sprite 0x41
      12'h411: dout <= 8'b00111000; // 1041 :  56 - 0x38
      12'h412: dout <= 8'b01111100; // 1042 : 124 - 0x7c
      12'h413: dout <= 8'b01111000; // 1043 : 120 - 0x78
      12'h414: dout <= 8'b00110000; // 1044 :  48 - 0x30
      12'h415: dout <= 8'b00000010; // 1045 :   2 - 0x2
      12'h416: dout <= 8'b00000101; // 1046 :   5 - 0x5
      12'h417: dout <= 8'b00000010; // 1047 :   2 - 0x2
      12'h418: dout <= 8'b11111111; // 1048 : 255 - 0xff -- plane 1
      12'h419: dout <= 8'b11111111; // 1049 : 255 - 0xff
      12'h41A: dout <= 8'b11111111; // 1050 : 255 - 0xff
      12'h41B: dout <= 8'b01111111; // 1051 : 127 - 0x7f
      12'h41C: dout <= 8'b01111111; // 1052 : 127 - 0x7f
      12'h41D: dout <= 8'b00111111; // 1053 :  63 - 0x3f
      12'h41E: dout <= 8'b10011111; // 1054 : 159 - 0x9f
      12'h41F: dout <= 8'b11000111; // 1055 : 199 - 0xc7
      12'h420: dout <= 8'b00010000; // 1056 :  16 - 0x10 -- Sprite 0x42
      12'h421: dout <= 8'b00111000; // 1057 :  56 - 0x38
      12'h422: dout <= 8'b01111100; // 1058 : 124 - 0x7c
      12'h423: dout <= 8'b11111000; // 1059 : 248 - 0xf8
      12'h424: dout <= 8'b01110000; // 1060 : 112 - 0x70
      12'h425: dout <= 8'b00100000; // 1061 :  32 - 0x20
      12'h426: dout <= 8'b00000001; // 1062 :   1 - 0x1
      12'h427: dout <= 8'b00000010; // 1063 :   2 - 0x2
      12'h428: dout <= 8'b11111111; // 1064 : 255 - 0xff -- plane 1
      12'h429: dout <= 8'b11111111; // 1065 : 255 - 0xff
      12'h42A: dout <= 8'b11111111; // 1066 : 255 - 0xff
      12'h42B: dout <= 8'b11111110; // 1067 : 254 - 0xfe
      12'h42C: dout <= 8'b11111110; // 1068 : 254 - 0xfe
      12'h42D: dout <= 8'b11111100; // 1069 : 252 - 0xfc
      12'h42E: dout <= 8'b11111001; // 1070 : 249 - 0xf9
      12'h42F: dout <= 8'b11100011; // 1071 : 227 - 0xe3
      12'h430: dout <= 8'b01000100; // 1072 :  68 - 0x44 -- Sprite 0x43
      12'h431: dout <= 8'b01000100; // 1073 :  68 - 0x44
      12'h432: dout <= 8'b01000100; // 1074 :  68 - 0x44
      12'h433: dout <= 8'b01000100; // 1075 :  68 - 0x44
      12'h434: dout <= 8'b10000100; // 1076 : 132 - 0x84
      12'h435: dout <= 8'b10000100; // 1077 : 132 - 0x84
      12'h436: dout <= 8'b00000100; // 1078 :   4 - 0x4
      12'h437: dout <= 8'b00001100; // 1079 :  12 - 0xc
      12'h438: dout <= 8'b01100110; // 1080 : 102 - 0x66 -- plane 1
      12'h439: dout <= 8'b01100110; // 1081 : 102 - 0x66
      12'h43A: dout <= 8'b01100110; // 1082 : 102 - 0x66
      12'h43B: dout <= 8'b01100110; // 1083 : 102 - 0x66
      12'h43C: dout <= 8'b11100110; // 1084 : 230 - 0xe6
      12'h43D: dout <= 8'b11000110; // 1085 : 198 - 0xc6
      12'h43E: dout <= 8'b11000110; // 1086 : 198 - 0xc6
      12'h43F: dout <= 8'b10000110; // 1087 : 134 - 0x86
      12'h440: dout <= 8'b00010000; // 1088 :  16 - 0x10 -- Sprite 0x44
      12'h441: dout <= 8'b00111000; // 1089 :  56 - 0x38
      12'h442: dout <= 8'b01111100; // 1090 : 124 - 0x7c
      12'h443: dout <= 8'b11111000; // 1091 : 248 - 0xf8
      12'h444: dout <= 8'b01110000; // 1092 : 112 - 0x70
      12'h445: dout <= 8'b00100010; // 1093 :  34 - 0x22
      12'h446: dout <= 8'b00000101; // 1094 :   5 - 0x5
      12'h447: dout <= 8'b00000010; // 1095 :   2 - 0x2
      12'h448: dout <= 8'b11111110; // 1096 : 254 - 0xfe -- plane 1
      12'h449: dout <= 8'b11111111; // 1097 : 255 - 0xff
      12'h44A: dout <= 8'b11111111; // 1098 : 255 - 0xff
      12'h44B: dout <= 8'b11111111; // 1099 : 255 - 0xff
      12'h44C: dout <= 8'b11111111; // 1100 : 255 - 0xff
      12'h44D: dout <= 8'b11111111; // 1101 : 255 - 0xff
      12'h44E: dout <= 8'b11111111; // 1102 : 255 - 0xff
      12'h44F: dout <= 8'b11111111; // 1103 : 255 - 0xff
      12'h450: dout <= 8'b01001111; // 1104 :  79 - 0x4f -- Sprite 0x45
      12'h451: dout <= 8'b01000111; // 1105 :  71 - 0x47
      12'h452: dout <= 8'b01000111; // 1106 :  71 - 0x47
      12'h453: dout <= 8'b01000111; // 1107 :  71 - 0x47
      12'h454: dout <= 8'b01000111; // 1108 :  71 - 0x47
      12'h455: dout <= 8'b01000111; // 1109 :  71 - 0x47
      12'h456: dout <= 8'b01000111; // 1110 :  71 - 0x47
      12'h457: dout <= 8'b01000111; // 1111 :  71 - 0x47
      12'h458: dout <= 8'b01100000; // 1112 :  96 - 0x60 -- plane 1
      12'h459: dout <= 8'b01100000; // 1113 :  96 - 0x60
      12'h45A: dout <= 8'b01100000; // 1114 :  96 - 0x60
      12'h45B: dout <= 8'b01100000; // 1115 :  96 - 0x60
      12'h45C: dout <= 8'b01100000; // 1116 :  96 - 0x60
      12'h45D: dout <= 8'b01100000; // 1117 :  96 - 0x60
      12'h45E: dout <= 8'b01100000; // 1118 :  96 - 0x60
      12'h45F: dout <= 8'b01100000; // 1119 :  96 - 0x60
      12'h460: dout <= 8'b10100000; // 1120 : 160 - 0xa0 -- Sprite 0x46
      12'h461: dout <= 8'b10011111; // 1121 : 159 - 0x9f
      12'h462: dout <= 8'b11000000; // 1122 : 192 - 0xc0
      12'h463: dout <= 8'b11100000; // 1123 : 224 - 0xe0
      12'h464: dout <= 8'b11111000; // 1124 : 248 - 0xf8
      12'h465: dout <= 8'b11111111; // 1125 : 255 - 0xff
      12'h466: dout <= 8'b11111111; // 1126 : 255 - 0xff
      12'h467: dout <= 8'b11111111; // 1127 : 255 - 0xff
      12'h468: dout <= 8'b11110000; // 1128 : 240 - 0xf0 -- plane 1
      12'h469: dout <= 8'b01111111; // 1129 : 127 - 0x7f
      12'h46A: dout <= 8'b00011111; // 1130 :  31 - 0x1f
      12'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      12'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      12'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      12'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      12'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      12'h470: dout <= 8'b00001100; // 1136 :  12 - 0xc -- Sprite 0x47
      12'h471: dout <= 8'b11110000; // 1137 : 240 - 0xf0
      12'h472: dout <= 8'b00000000; // 1138 :   0 - 0x0
      12'h473: dout <= 8'b00000000; // 1139 :   0 - 0x0
      12'h474: dout <= 8'b00000001; // 1140 :   1 - 0x1
      12'h475: dout <= 8'b11111111; // 1141 : 255 - 0xff
      12'h476: dout <= 8'b11111111; // 1142 : 255 - 0xff
      12'h477: dout <= 8'b11111111; // 1143 : 255 - 0xff
      12'h478: dout <= 8'b00001111; // 1144 :  15 - 0xf -- plane 1
      12'h479: dout <= 8'b11111110; // 1145 : 254 - 0xfe
      12'h47A: dout <= 8'b11111000; // 1146 : 248 - 0xf8
      12'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      12'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      12'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      12'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      12'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout <= 8'b00001100; // 1152 :  12 - 0xc -- Sprite 0x48
      12'h481: dout <= 8'b00011101; // 1153 :  29 - 0x1d
      12'h482: dout <= 8'b00111000; // 1154 :  56 - 0x38
      12'h483: dout <= 8'b01111110; // 1155 : 126 - 0x7e
      12'h484: dout <= 8'b11111110; // 1156 : 254 - 0xfe
      12'h485: dout <= 8'b11111111; // 1157 : 255 - 0xff
      12'h486: dout <= 8'b11111111; // 1158 : 255 - 0xff
      12'h487: dout <= 8'b11111111; // 1159 : 255 - 0xff
      12'h488: dout <= 8'b00000110; // 1160 :   6 - 0x6 -- plane 1
      12'h489: dout <= 8'b00000111; // 1161 :   7 - 0x7
      12'h48A: dout <= 8'b00000111; // 1162 :   7 - 0x7
      12'h48B: dout <= 8'b00000000; // 1163 :   0 - 0x0
      12'h48C: dout <= 8'b00000000; // 1164 :   0 - 0x0
      12'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      12'h48E: dout <= 8'b00000000; // 1166 :   0 - 0x0
      12'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout <= 8'b11111111; // 1168 : 255 - 0xff -- Sprite 0x49
      12'h491: dout <= 8'b11111111; // 1169 : 255 - 0xff
      12'h492: dout <= 8'b11111111; // 1170 : 255 - 0xff
      12'h493: dout <= 8'b11111111; // 1171 : 255 - 0xff
      12'h494: dout <= 8'b11111111; // 1172 : 255 - 0xff
      12'h495: dout <= 8'b11111111; // 1173 : 255 - 0xff
      12'h496: dout <= 8'b11111111; // 1174 : 255 - 0xff
      12'h497: dout <= 8'b11111111; // 1175 : 255 - 0xff
      12'h498: dout <= 8'b00000000; // 1176 :   0 - 0x0 -- plane 1
      12'h499: dout <= 8'b00000000; // 1177 :   0 - 0x0
      12'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      12'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      12'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      12'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      12'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      12'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      12'h4A0: dout <= 8'b11111111; // 1184 : 255 - 0xff -- Sprite 0x4a
      12'h4A1: dout <= 8'b11101111; // 1185 : 239 - 0xef
      12'h4A2: dout <= 8'b11111101; // 1186 : 253 - 0xfd
      12'h4A3: dout <= 8'b11111111; // 1187 : 255 - 0xff
      12'h4A4: dout <= 8'b11111111; // 1188 : 255 - 0xff
      12'h4A5: dout <= 8'b11101111; // 1189 : 239 - 0xef
      12'h4A6: dout <= 8'b11111110; // 1190 : 254 - 0xfe
      12'h4A7: dout <= 8'b11111111; // 1191 : 255 - 0xff
      12'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0 -- plane 1
      12'h4A9: dout <= 8'b01110110; // 1193 : 118 - 0x76
      12'h4AA: dout <= 8'b01010111; // 1194 :  87 - 0x57
      12'h4AB: dout <= 8'b01010101; // 1195 :  85 - 0x55
      12'h4AC: dout <= 8'b01010101; // 1196 :  85 - 0x55
      12'h4AD: dout <= 8'b01110101; // 1197 : 117 - 0x75
      12'h4AE: dout <= 8'b01000111; // 1198 :  71 - 0x47
      12'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      12'h4B0: dout <= 8'b11111111; // 1200 : 255 - 0xff -- Sprite 0x4b
      12'h4B1: dout <= 8'b11101010; // 1201 : 234 - 0xea
      12'h4B2: dout <= 8'b11111111; // 1202 : 255 - 0xff
      12'h4B3: dout <= 8'b10101111; // 1203 : 175 - 0xaf
      12'h4B4: dout <= 8'b11111111; // 1204 : 255 - 0xff
      12'h4B5: dout <= 8'b11111111; // 1205 : 255 - 0xff
      12'h4B6: dout <= 8'b11111010; // 1206 : 250 - 0xfa
      12'h4B7: dout <= 8'b11111111; // 1207 : 255 - 0xff
      12'h4B8: dout <= 8'b00000000; // 1208 :   0 - 0x0 -- plane 1
      12'h4B9: dout <= 8'b01110111; // 1209 : 119 - 0x77
      12'h4BA: dout <= 8'b00010101; // 1210 :  21 - 0x15
      12'h4BB: dout <= 8'b01110101; // 1211 : 117 - 0x75
      12'h4BC: dout <= 8'b01000101; // 1212 :  69 - 0x45
      12'h4BD: dout <= 8'b01000101; // 1213 :  69 - 0x45
      12'h4BE: dout <= 8'b01110111; // 1214 : 119 - 0x77
      12'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      12'h4C0: dout <= 8'b11111111; // 1216 : 255 - 0xff -- Sprite 0x4c
      12'h4C1: dout <= 8'b11111111; // 1217 : 255 - 0xff
      12'h4C2: dout <= 8'b11111111; // 1218 : 255 - 0xff
      12'h4C3: dout <= 8'b11111111; // 1219 : 255 - 0xff
      12'h4C4: dout <= 8'b11111111; // 1220 : 255 - 0xff
      12'h4C5: dout <= 8'b11111111; // 1221 : 255 - 0xff
      12'h4C6: dout <= 8'b11111110; // 1222 : 254 - 0xfe
      12'h4C7: dout <= 8'b11111111; // 1223 : 255 - 0xff
      12'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0 -- plane 1
      12'h4C9: dout <= 8'b00100100; // 1225 :  36 - 0x24
      12'h4CA: dout <= 8'b01101100; // 1226 : 108 - 0x6c
      12'h4CB: dout <= 8'b00100100; // 1227 :  36 - 0x24
      12'h4CC: dout <= 8'b00100100; // 1228 :  36 - 0x24
      12'h4CD: dout <= 8'b00100100; // 1229 :  36 - 0x24
      12'h4CE: dout <= 8'b00100101; // 1230 :  37 - 0x25
      12'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      12'h4D0: dout <= 8'b11111111; // 1232 : 255 - 0xff -- Sprite 0x4d
      12'h4D1: dout <= 8'b10111111; // 1233 : 191 - 0xbf
      12'h4D2: dout <= 8'b11111110; // 1234 : 254 - 0xfe
      12'h4D3: dout <= 8'b10101111; // 1235 : 175 - 0xaf
      12'h4D4: dout <= 8'b11111111; // 1236 : 255 - 0xff
      12'h4D5: dout <= 8'b11111111; // 1237 : 255 - 0xff
      12'h4D6: dout <= 8'b11101111; // 1238 : 239 - 0xef
      12'h4D7: dout <= 8'b11111111; // 1239 : 255 - 0xff
      12'h4D8: dout <= 8'b00000000; // 1240 :   0 - 0x0 -- plane 1
      12'h4D9: dout <= 8'b01110100; // 1241 : 116 - 0x74
      12'h4DA: dout <= 8'b01000111; // 1242 :  71 - 0x47
      12'h4DB: dout <= 8'b01110101; // 1243 : 117 - 0x75
      12'h4DC: dout <= 8'b00010101; // 1244 :  21 - 0x15
      12'h4DD: dout <= 8'b00010101; // 1245 :  21 - 0x15
      12'h4DE: dout <= 8'b01110101; // 1246 : 117 - 0x75
      12'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout <= 8'b11111111; // 1248 : 255 - 0xff -- Sprite 0x4e
      12'h4E1: dout <= 8'b11111111; // 1249 : 255 - 0xff
      12'h4E2: dout <= 8'b11111011; // 1250 : 251 - 0xfb
      12'h4E3: dout <= 8'b11111111; // 1251 : 255 - 0xff
      12'h4E4: dout <= 8'b11111111; // 1252 : 255 - 0xff
      12'h4E5: dout <= 8'b11111111; // 1253 : 255 - 0xff
      12'h4E6: dout <= 8'b11111110; // 1254 : 254 - 0xfe
      12'h4E7: dout <= 8'b11111111; // 1255 : 255 - 0xff
      12'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0 -- plane 1
      12'h4E9: dout <= 8'b01000000; // 1257 :  64 - 0x40
      12'h4EA: dout <= 8'b00011101; // 1258 :  29 - 0x1d
      12'h4EB: dout <= 8'b01010101; // 1259 :  85 - 0x55
      12'h4EC: dout <= 8'b01010001; // 1260 :  81 - 0x51
      12'h4ED: dout <= 8'b01010001; // 1261 :  81 - 0x51
      12'h4EE: dout <= 8'b01010001; // 1262 :  81 - 0x51
      12'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout <= 8'b11111111; // 1264 : 255 - 0xff -- Sprite 0x4f
      12'h4F1: dout <= 8'b11111111; // 1265 : 255 - 0xff
      12'h4F2: dout <= 8'b11110111; // 1266 : 247 - 0xf7
      12'h4F3: dout <= 8'b11111110; // 1267 : 254 - 0xfe
      12'h4F4: dout <= 8'b11111011; // 1268 : 251 - 0xfb
      12'h4F5: dout <= 8'b11111111; // 1269 : 255 - 0xff
      12'h4F6: dout <= 8'b11101111; // 1270 : 239 - 0xef
      12'h4F7: dout <= 8'b11111101; // 1271 : 253 - 0xfd
      12'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0 -- plane 1
      12'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout <= 8'b01001000; // 1274 :  72 - 0x48
      12'h4FB: dout <= 8'b01000001; // 1275 :  65 - 0x41
      12'h4FC: dout <= 8'b01000100; // 1276 :  68 - 0x44
      12'h4FD: dout <= 8'b01000000; // 1277 :  64 - 0x40
      12'h4FE: dout <= 8'b11010000; // 1278 : 208 - 0xd0
      12'h4FF: dout <= 8'b00000010; // 1279 :   2 - 0x2
      12'h500: dout <= 8'b11111111; // 1280 : 255 - 0xff -- Sprite 0x50
      12'h501: dout <= 8'b11111111; // 1281 : 255 - 0xff
      12'h502: dout <= 8'b00000011; // 1282 :   3 - 0x3
      12'h503: dout <= 8'b00000001; // 1283 :   1 - 0x1
      12'h504: dout <= 8'b11101110; // 1284 : 238 - 0xee
      12'h505: dout <= 8'b00000000; // 1285 :   0 - 0x0
      12'h506: dout <= 8'b11101110; // 1286 : 238 - 0xee
      12'h507: dout <= 8'b11101110; // 1287 : 238 - 0xee
      12'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0 -- plane 1
      12'h509: dout <= 8'b00000000; // 1289 :   0 - 0x0
      12'h50A: dout <= 8'b11111100; // 1290 : 252 - 0xfc
      12'h50B: dout <= 8'b11111110; // 1291 : 254 - 0xfe
      12'h50C: dout <= 8'b11101110; // 1292 : 238 - 0xee
      12'h50D: dout <= 8'b11101110; // 1293 : 238 - 0xee
      12'h50E: dout <= 8'b11101110; // 1294 : 238 - 0xee
      12'h50F: dout <= 8'b11101110; // 1295 : 238 - 0xee
      12'h510: dout <= 8'b11111111; // 1296 : 255 - 0xff -- Sprite 0x51
      12'h511: dout <= 8'b11111111; // 1297 : 255 - 0xff
      12'h512: dout <= 8'b00000011; // 1298 :   3 - 0x3
      12'h513: dout <= 8'b00000001; // 1299 :   1 - 0x1
      12'h514: dout <= 8'b11101110; // 1300 : 238 - 0xee
      12'h515: dout <= 8'b00000000; // 1301 :   0 - 0x0
      12'h516: dout <= 8'b11101110; // 1302 : 238 - 0xee
      12'h517: dout <= 8'b11101110; // 1303 : 238 - 0xee
      12'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0 -- plane 1
      12'h519: dout <= 8'b00000000; // 1305 :   0 - 0x0
      12'h51A: dout <= 8'b11111100; // 1306 : 252 - 0xfc
      12'h51B: dout <= 8'b11111110; // 1307 : 254 - 0xfe
      12'h51C: dout <= 8'b11101110; // 1308 : 238 - 0xee
      12'h51D: dout <= 8'b11101110; // 1309 : 238 - 0xee
      12'h51E: dout <= 8'b11101110; // 1310 : 238 - 0xee
      12'h51F: dout <= 8'b11101110; // 1311 : 238 - 0xee
      12'h520: dout <= 8'b11111111; // 1312 : 255 - 0xff -- Sprite 0x52
      12'h521: dout <= 8'b11111111; // 1313 : 255 - 0xff
      12'h522: dout <= 8'b00000001; // 1314 :   1 - 0x1
      12'h523: dout <= 8'b00000000; // 1315 :   0 - 0x0
      12'h524: dout <= 8'b11100000; // 1316 : 224 - 0xe0
      12'h525: dout <= 8'b00001111; // 1317 :  15 - 0xf
      12'h526: dout <= 8'b11111111; // 1318 : 255 - 0xff
      12'h527: dout <= 8'b11111011; // 1319 : 251 - 0xfb
      12'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0 -- plane 1
      12'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      12'h52A: dout <= 8'b11111110; // 1322 : 254 - 0xfe
      12'h52B: dout <= 8'b11111110; // 1323 : 254 - 0xfe
      12'h52C: dout <= 8'b11100000; // 1324 : 224 - 0xe0
      12'h52D: dout <= 8'b11100000; // 1325 : 224 - 0xe0
      12'h52E: dout <= 8'b11111000; // 1326 : 248 - 0xf8
      12'h52F: dout <= 8'b11111000; // 1327 : 248 - 0xf8
      12'h530: dout <= 8'b11111111; // 1328 : 255 - 0xff -- Sprite 0x53
      12'h531: dout <= 8'b11111111; // 1329 : 255 - 0xff
      12'h532: dout <= 8'b10000011; // 1330 : 131 - 0x83
      12'h533: dout <= 8'b00000001; // 1331 :   1 - 0x1
      12'h534: dout <= 8'b11101110; // 1332 : 238 - 0xee
      12'h535: dout <= 8'b00000000; // 1333 :   0 - 0x0
      12'h536: dout <= 8'b11111111; // 1334 : 255 - 0xff
      12'h537: dout <= 8'b11111111; // 1335 : 255 - 0xff
      12'h538: dout <= 8'b00000000; // 1336 :   0 - 0x0 -- plane 1
      12'h539: dout <= 8'b00000000; // 1337 :   0 - 0x0
      12'h53A: dout <= 8'b01111100; // 1338 : 124 - 0x7c
      12'h53B: dout <= 8'b11111110; // 1339 : 254 - 0xfe
      12'h53C: dout <= 8'b11101110; // 1340 : 238 - 0xee
      12'h53D: dout <= 8'b11100000; // 1341 : 224 - 0xe0
      12'h53E: dout <= 8'b11111100; // 1342 : 252 - 0xfc
      12'h53F: dout <= 8'b01111110; // 1343 : 126 - 0x7e
      12'h540: dout <= 8'b11111111; // 1344 : 255 - 0xff -- Sprite 0x54
      12'h541: dout <= 8'b11111111; // 1345 : 255 - 0xff
      12'h542: dout <= 8'b00000001; // 1346 :   1 - 0x1
      12'h543: dout <= 8'b00000000; // 1347 :   0 - 0x0
      12'h544: dout <= 8'b10111000; // 1348 : 184 - 0xb8
      12'h545: dout <= 8'b11000011; // 1349 : 195 - 0xc3
      12'h546: dout <= 8'b11111011; // 1350 : 251 - 0xfb
      12'h547: dout <= 8'b11111011; // 1351 : 251 - 0xfb
      12'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0 -- plane 1
      12'h549: dout <= 8'b00000000; // 1353 :   0 - 0x0
      12'h54A: dout <= 8'b11111110; // 1354 : 254 - 0xfe
      12'h54B: dout <= 8'b11111110; // 1355 : 254 - 0xfe
      12'h54C: dout <= 8'b00111000; // 1356 :  56 - 0x38
      12'h54D: dout <= 8'b00111000; // 1357 :  56 - 0x38
      12'h54E: dout <= 8'b00111000; // 1358 :  56 - 0x38
      12'h54F: dout <= 8'b00111000; // 1359 :  56 - 0x38
      12'h550: dout <= 8'b11111111; // 1360 : 255 - 0xff -- Sprite 0x55
      12'h551: dout <= 8'b11111111; // 1361 : 255 - 0xff
      12'h552: dout <= 8'b10000011; // 1362 : 131 - 0x83
      12'h553: dout <= 8'b00000001; // 1363 :   1 - 0x1
      12'h554: dout <= 8'b11101110; // 1364 : 238 - 0xee
      12'h555: dout <= 8'b00000000; // 1365 :   0 - 0x0
      12'h556: dout <= 8'b11101110; // 1366 : 238 - 0xee
      12'h557: dout <= 8'b11101110; // 1367 : 238 - 0xee
      12'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0 -- plane 1
      12'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout <= 8'b01111100; // 1370 : 124 - 0x7c
      12'h55B: dout <= 8'b11111110; // 1371 : 254 - 0xfe
      12'h55C: dout <= 8'b11101110; // 1372 : 238 - 0xee
      12'h55D: dout <= 8'b11101110; // 1373 : 238 - 0xee
      12'h55E: dout <= 8'b11101110; // 1374 : 238 - 0xee
      12'h55F: dout <= 8'b11101110; // 1375 : 238 - 0xee
      12'h560: dout <= 8'b11111111; // 1376 : 255 - 0xff -- Sprite 0x56
      12'h561: dout <= 8'b11111111; // 1377 : 255 - 0xff
      12'h562: dout <= 8'b00011111; // 1378 :  31 - 0x1f
      12'h563: dout <= 8'b00001111; // 1379 :  15 - 0xf
      12'h564: dout <= 8'b11101111; // 1380 : 239 - 0xef
      12'h565: dout <= 8'b00001111; // 1381 :  15 - 0xf
      12'h566: dout <= 8'b11101111; // 1382 : 239 - 0xef
      12'h567: dout <= 8'b11101111; // 1383 : 239 - 0xef
      12'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0 -- plane 1
      12'h569: dout <= 8'b00000000; // 1385 :   0 - 0x0
      12'h56A: dout <= 8'b11100000; // 1386 : 224 - 0xe0
      12'h56B: dout <= 8'b11100000; // 1387 : 224 - 0xe0
      12'h56C: dout <= 8'b11100000; // 1388 : 224 - 0xe0
      12'h56D: dout <= 8'b11100000; // 1389 : 224 - 0xe0
      12'h56E: dout <= 8'b11100000; // 1390 : 224 - 0xe0
      12'h56F: dout <= 8'b11100000; // 1391 : 224 - 0xe0
      12'h570: dout <= 8'b11111111; // 1392 : 255 - 0xff -- Sprite 0x57
      12'h571: dout <= 8'b11111111; // 1393 : 255 - 0xff
      12'h572: dout <= 8'b00010001; // 1394 :  17 - 0x11
      12'h573: dout <= 8'b00000000; // 1395 :   0 - 0x0
      12'h574: dout <= 8'b11101110; // 1396 : 238 - 0xee
      12'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      12'h576: dout <= 8'b11101110; // 1398 : 238 - 0xee
      12'h577: dout <= 8'b11101110; // 1399 : 238 - 0xee
      12'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0 -- plane 1
      12'h579: dout <= 8'b00000000; // 1401 :   0 - 0x0
      12'h57A: dout <= 8'b11101110; // 1402 : 238 - 0xee
      12'h57B: dout <= 8'b11101110; // 1403 : 238 - 0xee
      12'h57C: dout <= 8'b11101110; // 1404 : 238 - 0xee
      12'h57D: dout <= 8'b11101110; // 1405 : 238 - 0xee
      12'h57E: dout <= 8'b11101110; // 1406 : 238 - 0xee
      12'h57F: dout <= 8'b11101110; // 1407 : 238 - 0xee
      12'h580: dout <= 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0x58
      12'h581: dout <= 8'b11111111; // 1409 : 255 - 0xff
      12'h582: dout <= 8'b01110001; // 1410 : 113 - 0x71
      12'h583: dout <= 8'b00110000; // 1411 :  48 - 0x30
      12'h584: dout <= 8'b11111110; // 1412 : 254 - 0xfe
      12'h585: dout <= 8'b00000000; // 1413 :   0 - 0x0
      12'h586: dout <= 8'b11111110; // 1414 : 254 - 0xfe
      12'h587: dout <= 8'b11101110; // 1415 : 238 - 0xee
      12'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0 -- plane 1
      12'h589: dout <= 8'b00000000; // 1417 :   0 - 0x0
      12'h58A: dout <= 8'b10001110; // 1418 : 142 - 0x8e
      12'h58B: dout <= 8'b11001110; // 1419 : 206 - 0xce
      12'h58C: dout <= 8'b11101110; // 1420 : 238 - 0xee
      12'h58D: dout <= 8'b11111110; // 1421 : 254 - 0xfe
      12'h58E: dout <= 8'b11111110; // 1422 : 254 - 0xfe
      12'h58F: dout <= 8'b11101110; // 1423 : 238 - 0xee
      12'h590: dout <= 8'b11111111; // 1424 : 255 - 0xff -- Sprite 0x59
      12'h591: dout <= 8'b11111111; // 1425 : 255 - 0xff
      12'h592: dout <= 8'b00000011; // 1426 :   3 - 0x3
      12'h593: dout <= 8'b00000001; // 1427 :   1 - 0x1
      12'h594: dout <= 8'b11101110; // 1428 : 238 - 0xee
      12'h595: dout <= 8'b00000000; // 1429 :   0 - 0x0
      12'h596: dout <= 8'b11101110; // 1430 : 238 - 0xee
      12'h597: dout <= 8'b11101110; // 1431 : 238 - 0xee
      12'h598: dout <= 8'b00000000; // 1432 :   0 - 0x0 -- plane 1
      12'h599: dout <= 8'b00000000; // 1433 :   0 - 0x0
      12'h59A: dout <= 8'b11111100; // 1434 : 252 - 0xfc
      12'h59B: dout <= 8'b11111110; // 1435 : 254 - 0xfe
      12'h59C: dout <= 8'b11101110; // 1436 : 238 - 0xee
      12'h59D: dout <= 8'b11101110; // 1437 : 238 - 0xee
      12'h59E: dout <= 8'b11101110; // 1438 : 238 - 0xee
      12'h59F: dout <= 8'b11101110; // 1439 : 238 - 0xee
      12'h5A0: dout <= 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0x5a
      12'h5A1: dout <= 8'b11111111; // 1441 : 255 - 0xff
      12'h5A2: dout <= 8'b10000011; // 1442 : 131 - 0x83
      12'h5A3: dout <= 8'b00000001; // 1443 :   1 - 0x1
      12'h5A4: dout <= 8'b11101110; // 1444 : 238 - 0xee
      12'h5A5: dout <= 8'b00000000; // 1445 :   0 - 0x0
      12'h5A6: dout <= 8'b11101110; // 1446 : 238 - 0xee
      12'h5A7: dout <= 8'b11101110; // 1447 : 238 - 0xee
      12'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0 -- plane 1
      12'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      12'h5AA: dout <= 8'b01111100; // 1450 : 124 - 0x7c
      12'h5AB: dout <= 8'b11111110; // 1451 : 254 - 0xfe
      12'h5AC: dout <= 8'b11101110; // 1452 : 238 - 0xee
      12'h5AD: dout <= 8'b11101110; // 1453 : 238 - 0xee
      12'h5AE: dout <= 8'b11101110; // 1454 : 238 - 0xee
      12'h5AF: dout <= 8'b11101110; // 1455 : 238 - 0xee
      12'h5B0: dout <= 8'b11111111; // 1456 : 255 - 0xff -- Sprite 0x5b
      12'h5B1: dout <= 8'b11111111; // 1457 : 255 - 0xff
      12'h5B2: dout <= 8'b00000001; // 1458 :   1 - 0x1
      12'h5B3: dout <= 8'b00000000; // 1459 :   0 - 0x0
      12'h5B4: dout <= 8'b11100000; // 1460 : 224 - 0xe0
      12'h5B5: dout <= 8'b00001111; // 1461 :  15 - 0xf
      12'h5B6: dout <= 8'b11111111; // 1462 : 255 - 0xff
      12'h5B7: dout <= 8'b11111011; // 1463 : 251 - 0xfb
      12'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0 -- plane 1
      12'h5B9: dout <= 8'b00000000; // 1465 :   0 - 0x0
      12'h5BA: dout <= 8'b11111110; // 1466 : 254 - 0xfe
      12'h5BB: dout <= 8'b11111110; // 1467 : 254 - 0xfe
      12'h5BC: dout <= 8'b11100000; // 1468 : 224 - 0xe0
      12'h5BD: dout <= 8'b11100000; // 1469 : 224 - 0xe0
      12'h5BE: dout <= 8'b11111000; // 1470 : 248 - 0xf8
      12'h5BF: dout <= 8'b11111000; // 1471 : 248 - 0xf8
      12'h5C0: dout <= 8'b11111111; // 1472 : 255 - 0xff -- Sprite 0x5c
      12'h5C1: dout <= 8'b11111111; // 1473 : 255 - 0xff
      12'h5C2: dout <= 8'b11111111; // 1474 : 255 - 0xff
      12'h5C3: dout <= 8'b11111111; // 1475 : 255 - 0xff
      12'h5C4: dout <= 8'b11111111; // 1476 : 255 - 0xff
      12'h5C5: dout <= 8'b11111111; // 1477 : 255 - 0xff
      12'h5C6: dout <= 8'b11111111; // 1478 : 255 - 0xff
      12'h5C7: dout <= 8'b11011101; // 1479 : 221 - 0xdd
      12'h5C8: dout <= 8'b00000000; // 1480 :   0 - 0x0 -- plane 1
      12'h5C9: dout <= 8'b00000000; // 1481 :   0 - 0x0
      12'h5CA: dout <= 8'b00000000; // 1482 :   0 - 0x0
      12'h5CB: dout <= 8'b00000000; // 1483 :   0 - 0x0
      12'h5CC: dout <= 8'b00000000; // 1484 :   0 - 0x0
      12'h5CD: dout <= 8'b00000000; // 1485 :   0 - 0x0
      12'h5CE: dout <= 8'b11001100; // 1486 : 204 - 0xcc
      12'h5CF: dout <= 8'b11001100; // 1487 : 204 - 0xcc
      12'h5D0: dout <= 8'b11111111; // 1488 : 255 - 0xff -- Sprite 0x5d
      12'h5D1: dout <= 8'b11111111; // 1489 : 255 - 0xff
      12'h5D2: dout <= 8'b00000001; // 1490 :   1 - 0x1
      12'h5D3: dout <= 8'b00000000; // 1491 :   0 - 0x0
      12'h5D4: dout <= 8'b11100000; // 1492 : 224 - 0xe0
      12'h5D5: dout <= 8'b00001111; // 1493 :  15 - 0xf
      12'h5D6: dout <= 8'b11111111; // 1494 : 255 - 0xff
      12'h5D7: dout <= 8'b11111011; // 1495 : 251 - 0xfb
      12'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0 -- plane 1
      12'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout <= 8'b11111110; // 1498 : 254 - 0xfe
      12'h5DB: dout <= 8'b11111110; // 1499 : 254 - 0xfe
      12'h5DC: dout <= 8'b11100000; // 1500 : 224 - 0xe0
      12'h5DD: dout <= 8'b11100000; // 1501 : 224 - 0xe0
      12'h5DE: dout <= 8'b11111000; // 1502 : 248 - 0xf8
      12'h5DF: dout <= 8'b11111000; // 1503 : 248 - 0xf8
      12'h5E0: dout <= 8'b11111111; // 1504 : 255 - 0xff -- Sprite 0x5e
      12'h5E1: dout <= 8'b11111111; // 1505 : 255 - 0xff
      12'h5E2: dout <= 8'b00010001; // 1506 :  17 - 0x11
      12'h5E3: dout <= 8'b00000000; // 1507 :   0 - 0x0
      12'h5E4: dout <= 8'b11101110; // 1508 : 238 - 0xee
      12'h5E5: dout <= 8'b00000000; // 1509 :   0 - 0x0
      12'h5E6: dout <= 8'b11101110; // 1510 : 238 - 0xee
      12'h5E7: dout <= 8'b11101110; // 1511 : 238 - 0xee
      12'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0 -- plane 1
      12'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      12'h5EA: dout <= 8'b11101110; // 1514 : 238 - 0xee
      12'h5EB: dout <= 8'b11101110; // 1515 : 238 - 0xee
      12'h5EC: dout <= 8'b11101110; // 1516 : 238 - 0xee
      12'h5ED: dout <= 8'b11101110; // 1517 : 238 - 0xee
      12'h5EE: dout <= 8'b11101110; // 1518 : 238 - 0xee
      12'h5EF: dout <= 8'b11101110; // 1519 : 238 - 0xee
      12'h5F0: dout <= 8'b10111101; // 1520 : 189 - 0xbd -- Sprite 0x5f
      12'h5F1: dout <= 8'b11111111; // 1521 : 255 - 0xff
      12'h5F2: dout <= 8'b11111111; // 1522 : 255 - 0xff
      12'h5F3: dout <= 8'b11111111; // 1523 : 255 - 0xff
      12'h5F4: dout <= 8'b11111111; // 1524 : 255 - 0xff
      12'h5F5: dout <= 8'b11111111; // 1525 : 255 - 0xff
      12'h5F6: dout <= 8'b11111111; // 1526 : 255 - 0xff
      12'h5F7: dout <= 8'b11111111; // 1527 : 255 - 0xff
      12'h5F8: dout <= 8'b01111110; // 1528 : 126 - 0x7e -- plane 1
      12'h5F9: dout <= 8'b01111110; // 1529 : 126 - 0x7e
      12'h5FA: dout <= 8'b01111110; // 1530 : 126 - 0x7e
      12'h5FB: dout <= 8'b01111110; // 1531 : 126 - 0x7e
      12'h5FC: dout <= 8'b01111110; // 1532 : 126 - 0x7e
      12'h5FD: dout <= 8'b01111110; // 1533 : 126 - 0x7e
      12'h5FE: dout <= 8'b01111110; // 1534 : 126 - 0x7e
      12'h5FF: dout <= 8'b01111110; // 1535 : 126 - 0x7e
      12'h600: dout <= 8'b11101110; // 1536 : 238 - 0xee -- Sprite 0x60
      12'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout <= 8'b11111110; // 1538 : 254 - 0xfe
      12'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      12'h604: dout <= 8'b00000001; // 1540 :   1 - 0x1
      12'h605: dout <= 8'b00001111; // 1541 :  15 - 0xf
      12'h606: dout <= 8'b10001111; // 1542 : 143 - 0x8f
      12'h607: dout <= 8'b11111111; // 1543 : 255 - 0xff
      12'h608: dout <= 8'b11101110; // 1544 : 238 - 0xee -- plane 1
      12'h609: dout <= 8'b11101110; // 1545 : 238 - 0xee
      12'h60A: dout <= 8'b11111110; // 1546 : 254 - 0xfe
      12'h60B: dout <= 8'b11111100; // 1547 : 252 - 0xfc
      12'h60C: dout <= 8'b11100000; // 1548 : 224 - 0xe0
      12'h60D: dout <= 8'b11100000; // 1549 : 224 - 0xe0
      12'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      12'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout <= 8'b11101110; // 1552 : 238 - 0xee -- Sprite 0x61
      12'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      12'h612: dout <= 8'b11111100; // 1554 : 252 - 0xfc
      12'h613: dout <= 8'b00000001; // 1555 :   1 - 0x1
      12'h614: dout <= 8'b00000001; // 1556 :   1 - 0x1
      12'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      12'h616: dout <= 8'b10001000; // 1558 : 136 - 0x88
      12'h617: dout <= 8'b11111111; // 1559 : 255 - 0xff
      12'h618: dout <= 8'b11101110; // 1560 : 238 - 0xee -- plane 1
      12'h619: dout <= 8'b11101110; // 1561 : 238 - 0xee
      12'h61A: dout <= 8'b11111100; // 1562 : 252 - 0xfc
      12'h61B: dout <= 8'b11111100; // 1563 : 252 - 0xfc
      12'h61C: dout <= 8'b11101110; // 1564 : 238 - 0xee
      12'h61D: dout <= 8'b11101110; // 1565 : 238 - 0xee
      12'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      12'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout <= 8'b11100011; // 1568 : 227 - 0xe3 -- Sprite 0x62
      12'h621: dout <= 8'b00001111; // 1569 :  15 - 0xf
      12'h622: dout <= 8'b11101111; // 1570 : 239 - 0xef
      12'h623: dout <= 8'b00001111; // 1571 :  15 - 0xf
      12'h624: dout <= 8'b00000001; // 1572 :   1 - 0x1
      12'h625: dout <= 8'b00000000; // 1573 :   0 - 0x0
      12'h626: dout <= 8'b10000000; // 1574 : 128 - 0x80
      12'h627: dout <= 8'b11111111; // 1575 : 255 - 0xff
      12'h628: dout <= 8'b11100000; // 1576 : 224 - 0xe0 -- plane 1
      12'h629: dout <= 8'b11100000; // 1577 : 224 - 0xe0
      12'h62A: dout <= 8'b11100000; // 1578 : 224 - 0xe0
      12'h62B: dout <= 8'b11100000; // 1579 : 224 - 0xe0
      12'h62C: dout <= 8'b11111110; // 1580 : 254 - 0xfe
      12'h62D: dout <= 8'b11111110; // 1581 : 254 - 0xfe
      12'h62E: dout <= 8'b00000000; // 1582 :   0 - 0x0
      12'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout <= 8'b11001110; // 1584 : 206 - 0xce -- Sprite 0x63
      12'h631: dout <= 8'b11110000; // 1585 : 240 - 0xf0
      12'h632: dout <= 8'b11111110; // 1586 : 254 - 0xfe
      12'h633: dout <= 8'b00010000; // 1587 :  16 - 0x10
      12'h634: dout <= 8'b00000000; // 1588 :   0 - 0x0
      12'h635: dout <= 8'b10000000; // 1589 : 128 - 0x80
      12'h636: dout <= 8'b11000001; // 1590 : 193 - 0xc1
      12'h637: dout <= 8'b11111111; // 1591 : 255 - 0xff
      12'h638: dout <= 8'b00001110; // 1592 :  14 - 0xe -- plane 1
      12'h639: dout <= 8'b00001110; // 1593 :  14 - 0xe
      12'h63A: dout <= 8'b00001110; // 1594 :  14 - 0xe
      12'h63B: dout <= 8'b11101110; // 1595 : 238 - 0xee
      12'h63C: dout <= 8'b11111110; // 1596 : 254 - 0xfe
      12'h63D: dout <= 8'b01111100; // 1597 : 124 - 0x7c
      12'h63E: dout <= 8'b00000000; // 1598 :   0 - 0x0
      12'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout <= 8'b11111011; // 1600 : 251 - 0xfb -- Sprite 0x64
      12'h641: dout <= 8'b11000011; // 1601 : 195 - 0xc3
      12'h642: dout <= 8'b11111011; // 1602 : 251 - 0xfb
      12'h643: dout <= 8'b11000011; // 1603 : 195 - 0xc3
      12'h644: dout <= 8'b11000011; // 1604 : 195 - 0xc3
      12'h645: dout <= 8'b11000011; // 1605 : 195 - 0xc3
      12'h646: dout <= 8'b11100011; // 1606 : 227 - 0xe3
      12'h647: dout <= 8'b11111111; // 1607 : 255 - 0xff
      12'h648: dout <= 8'b00111000; // 1608 :  56 - 0x38 -- plane 1
      12'h649: dout <= 8'b00111000; // 1609 :  56 - 0x38
      12'h64A: dout <= 8'b00111000; // 1610 :  56 - 0x38
      12'h64B: dout <= 8'b00111000; // 1611 :  56 - 0x38
      12'h64C: dout <= 8'b00111000; // 1612 :  56 - 0x38
      12'h64D: dout <= 8'b00111000; // 1613 :  56 - 0x38
      12'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout <= 8'b11101110; // 1616 : 238 - 0xee -- Sprite 0x65
      12'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      12'h652: dout <= 8'b11111110; // 1618 : 254 - 0xfe
      12'h653: dout <= 8'b00000000; // 1619 :   0 - 0x0
      12'h654: dout <= 8'b00000000; // 1620 :   0 - 0x0
      12'h655: dout <= 8'b00000000; // 1621 :   0 - 0x0
      12'h656: dout <= 8'b10001000; // 1622 : 136 - 0x88
      12'h657: dout <= 8'b11111111; // 1623 : 255 - 0xff
      12'h658: dout <= 8'b11101110; // 1624 : 238 - 0xee -- plane 1
      12'h659: dout <= 8'b11101110; // 1625 : 238 - 0xee
      12'h65A: dout <= 8'b11111110; // 1626 : 254 - 0xfe
      12'h65B: dout <= 8'b11111110; // 1627 : 254 - 0xfe
      12'h65C: dout <= 8'b11101110; // 1628 : 238 - 0xee
      12'h65D: dout <= 8'b11101110; // 1629 : 238 - 0xee
      12'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout <= 8'b11101111; // 1632 : 239 - 0xef -- Sprite 0x66
      12'h661: dout <= 8'b00001111; // 1633 :  15 - 0xf
      12'h662: dout <= 8'b11101111; // 1634 : 239 - 0xef
      12'h663: dout <= 8'b00000001; // 1635 :   1 - 0x1
      12'h664: dout <= 8'b00000000; // 1636 :   0 - 0x0
      12'h665: dout <= 8'b00000000; // 1637 :   0 - 0x0
      12'h666: dout <= 8'b10000000; // 1638 : 128 - 0x80
      12'h667: dout <= 8'b11111111; // 1639 : 255 - 0xff
      12'h668: dout <= 8'b11100000; // 1640 : 224 - 0xe0 -- plane 1
      12'h669: dout <= 8'b11100000; // 1641 : 224 - 0xe0
      12'h66A: dout <= 8'b11100000; // 1642 : 224 - 0xe0
      12'h66B: dout <= 8'b11101110; // 1643 : 238 - 0xee
      12'h66C: dout <= 8'b11111110; // 1644 : 254 - 0xfe
      12'h66D: dout <= 8'b11111110; // 1645 : 254 - 0xfe
      12'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      12'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      12'h670: dout <= 8'b11101110; // 1648 : 238 - 0xee -- Sprite 0x67
      12'h671: dout <= 8'b00000000; // 1649 :   0 - 0x0
      12'h672: dout <= 8'b11111110; // 1650 : 254 - 0xfe
      12'h673: dout <= 8'b00000000; // 1651 :   0 - 0x0
      12'h674: dout <= 8'b00000000; // 1652 :   0 - 0x0
      12'h675: dout <= 8'b00001000; // 1653 :   8 - 0x8
      12'h676: dout <= 8'b10011100; // 1654 : 156 - 0x9c
      12'h677: dout <= 8'b11111111; // 1655 : 255 - 0xff
      12'h678: dout <= 8'b11101110; // 1656 : 238 - 0xee -- plane 1
      12'h679: dout <= 8'b11101110; // 1657 : 238 - 0xee
      12'h67A: dout <= 8'b11111110; // 1658 : 254 - 0xfe
      12'h67B: dout <= 8'b11111110; // 1659 : 254 - 0xfe
      12'h67C: dout <= 8'b11101110; // 1660 : 238 - 0xee
      12'h67D: dout <= 8'b11000110; // 1661 : 198 - 0xc6
      12'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout <= 8'b11101110; // 1664 : 238 - 0xee -- Sprite 0x68
      12'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout <= 8'b11101110; // 1666 : 238 - 0xee
      12'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      12'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      12'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      12'h686: dout <= 8'b10001000; // 1670 : 136 - 0x88
      12'h687: dout <= 8'b11111111; // 1671 : 255 - 0xff
      12'h688: dout <= 8'b11101110; // 1672 : 238 - 0xee -- plane 1
      12'h689: dout <= 8'b11101110; // 1673 : 238 - 0xee
      12'h68A: dout <= 8'b11101110; // 1674 : 238 - 0xee
      12'h68B: dout <= 8'b11101110; // 1675 : 238 - 0xee
      12'h68C: dout <= 8'b11101110; // 1676 : 238 - 0xee
      12'h68D: dout <= 8'b11101110; // 1677 : 238 - 0xee
      12'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      12'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout <= 8'b11101110; // 1680 : 238 - 0xee -- Sprite 0x69
      12'h691: dout <= 8'b00000000; // 1681 :   0 - 0x0
      12'h692: dout <= 8'b11101110; // 1682 : 238 - 0xee
      12'h693: dout <= 8'b00000000; // 1683 :   0 - 0x0
      12'h694: dout <= 8'b00000000; // 1684 :   0 - 0x0
      12'h695: dout <= 8'b00000000; // 1685 :   0 - 0x0
      12'h696: dout <= 8'b10000001; // 1686 : 129 - 0x81
      12'h697: dout <= 8'b11111111; // 1687 : 255 - 0xff
      12'h698: dout <= 8'b11101110; // 1688 : 238 - 0xee -- plane 1
      12'h699: dout <= 8'b11101110; // 1689 : 238 - 0xee
      12'h69A: dout <= 8'b11101110; // 1690 : 238 - 0xee
      12'h69B: dout <= 8'b11101110; // 1691 : 238 - 0xee
      12'h69C: dout <= 8'b11111110; // 1692 : 254 - 0xfe
      12'h69D: dout <= 8'b11111100; // 1693 : 252 - 0xfc
      12'h69E: dout <= 8'b00000000; // 1694 :   0 - 0x0
      12'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      12'h6A0: dout <= 8'b11101110; // 1696 : 238 - 0xee -- Sprite 0x6a
      12'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout <= 8'b11101110; // 1698 : 238 - 0xee
      12'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      12'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      12'h6A5: dout <= 8'b10000000; // 1701 : 128 - 0x80
      12'h6A6: dout <= 8'b11000001; // 1702 : 193 - 0xc1
      12'h6A7: dout <= 8'b11111111; // 1703 : 255 - 0xff
      12'h6A8: dout <= 8'b11101110; // 1704 : 238 - 0xee -- plane 1
      12'h6A9: dout <= 8'b11101110; // 1705 : 238 - 0xee
      12'h6AA: dout <= 8'b11101110; // 1706 : 238 - 0xee
      12'h6AB: dout <= 8'b11101110; // 1707 : 238 - 0xee
      12'h6AC: dout <= 8'b11111110; // 1708 : 254 - 0xfe
      12'h6AD: dout <= 8'b01111100; // 1709 : 124 - 0x7c
      12'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      12'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout <= 8'b11100011; // 1712 : 227 - 0xe3 -- Sprite 0x6b
      12'h6B1: dout <= 8'b00001111; // 1713 :  15 - 0xf
      12'h6B2: dout <= 8'b11101111; // 1714 : 239 - 0xef
      12'h6B3: dout <= 8'b00001111; // 1715 :  15 - 0xf
      12'h6B4: dout <= 8'b00000001; // 1716 :   1 - 0x1
      12'h6B5: dout <= 8'b00000000; // 1717 :   0 - 0x0
      12'h6B6: dout <= 8'b10000000; // 1718 : 128 - 0x80
      12'h6B7: dout <= 8'b11111111; // 1719 : 255 - 0xff
      12'h6B8: dout <= 8'b11100000; // 1720 : 224 - 0xe0 -- plane 1
      12'h6B9: dout <= 8'b11100000; // 1721 : 224 - 0xe0
      12'h6BA: dout <= 8'b11100000; // 1722 : 224 - 0xe0
      12'h6BB: dout <= 8'b11100000; // 1723 : 224 - 0xe0
      12'h6BC: dout <= 8'b11111110; // 1724 : 254 - 0xfe
      12'h6BD: dout <= 8'b11111110; // 1725 : 254 - 0xfe
      12'h6BE: dout <= 8'b00000000; // 1726 :   0 - 0x0
      12'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout <= 8'b10011001; // 1728 : 153 - 0x99 -- Sprite 0x6c
      12'h6C1: dout <= 8'b11100011; // 1729 : 227 - 0xe3
      12'h6C2: dout <= 8'b11110011; // 1730 : 243 - 0xf3
      12'h6C3: dout <= 8'b11000111; // 1731 : 199 - 0xc7
      12'h6C4: dout <= 8'b10000001; // 1732 : 129 - 0x81
      12'h6C5: dout <= 8'b10001000; // 1733 : 136 - 0x88
      12'h6C6: dout <= 8'b11001100; // 1734 : 204 - 0xcc
      12'h6C7: dout <= 8'b11111111; // 1735 : 255 - 0xff
      12'h6C8: dout <= 8'b00011000; // 1736 :  24 - 0x18 -- plane 1
      12'h6C9: dout <= 8'b00011000; // 1737 :  24 - 0x18
      12'h6CA: dout <= 8'b00110000; // 1738 :  48 - 0x30
      12'h6CB: dout <= 8'b00110000; // 1739 :  48 - 0x30
      12'h6CC: dout <= 8'b01100110; // 1740 : 102 - 0x66
      12'h6CD: dout <= 8'b01100110; // 1741 : 102 - 0x66
      12'h6CE: dout <= 8'b00000000; // 1742 :   0 - 0x0
      12'h6CF: dout <= 8'b00000000; // 1743 :   0 - 0x0
      12'h6D0: dout <= 8'b11100011; // 1744 : 227 - 0xe3 -- Sprite 0x6d
      12'h6D1: dout <= 8'b00001111; // 1745 :  15 - 0xf
      12'h6D2: dout <= 8'b11101111; // 1746 : 239 - 0xef
      12'h6D3: dout <= 8'b00001111; // 1747 :  15 - 0xf
      12'h6D4: dout <= 8'b00001111; // 1748 :  15 - 0xf
      12'h6D5: dout <= 8'b00001111; // 1749 :  15 - 0xf
      12'h6D6: dout <= 8'b10001111; // 1750 : 143 - 0x8f
      12'h6D7: dout <= 8'b11111111; // 1751 : 255 - 0xff
      12'h6D8: dout <= 8'b11100000; // 1752 : 224 - 0xe0 -- plane 1
      12'h6D9: dout <= 8'b11100000; // 1753 : 224 - 0xe0
      12'h6DA: dout <= 8'b11100000; // 1754 : 224 - 0xe0
      12'h6DB: dout <= 8'b11100000; // 1755 : 224 - 0xe0
      12'h6DC: dout <= 8'b11100000; // 1756 : 224 - 0xe0
      12'h6DD: dout <= 8'b11100000; // 1757 : 224 - 0xe0
      12'h6DE: dout <= 8'b00000000; // 1758 :   0 - 0x0
      12'h6DF: dout <= 8'b00000000; // 1759 :   0 - 0x0
      12'h6E0: dout <= 8'b11101110; // 1760 : 238 - 0xee -- Sprite 0x6e
      12'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout <= 8'b11101110; // 1762 : 238 - 0xee
      12'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      12'h6E5: dout <= 8'b10000000; // 1765 : 128 - 0x80
      12'h6E6: dout <= 8'b11000001; // 1766 : 193 - 0xc1
      12'h6E7: dout <= 8'b11111111; // 1767 : 255 - 0xff
      12'h6E8: dout <= 8'b11101110; // 1768 : 238 - 0xee -- plane 1
      12'h6E9: dout <= 8'b11101110; // 1769 : 238 - 0xee
      12'h6EA: dout <= 8'b11101110; // 1770 : 238 - 0xee
      12'h6EB: dout <= 8'b11101110; // 1771 : 238 - 0xee
      12'h6EC: dout <= 8'b11111110; // 1772 : 254 - 0xfe
      12'h6ED: dout <= 8'b01111100; // 1773 : 124 - 0x7c
      12'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      12'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      12'h6F0: dout <= 8'b11111111; // 1776 : 255 - 0xff -- Sprite 0x6f
      12'h6F1: dout <= 8'b11111111; // 1777 : 255 - 0xff
      12'h6F2: dout <= 8'b11111111; // 1778 : 255 - 0xff
      12'h6F3: dout <= 8'b10111101; // 1779 : 189 - 0xbd
      12'h6F4: dout <= 8'b11111111; // 1780 : 255 - 0xff
      12'h6F5: dout <= 8'b11011011; // 1781 : 219 - 0xdb
      12'h6F6: dout <= 8'b11111111; // 1782 : 255 - 0xff
      12'h6F7: dout <= 8'b11111111; // 1783 : 255 - 0xff
      12'h6F8: dout <= 8'b01111110; // 1784 : 126 - 0x7e -- plane 1
      12'h6F9: dout <= 8'b01111110; // 1785 : 126 - 0x7e
      12'h6FA: dout <= 8'b01111110; // 1786 : 126 - 0x7e
      12'h6FB: dout <= 8'b01111110; // 1787 : 126 - 0x7e
      12'h6FC: dout <= 8'b00111100; // 1788 :  60 - 0x3c
      12'h6FD: dout <= 8'b00111100; // 1789 :  60 - 0x3c
      12'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      12'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout <= 8'b11111011; // 1792 : 251 - 0xfb -- Sprite 0x70
      12'h701: dout <= 8'b11101111; // 1793 : 239 - 0xef
      12'h702: dout <= 8'b11011111; // 1794 : 223 - 0xdf
      12'h703: dout <= 8'b11111111; // 1795 : 255 - 0xff
      12'h704: dout <= 8'b10111111; // 1796 : 191 - 0xbf
      12'h705: dout <= 8'b10111111; // 1797 : 191 - 0xbf
      12'h706: dout <= 8'b11111110; // 1798 : 254 - 0xfe
      12'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      12'h708: dout <= 8'b00000111; // 1800 :   7 - 0x7 -- plane 1
      12'h709: dout <= 8'b00011111; // 1801 :  31 - 0x1f
      12'h70A: dout <= 8'b00111111; // 1802 :  63 - 0x3f
      12'h70B: dout <= 8'b00111111; // 1803 :  63 - 0x3f
      12'h70C: dout <= 8'b01111111; // 1804 : 127 - 0x7f
      12'h70D: dout <= 8'b01111111; // 1805 : 127 - 0x7f
      12'h70E: dout <= 8'b01111111; // 1806 : 127 - 0x7f
      12'h70F: dout <= 8'b01111110; // 1807 : 126 - 0x7e
      12'h710: dout <= 8'b11011111; // 1808 : 223 - 0xdf -- Sprite 0x71
      12'h711: dout <= 8'b11110111; // 1809 : 247 - 0xf7
      12'h712: dout <= 8'b11111011; // 1810 : 251 - 0xfb
      12'h713: dout <= 8'b11111111; // 1811 : 255 - 0xff
      12'h714: dout <= 8'b11111101; // 1812 : 253 - 0xfd
      12'h715: dout <= 8'b11111101; // 1813 : 253 - 0xfd
      12'h716: dout <= 8'b01111111; // 1814 : 127 - 0x7f
      12'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      12'h718: dout <= 8'b11100000; // 1816 : 224 - 0xe0 -- plane 1
      12'h719: dout <= 8'b11111000; // 1817 : 248 - 0xf8
      12'h71A: dout <= 8'b11111100; // 1818 : 252 - 0xfc
      12'h71B: dout <= 8'b11111100; // 1819 : 252 - 0xfc
      12'h71C: dout <= 8'b11111110; // 1820 : 254 - 0xfe
      12'h71D: dout <= 8'b11111110; // 1821 : 254 - 0xfe
      12'h71E: dout <= 8'b11111110; // 1822 : 254 - 0xfe
      12'h71F: dout <= 8'b01111110; // 1823 : 126 - 0x7e
      12'h720: dout <= 8'b11111111; // 1824 : 255 - 0xff -- Sprite 0x72
      12'h721: dout <= 8'b11111111; // 1825 : 255 - 0xff
      12'h722: dout <= 8'b11111111; // 1826 : 255 - 0xff
      12'h723: dout <= 8'b11111111; // 1827 : 255 - 0xff
      12'h724: dout <= 8'b11111111; // 1828 : 255 - 0xff
      12'h725: dout <= 8'b11111111; // 1829 : 255 - 0xff
      12'h726: dout <= 8'b11111111; // 1830 : 255 - 0xff
      12'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      12'h728: dout <= 8'b01111110; // 1832 : 126 - 0x7e -- plane 1
      12'h729: dout <= 8'b01111110; // 1833 : 126 - 0x7e
      12'h72A: dout <= 8'b01111110; // 1834 : 126 - 0x7e
      12'h72B: dout <= 8'b01111110; // 1835 : 126 - 0x7e
      12'h72C: dout <= 8'b01111110; // 1836 : 126 - 0x7e
      12'h72D: dout <= 8'b01111110; // 1837 : 126 - 0x7e
      12'h72E: dout <= 8'b01111110; // 1838 : 126 - 0x7e
      12'h72F: dout <= 8'b01111110; // 1839 : 126 - 0x7e
      12'h730: dout <= 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0x73
      12'h731: dout <= 8'b11111110; // 1841 : 254 - 0xfe
      12'h732: dout <= 8'b10111111; // 1842 : 191 - 0xbf
      12'h733: dout <= 8'b10111111; // 1843 : 191 - 0xbf
      12'h734: dout <= 8'b11111111; // 1844 : 255 - 0xff
      12'h735: dout <= 8'b11011111; // 1845 : 223 - 0xdf
      12'h736: dout <= 8'b11101111; // 1846 : 239 - 0xef
      12'h737: dout <= 8'b11111011; // 1847 : 251 - 0xfb
      12'h738: dout <= 8'b01111110; // 1848 : 126 - 0x7e -- plane 1
      12'h739: dout <= 8'b01111111; // 1849 : 127 - 0x7f
      12'h73A: dout <= 8'b01111111; // 1850 : 127 - 0x7f
      12'h73B: dout <= 8'b01111111; // 1851 : 127 - 0x7f
      12'h73C: dout <= 8'b00111111; // 1852 :  63 - 0x3f
      12'h73D: dout <= 8'b00111111; // 1853 :  63 - 0x3f
      12'h73E: dout <= 8'b00011111; // 1854 :  31 - 0x1f
      12'h73F: dout <= 8'b00000111; // 1855 :   7 - 0x7
      12'h740: dout <= 8'b11111111; // 1856 : 255 - 0xff -- Sprite 0x74
      12'h741: dout <= 8'b01111111; // 1857 : 127 - 0x7f
      12'h742: dout <= 8'b11111101; // 1858 : 253 - 0xfd
      12'h743: dout <= 8'b11111101; // 1859 : 253 - 0xfd
      12'h744: dout <= 8'b11111111; // 1860 : 255 - 0xff
      12'h745: dout <= 8'b11111011; // 1861 : 251 - 0xfb
      12'h746: dout <= 8'b11110111; // 1862 : 247 - 0xf7
      12'h747: dout <= 8'b11011111; // 1863 : 223 - 0xdf
      12'h748: dout <= 8'b01111110; // 1864 : 126 - 0x7e -- plane 1
      12'h749: dout <= 8'b11111110; // 1865 : 254 - 0xfe
      12'h74A: dout <= 8'b11111110; // 1866 : 254 - 0xfe
      12'h74B: dout <= 8'b11111110; // 1867 : 254 - 0xfe
      12'h74C: dout <= 8'b11111100; // 1868 : 252 - 0xfc
      12'h74D: dout <= 8'b11111100; // 1869 : 252 - 0xfc
      12'h74E: dout <= 8'b11111000; // 1870 : 248 - 0xf8
      12'h74F: dout <= 8'b11100000; // 1871 : 224 - 0xe0
      12'h750: dout <= 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0x75
      12'h751: dout <= 8'b11111111; // 1873 : 255 - 0xff
      12'h752: dout <= 8'b11111111; // 1874 : 255 - 0xff
      12'h753: dout <= 8'b11111111; // 1875 : 255 - 0xff
      12'h754: dout <= 8'b11111111; // 1876 : 255 - 0xff
      12'h755: dout <= 8'b11111111; // 1877 : 255 - 0xff
      12'h756: dout <= 8'b11111111; // 1878 : 255 - 0xff
      12'h757: dout <= 8'b11111111; // 1879 : 255 - 0xff
      12'h758: dout <= 8'b01111111; // 1880 : 127 - 0x7f -- plane 1
      12'h759: dout <= 8'b01111111; // 1881 : 127 - 0x7f
      12'h75A: dout <= 8'b01111111; // 1882 : 127 - 0x7f
      12'h75B: dout <= 8'b01111111; // 1883 : 127 - 0x7f
      12'h75C: dout <= 8'b01111111; // 1884 : 127 - 0x7f
      12'h75D: dout <= 8'b01111111; // 1885 : 127 - 0x7f
      12'h75E: dout <= 8'b00000111; // 1886 :   7 - 0x7
      12'h75F: dout <= 8'b00000111; // 1887 :   7 - 0x7
      12'h760: dout <= 8'b11111111; // 1888 : 255 - 0xff -- Sprite 0x76
      12'h761: dout <= 8'b11111111; // 1889 : 255 - 0xff
      12'h762: dout <= 8'b11111111; // 1890 : 255 - 0xff
      12'h763: dout <= 8'b11111111; // 1891 : 255 - 0xff
      12'h764: dout <= 8'b11111111; // 1892 : 255 - 0xff
      12'h765: dout <= 8'b11111111; // 1893 : 255 - 0xff
      12'h766: dout <= 8'b11111111; // 1894 : 255 - 0xff
      12'h767: dout <= 8'b11111111; // 1895 : 255 - 0xff
      12'h768: dout <= 8'b11111110; // 1896 : 254 - 0xfe -- plane 1
      12'h769: dout <= 8'b11111110; // 1897 : 254 - 0xfe
      12'h76A: dout <= 8'b11111110; // 1898 : 254 - 0xfe
      12'h76B: dout <= 8'b11111110; // 1899 : 254 - 0xfe
      12'h76C: dout <= 8'b11111110; // 1900 : 254 - 0xfe
      12'h76D: dout <= 8'b11111110; // 1901 : 254 - 0xfe
      12'h76E: dout <= 8'b11100000; // 1902 : 224 - 0xe0
      12'h76F: dout <= 8'b11100000; // 1903 : 224 - 0xe0
      12'h770: dout <= 8'b11111111; // 1904 : 255 - 0xff -- Sprite 0x77
      12'h771: dout <= 8'b11111111; // 1905 : 255 - 0xff
      12'h772: dout <= 8'b11111111; // 1906 : 255 - 0xff
      12'h773: dout <= 8'b11111111; // 1907 : 255 - 0xff
      12'h774: dout <= 8'b11111111; // 1908 : 255 - 0xff
      12'h775: dout <= 8'b11111111; // 1909 : 255 - 0xff
      12'h776: dout <= 8'b11111111; // 1910 : 255 - 0xff
      12'h777: dout <= 8'b11111111; // 1911 : 255 - 0xff
      12'h778: dout <= 8'b00000111; // 1912 :   7 - 0x7 -- plane 1
      12'h779: dout <= 8'b00000111; // 1913 :   7 - 0x7
      12'h77A: dout <= 8'b00000111; // 1914 :   7 - 0x7
      12'h77B: dout <= 8'b00000111; // 1915 :   7 - 0x7
      12'h77C: dout <= 8'b00000111; // 1916 :   7 - 0x7
      12'h77D: dout <= 8'b00000111; // 1917 :   7 - 0x7
      12'h77E: dout <= 8'b00000111; // 1918 :   7 - 0x7
      12'h77F: dout <= 8'b00000111; // 1919 :   7 - 0x7
      12'h780: dout <= 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0x78
      12'h781: dout <= 8'b11111111; // 1921 : 255 - 0xff
      12'h782: dout <= 8'b11111111; // 1922 : 255 - 0xff
      12'h783: dout <= 8'b11111111; // 1923 : 255 - 0xff
      12'h784: dout <= 8'b11111111; // 1924 : 255 - 0xff
      12'h785: dout <= 8'b11111111; // 1925 : 255 - 0xff
      12'h786: dout <= 8'b11111111; // 1926 : 255 - 0xff
      12'h787: dout <= 8'b11111111; // 1927 : 255 - 0xff
      12'h788: dout <= 8'b11100000; // 1928 : 224 - 0xe0 -- plane 1
      12'h789: dout <= 8'b11100000; // 1929 : 224 - 0xe0
      12'h78A: dout <= 8'b11100000; // 1930 : 224 - 0xe0
      12'h78B: dout <= 8'b11100000; // 1931 : 224 - 0xe0
      12'h78C: dout <= 8'b11100000; // 1932 : 224 - 0xe0
      12'h78D: dout <= 8'b11100000; // 1933 : 224 - 0xe0
      12'h78E: dout <= 8'b11100000; // 1934 : 224 - 0xe0
      12'h78F: dout <= 8'b11100000; // 1935 : 224 - 0xe0
      12'h790: dout <= 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0x79
      12'h791: dout <= 8'b11111111; // 1937 : 255 - 0xff
      12'h792: dout <= 8'b11111111; // 1938 : 255 - 0xff
      12'h793: dout <= 8'b11111111; // 1939 : 255 - 0xff
      12'h794: dout <= 8'b11111111; // 1940 : 255 - 0xff
      12'h795: dout <= 8'b11111111; // 1941 : 255 - 0xff
      12'h796: dout <= 8'b11111111; // 1942 : 255 - 0xff
      12'h797: dout <= 8'b11111111; // 1943 : 255 - 0xff
      12'h798: dout <= 8'b01111111; // 1944 : 127 - 0x7f -- plane 1
      12'h799: dout <= 8'b01111111; // 1945 : 127 - 0x7f
      12'h79A: dout <= 8'b01111111; // 1946 : 127 - 0x7f
      12'h79B: dout <= 8'b01111111; // 1947 : 127 - 0x7f
      12'h79C: dout <= 8'b01111111; // 1948 : 127 - 0x7f
      12'h79D: dout <= 8'b01111111; // 1949 : 127 - 0x7f
      12'h79E: dout <= 8'b01111110; // 1950 : 126 - 0x7e
      12'h79F: dout <= 8'b01111110; // 1951 : 126 - 0x7e
      12'h7A0: dout <= 8'b11111111; // 1952 : 255 - 0xff -- Sprite 0x7a
      12'h7A1: dout <= 8'b11111111; // 1953 : 255 - 0xff
      12'h7A2: dout <= 8'b11111111; // 1954 : 255 - 0xff
      12'h7A3: dout <= 8'b11111111; // 1955 : 255 - 0xff
      12'h7A4: dout <= 8'b11111111; // 1956 : 255 - 0xff
      12'h7A5: dout <= 8'b11111111; // 1957 : 255 - 0xff
      12'h7A6: dout <= 8'b11111111; // 1958 : 255 - 0xff
      12'h7A7: dout <= 8'b11111111; // 1959 : 255 - 0xff
      12'h7A8: dout <= 8'b11111110; // 1960 : 254 - 0xfe -- plane 1
      12'h7A9: dout <= 8'b11111110; // 1961 : 254 - 0xfe
      12'h7AA: dout <= 8'b11111110; // 1962 : 254 - 0xfe
      12'h7AB: dout <= 8'b11111110; // 1963 : 254 - 0xfe
      12'h7AC: dout <= 8'b11111110; // 1964 : 254 - 0xfe
      12'h7AD: dout <= 8'b11111110; // 1965 : 254 - 0xfe
      12'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      12'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout <= 8'b11111111; // 1968 : 255 - 0xff -- Sprite 0x7b
      12'h7B1: dout <= 8'b11111111; // 1969 : 255 - 0xff
      12'h7B2: dout <= 8'b11111111; // 1970 : 255 - 0xff
      12'h7B3: dout <= 8'b11111111; // 1971 : 255 - 0xff
      12'h7B4: dout <= 8'b11111111; // 1972 : 255 - 0xff
      12'h7B5: dout <= 8'b11111111; // 1973 : 255 - 0xff
      12'h7B6: dout <= 8'b11111111; // 1974 : 255 - 0xff
      12'h7B7: dout <= 8'b11111111; // 1975 : 255 - 0xff
      12'h7B8: dout <= 8'b01111110; // 1976 : 126 - 0x7e -- plane 1
      12'h7B9: dout <= 8'b01111111; // 1977 : 127 - 0x7f
      12'h7BA: dout <= 8'b01111111; // 1978 : 127 - 0x7f
      12'h7BB: dout <= 8'b01111111; // 1979 : 127 - 0x7f
      12'h7BC: dout <= 8'b01111111; // 1980 : 127 - 0x7f
      12'h7BD: dout <= 8'b01111111; // 1981 : 127 - 0x7f
      12'h7BE: dout <= 8'b01111111; // 1982 : 127 - 0x7f
      12'h7BF: dout <= 8'b01111110; // 1983 : 126 - 0x7e
      12'h7C0: dout <= 8'b11111111; // 1984 : 255 - 0xff -- Sprite 0x7c
      12'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      12'h7C2: dout <= 8'b11111111; // 1986 : 255 - 0xff
      12'h7C3: dout <= 8'b11111111; // 1987 : 255 - 0xff
      12'h7C4: dout <= 8'b11111111; // 1988 : 255 - 0xff
      12'h7C5: dout <= 8'b11111111; // 1989 : 255 - 0xff
      12'h7C6: dout <= 8'b11111111; // 1990 : 255 - 0xff
      12'h7C7: dout <= 8'b11111111; // 1991 : 255 - 0xff
      12'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0 -- plane 1
      12'h7C9: dout <= 8'b11110000; // 1993 : 240 - 0xf0
      12'h7CA: dout <= 8'b11110000; // 1994 : 240 - 0xf0
      12'h7CB: dout <= 8'b11110000; // 1995 : 240 - 0xf0
      12'h7CC: dout <= 8'b11110000; // 1996 : 240 - 0xf0
      12'h7CD: dout <= 8'b11110000; // 1997 : 240 - 0xf0
      12'h7CE: dout <= 8'b11110000; // 1998 : 240 - 0xf0
      12'h7CF: dout <= 8'b00000000; // 1999 :   0 - 0x0
      12'h7D0: dout <= 8'b11111111; // 2000 : 255 - 0xff -- Sprite 0x7d
      12'h7D1: dout <= 8'b11111111; // 2001 : 255 - 0xff
      12'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      12'h7D3: dout <= 8'b11111111; // 2003 : 255 - 0xff
      12'h7D4: dout <= 8'b11111111; // 2004 : 255 - 0xff
      12'h7D5: dout <= 8'b11111111; // 2005 : 255 - 0xff
      12'h7D6: dout <= 8'b11111111; // 2006 : 255 - 0xff
      12'h7D7: dout <= 8'b11111111; // 2007 : 255 - 0xff
      12'h7D8: dout <= 8'b01111110; // 2008 : 126 - 0x7e -- plane 1
      12'h7D9: dout <= 8'b01111110; // 2009 : 126 - 0x7e
      12'h7DA: dout <= 8'b01111111; // 2010 : 127 - 0x7f
      12'h7DB: dout <= 8'b01111111; // 2011 : 127 - 0x7f
      12'h7DC: dout <= 8'b01111111; // 2012 : 127 - 0x7f
      12'h7DD: dout <= 8'b01111111; // 2013 : 127 - 0x7f
      12'h7DE: dout <= 8'b01111111; // 2014 : 127 - 0x7f
      12'h7DF: dout <= 8'b01111111; // 2015 : 127 - 0x7f
      12'h7E0: dout <= 8'b11111111; // 2016 : 255 - 0xff -- Sprite 0x7e
      12'h7E1: dout <= 8'b11111111; // 2017 : 255 - 0xff
      12'h7E2: dout <= 8'b11111111; // 2018 : 255 - 0xff
      12'h7E3: dout <= 8'b11111111; // 2019 : 255 - 0xff
      12'h7E4: dout <= 8'b11111111; // 2020 : 255 - 0xff
      12'h7E5: dout <= 8'b11111111; // 2021 : 255 - 0xff
      12'h7E6: dout <= 8'b11111111; // 2022 : 255 - 0xff
      12'h7E7: dout <= 8'b11111111; // 2023 : 255 - 0xff
      12'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0 -- plane 1
      12'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout <= 8'b11111110; // 2026 : 254 - 0xfe
      12'h7EB: dout <= 8'b11111110; // 2027 : 254 - 0xfe
      12'h7EC: dout <= 8'b11111110; // 2028 : 254 - 0xfe
      12'h7ED: dout <= 8'b11111110; // 2029 : 254 - 0xfe
      12'h7EE: dout <= 8'b11111110; // 2030 : 254 - 0xfe
      12'h7EF: dout <= 8'b11111110; // 2031 : 254 - 0xfe
      12'h7F0: dout <= 8'b11111111; // 2032 : 255 - 0xff -- Sprite 0x7f
      12'h7F1: dout <= 8'b11111111; // 2033 : 255 - 0xff
      12'h7F2: dout <= 8'b11111111; // 2034 : 255 - 0xff
      12'h7F3: dout <= 8'b11111111; // 2035 : 255 - 0xff
      12'h7F4: dout <= 8'b11111111; // 2036 : 255 - 0xff
      12'h7F5: dout <= 8'b11111111; // 2037 : 255 - 0xff
      12'h7F6: dout <= 8'b11111111; // 2038 : 255 - 0xff
      12'h7F7: dout <= 8'b11111111; // 2039 : 255 - 0xff
      12'h7F8: dout <= 8'b01111110; // 2040 : 126 - 0x7e -- plane 1
      12'h7F9: dout <= 8'b11111110; // 2041 : 254 - 0xfe
      12'h7FA: dout <= 8'b11111110; // 2042 : 254 - 0xfe
      12'h7FB: dout <= 8'b11111110; // 2043 : 254 - 0xfe
      12'h7FC: dout <= 8'b11111110; // 2044 : 254 - 0xfe
      12'h7FD: dout <= 8'b11111110; // 2045 : 254 - 0xfe
      12'h7FE: dout <= 8'b11111110; // 2046 : 254 - 0xfe
      12'h7FF: dout <= 8'b01111110; // 2047 : 126 - 0x7e
      12'h800: dout <= 8'b10111111; // 2048 : 191 - 0xbf -- Sprite 0x80
      12'h801: dout <= 8'b11110111; // 2049 : 247 - 0xf7
      12'h802: dout <= 8'b11111101; // 2050 : 253 - 0xfd
      12'h803: dout <= 8'b11011111; // 2051 : 223 - 0xdf
      12'h804: dout <= 8'b11111011; // 2052 : 251 - 0xfb
      12'h805: dout <= 8'b10111111; // 2053 : 191 - 0xbf
      12'h806: dout <= 8'b11111110; // 2054 : 254 - 0xfe
      12'h807: dout <= 8'b11101111; // 2055 : 239 - 0xef
      12'h808: dout <= 8'b01000000; // 2056 :  64 - 0x40 -- plane 1
      12'h809: dout <= 8'b00001000; // 2057 :   8 - 0x8
      12'h80A: dout <= 8'b00000010; // 2058 :   2 - 0x2
      12'h80B: dout <= 8'b00100000; // 2059 :  32 - 0x20
      12'h80C: dout <= 8'b00000100; // 2060 :   4 - 0x4
      12'h80D: dout <= 8'b01000000; // 2061 :  64 - 0x40
      12'h80E: dout <= 8'b00000001; // 2062 :   1 - 0x1
      12'h80F: dout <= 8'b00010000; // 2063 :  16 - 0x10
      12'h810: dout <= 8'b11111111; // 2064 : 255 - 0xff -- Sprite 0x81
      12'h811: dout <= 8'b11101110; // 2065 : 238 - 0xee
      12'h812: dout <= 8'b11111111; // 2066 : 255 - 0xff
      12'h813: dout <= 8'b11011111; // 2067 : 223 - 0xdf
      12'h814: dout <= 8'b01110111; // 2068 : 119 - 0x77
      12'h815: dout <= 8'b11111101; // 2069 : 253 - 0xfd
      12'h816: dout <= 8'b11011111; // 2070 : 223 - 0xdf
      12'h817: dout <= 8'b10111111; // 2071 : 191 - 0xbf
      12'h818: dout <= 8'b00000000; // 2072 :   0 - 0x0 -- plane 1
      12'h819: dout <= 8'b00010001; // 2073 :  17 - 0x11
      12'h81A: dout <= 8'b00000000; // 2074 :   0 - 0x0
      12'h81B: dout <= 8'b00100000; // 2075 :  32 - 0x20
      12'h81C: dout <= 8'b10001000; // 2076 : 136 - 0x88
      12'h81D: dout <= 8'b00000010; // 2077 :   2 - 0x2
      12'h81E: dout <= 8'b00100000; // 2078 :  32 - 0x20
      12'h81F: dout <= 8'b01000000; // 2079 :  64 - 0x40
      12'h820: dout <= 8'b11111110; // 2080 : 254 - 0xfe -- Sprite 0x82
      12'h821: dout <= 8'b11101111; // 2081 : 239 - 0xef
      12'h822: dout <= 8'b10111111; // 2082 : 191 - 0xbf
      12'h823: dout <= 8'b11110111; // 2083 : 247 - 0xf7
      12'h824: dout <= 8'b11111101; // 2084 : 253 - 0xfd
      12'h825: dout <= 8'b11011111; // 2085 : 223 - 0xdf
      12'h826: dout <= 8'b11111011; // 2086 : 251 - 0xfb
      12'h827: dout <= 8'b10111111; // 2087 : 191 - 0xbf
      12'h828: dout <= 8'b00000001; // 2088 :   1 - 0x1 -- plane 1
      12'h829: dout <= 8'b00010000; // 2089 :  16 - 0x10
      12'h82A: dout <= 8'b01000000; // 2090 :  64 - 0x40
      12'h82B: dout <= 8'b00001000; // 2091 :   8 - 0x8
      12'h82C: dout <= 8'b00000010; // 2092 :   2 - 0x2
      12'h82D: dout <= 8'b00100000; // 2093 :  32 - 0x20
      12'h82E: dout <= 8'b00000100; // 2094 :   4 - 0x4
      12'h82F: dout <= 8'b01000000; // 2095 :  64 - 0x40
      12'h830: dout <= 8'b11101111; // 2096 : 239 - 0xef -- Sprite 0x83
      12'h831: dout <= 8'b11111111; // 2097 : 255 - 0xff
      12'h832: dout <= 8'b10111011; // 2098 : 187 - 0xbb
      12'h833: dout <= 8'b11111111; // 2099 : 255 - 0xff
      12'h834: dout <= 8'b11110111; // 2100 : 247 - 0xf7
      12'h835: dout <= 8'b11011101; // 2101 : 221 - 0xdd
      12'h836: dout <= 8'b01111111; // 2102 : 127 - 0x7f
      12'h837: dout <= 8'b11110111; // 2103 : 247 - 0xf7
      12'h838: dout <= 8'b00010000; // 2104 :  16 - 0x10 -- plane 1
      12'h839: dout <= 8'b00000000; // 2105 :   0 - 0x0
      12'h83A: dout <= 8'b01000100; // 2106 :  68 - 0x44
      12'h83B: dout <= 8'b00000000; // 2107 :   0 - 0x0
      12'h83C: dout <= 8'b00001000; // 2108 :   8 - 0x8
      12'h83D: dout <= 8'b00100010; // 2109 :  34 - 0x22
      12'h83E: dout <= 8'b10000000; // 2110 : 128 - 0x80
      12'h83F: dout <= 8'b00001000; // 2111 :   8 - 0x8
      12'h840: dout <= 8'b11111111; // 2112 : 255 - 0xff -- Sprite 0x84
      12'h841: dout <= 8'b11101110; // 2113 : 238 - 0xee
      12'h842: dout <= 8'b11111011; // 2114 : 251 - 0xfb
      12'h843: dout <= 8'b10111111; // 2115 : 191 - 0xbf
      12'h844: dout <= 8'b01111111; // 2116 : 127 - 0x7f
      12'h845: dout <= 8'b11101101; // 2117 : 237 - 0xed
      12'h846: dout <= 8'b11111111; // 2118 : 255 - 0xff
      12'h847: dout <= 8'b10111111; // 2119 : 191 - 0xbf
      12'h848: dout <= 8'b00010100; // 2120 :  20 - 0x14 -- plane 1
      12'h849: dout <= 8'b10110101; // 2121 : 181 - 0xb5
      12'h84A: dout <= 8'b01000100; // 2122 :  68 - 0x44
      12'h84B: dout <= 8'b01001010; // 2123 :  74 - 0x4a
      12'h84C: dout <= 8'b10010010; // 2124 : 146 - 0x92
      12'h84D: dout <= 8'b10010010; // 2125 : 146 - 0x92
      12'h84E: dout <= 8'b01000100; // 2126 :  68 - 0x44
      12'h84F: dout <= 8'b01001001; // 2127 :  73 - 0x49
      12'h850: dout <= 8'b11111111; // 2128 : 255 - 0xff -- Sprite 0x85
      12'h851: dout <= 8'b10111111; // 2129 : 191 - 0xbf
      12'h852: dout <= 8'b01111101; // 2130 : 125 - 0x7d
      12'h853: dout <= 8'b11110111; // 2131 : 247 - 0xf7
      12'h854: dout <= 8'b11011011; // 2132 : 219 - 0xdb
      12'h855: dout <= 8'b11111101; // 2133 : 253 - 0xfd
      12'h856: dout <= 8'b01111110; // 2134 : 126 - 0x7e
      12'h857: dout <= 8'b11111011; // 2135 : 251 - 0xfb
      12'h858: dout <= 8'b01000010; // 2136 :  66 - 0x42 -- plane 1
      12'h859: dout <= 8'b01001010; // 2137 :  74 - 0x4a
      12'h85A: dout <= 8'b11001010; // 2138 : 202 - 0xca
      12'h85B: dout <= 8'b00101001; // 2139 :  41 - 0x29
      12'h85C: dout <= 8'b10100110; // 2140 : 166 - 0xa6
      12'h85D: dout <= 8'b10010010; // 2141 : 146 - 0x92
      12'h85E: dout <= 8'b10001001; // 2142 : 137 - 0x89
      12'h85F: dout <= 8'b00101101; // 2143 :  45 - 0x2d
      12'h860: dout <= 8'b11111111; // 2144 : 255 - 0xff -- Sprite 0x86
      12'h861: dout <= 8'b11110111; // 2145 : 247 - 0xf7
      12'h862: dout <= 8'b11111111; // 2146 : 255 - 0xff
      12'h863: dout <= 8'b11011101; // 2147 : 221 - 0xdd
      12'h864: dout <= 8'b01111111; // 2148 : 127 - 0x7f
      12'h865: dout <= 8'b11110111; // 2149 : 247 - 0xf7
      12'h866: dout <= 8'b11101111; // 2150 : 239 - 0xef
      12'h867: dout <= 8'b10111101; // 2151 : 189 - 0xbd
      12'h868: dout <= 8'b10001000; // 2152 : 136 - 0x88 -- plane 1
      12'h869: dout <= 8'b00101001; // 2153 :  41 - 0x29
      12'h86A: dout <= 8'b10000010; // 2154 : 130 - 0x82
      12'h86B: dout <= 8'b10110110; // 2155 : 182 - 0xb6
      12'h86C: dout <= 8'b10001000; // 2156 : 136 - 0x88
      12'h86D: dout <= 8'b01001001; // 2157 :  73 - 0x49
      12'h86E: dout <= 8'b01010010; // 2158 :  82 - 0x52
      12'h86F: dout <= 8'b01010010; // 2159 :  82 - 0x52
      12'h870: dout <= 8'b01011111; // 2160 :  95 - 0x5f -- Sprite 0x87
      12'h871: dout <= 8'b11111101; // 2161 : 253 - 0xfd
      12'h872: dout <= 8'b11110110; // 2162 : 246 - 0xf6
      12'h873: dout <= 8'b01111111; // 2163 : 127 - 0x7f
      12'h874: dout <= 8'b10011111; // 2164 : 159 - 0x9f
      12'h875: dout <= 8'b11111110; // 2165 : 254 - 0xfe
      12'h876: dout <= 8'b11111111; // 2166 : 255 - 0xff
      12'h877: dout <= 8'b11101111; // 2167 : 239 - 0xef
      12'h878: dout <= 8'b10110010; // 2168 : 178 - 0xb2 -- plane 1
      12'h879: dout <= 8'b01001010; // 2169 :  74 - 0x4a
      12'h87A: dout <= 8'b10101001; // 2170 : 169 - 0xa9
      12'h87B: dout <= 8'b10100100; // 2171 : 164 - 0xa4
      12'h87C: dout <= 8'b01100010; // 2172 :  98 - 0x62
      12'h87D: dout <= 8'b01001011; // 2173 :  75 - 0x4b
      12'h87E: dout <= 8'b10010000; // 2174 : 144 - 0x90
      12'h87F: dout <= 8'b10010010; // 2175 : 146 - 0x92
      12'h880: dout <= 8'b11111111; // 2176 : 255 - 0xff -- Sprite 0x88
      12'h881: dout <= 8'b11111111; // 2177 : 255 - 0xff
      12'h882: dout <= 8'b10011111; // 2178 : 159 - 0x9f
      12'h883: dout <= 8'b10110011; // 2179 : 179 - 0xb3
      12'h884: dout <= 8'b11110011; // 2180 : 243 - 0xf3
      12'h885: dout <= 8'b11111111; // 2181 : 255 - 0xff
      12'h886: dout <= 8'b11111111; // 2182 : 255 - 0xff
      12'h887: dout <= 8'b11111111; // 2183 : 255 - 0xff
      12'h888: dout <= 8'b00000000; // 2184 :   0 - 0x0 -- plane 1
      12'h889: dout <= 8'b01100000; // 2185 :  96 - 0x60
      12'h88A: dout <= 8'b11111110; // 2186 : 254 - 0xfe
      12'h88B: dout <= 8'b11111111; // 2187 : 255 - 0xff
      12'h88C: dout <= 8'b01111111; // 2188 : 127 - 0x7f
      12'h88D: dout <= 8'b00011111; // 2189 :  31 - 0x1f
      12'h88E: dout <= 8'b00001110; // 2190 :  14 - 0xe
      12'h88F: dout <= 8'b00000000; // 2191 :   0 - 0x0
      12'h890: dout <= 8'b11111111; // 2192 : 255 - 0xff -- Sprite 0x89
      12'h891: dout <= 8'b11001111; // 2193 : 207 - 0xcf
      12'h892: dout <= 8'b11011111; // 2194 : 223 - 0xdf
      12'h893: dout <= 8'b11111111; // 2195 : 255 - 0xff
      12'h894: dout <= 8'b11110011; // 2196 : 243 - 0xf3
      12'h895: dout <= 8'b11110011; // 2197 : 243 - 0xf3
      12'h896: dout <= 8'b11111111; // 2198 : 255 - 0xff
      12'h897: dout <= 8'b11111111; // 2199 : 255 - 0xff
      12'h898: dout <= 8'b00110000; // 2200 :  48 - 0x30 -- plane 1
      12'h899: dout <= 8'b01111000; // 2201 : 120 - 0x78
      12'h89A: dout <= 8'b01111000; // 2202 : 120 - 0x78
      12'h89B: dout <= 8'b00111110; // 2203 :  62 - 0x3e
      12'h89C: dout <= 8'b00011111; // 2204 :  31 - 0x1f
      12'h89D: dout <= 8'b00011111; // 2205 :  31 - 0x1f
      12'h89E: dout <= 8'b00011111; // 2206 :  31 - 0x1f
      12'h89F: dout <= 8'b00001110; // 2207 :  14 - 0xe
      12'h8A0: dout <= 8'b10111111; // 2208 : 191 - 0xbf -- Sprite 0x8a
      12'h8A1: dout <= 8'b11110111; // 2209 : 247 - 0xf7
      12'h8A2: dout <= 8'b11111101; // 2210 : 253 - 0xfd
      12'h8A3: dout <= 8'b11111111; // 2211 : 255 - 0xff
      12'h8A4: dout <= 8'b11111011; // 2212 : 251 - 0xfb
      12'h8A5: dout <= 8'b10111111; // 2213 : 191 - 0xbf
      12'h8A6: dout <= 8'b11111110; // 2214 : 254 - 0xfe
      12'h8A7: dout <= 8'b11101111; // 2215 : 239 - 0xef
      12'h8A8: dout <= 8'b01000000; // 2216 :  64 - 0x40 -- plane 1
      12'h8A9: dout <= 8'b00001000; // 2217 :   8 - 0x8
      12'h8AA: dout <= 8'b00000010; // 2218 :   2 - 0x2
      12'h8AB: dout <= 8'b00101000; // 2219 :  40 - 0x28
      12'h8AC: dout <= 8'b00010100; // 2220 :  20 - 0x14
      12'h8AD: dout <= 8'b01010100; // 2221 :  84 - 0x54
      12'h8AE: dout <= 8'b00000001; // 2222 :   1 - 0x1
      12'h8AF: dout <= 8'b00010000; // 2223 :  16 - 0x10
      12'h8B0: dout <= 8'b10111111; // 2224 : 191 - 0xbf -- Sprite 0x8b
      12'h8B1: dout <= 8'b11111111; // 2225 : 255 - 0xff
      12'h8B2: dout <= 8'b11101110; // 2226 : 238 - 0xee
      12'h8B3: dout <= 8'b11111111; // 2227 : 255 - 0xff
      12'h8B4: dout <= 8'b11011111; // 2228 : 223 - 0xdf
      12'h8B5: dout <= 8'b01111101; // 2229 : 125 - 0x7d
      12'h8B6: dout <= 8'b11111111; // 2230 : 255 - 0xff
      12'h8B7: dout <= 8'b11011111; // 2231 : 223 - 0xdf
      12'h8B8: dout <= 8'b01000000; // 2232 :  64 - 0x40 -- plane 1
      12'h8B9: dout <= 8'b00000000; // 2233 :   0 - 0x0
      12'h8BA: dout <= 8'b10010001; // 2234 : 145 - 0x91
      12'h8BB: dout <= 8'b00010100; // 2235 :  20 - 0x14
      12'h8BC: dout <= 8'b00101000; // 2236 :  40 - 0x28
      12'h8BD: dout <= 8'b10001010; // 2237 : 138 - 0x8a
      12'h8BE: dout <= 8'b01000000; // 2238 :  64 - 0x40
      12'h8BF: dout <= 8'b00100000; // 2239 :  32 - 0x20
      12'h8C0: dout <= 8'b11111111; // 2240 : 255 - 0xff -- Sprite 0x8c
      12'h8C1: dout <= 8'b11111000; // 2241 : 248 - 0xf8
      12'h8C2: dout <= 8'b11100010; // 2242 : 226 - 0xe2
      12'h8C3: dout <= 8'b11010111; // 2243 : 215 - 0xd7
      12'h8C4: dout <= 8'b11001111; // 2244 : 207 - 0xcf
      12'h8C5: dout <= 8'b10011111; // 2245 : 159 - 0x9f
      12'h8C6: dout <= 8'b10111110; // 2246 : 190 - 0xbe
      12'h8C7: dout <= 8'b10011101; // 2247 : 157 - 0x9d
      12'h8C8: dout <= 8'b00000000; // 2248 :   0 - 0x0 -- plane 1
      12'h8C9: dout <= 8'b00000111; // 2249 :   7 - 0x7
      12'h8CA: dout <= 8'b00011111; // 2250 :  31 - 0x1f
      12'h8CB: dout <= 8'b00111111; // 2251 :  63 - 0x3f
      12'h8CC: dout <= 8'b00111111; // 2252 :  63 - 0x3f
      12'h8CD: dout <= 8'b01111111; // 2253 : 127 - 0x7f
      12'h8CE: dout <= 8'b01111111; // 2254 : 127 - 0x7f
      12'h8CF: dout <= 8'b01111111; // 2255 : 127 - 0x7f
      12'h8D0: dout <= 8'b11111111; // 2256 : 255 - 0xff -- Sprite 0x8d
      12'h8D1: dout <= 8'b00011111; // 2257 :  31 - 0x1f
      12'h8D2: dout <= 8'b10100111; // 2258 : 167 - 0xa7
      12'h8D3: dout <= 8'b11000011; // 2259 : 195 - 0xc3
      12'h8D4: dout <= 8'b11100011; // 2260 : 227 - 0xe3
      12'h8D5: dout <= 8'b01000001; // 2261 :  65 - 0x41
      12'h8D6: dout <= 8'b10100001; // 2262 : 161 - 0xa1
      12'h8D7: dout <= 8'b00000001; // 2263 :   1 - 0x1
      12'h8D8: dout <= 8'b00000000; // 2264 :   0 - 0x0 -- plane 1
      12'h8D9: dout <= 8'b11100000; // 2265 : 224 - 0xe0
      12'h8DA: dout <= 8'b11111000; // 2266 : 248 - 0xf8
      12'h8DB: dout <= 8'b11111000; // 2267 : 248 - 0xf8
      12'h8DC: dout <= 8'b11110000; // 2268 : 240 - 0xf0
      12'h8DD: dout <= 8'b11111000; // 2269 : 248 - 0xf8
      12'h8DE: dout <= 8'b11110100; // 2270 : 244 - 0xf4
      12'h8DF: dout <= 8'b11111000; // 2271 : 248 - 0xf8
      12'h8E0: dout <= 8'b10111110; // 2272 : 190 - 0xbe -- Sprite 0x8e
      12'h8E1: dout <= 8'b11111111; // 2273 : 255 - 0xff
      12'h8E2: dout <= 8'b11011111; // 2274 : 223 - 0xdf
      12'h8E3: dout <= 8'b11111111; // 2275 : 255 - 0xff
      12'h8E4: dout <= 8'b11101111; // 2276 : 239 - 0xef
      12'h8E5: dout <= 8'b11111111; // 2277 : 255 - 0xff
      12'h8E6: dout <= 8'b11110111; // 2278 : 247 - 0xf7
      12'h8E7: dout <= 8'b11111111; // 2279 : 255 - 0xff
      12'h8E8: dout <= 8'b01111111; // 2280 : 127 - 0x7f -- plane 1
      12'h8E9: dout <= 8'b00111111; // 2281 :  63 - 0x3f
      12'h8EA: dout <= 8'b00111111; // 2282 :  63 - 0x3f
      12'h8EB: dout <= 8'b00011111; // 2283 :  31 - 0x1f
      12'h8EC: dout <= 8'b00011111; // 2284 :  31 - 0x1f
      12'h8ED: dout <= 8'b00001111; // 2285 :  15 - 0xf
      12'h8EE: dout <= 8'b00001111; // 2286 :  15 - 0xf
      12'h8EF: dout <= 8'b00000111; // 2287 :   7 - 0x7
      12'h8F0: dout <= 8'b01111101; // 2288 : 125 - 0x7d -- Sprite 0x8f
      12'h8F1: dout <= 8'b11111111; // 2289 : 255 - 0xff
      12'h8F2: dout <= 8'b11111011; // 2290 : 251 - 0xfb
      12'h8F3: dout <= 8'b11111111; // 2291 : 255 - 0xff
      12'h8F4: dout <= 8'b11110111; // 2292 : 247 - 0xf7
      12'h8F5: dout <= 8'b11111111; // 2293 : 255 - 0xff
      12'h8F6: dout <= 8'b11101111; // 2294 : 239 - 0xef
      12'h8F7: dout <= 8'b11111111; // 2295 : 255 - 0xff
      12'h8F8: dout <= 8'b11111110; // 2296 : 254 - 0xfe -- plane 1
      12'h8F9: dout <= 8'b11111100; // 2297 : 252 - 0xfc
      12'h8FA: dout <= 8'b11111100; // 2298 : 252 - 0xfc
      12'h8FB: dout <= 8'b11111000; // 2299 : 248 - 0xf8
      12'h8FC: dout <= 8'b11111000; // 2300 : 248 - 0xf8
      12'h8FD: dout <= 8'b11110000; // 2301 : 240 - 0xf0
      12'h8FE: dout <= 8'b11110000; // 2302 : 240 - 0xf0
      12'h8FF: dout <= 8'b11100000; // 2303 : 224 - 0xe0
      12'h900: dout <= 8'b10111110; // 2304 : 190 - 0xbe -- Sprite 0x90
      12'h901: dout <= 8'b11110111; // 2305 : 247 - 0xf7
      12'h902: dout <= 8'b11111111; // 2306 : 255 - 0xff
      12'h903: dout <= 8'b11011111; // 2307 : 223 - 0xdf
      12'h904: dout <= 8'b11111011; // 2308 : 251 - 0xfb
      12'h905: dout <= 8'b11111110; // 2309 : 254 - 0xfe
      12'h906: dout <= 8'b10111111; // 2310 : 191 - 0xbf
      12'h907: dout <= 8'b11110111; // 2311 : 247 - 0xf7
      12'h908: dout <= 8'b01000001; // 2312 :  65 - 0x41 -- plane 1
      12'h909: dout <= 8'b00001000; // 2313 :   8 - 0x8
      12'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout <= 8'b00100000; // 2315 :  32 - 0x20
      12'h90C: dout <= 8'b00000100; // 2316 :   4 - 0x4
      12'h90D: dout <= 8'b00000001; // 2317 :   1 - 0x1
      12'h90E: dout <= 8'b01000000; // 2318 :  64 - 0x40
      12'h90F: dout <= 8'b00001000; // 2319 :   8 - 0x8
      12'h910: dout <= 8'b11101110; // 2320 : 238 - 0xee -- Sprite 0x91
      12'h911: dout <= 8'b11111111; // 2321 : 255 - 0xff
      12'h912: dout <= 8'b01111011; // 2322 : 123 - 0x7b
      12'h913: dout <= 8'b11111101; // 2323 : 253 - 0xfd
      12'h914: dout <= 8'b11101111; // 2324 : 239 - 0xef
      12'h915: dout <= 8'b11111111; // 2325 : 255 - 0xff
      12'h916: dout <= 8'b10111101; // 2326 : 189 - 0xbd
      12'h917: dout <= 8'b11111111; // 2327 : 255 - 0xff
      12'h918: dout <= 8'b00010001; // 2328 :  17 - 0x11 -- plane 1
      12'h919: dout <= 8'b00000000; // 2329 :   0 - 0x0
      12'h91A: dout <= 8'b10000100; // 2330 : 132 - 0x84
      12'h91B: dout <= 8'b00000010; // 2331 :   2 - 0x2
      12'h91C: dout <= 8'b00010000; // 2332 :  16 - 0x10
      12'h91D: dout <= 8'b00000000; // 2333 :   0 - 0x0
      12'h91E: dout <= 8'b01000010; // 2334 :  66 - 0x42
      12'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout <= 8'b11111011; // 2336 : 251 - 0xfb -- Sprite 0x92
      12'h921: dout <= 8'b10111111; // 2337 : 191 - 0xbf
      12'h922: dout <= 8'b11101111; // 2338 : 239 - 0xef
      12'h923: dout <= 8'b11111101; // 2339 : 253 - 0xfd
      12'h924: dout <= 8'b11111111; // 2340 : 255 - 0xff
      12'h925: dout <= 8'b10111111; // 2341 : 191 - 0xbf
      12'h926: dout <= 8'b11111011; // 2342 : 251 - 0xfb
      12'h927: dout <= 8'b11011111; // 2343 : 223 - 0xdf
      12'h928: dout <= 8'b00000100; // 2344 :   4 - 0x4 -- plane 1
      12'h929: dout <= 8'b01000000; // 2345 :  64 - 0x40
      12'h92A: dout <= 8'b00010000; // 2346 :  16 - 0x10
      12'h92B: dout <= 8'b00000010; // 2347 :   2 - 0x2
      12'h92C: dout <= 8'b00000000; // 2348 :   0 - 0x0
      12'h92D: dout <= 8'b01000000; // 2349 :  64 - 0x40
      12'h92E: dout <= 8'b00000100; // 2350 :   4 - 0x4
      12'h92F: dout <= 8'b00100000; // 2351 :  32 - 0x20
      12'h930: dout <= 8'b10111101; // 2352 : 189 - 0xbd -- Sprite 0x93
      12'h931: dout <= 8'b11111111; // 2353 : 255 - 0xff
      12'h932: dout <= 8'b01110111; // 2354 : 119 - 0x77
      12'h933: dout <= 8'b11111110; // 2355 : 254 - 0xfe
      12'h934: dout <= 8'b11011111; // 2356 : 223 - 0xdf
      12'h935: dout <= 8'b11111011; // 2357 : 251 - 0xfb
      12'h936: dout <= 8'b11101111; // 2358 : 239 - 0xef
      12'h937: dout <= 8'b01111111; // 2359 : 127 - 0x7f
      12'h938: dout <= 8'b01000010; // 2360 :  66 - 0x42 -- plane 1
      12'h939: dout <= 8'b00000000; // 2361 :   0 - 0x0
      12'h93A: dout <= 8'b10001000; // 2362 : 136 - 0x88
      12'h93B: dout <= 8'b00000001; // 2363 :   1 - 0x1
      12'h93C: dout <= 8'b00100000; // 2364 :  32 - 0x20
      12'h93D: dout <= 8'b00000100; // 2365 :   4 - 0x4
      12'h93E: dout <= 8'b00010000; // 2366 :  16 - 0x10
      12'h93F: dout <= 8'b10000000; // 2367 : 128 - 0x80
      12'h940: dout <= 8'b01111111; // 2368 : 127 - 0x7f -- Sprite 0x94
      12'h941: dout <= 8'b11110111; // 2369 : 247 - 0xf7
      12'h942: dout <= 8'b11011101; // 2370 : 221 - 0xdd
      12'h943: dout <= 8'b01111011; // 2371 : 123 - 0x7b
      12'h944: dout <= 8'b11111111; // 2372 : 255 - 0xff
      12'h945: dout <= 8'b11101110; // 2373 : 238 - 0xee
      12'h946: dout <= 8'b10111011; // 2374 : 187 - 0xbb
      12'h947: dout <= 8'b11111101; // 2375 : 253 - 0xfd
      12'h948: dout <= 8'b11001000; // 2376 : 200 - 0xc8 -- plane 1
      12'h949: dout <= 8'b00101010; // 2377 :  42 - 0x2a
      12'h94A: dout <= 8'b10100010; // 2378 : 162 - 0xa2
      12'h94B: dout <= 8'b10010100; // 2379 : 148 - 0x94
      12'h94C: dout <= 8'b10010001; // 2380 : 145 - 0x91
      12'h94D: dout <= 8'b01010101; // 2381 :  85 - 0x55
      12'h94E: dout <= 8'b01000100; // 2382 :  68 - 0x44
      12'h94F: dout <= 8'b00010010; // 2383 :  18 - 0x12
      12'h950: dout <= 8'b11010111; // 2384 : 215 - 0xd7 -- Sprite 0x95
      12'h951: dout <= 8'b01111111; // 2385 : 127 - 0x7f
      12'h952: dout <= 8'b11111101; // 2386 : 253 - 0xfd
      12'h953: dout <= 8'b11101110; // 2387 : 238 - 0xee
      12'h954: dout <= 8'b11110111; // 2388 : 247 - 0xf7
      12'h955: dout <= 8'b10111011; // 2389 : 187 - 0xbb
      12'h956: dout <= 8'b11101111; // 2390 : 239 - 0xef
      12'h957: dout <= 8'b11110111; // 2391 : 247 - 0xf7
      12'h958: dout <= 8'b10101010; // 2392 : 170 - 0xaa -- plane 1
      12'h959: dout <= 8'b10100010; // 2393 : 162 - 0xa2
      12'h95A: dout <= 8'b00010010; // 2394 :  18 - 0x12
      12'h95B: dout <= 8'b01010011; // 2395 :  83 - 0x53
      12'h95C: dout <= 8'b01001100; // 2396 :  76 - 0x4c
      12'h95D: dout <= 8'b01010101; // 2397 :  85 - 0x55
      12'h95E: dout <= 8'b10010001; // 2398 : 145 - 0x91
      12'h95F: dout <= 8'b01001000; // 2399 :  72 - 0x48
      12'h960: dout <= 8'b10111111; // 2400 : 191 - 0xbf -- Sprite 0x96
      12'h961: dout <= 8'b11101110; // 2401 : 238 - 0xee
      12'h962: dout <= 8'b11011011; // 2402 : 219 - 0xdb
      12'h963: dout <= 8'b11111111; // 2403 : 255 - 0xff
      12'h964: dout <= 8'b01110111; // 2404 : 119 - 0x77
      12'h965: dout <= 8'b11011101; // 2405 : 221 - 0xdd
      12'h966: dout <= 8'b11101111; // 2406 : 239 - 0xef
      12'h967: dout <= 8'b11111011; // 2407 : 251 - 0xfb
      12'h968: dout <= 8'b01010001; // 2408 :  81 - 0x51 -- plane 1
      12'h969: dout <= 8'b00010101; // 2409 :  21 - 0x15
      12'h96A: dout <= 8'b10100100; // 2410 : 164 - 0xa4
      12'h96B: dout <= 8'b10001100; // 2411 : 140 - 0x8c
      12'h96C: dout <= 8'b10101010; // 2412 : 170 - 0xaa
      12'h96D: dout <= 8'b00100010; // 2413 :  34 - 0x22
      12'h96E: dout <= 8'b10010000; // 2414 : 144 - 0x90
      12'h96F: dout <= 8'b01000110; // 2415 :  70 - 0x46
      12'h970: dout <= 8'b11111101; // 2416 : 253 - 0xfd -- Sprite 0x97
      12'h971: dout <= 8'b11101110; // 2417 : 238 - 0xee
      12'h972: dout <= 8'b11111011; // 2418 : 251 - 0xfb
      12'h973: dout <= 8'b11111101; // 2419 : 253 - 0xfd
      12'h974: dout <= 8'b11110101; // 2420 : 245 - 0xf5
      12'h975: dout <= 8'b11011111; // 2421 : 223 - 0xdf
      12'h976: dout <= 8'b01111111; // 2422 : 127 - 0x7f
      12'h977: dout <= 8'b10111011; // 2423 : 187 - 0xbb
      12'h978: dout <= 8'b00010011; // 2424 :  19 - 0x13 -- plane 1
      12'h979: dout <= 8'b01010101; // 2425 :  85 - 0x55
      12'h97A: dout <= 8'b01100100; // 2426 : 100 - 0x64
      12'h97B: dout <= 8'b00010010; // 2427 :  18 - 0x12
      12'h97C: dout <= 8'b10101010; // 2428 : 170 - 0xaa
      12'h97D: dout <= 8'b10101000; // 2429 : 168 - 0xa8
      12'h97E: dout <= 8'b10000100; // 2430 : 132 - 0x84
      12'h97F: dout <= 8'b11010100; // 2431 : 212 - 0xd4
      12'h980: dout <= 8'b11111111; // 2432 : 255 - 0xff -- Sprite 0x98
      12'h981: dout <= 8'b11001111; // 2433 : 207 - 0xcf
      12'h982: dout <= 8'b11011111; // 2434 : 223 - 0xdf
      12'h983: dout <= 8'b11111111; // 2435 : 255 - 0xff
      12'h984: dout <= 8'b11110011; // 2436 : 243 - 0xf3
      12'h985: dout <= 8'b11110011; // 2437 : 243 - 0xf3
      12'h986: dout <= 8'b11111111; // 2438 : 255 - 0xff
      12'h987: dout <= 8'b11111111; // 2439 : 255 - 0xff
      12'h988: dout <= 8'b00110000; // 2440 :  48 - 0x30 -- plane 1
      12'h989: dout <= 8'b01111000; // 2441 : 120 - 0x78
      12'h98A: dout <= 8'b01111000; // 2442 : 120 - 0x78
      12'h98B: dout <= 8'b00111110; // 2443 :  62 - 0x3e
      12'h98C: dout <= 8'b00011111; // 2444 :  31 - 0x1f
      12'h98D: dout <= 8'b00011111; // 2445 :  31 - 0x1f
      12'h98E: dout <= 8'b00011111; // 2446 :  31 - 0x1f
      12'h98F: dout <= 8'b00001110; // 2447 :  14 - 0xe
      12'h990: dout <= 8'b11111111; // 2448 : 255 - 0xff -- Sprite 0x99
      12'h991: dout <= 8'b11111111; // 2449 : 255 - 0xff
      12'h992: dout <= 8'b10011111; // 2450 : 159 - 0x9f
      12'h993: dout <= 8'b10110011; // 2451 : 179 - 0xb3
      12'h994: dout <= 8'b11110011; // 2452 : 243 - 0xf3
      12'h995: dout <= 8'b11111111; // 2453 : 255 - 0xff
      12'h996: dout <= 8'b11111111; // 2454 : 255 - 0xff
      12'h997: dout <= 8'b11111111; // 2455 : 255 - 0xff
      12'h998: dout <= 8'b00000000; // 2456 :   0 - 0x0 -- plane 1
      12'h999: dout <= 8'b01100000; // 2457 :  96 - 0x60
      12'h99A: dout <= 8'b11111110; // 2458 : 254 - 0xfe
      12'h99B: dout <= 8'b11111111; // 2459 : 255 - 0xff
      12'h99C: dout <= 8'b01111111; // 2460 : 127 - 0x7f
      12'h99D: dout <= 8'b00011111; // 2461 :  31 - 0x1f
      12'h99E: dout <= 8'b00001110; // 2462 :  14 - 0xe
      12'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout <= 8'b10111111; // 2464 : 191 - 0xbf -- Sprite 0x9a
      12'h9A1: dout <= 8'b11110111; // 2465 : 247 - 0xf7
      12'h9A2: dout <= 8'b11111111; // 2466 : 255 - 0xff
      12'h9A3: dout <= 8'b11011111; // 2467 : 223 - 0xdf
      12'h9A4: dout <= 8'b11111011; // 2468 : 251 - 0xfb
      12'h9A5: dout <= 8'b11111111; // 2469 : 255 - 0xff
      12'h9A6: dout <= 8'b10111111; // 2470 : 191 - 0xbf
      12'h9A7: dout <= 8'b11110111; // 2471 : 247 - 0xf7
      12'h9A8: dout <= 8'b01000000; // 2472 :  64 - 0x40 -- plane 1
      12'h9A9: dout <= 8'b00001100; // 2473 :  12 - 0xc
      12'h9AA: dout <= 8'b00000000; // 2474 :   0 - 0x0
      12'h9AB: dout <= 8'b00101000; // 2475 :  40 - 0x28
      12'h9AC: dout <= 8'b00101100; // 2476 :  44 - 0x2c
      12'h9AD: dout <= 8'b00010001; // 2477 :  17 - 0x11
      12'h9AE: dout <= 8'b01000000; // 2478 :  64 - 0x40
      12'h9AF: dout <= 8'b00001000; // 2479 :   8 - 0x8
      12'h9B0: dout <= 8'b11011111; // 2480 : 223 - 0xdf -- Sprite 0x9b
      12'h9B1: dout <= 8'b11111111; // 2481 : 255 - 0xff
      12'h9B2: dout <= 8'b01111011; // 2482 : 123 - 0x7b
      12'h9B3: dout <= 8'b11111111; // 2483 : 255 - 0xff
      12'h9B4: dout <= 8'b11101111; // 2484 : 239 - 0xef
      12'h9B5: dout <= 8'b11111101; // 2485 : 253 - 0xfd
      12'h9B6: dout <= 8'b10111111; // 2486 : 191 - 0xbf
      12'h9B7: dout <= 8'b11111111; // 2487 : 255 - 0xff
      12'h9B8: dout <= 8'b00100000; // 2488 :  32 - 0x20 -- plane 1
      12'h9B9: dout <= 8'b00000000; // 2489 :   0 - 0x0
      12'h9BA: dout <= 8'b10010100; // 2490 : 148 - 0x94
      12'h9BB: dout <= 8'b01001000; // 2491 :  72 - 0x48
      12'h9BC: dout <= 8'b00011000; // 2492 :  24 - 0x18
      12'h9BD: dout <= 8'b00000110; // 2493 :   6 - 0x6
      12'h9BE: dout <= 8'b01000000; // 2494 :  64 - 0x40
      12'h9BF: dout <= 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout <= 8'b10111010; // 2496 : 186 - 0xba -- Sprite 0x9c
      12'h9C1: dout <= 8'b10011100; // 2497 : 156 - 0x9c
      12'h9C2: dout <= 8'b10101010; // 2498 : 170 - 0xaa
      12'h9C3: dout <= 8'b11000000; // 2499 : 192 - 0xc0
      12'h9C4: dout <= 8'b11000000; // 2500 : 192 - 0xc0
      12'h9C5: dout <= 8'b11100000; // 2501 : 224 - 0xe0
      12'h9C6: dout <= 8'b11111000; // 2502 : 248 - 0xf8
      12'h9C7: dout <= 8'b11111111; // 2503 : 255 - 0xff
      12'h9C8: dout <= 8'b01111111; // 2504 : 127 - 0x7f -- plane 1
      12'h9C9: dout <= 8'b01111111; // 2505 : 127 - 0x7f
      12'h9CA: dout <= 8'b01111111; // 2506 : 127 - 0x7f
      12'h9CB: dout <= 8'b00111111; // 2507 :  63 - 0x3f
      12'h9CC: dout <= 8'b00110101; // 2508 :  53 - 0x35
      12'h9CD: dout <= 8'b00000010; // 2509 :   2 - 0x2
      12'h9CE: dout <= 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout <= 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout <= 8'b00000001; // 2512 :   1 - 0x1 -- Sprite 0x9d
      12'h9D1: dout <= 8'b00000001; // 2513 :   1 - 0x1
      12'h9D2: dout <= 8'b00000001; // 2514 :   1 - 0x1
      12'h9D3: dout <= 8'b00000011; // 2515 :   3 - 0x3
      12'h9D4: dout <= 8'b00000011; // 2516 :   3 - 0x3
      12'h9D5: dout <= 8'b00000111; // 2517 :   7 - 0x7
      12'h9D6: dout <= 8'b00011111; // 2518 :  31 - 0x1f
      12'h9D7: dout <= 8'b11111111; // 2519 : 255 - 0xff
      12'h9D8: dout <= 8'b11110100; // 2520 : 244 - 0xf4 -- plane 1
      12'h9D9: dout <= 8'b11111000; // 2521 : 248 - 0xf8
      12'h9DA: dout <= 8'b11110000; // 2522 : 240 - 0xf0
      12'h9DB: dout <= 8'b11101000; // 2523 : 232 - 0xe8
      12'h9DC: dout <= 8'b01010000; // 2524 :  80 - 0x50
      12'h9DD: dout <= 8'b10000000; // 2525 : 128 - 0x80
      12'h9DE: dout <= 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout <= 8'b01111101; // 2528 : 125 - 0x7d -- Sprite 0x9e
      12'h9E1: dout <= 8'b11111111; // 2529 : 255 - 0xff
      12'h9E2: dout <= 8'b11111011; // 2530 : 251 - 0xfb
      12'h9E3: dout <= 8'b11111111; // 2531 : 255 - 0xff
      12'h9E4: dout <= 8'b11111111; // 2532 : 255 - 0xff
      12'h9E5: dout <= 8'b11111011; // 2533 : 251 - 0xfb
      12'h9E6: dout <= 8'b11111111; // 2534 : 255 - 0xff
      12'h9E7: dout <= 8'b01111101; // 2535 : 125 - 0x7d
      12'h9E8: dout <= 8'b11111110; // 2536 : 254 - 0xfe -- plane 1
      12'h9E9: dout <= 8'b11111100; // 2537 : 252 - 0xfc
      12'h9EA: dout <= 8'b11111100; // 2538 : 252 - 0xfc
      12'h9EB: dout <= 8'b11111000; // 2539 : 248 - 0xf8
      12'h9EC: dout <= 8'b11111000; // 2540 : 248 - 0xf8
      12'h9ED: dout <= 8'b11111100; // 2541 : 252 - 0xfc
      12'h9EE: dout <= 8'b11111100; // 2542 : 252 - 0xfc
      12'h9EF: dout <= 8'b11111110; // 2543 : 254 - 0xfe
      12'h9F0: dout <= 8'b11111111; // 2544 : 255 - 0xff -- Sprite 0x9f
      12'h9F1: dout <= 8'b11111111; // 2545 : 255 - 0xff
      12'h9F2: dout <= 8'b10111101; // 2546 : 189 - 0xbd
      12'h9F3: dout <= 8'b11111111; // 2547 : 255 - 0xff
      12'h9F4: dout <= 8'b11111111; // 2548 : 255 - 0xff
      12'h9F5: dout <= 8'b11111111; // 2549 : 255 - 0xff
      12'h9F6: dout <= 8'b11111111; // 2550 : 255 - 0xff
      12'h9F7: dout <= 8'b10111101; // 2551 : 189 - 0xbd
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- plane 1
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b01111110; // 2554 : 126 - 0x7e
      12'h9FB: dout <= 8'b01111110; // 2555 : 126 - 0x7e
      12'h9FC: dout <= 8'b01111110; // 2556 : 126 - 0x7e
      12'h9FD: dout <= 8'b01111110; // 2557 : 126 - 0x7e
      12'h9FE: dout <= 8'b01111110; // 2558 : 126 - 0x7e
      12'h9FF: dout <= 8'b01111110; // 2559 : 126 - 0x7e
      12'hA00: dout <= 8'b11101111; // 2560 : 239 - 0xef -- Sprite 0xa0
      12'hA01: dout <= 8'b11000111; // 2561 : 199 - 0xc7
      12'hA02: dout <= 8'b10000011; // 2562 : 131 - 0x83
      12'hA03: dout <= 8'b00000111; // 2563 :   7 - 0x7
      12'hA04: dout <= 8'b10001111; // 2564 : 143 - 0x8f
      12'hA05: dout <= 8'b11011101; // 2565 : 221 - 0xdd
      12'hA06: dout <= 8'b11111010; // 2566 : 250 - 0xfa
      12'hA07: dout <= 8'b11111101; // 2567 : 253 - 0xfd
      12'hA08: dout <= 8'b00010000; // 2568 :  16 - 0x10 -- plane 1
      12'hA09: dout <= 8'b00111000; // 2569 :  56 - 0x38
      12'hA0A: dout <= 8'b01111100; // 2570 : 124 - 0x7c
      12'hA0B: dout <= 8'b11111000; // 2571 : 248 - 0xf8
      12'hA0C: dout <= 8'b01110000; // 2572 : 112 - 0x70
      12'hA0D: dout <= 8'b00100010; // 2573 :  34 - 0x22
      12'hA0E: dout <= 8'b00000101; // 2574 :   5 - 0x5
      12'hA0F: dout <= 8'b00000010; // 2575 :   2 - 0x2
      12'hA10: dout <= 8'b11101111; // 2576 : 239 - 0xef -- Sprite 0xa1
      12'hA11: dout <= 8'b11000111; // 2577 : 199 - 0xc7
      12'hA12: dout <= 8'b10000011; // 2578 : 131 - 0x83
      12'hA13: dout <= 8'b00011111; // 2579 :  31 - 0x1f
      12'hA14: dout <= 8'b10010000; // 2580 : 144 - 0x90
      12'hA15: dout <= 8'b11010100; // 2581 : 212 - 0xd4
      12'hA16: dout <= 8'b11110011; // 2582 : 243 - 0xf3
      12'hA17: dout <= 8'b11110010; // 2583 : 242 - 0xf2
      12'hA18: dout <= 8'b00010000; // 2584 :  16 - 0x10 -- plane 1
      12'hA19: dout <= 8'b00111000; // 2585 :  56 - 0x38
      12'hA1A: dout <= 8'b01111100; // 2586 : 124 - 0x7c
      12'hA1B: dout <= 8'b11100000; // 2587 : 224 - 0xe0
      12'hA1C: dout <= 8'b01100000; // 2588 :  96 - 0x60
      12'hA1D: dout <= 8'b00100000; // 2589 :  32 - 0x20
      12'hA1E: dout <= 8'b00000000; // 2590 :   0 - 0x0
      12'hA1F: dout <= 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout <= 8'b11101111; // 2592 : 239 - 0xef -- Sprite 0xa2
      12'hA21: dout <= 8'b11000111; // 2593 : 199 - 0xc7
      12'hA22: dout <= 8'b10000011; // 2594 : 131 - 0x83
      12'hA23: dout <= 8'b11111111; // 2595 : 255 - 0xff
      12'hA24: dout <= 8'b00000000; // 2596 :   0 - 0x0
      12'hA25: dout <= 8'b00000000; // 2597 :   0 - 0x0
      12'hA26: dout <= 8'b01010101; // 2598 :  85 - 0x55
      12'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout <= 8'b00010000; // 2600 :  16 - 0x10 -- plane 1
      12'hA29: dout <= 8'b00111000; // 2601 :  56 - 0x38
      12'hA2A: dout <= 8'b01111100; // 2602 : 124 - 0x7c
      12'hA2B: dout <= 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout <= 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout <= 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout <= 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout <= 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout <= 8'b11110000; // 2608 : 240 - 0xf0 -- Sprite 0xa3
      12'hA31: dout <= 8'b11010010; // 2609 : 210 - 0xd2
      12'hA32: dout <= 8'b10010000; // 2610 : 144 - 0x90
      12'hA33: dout <= 8'b00010010; // 2611 :  18 - 0x12
      12'hA34: dout <= 8'b10010000; // 2612 : 144 - 0x90
      12'hA35: dout <= 8'b11010010; // 2613 : 210 - 0xd2
      12'hA36: dout <= 8'b11110000; // 2614 : 240 - 0xf0
      12'hA37: dout <= 8'b11110010; // 2615 : 242 - 0xf2
      12'hA38: dout <= 8'b00000000; // 2616 :   0 - 0x0 -- plane 1
      12'hA39: dout <= 8'b00100000; // 2617 :  32 - 0x20
      12'hA3A: dout <= 8'b01100000; // 2618 :  96 - 0x60
      12'hA3B: dout <= 8'b11100000; // 2619 : 224 - 0xe0
      12'hA3C: dout <= 8'b01100000; // 2620 :  96 - 0x60
      12'hA3D: dout <= 8'b00100000; // 2621 :  32 - 0x20
      12'hA3E: dout <= 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout <= 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout <= 8'b11110000; // 2624 : 240 - 0xf0 -- Sprite 0xa4
      12'hA41: dout <= 8'b11010011; // 2625 : 211 - 0xd3
      12'hA42: dout <= 8'b10010100; // 2626 : 148 - 0x94
      12'hA43: dout <= 8'b00011000; // 2627 :  24 - 0x18
      12'hA44: dout <= 8'b10011111; // 2628 : 159 - 0x9f
      12'hA45: dout <= 8'b11011101; // 2629 : 221 - 0xdd
      12'hA46: dout <= 8'b11111010; // 2630 : 250 - 0xfa
      12'hA47: dout <= 8'b11111101; // 2631 : 253 - 0xfd
      12'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0 -- plane 1
      12'hA49: dout <= 8'b00100000; // 2633 :  32 - 0x20
      12'hA4A: dout <= 8'b01100011; // 2634 :  99 - 0x63
      12'hA4B: dout <= 8'b11100111; // 2635 : 231 - 0xe7
      12'hA4C: dout <= 8'b01100000; // 2636 :  96 - 0x60
      12'hA4D: dout <= 8'b00100010; // 2637 :  34 - 0x22
      12'hA4E: dout <= 8'b00000101; // 2638 :   5 - 0x5
      12'hA4F: dout <= 8'b00000010; // 2639 :   2 - 0x2
      12'hA50: dout <= 8'b00000000; // 2640 :   0 - 0x0 -- Sprite 0xa5
      12'hA51: dout <= 8'b11111111; // 2641 : 255 - 0xff
      12'hA52: dout <= 8'b00000000; // 2642 :   0 - 0x0
      12'hA53: dout <= 8'b00000000; // 2643 :   0 - 0x0
      12'hA54: dout <= 8'b11111111; // 2644 : 255 - 0xff
      12'hA55: dout <= 8'b11011101; // 2645 : 221 - 0xdd
      12'hA56: dout <= 8'b11111010; // 2646 : 250 - 0xfa
      12'hA57: dout <= 8'b11111101; // 2647 : 253 - 0xfd
      12'hA58: dout <= 8'b00000000; // 2648 :   0 - 0x0 -- plane 1
      12'hA59: dout <= 8'b00000000; // 2649 :   0 - 0x0
      12'hA5A: dout <= 8'b11111111; // 2650 : 255 - 0xff
      12'hA5B: dout <= 8'b11111111; // 2651 : 255 - 0xff
      12'hA5C: dout <= 8'b00000000; // 2652 :   0 - 0x0
      12'hA5D: dout <= 8'b00100010; // 2653 :  34 - 0x22
      12'hA5E: dout <= 8'b00000101; // 2654 :   5 - 0x5
      12'hA5F: dout <= 8'b00000010; // 2655 :   2 - 0x2
      12'hA60: dout <= 8'b11101111; // 2656 : 239 - 0xef -- Sprite 0xa6
      12'hA61: dout <= 8'b11000111; // 2657 : 199 - 0xc7
      12'hA62: dout <= 8'b10000011; // 2658 : 131 - 0x83
      12'hA63: dout <= 8'b11111111; // 2659 : 255 - 0xff
      12'hA64: dout <= 8'b00011111; // 2660 :  31 - 0x1f
      12'hA65: dout <= 8'b00101101; // 2661 :  45 - 0x2d
      12'hA66: dout <= 8'b01001010; // 2662 :  74 - 0x4a
      12'hA67: dout <= 8'b01001101; // 2663 :  77 - 0x4d
      12'hA68: dout <= 8'b00010000; // 2664 :  16 - 0x10 -- plane 1
      12'hA69: dout <= 8'b00111000; // 2665 :  56 - 0x38
      12'hA6A: dout <= 8'b01111100; // 2666 : 124 - 0x7c
      12'hA6B: dout <= 8'b00000000; // 2667 :   0 - 0x0
      12'hA6C: dout <= 8'b00000000; // 2668 :   0 - 0x0
      12'hA6D: dout <= 8'b00010010; // 2669 :  18 - 0x12
      12'hA6E: dout <= 8'b00110101; // 2670 :  53 - 0x35
      12'hA6F: dout <= 8'b00110010; // 2671 :  50 - 0x32
      12'hA70: dout <= 8'b01001111; // 2672 :  79 - 0x4f -- Sprite 0xa7
      12'hA71: dout <= 8'b01001111; // 2673 :  79 - 0x4f
      12'hA72: dout <= 8'b01001011; // 2674 :  75 - 0x4b
      12'hA73: dout <= 8'b01001111; // 2675 :  79 - 0x4f
      12'hA74: dout <= 8'b01001111; // 2676 :  79 - 0x4f
      12'hA75: dout <= 8'b01001101; // 2677 :  77 - 0x4d
      12'hA76: dout <= 8'b01001010; // 2678 :  74 - 0x4a
      12'hA77: dout <= 8'b01001101; // 2679 :  77 - 0x4d
      12'hA78: dout <= 8'b00110000; // 2680 :  48 - 0x30 -- plane 1
      12'hA79: dout <= 8'b00110000; // 2681 :  48 - 0x30
      12'hA7A: dout <= 8'b00110100; // 2682 :  52 - 0x34
      12'hA7B: dout <= 8'b00110000; // 2683 :  48 - 0x30
      12'hA7C: dout <= 8'b00110000; // 2684 :  48 - 0x30
      12'hA7D: dout <= 8'b00110010; // 2685 :  50 - 0x32
      12'hA7E: dout <= 8'b00110101; // 2686 :  53 - 0x35
      12'hA7F: dout <= 8'b00110010; // 2687 :  50 - 0x32
      12'hA80: dout <= 8'b01001111; // 2688 :  79 - 0x4f -- Sprite 0xa8
      12'hA81: dout <= 8'b11001111; // 2689 : 207 - 0xcf
      12'hA82: dout <= 8'b00001011; // 2690 :  11 - 0xb
      12'hA83: dout <= 8'b00001111; // 2691 :  15 - 0xf
      12'hA84: dout <= 8'b11111111; // 2692 : 255 - 0xff
      12'hA85: dout <= 8'b11011101; // 2693 : 221 - 0xdd
      12'hA86: dout <= 8'b11111010; // 2694 : 250 - 0xfa
      12'hA87: dout <= 8'b11111101; // 2695 : 253 - 0xfd
      12'hA88: dout <= 8'b00110000; // 2696 :  48 - 0x30 -- plane 1
      12'hA89: dout <= 8'b00110000; // 2697 :  48 - 0x30
      12'hA8A: dout <= 8'b11110100; // 2698 : 244 - 0xf4
      12'hA8B: dout <= 8'b11110000; // 2699 : 240 - 0xf0
      12'hA8C: dout <= 8'b00000000; // 2700 :   0 - 0x0
      12'hA8D: dout <= 8'b00100010; // 2701 :  34 - 0x22
      12'hA8E: dout <= 8'b00000101; // 2702 :   5 - 0x5
      12'hA8F: dout <= 8'b00000010; // 2703 :   2 - 0x2
      12'hA90: dout <= 8'b11111111; // 2704 : 255 - 0xff -- Sprite 0xa9
      12'hA91: dout <= 8'b11111111; // 2705 : 255 - 0xff
      12'hA92: dout <= 8'b11111111; // 2706 : 255 - 0xff
      12'hA93: dout <= 8'b11111111; // 2707 : 255 - 0xff
      12'hA94: dout <= 8'b11111111; // 2708 : 255 - 0xff
      12'hA95: dout <= 8'b11111111; // 2709 : 255 - 0xff
      12'hA96: dout <= 8'b11111111; // 2710 : 255 - 0xff
      12'hA97: dout <= 8'b11111111; // 2711 : 255 - 0xff
      12'hA98: dout <= 8'b00000000; // 2712 :   0 - 0x0 -- plane 1
      12'hA99: dout <= 8'b00000000; // 2713 :   0 - 0x0
      12'hA9A: dout <= 8'b00000000; // 2714 :   0 - 0x0
      12'hA9B: dout <= 8'b00000000; // 2715 :   0 - 0x0
      12'hA9C: dout <= 8'b00000000; // 2716 :   0 - 0x0
      12'hA9D: dout <= 8'b00000000; // 2717 :   0 - 0x0
      12'hA9E: dout <= 8'b00000000; // 2718 :   0 - 0x0
      12'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout <= 8'b11111111; // 2720 : 255 - 0xff -- Sprite 0xaa
      12'hAA1: dout <= 8'b11111111; // 2721 : 255 - 0xff
      12'hAA2: dout <= 8'b10101111; // 2722 : 175 - 0xaf
      12'hAA3: dout <= 8'b01010111; // 2723 :  87 - 0x57
      12'hAA4: dout <= 8'b10001111; // 2724 : 143 - 0x8f
      12'hAA5: dout <= 8'b11011101; // 2725 : 221 - 0xdd
      12'hAA6: dout <= 8'b11111010; // 2726 : 250 - 0xfa
      12'hAA7: dout <= 8'b11111101; // 2727 : 253 - 0xfd
      12'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0 -- plane 1
      12'hAA9: dout <= 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout <= 8'b01010000; // 2730 :  80 - 0x50
      12'hAAB: dout <= 8'b10101000; // 2731 : 168 - 0xa8
      12'hAAC: dout <= 8'b01110000; // 2732 : 112 - 0x70
      12'hAAD: dout <= 8'b00100010; // 2733 :  34 - 0x22
      12'hAAE: dout <= 8'b00000101; // 2734 :   5 - 0x5
      12'hAAF: dout <= 8'b00000010; // 2735 :   2 - 0x2
      12'hAB0: dout <= 8'b11111111; // 2736 : 255 - 0xff -- Sprite 0xab
      12'hAB1: dout <= 8'b00000000; // 2737 :   0 - 0x0
      12'hAB2: dout <= 8'b00000000; // 2738 :   0 - 0x0
      12'hAB3: dout <= 8'b00000000; // 2739 :   0 - 0x0
      12'hAB4: dout <= 8'b00000000; // 2740 :   0 - 0x0
      12'hAB5: dout <= 8'b00000000; // 2741 :   0 - 0x0
      12'hAB6: dout <= 8'b00000000; // 2742 :   0 - 0x0
      12'hAB7: dout <= 8'b00000000; // 2743 :   0 - 0x0
      12'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0 -- plane 1
      12'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout <= 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout <= 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout <= 8'b00000000; // 2752 :   0 - 0x0 -- Sprite 0xac
      12'hAC1: dout <= 8'b00000000; // 2753 :   0 - 0x0
      12'hAC2: dout <= 8'b00000000; // 2754 :   0 - 0x0
      12'hAC3: dout <= 8'b00000000; // 2755 :   0 - 0x0
      12'hAC4: dout <= 8'b00000000; // 2756 :   0 - 0x0
      12'hAC5: dout <= 8'b00000000; // 2757 :   0 - 0x0
      12'hAC6: dout <= 8'b00000000; // 2758 :   0 - 0x0
      12'hAC7: dout <= 8'b00000000; // 2759 :   0 - 0x0
      12'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0 -- plane 1
      12'hAC9: dout <= 8'b00000000; // 2761 :   0 - 0x0
      12'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout <= 8'b00000000; // 2763 :   0 - 0x0
      12'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      12'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout <= 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout <= 8'b00000000; // 2768 :   0 - 0x0 -- Sprite 0xad
      12'hAD1: dout <= 8'b11111111; // 2769 : 255 - 0xff
      12'hAD2: dout <= 8'b00000000; // 2770 :   0 - 0x0
      12'hAD3: dout <= 8'b11111111; // 2771 : 255 - 0xff
      12'hAD4: dout <= 8'b11111111; // 2772 : 255 - 0xff
      12'hAD5: dout <= 8'b11111111; // 2773 : 255 - 0xff
      12'hAD6: dout <= 8'b11111111; // 2774 : 255 - 0xff
      12'hAD7: dout <= 8'b11111111; // 2775 : 255 - 0xff
      12'hAD8: dout <= 8'b00000000; // 2776 :   0 - 0x0 -- plane 1
      12'hAD9: dout <= 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout <= 8'b11111111; // 2778 : 255 - 0xff
      12'hADB: dout <= 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout <= 8'b00000000; // 2780 :   0 - 0x0
      12'hADD: dout <= 8'b00000000; // 2781 :   0 - 0x0
      12'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      12'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout <= 8'b11111111; // 2784 : 255 - 0xff -- Sprite 0xae
      12'hAE1: dout <= 8'b11111111; // 2785 : 255 - 0xff
      12'hAE2: dout <= 8'b11111111; // 2786 : 255 - 0xff
      12'hAE3: dout <= 8'b11111111; // 2787 : 255 - 0xff
      12'hAE4: dout <= 8'b11111111; // 2788 : 255 - 0xff
      12'hAE5: dout <= 8'b00000000; // 2789 :   0 - 0x0
      12'hAE6: dout <= 8'b11111111; // 2790 : 255 - 0xff
      12'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0 -- plane 1
      12'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout <= 8'b00000000; // 2794 :   0 - 0x0
      12'hAEB: dout <= 8'b00000000; // 2795 :   0 - 0x0
      12'hAEC: dout <= 8'b00000000; // 2796 :   0 - 0x0
      12'hAED: dout <= 8'b11111111; // 2797 : 255 - 0xff
      12'hAEE: dout <= 8'b00000000; // 2798 :   0 - 0x0
      12'hAEF: dout <= 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout <= 8'b11111111; // 2800 : 255 - 0xff -- Sprite 0xaf
      12'hAF1: dout <= 8'b11111111; // 2801 : 255 - 0xff
      12'hAF2: dout <= 8'b11111111; // 2802 : 255 - 0xff
      12'hAF3: dout <= 8'b11111111; // 2803 : 255 - 0xff
      12'hAF4: dout <= 8'b11111111; // 2804 : 255 - 0xff
      12'hAF5: dout <= 8'b11111111; // 2805 : 255 - 0xff
      12'hAF6: dout <= 8'b11111111; // 2806 : 255 - 0xff
      12'hAF7: dout <= 8'b11111111; // 2807 : 255 - 0xff
      12'hAF8: dout <= 8'b00000000; // 2808 :   0 - 0x0 -- plane 1
      12'hAF9: dout <= 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout <= 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout <= 8'b00000000; // 2811 :   0 - 0x0
      12'hAFC: dout <= 8'b00000000; // 2812 :   0 - 0x0
      12'hAFD: dout <= 8'b00000000; // 2813 :   0 - 0x0
      12'hAFE: dout <= 8'b00000000; // 2814 :   0 - 0x0
      12'hAFF: dout <= 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout <= 8'b00000000; // 2816 :   0 - 0x0 -- Sprite 0xb0
      12'hB01: dout <= 8'b00011111; // 2817 :  31 - 0x1f
      12'hB02: dout <= 8'b00010000; // 2818 :  16 - 0x10
      12'hB03: dout <= 8'b00010000; // 2819 :  16 - 0x10
      12'hB04: dout <= 8'b00010000; // 2820 :  16 - 0x10
      12'hB05: dout <= 8'b00010000; // 2821 :  16 - 0x10
      12'hB06: dout <= 8'b00010000; // 2822 :  16 - 0x10
      12'hB07: dout <= 8'b00010000; // 2823 :  16 - 0x10
      12'hB08: dout <= 8'b00000000; // 2824 :   0 - 0x0 -- plane 1
      12'hB09: dout <= 8'b00011111; // 2825 :  31 - 0x1f
      12'hB0A: dout <= 8'b00011111; // 2826 :  31 - 0x1f
      12'hB0B: dout <= 8'b00011111; // 2827 :  31 - 0x1f
      12'hB0C: dout <= 8'b00011111; // 2828 :  31 - 0x1f
      12'hB0D: dout <= 8'b00011111; // 2829 :  31 - 0x1f
      12'hB0E: dout <= 8'b00011111; // 2830 :  31 - 0x1f
      12'hB0F: dout <= 8'b00011111; // 2831 :  31 - 0x1f
      12'hB10: dout <= 8'b00000000; // 2832 :   0 - 0x0 -- Sprite 0xb1
      12'hB11: dout <= 8'b11111000; // 2833 : 248 - 0xf8
      12'hB12: dout <= 8'b00001000; // 2834 :   8 - 0x8
      12'hB13: dout <= 8'b00001000; // 2835 :   8 - 0x8
      12'hB14: dout <= 8'b00001000; // 2836 :   8 - 0x8
      12'hB15: dout <= 8'b00001000; // 2837 :   8 - 0x8
      12'hB16: dout <= 8'b00001000; // 2838 :   8 - 0x8
      12'hB17: dout <= 8'b00001000; // 2839 :   8 - 0x8
      12'hB18: dout <= 8'b00000000; // 2840 :   0 - 0x0 -- plane 1
      12'hB19: dout <= 8'b11110000; // 2841 : 240 - 0xf0
      12'hB1A: dout <= 8'b11110000; // 2842 : 240 - 0xf0
      12'hB1B: dout <= 8'b11110000; // 2843 : 240 - 0xf0
      12'hB1C: dout <= 8'b11110000; // 2844 : 240 - 0xf0
      12'hB1D: dout <= 8'b11110000; // 2845 : 240 - 0xf0
      12'hB1E: dout <= 8'b11110000; // 2846 : 240 - 0xf0
      12'hB1F: dout <= 8'b11110000; // 2847 : 240 - 0xf0
      12'hB20: dout <= 8'b00010000; // 2848 :  16 - 0x10 -- Sprite 0xb2
      12'hB21: dout <= 8'b00010000; // 2849 :  16 - 0x10
      12'hB22: dout <= 8'b00010000; // 2850 :  16 - 0x10
      12'hB23: dout <= 8'b00010000; // 2851 :  16 - 0x10
      12'hB24: dout <= 8'b00011111; // 2852 :  31 - 0x1f
      12'hB25: dout <= 8'b00011111; // 2853 :  31 - 0x1f
      12'hB26: dout <= 8'b00001111; // 2854 :  15 - 0xf
      12'hB27: dout <= 8'b00000000; // 2855 :   0 - 0x0
      12'hB28: dout <= 8'b00011111; // 2856 :  31 - 0x1f -- plane 1
      12'hB29: dout <= 8'b00011111; // 2857 :  31 - 0x1f
      12'hB2A: dout <= 8'b00011111; // 2858 :  31 - 0x1f
      12'hB2B: dout <= 8'b00011111; // 2859 :  31 - 0x1f
      12'hB2C: dout <= 8'b00000000; // 2860 :   0 - 0x0
      12'hB2D: dout <= 8'b00000000; // 2861 :   0 - 0x0
      12'hB2E: dout <= 8'b00000000; // 2862 :   0 - 0x0
      12'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout <= 8'b00001000; // 2864 :   8 - 0x8 -- Sprite 0xb3
      12'hB31: dout <= 8'b00001000; // 2865 :   8 - 0x8
      12'hB32: dout <= 8'b00001000; // 2866 :   8 - 0x8
      12'hB33: dout <= 8'b00001000; // 2867 :   8 - 0x8
      12'hB34: dout <= 8'b11111000; // 2868 : 248 - 0xf8
      12'hB35: dout <= 8'b11111000; // 2869 : 248 - 0xf8
      12'hB36: dout <= 8'b11110000; // 2870 : 240 - 0xf0
      12'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      12'hB38: dout <= 8'b11110000; // 2872 : 240 - 0xf0 -- plane 1
      12'hB39: dout <= 8'b11110000; // 2873 : 240 - 0xf0
      12'hB3A: dout <= 8'b11110000; // 2874 : 240 - 0xf0
      12'hB3B: dout <= 8'b11110000; // 2875 : 240 - 0xf0
      12'hB3C: dout <= 8'b00000000; // 2876 :   0 - 0x0
      12'hB3D: dout <= 8'b00000000; // 2877 :   0 - 0x0
      12'hB3E: dout <= 8'b00000000; // 2878 :   0 - 0x0
      12'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout <= 8'b00000000; // 2880 :   0 - 0x0 -- Sprite 0xb4
      12'hB41: dout <= 8'b00000000; // 2881 :   0 - 0x0
      12'hB42: dout <= 8'b00111111; // 2882 :  63 - 0x3f
      12'hB43: dout <= 8'b01100000; // 2883 :  96 - 0x60
      12'hB44: dout <= 8'b01100000; // 2884 :  96 - 0x60
      12'hB45: dout <= 8'b01100000; // 2885 :  96 - 0x60
      12'hB46: dout <= 8'b01100000; // 2886 :  96 - 0x60
      12'hB47: dout <= 8'b01100000; // 2887 :  96 - 0x60
      12'hB48: dout <= 8'b00000000; // 2888 :   0 - 0x0 -- plane 1
      12'hB49: dout <= 8'b00000000; // 2889 :   0 - 0x0
      12'hB4A: dout <= 8'b00111111; // 2890 :  63 - 0x3f
      12'hB4B: dout <= 8'b01111111; // 2891 : 127 - 0x7f
      12'hB4C: dout <= 8'b01111111; // 2892 : 127 - 0x7f
      12'hB4D: dout <= 8'b01111111; // 2893 : 127 - 0x7f
      12'hB4E: dout <= 8'b01111111; // 2894 : 127 - 0x7f
      12'hB4F: dout <= 8'b01111111; // 2895 : 127 - 0x7f
      12'hB50: dout <= 8'b00000000; // 2896 :   0 - 0x0 -- Sprite 0xb5
      12'hB51: dout <= 8'b00000000; // 2897 :   0 - 0x0
      12'hB52: dout <= 8'b11111100; // 2898 : 252 - 0xfc
      12'hB53: dout <= 8'b00000110; // 2899 :   6 - 0x6
      12'hB54: dout <= 8'b00000110; // 2900 :   6 - 0x6
      12'hB55: dout <= 8'b00000110; // 2901 :   6 - 0x6
      12'hB56: dout <= 8'b00000110; // 2902 :   6 - 0x6
      12'hB57: dout <= 8'b00000110; // 2903 :   6 - 0x6
      12'hB58: dout <= 8'b00000000; // 2904 :   0 - 0x0 -- plane 1
      12'hB59: dout <= 8'b00000000; // 2905 :   0 - 0x0
      12'hB5A: dout <= 8'b11111000; // 2906 : 248 - 0xf8
      12'hB5B: dout <= 8'b11111000; // 2907 : 248 - 0xf8
      12'hB5C: dout <= 8'b11111000; // 2908 : 248 - 0xf8
      12'hB5D: dout <= 8'b11111000; // 2909 : 248 - 0xf8
      12'hB5E: dout <= 8'b11111000; // 2910 : 248 - 0xf8
      12'hB5F: dout <= 8'b11111000; // 2911 : 248 - 0xf8
      12'hB60: dout <= 8'b01100000; // 2912 :  96 - 0x60 -- Sprite 0xb6
      12'hB61: dout <= 8'b01100000; // 2913 :  96 - 0x60
      12'hB62: dout <= 8'b01100000; // 2914 :  96 - 0x60
      12'hB63: dout <= 8'b01111111; // 2915 : 127 - 0x7f
      12'hB64: dout <= 8'b01111111; // 2916 : 127 - 0x7f
      12'hB65: dout <= 8'b00111111; // 2917 :  63 - 0x3f
      12'hB66: dout <= 8'b00000000; // 2918 :   0 - 0x0
      12'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout <= 8'b01111111; // 2920 : 127 - 0x7f -- plane 1
      12'hB69: dout <= 8'b01111111; // 2921 : 127 - 0x7f
      12'hB6A: dout <= 8'b01111111; // 2922 : 127 - 0x7f
      12'hB6B: dout <= 8'b01000000; // 2923 :  64 - 0x40
      12'hB6C: dout <= 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout <= 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout <= 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout <= 8'b00000110; // 2928 :   6 - 0x6 -- Sprite 0xb7
      12'hB71: dout <= 8'b00000110; // 2929 :   6 - 0x6
      12'hB72: dout <= 8'b00000110; // 2930 :   6 - 0x6
      12'hB73: dout <= 8'b11111110; // 2931 : 254 - 0xfe
      12'hB74: dout <= 8'b11111110; // 2932 : 254 - 0xfe
      12'hB75: dout <= 8'b11111100; // 2933 : 252 - 0xfc
      12'hB76: dout <= 8'b00000000; // 2934 :   0 - 0x0
      12'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout <= 8'b11111000; // 2936 : 248 - 0xf8 -- plane 1
      12'hB79: dout <= 8'b11111000; // 2937 : 248 - 0xf8
      12'hB7A: dout <= 8'b11111000; // 2938 : 248 - 0xf8
      12'hB7B: dout <= 8'b00000000; // 2939 :   0 - 0x0
      12'hB7C: dout <= 8'b00000000; // 2940 :   0 - 0x0
      12'hB7D: dout <= 8'b00000000; // 2941 :   0 - 0x0
      12'hB7E: dout <= 8'b00000000; // 2942 :   0 - 0x0
      12'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout <= 8'b01100000; // 2944 :  96 - 0x60 -- Sprite 0xb8
      12'hB81: dout <= 8'b11110011; // 2945 : 243 - 0xf3
      12'hB82: dout <= 8'b11000111; // 2946 : 199 - 0xc7
      12'hB83: dout <= 8'b10000110; // 2947 : 134 - 0x86
      12'hB84: dout <= 8'b00000100; // 2948 :   4 - 0x4
      12'hB85: dout <= 8'b00000100; // 2949 :   4 - 0x4
      12'hB86: dout <= 8'b00000111; // 2950 :   7 - 0x7
      12'hB87: dout <= 8'b00000111; // 2951 :   7 - 0x7
      12'hB88: dout <= 8'b00000000; // 2952 :   0 - 0x0 -- plane 1
      12'hB89: dout <= 8'b00000011; // 2953 :   3 - 0x3
      12'hB8A: dout <= 8'b00000111; // 2954 :   7 - 0x7
      12'hB8B: dout <= 8'b00000111; // 2955 :   7 - 0x7
      12'hB8C: dout <= 8'b00000111; // 2956 :   7 - 0x7
      12'hB8D: dout <= 8'b00000011; // 2957 :   3 - 0x3
      12'hB8E: dout <= 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b00000110; // 2960 :   6 - 0x6 -- Sprite 0xb9
      12'hB91: dout <= 8'b10001111; // 2961 : 143 - 0x8f
      12'hB92: dout <= 8'b11000101; // 2962 : 197 - 0xc5
      12'hB93: dout <= 8'b00100011; // 2963 :  35 - 0x23
      12'hB94: dout <= 8'b00101110; // 2964 :  46 - 0x2e
      12'hB95: dout <= 8'b01100000; // 2965 :  96 - 0x60
      12'hB96: dout <= 8'b11100001; // 2966 : 225 - 0xe1
      12'hB97: dout <= 8'b11100001; // 2967 : 225 - 0xe1
      12'hB98: dout <= 8'b00000000; // 2968 :   0 - 0x0 -- plane 1
      12'hB99: dout <= 8'b11000001; // 2969 : 193 - 0xc1
      12'hB9A: dout <= 8'b11100010; // 2970 : 226 - 0xe2
      12'hB9B: dout <= 8'b11001100; // 2971 : 204 - 0xcc
      12'hB9C: dout <= 8'b11000000; // 2972 : 192 - 0xc0
      12'hB9D: dout <= 8'b10000000; // 2973 : 128 - 0x80
      12'hB9E: dout <= 8'b00000001; // 2974 :   1 - 0x1
      12'hB9F: dout <= 8'b00000010; // 2975 :   2 - 0x2
      12'hBA0: dout <= 8'b11001000; // 2976 : 200 - 0xc8 -- Sprite 0xba
      12'hBA1: dout <= 8'b11111000; // 2977 : 248 - 0xf8
      12'hBA2: dout <= 8'b10110000; // 2978 : 176 - 0xb0
      12'hBA3: dout <= 8'b00010000; // 2979 :  16 - 0x10
      12'hBA4: dout <= 8'b00110000; // 2980 :  48 - 0x30
      12'hBA5: dout <= 8'b11001000; // 2981 : 200 - 0xc8
      12'hBA6: dout <= 8'b11111000; // 2982 : 248 - 0xf8
      12'hBA7: dout <= 8'b10000000; // 2983 : 128 - 0x80
      12'hBA8: dout <= 8'b11110000; // 2984 : 240 - 0xf0 -- plane 1
      12'hBA9: dout <= 8'b00000000; // 2985 :   0 - 0x0
      12'hBAA: dout <= 8'b00100000; // 2986 :  32 - 0x20
      12'hBAB: dout <= 8'b00100000; // 2987 :  32 - 0x20
      12'hBAC: dout <= 8'b00000000; // 2988 :   0 - 0x0
      12'hBAD: dout <= 8'b11110000; // 2989 : 240 - 0xf0
      12'hBAE: dout <= 8'b00000000; // 2990 :   0 - 0x0
      12'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout <= 8'b00000011; // 2992 :   3 - 0x3 -- Sprite 0xbb
      12'hBB1: dout <= 8'b00000000; // 2993 :   0 - 0x0
      12'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      12'hBB3: dout <= 8'b01100000; // 2995 :  96 - 0x60
      12'hBB4: dout <= 8'b11110000; // 2996 : 240 - 0xf0
      12'hBB5: dout <= 8'b11010000; // 2997 : 208 - 0xd0
      12'hBB6: dout <= 8'b10010000; // 2998 : 144 - 0x90
      12'hBB7: dout <= 8'b01100000; // 2999 :  96 - 0x60
      12'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0 -- plane 1
      12'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      12'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      12'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      12'hBBD: dout <= 8'b01100000; // 3005 :  96 - 0x60
      12'hBBE: dout <= 8'b01100000; // 3006 :  96 - 0x60
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b11000011; // 3008 : 195 - 0xc3 -- Sprite 0xbc
      12'hBC1: dout <= 8'b00001110; // 3009 :  14 - 0xe
      12'hBC2: dout <= 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout <= 8'b00000110; // 3011 :   6 - 0x6
      12'hBC4: dout <= 8'b00001111; // 3012 :  15 - 0xf
      12'hBC5: dout <= 8'b00001101; // 3013 :  13 - 0xd
      12'hBC6: dout <= 8'b00001001; // 3014 :   9 - 0x9
      12'hBC7: dout <= 8'b00000110; // 3015 :   6 - 0x6
      12'hBC8: dout <= 8'b00001100; // 3016 :  12 - 0xc -- plane 1
      12'hBC9: dout <= 8'b00000000; // 3017 :   0 - 0x0
      12'hBCA: dout <= 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout <= 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout <= 8'b00000110; // 3021 :   6 - 0x6
      12'hBCE: dout <= 8'b00000110; // 3022 :   6 - 0x6
      12'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout <= 8'b11100000; // 3024 : 224 - 0xe0 -- Sprite 0xbd
      12'hBD1: dout <= 8'b01100011; // 3025 :  99 - 0x63
      12'hBD2: dout <= 8'b11100111; // 3026 : 231 - 0xe7
      12'hBD3: dout <= 8'b11100110; // 3027 : 230 - 0xe6
      12'hBD4: dout <= 8'b00000100; // 3028 :   4 - 0x4
      12'hBD5: dout <= 8'b00000100; // 3029 :   4 - 0x4
      12'hBD6: dout <= 8'b00000111; // 3030 :   7 - 0x7
      12'hBD7: dout <= 8'b00000111; // 3031 :   7 - 0x7
      12'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0 -- plane 1
      12'hBD9: dout <= 8'b10000011; // 3033 : 131 - 0x83
      12'hBDA: dout <= 8'b00000111; // 3034 :   7 - 0x7
      12'hBDB: dout <= 8'b00000111; // 3035 :   7 - 0x7
      12'hBDC: dout <= 8'b00000111; // 3036 :   7 - 0x7
      12'hBDD: dout <= 8'b00000011; // 3037 :   3 - 0x3
      12'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout <= 8'b00000111; // 3040 :   7 - 0x7 -- Sprite 0xbe
      12'hBE1: dout <= 8'b10000011; // 3041 : 131 - 0x83
      12'hBE2: dout <= 8'b11000111; // 3042 : 199 - 0xc7
      12'hBE3: dout <= 8'b00100111; // 3043 :  39 - 0x27
      12'hBE4: dout <= 8'b00100000; // 3044 :  32 - 0x20
      12'hBE5: dout <= 8'b01100000; // 3045 :  96 - 0x60
      12'hBE6: dout <= 8'b11100000; // 3046 : 224 - 0xe0
      12'hBE7: dout <= 8'b11100000; // 3047 : 224 - 0xe0
      12'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0 -- plane 1
      12'hBE9: dout <= 8'b11000100; // 3049 : 196 - 0xc4
      12'hBEA: dout <= 8'b11100000; // 3050 : 224 - 0xe0
      12'hBEB: dout <= 8'b11000000; // 3051 : 192 - 0xc0
      12'hBEC: dout <= 8'b11000000; // 3052 : 192 - 0xc0
      12'hBED: dout <= 8'b10000000; // 3053 : 128 - 0x80
      12'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      12'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout <= 8'b00000011; // 3056 :   3 - 0x3 -- Sprite 0xbf
      12'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout <= 8'b00001100; // 3058 :  12 - 0xc
      12'hBF3: dout <= 8'b00001100; // 3059 :  12 - 0xc
      12'hBF4: dout <= 8'b11100100; // 3060 : 228 - 0xe4
      12'hBF5: dout <= 8'b01101100; // 3061 : 108 - 0x6c
      12'hBF6: dout <= 8'b11101101; // 3062 : 237 - 0xed
      12'hBF7: dout <= 8'b11100111; // 3063 : 231 - 0xe7
      12'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0 -- plane 1
      12'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      12'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout <= 8'b00001000; // 3068 :   8 - 0x8
      12'hBFD: dout <= 8'b10001000; // 3069 : 136 - 0x88
      12'hBFE: dout <= 8'b00001011; // 3070 :  11 - 0xb
      12'hBFF: dout <= 8'b00001000; // 3071 :   8 - 0x8
      12'hC00: dout <= 8'b11000000; // 3072 : 192 - 0xc0 -- Sprite 0xc0
      12'hC01: dout <= 8'b00000000; // 3073 :   0 - 0x0
      12'hC02: dout <= 8'b00110000; // 3074 :  48 - 0x30
      12'hC03: dout <= 8'b00110000; // 3075 :  48 - 0x30
      12'hC04: dout <= 8'b00010111; // 3076 :  23 - 0x17
      12'hC05: dout <= 8'b00110011; // 3077 :  51 - 0x33
      12'hC06: dout <= 8'b01110111; // 3078 : 119 - 0x77
      12'hC07: dout <= 8'b11010111; // 3079 : 215 - 0xd7
      12'hC08: dout <= 8'b00000000; // 3080 :   0 - 0x0 -- plane 1
      12'hC09: dout <= 8'b00000000; // 3081 :   0 - 0x0
      12'hC0A: dout <= 8'b00000000; // 3082 :   0 - 0x0
      12'hC0B: dout <= 8'b00000000; // 3083 :   0 - 0x0
      12'hC0C: dout <= 8'b00100000; // 3084 :  32 - 0x20
      12'hC0D: dout <= 8'b00100100; // 3085 :  36 - 0x24
      12'hC0E: dout <= 8'b10100000; // 3086 : 160 - 0xa0
      12'hC0F: dout <= 8'b00100000; // 3087 :  32 - 0x20
      12'hC10: dout <= 8'b00001100; // 3088 :  12 - 0xc -- Sprite 0xc1
      12'hC11: dout <= 8'b00000000; // 3089 :   0 - 0x0
      12'hC12: dout <= 8'b00000000; // 3090 :   0 - 0x0
      12'hC13: dout <= 8'b00000000; // 3091 :   0 - 0x0
      12'hC14: dout <= 8'b00000000; // 3092 :   0 - 0x0
      12'hC15: dout <= 8'b00000000; // 3093 :   0 - 0x0
      12'hC16: dout <= 8'b00000000; // 3094 :   0 - 0x0
      12'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      12'hC18: dout <= 8'b00000000; // 3096 :   0 - 0x0 -- plane 1
      12'hC19: dout <= 8'b00000000; // 3097 :   0 - 0x0
      12'hC1A: dout <= 8'b00000000; // 3098 :   0 - 0x0
      12'hC1B: dout <= 8'b00000000; // 3099 :   0 - 0x0
      12'hC1C: dout <= 8'b00000000; // 3100 :   0 - 0x0
      12'hC1D: dout <= 8'b00000000; // 3101 :   0 - 0x0
      12'hC1E: dout <= 8'b00000000; // 3102 :   0 - 0x0
      12'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout <= 8'b00110000; // 3104 :  48 - 0x30 -- Sprite 0xc2
      12'hC21: dout <= 8'b00000000; // 3105 :   0 - 0x0
      12'hC22: dout <= 8'b00000000; // 3106 :   0 - 0x0
      12'hC23: dout <= 8'b00000000; // 3107 :   0 - 0x0
      12'hC24: dout <= 8'b00000000; // 3108 :   0 - 0x0
      12'hC25: dout <= 8'b00000000; // 3109 :   0 - 0x0
      12'hC26: dout <= 8'b00000000; // 3110 :   0 - 0x0
      12'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      12'hC28: dout <= 8'b00000000; // 3112 :   0 - 0x0 -- plane 1
      12'hC29: dout <= 8'b00000000; // 3113 :   0 - 0x0
      12'hC2A: dout <= 8'b00000000; // 3114 :   0 - 0x0
      12'hC2B: dout <= 8'b00000000; // 3115 :   0 - 0x0
      12'hC2C: dout <= 8'b00000000; // 3116 :   0 - 0x0
      12'hC2D: dout <= 8'b00000000; // 3117 :   0 - 0x0
      12'hC2E: dout <= 8'b00000000; // 3118 :   0 - 0x0
      12'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      12'hC30: dout <= 8'b00000000; // 3120 :   0 - 0x0 -- Sprite 0xc3
      12'hC31: dout <= 8'b00000000; // 3121 :   0 - 0x0
      12'hC32: dout <= 8'b00000100; // 3122 :   4 - 0x4
      12'hC33: dout <= 8'b00001101; // 3123 :  13 - 0xd
      12'hC34: dout <= 8'b00001111; // 3124 :  15 - 0xf
      12'hC35: dout <= 8'b00001100; // 3125 :  12 - 0xc
      12'hC36: dout <= 8'b00001100; // 3126 :  12 - 0xc
      12'hC37: dout <= 8'b00000100; // 3127 :   4 - 0x4
      12'hC38: dout <= 8'b00000000; // 3128 :   0 - 0x0 -- plane 1
      12'hC39: dout <= 8'b00000000; // 3129 :   0 - 0x0
      12'hC3A: dout <= 8'b00001000; // 3130 :   8 - 0x8
      12'hC3B: dout <= 8'b00001011; // 3131 :  11 - 0xb
      12'hC3C: dout <= 8'b00001000; // 3132 :   8 - 0x8
      12'hC3D: dout <= 8'b00001000; // 3133 :   8 - 0x8
      12'hC3E: dout <= 8'b00001000; // 3134 :   8 - 0x8
      12'hC3F: dout <= 8'b00001000; // 3135 :   8 - 0x8
      12'hC40: dout <= 8'b00000000; // 3136 :   0 - 0x0 -- Sprite 0xc4
      12'hC41: dout <= 8'b00000000; // 3137 :   0 - 0x0
      12'hC42: dout <= 8'b00010000; // 3138 :  16 - 0x10
      12'hC43: dout <= 8'b01110000; // 3139 : 112 - 0x70
      12'hC44: dout <= 8'b11110000; // 3140 : 240 - 0xf0
      12'hC45: dout <= 8'b00110000; // 3141 :  48 - 0x30
      12'hC46: dout <= 8'b00110000; // 3142 :  48 - 0x30
      12'hC47: dout <= 8'b00010000; // 3143 :  16 - 0x10
      12'hC48: dout <= 8'b00000000; // 3144 :   0 - 0x0 -- plane 1
      12'hC49: dout <= 8'b00000000; // 3145 :   0 - 0x0
      12'hC4A: dout <= 8'b00100000; // 3146 :  32 - 0x20
      12'hC4B: dout <= 8'b10100000; // 3147 : 160 - 0xa0
      12'hC4C: dout <= 8'b00100000; // 3148 :  32 - 0x20
      12'hC4D: dout <= 8'b00100000; // 3149 :  32 - 0x20
      12'hC4E: dout <= 8'b00100000; // 3150 :  32 - 0x20
      12'hC4F: dout <= 8'b00100000; // 3151 :  32 - 0x20
      12'hC50: dout <= 8'b11100100; // 3152 : 228 - 0xe4 -- Sprite 0xc5
      12'hC51: dout <= 8'b00100100; // 3153 :  36 - 0x24
      12'hC52: dout <= 8'b11101111; // 3154 : 239 - 0xef
      12'hC53: dout <= 8'b11100111; // 3155 : 231 - 0xe7
      12'hC54: dout <= 8'b00000110; // 3156 :   6 - 0x6
      12'hC55: dout <= 8'b00000100; // 3157 :   4 - 0x4
      12'hC56: dout <= 8'b00000100; // 3158 :   4 - 0x4
      12'hC57: dout <= 8'b00000111; // 3159 :   7 - 0x7
      12'hC58: dout <= 8'b00001000; // 3160 :   8 - 0x8 -- plane 1
      12'hC59: dout <= 8'b11001000; // 3161 : 200 - 0xc8
      12'hC5A: dout <= 8'b00000011; // 3162 :   3 - 0x3
      12'hC5B: dout <= 8'b00000111; // 3163 :   7 - 0x7
      12'hC5C: dout <= 8'b00000111; // 3164 :   7 - 0x7
      12'hC5D: dout <= 8'b00000111; // 3165 :   7 - 0x7
      12'hC5E: dout <= 8'b00000011; // 3166 :   3 - 0x3
      12'hC5F: dout <= 8'b00000000; // 3167 :   0 - 0x0
      12'hC60: dout <= 8'b00010111; // 3168 :  23 - 0x17 -- Sprite 0xc6
      12'hC61: dout <= 8'b00010001; // 3169 :  17 - 0x11
      12'hC62: dout <= 8'b10110111; // 3170 : 183 - 0xb7
      12'hC63: dout <= 8'b11000111; // 3171 : 199 - 0xc7
      12'hC64: dout <= 8'b00100000; // 3172 :  32 - 0x20
      12'hC65: dout <= 8'b00100000; // 3173 :  32 - 0x20
      12'hC66: dout <= 8'b01100000; // 3174 :  96 - 0x60
      12'hC67: dout <= 8'b11100000; // 3175 : 224 - 0xe0
      12'hC68: dout <= 8'b00100000; // 3176 :  32 - 0x20 -- plane 1
      12'hC69: dout <= 8'b00100110; // 3177 :  38 - 0x26
      12'hC6A: dout <= 8'b11000000; // 3178 : 192 - 0xc0
      12'hC6B: dout <= 8'b11100000; // 3179 : 224 - 0xe0
      12'hC6C: dout <= 8'b11000000; // 3180 : 192 - 0xc0
      12'hC6D: dout <= 8'b11000000; // 3181 : 192 - 0xc0
      12'hC6E: dout <= 8'b10000000; // 3182 : 128 - 0x80
      12'hC6F: dout <= 8'b00000000; // 3183 :   0 - 0x0
      12'hC70: dout <= 8'b00000111; // 3184 :   7 - 0x7 -- Sprite 0xc7
      12'hC71: dout <= 8'b00000011; // 3185 :   3 - 0x3
      12'hC72: dout <= 8'b00000000; // 3186 :   0 - 0x0
      12'hC73: dout <= 8'b00000000; // 3187 :   0 - 0x0
      12'hC74: dout <= 8'b11100000; // 3188 : 224 - 0xe0
      12'hC75: dout <= 8'b00100000; // 3189 :  32 - 0x20
      12'hC76: dout <= 8'b11100000; // 3190 : 224 - 0xe0
      12'hC77: dout <= 8'b11100000; // 3191 : 224 - 0xe0
      12'hC78: dout <= 8'b00000000; // 3192 :   0 - 0x0 -- plane 1
      12'hC79: dout <= 8'b00000000; // 3193 :   0 - 0x0
      12'hC7A: dout <= 8'b00000000; // 3194 :   0 - 0x0
      12'hC7B: dout <= 8'b00000000; // 3195 :   0 - 0x0
      12'hC7C: dout <= 8'b00000000; // 3196 :   0 - 0x0
      12'hC7D: dout <= 8'b11000000; // 3197 : 192 - 0xc0
      12'hC7E: dout <= 8'b00000000; // 3198 :   0 - 0x0
      12'hC7F: dout <= 8'b00000000; // 3199 :   0 - 0x0
      12'hC80: dout <= 8'b11100000; // 3200 : 224 - 0xe0 -- Sprite 0xc8
      12'hC81: dout <= 8'b11000000; // 3201 : 192 - 0xc0
      12'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      12'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      12'hC84: dout <= 8'b00000111; // 3204 :   7 - 0x7
      12'hC85: dout <= 8'b00000001; // 3205 :   1 - 0x1
      12'hC86: dout <= 8'b00000111; // 3206 :   7 - 0x7
      12'hC87: dout <= 8'b00000111; // 3207 :   7 - 0x7
      12'hC88: dout <= 8'b00000000; // 3208 :   0 - 0x0 -- plane 1
      12'hC89: dout <= 8'b00000000; // 3209 :   0 - 0x0
      12'hC8A: dout <= 8'b00000000; // 3210 :   0 - 0x0
      12'hC8B: dout <= 8'b00000000; // 3211 :   0 - 0x0
      12'hC8C: dout <= 8'b00000000; // 3212 :   0 - 0x0
      12'hC8D: dout <= 8'b00000110; // 3213 :   6 - 0x6
      12'hC8E: dout <= 8'b00000000; // 3214 :   0 - 0x0
      12'hC8F: dout <= 8'b00000000; // 3215 :   0 - 0x0
      12'hC90: dout <= 8'b00010011; // 3216 :  19 - 0x13 -- Sprite 0xc9
      12'hC91: dout <= 8'b00011111; // 3217 :  31 - 0x1f
      12'hC92: dout <= 8'b00001101; // 3218 :  13 - 0xd
      12'hC93: dout <= 8'b00000100; // 3219 :   4 - 0x4
      12'hC94: dout <= 8'b00001100; // 3220 :  12 - 0xc
      12'hC95: dout <= 8'b00010011; // 3221 :  19 - 0x13
      12'hC96: dout <= 8'b00011111; // 3222 :  31 - 0x1f
      12'hC97: dout <= 8'b00000001; // 3223 :   1 - 0x1
      12'hC98: dout <= 8'b00001111; // 3224 :  15 - 0xf -- plane 1
      12'hC99: dout <= 8'b00000000; // 3225 :   0 - 0x0
      12'hC9A: dout <= 8'b00001000; // 3226 :   8 - 0x8
      12'hC9B: dout <= 8'b00001000; // 3227 :   8 - 0x8
      12'hC9C: dout <= 8'b00000000; // 3228 :   0 - 0x0
      12'hC9D: dout <= 8'b00001111; // 3229 :  15 - 0xf
      12'hC9E: dout <= 8'b00000000; // 3230 :   0 - 0x0
      12'hC9F: dout <= 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout <= 8'b01100000; // 3232 :  96 - 0x60 -- Sprite 0xca
      12'hCA1: dout <= 8'b11110011; // 3233 : 243 - 0xf3
      12'hCA2: dout <= 8'b10100111; // 3234 : 167 - 0xa7
      12'hCA3: dout <= 8'b11000110; // 3235 : 198 - 0xc6
      12'hCA4: dout <= 8'b01110100; // 3236 : 116 - 0x74
      12'hCA5: dout <= 8'b00000100; // 3237 :   4 - 0x4
      12'hCA6: dout <= 8'b10000111; // 3238 : 135 - 0x87
      12'hCA7: dout <= 8'b10000111; // 3239 : 135 - 0x87
      12'hCA8: dout <= 8'b00000000; // 3240 :   0 - 0x0 -- plane 1
      12'hCA9: dout <= 8'b10000011; // 3241 : 131 - 0x83
      12'hCAA: dout <= 8'b01000111; // 3242 :  71 - 0x47
      12'hCAB: dout <= 8'b00110111; // 3243 :  55 - 0x37
      12'hCAC: dout <= 8'b00000111; // 3244 :   7 - 0x7
      12'hCAD: dout <= 8'b00000011; // 3245 :   3 - 0x3
      12'hCAE: dout <= 8'b10000000; // 3246 : 128 - 0x80
      12'hCAF: dout <= 8'b01000000; // 3247 :  64 - 0x40
      12'hCB0: dout <= 8'b00000110; // 3248 :   6 - 0x6 -- Sprite 0xcb
      12'hCB1: dout <= 8'b10001111; // 3249 : 143 - 0x8f
      12'hCB2: dout <= 8'b11000011; // 3250 : 195 - 0xc3
      12'hCB3: dout <= 8'b00100001; // 3251 :  33 - 0x21
      12'hCB4: dout <= 8'b00100000; // 3252 :  32 - 0x20
      12'hCB5: dout <= 8'b01100000; // 3253 :  96 - 0x60
      12'hCB6: dout <= 8'b11100000; // 3254 : 224 - 0xe0
      12'hCB7: dout <= 8'b11100000; // 3255 : 224 - 0xe0
      12'hCB8: dout <= 8'b00000000; // 3256 :   0 - 0x0 -- plane 1
      12'hCB9: dout <= 8'b11000000; // 3257 : 192 - 0xc0
      12'hCBA: dout <= 8'b11100000; // 3258 : 224 - 0xe0
      12'hCBB: dout <= 8'b11000000; // 3259 : 192 - 0xc0
      12'hCBC: dout <= 8'b11000000; // 3260 : 192 - 0xc0
      12'hCBD: dout <= 8'b10000000; // 3261 : 128 - 0x80
      12'hCBE: dout <= 8'b00000000; // 3262 :   0 - 0x0
      12'hCBF: dout <= 8'b00000000; // 3263 :   0 - 0x0
      12'hCC0: dout <= 8'b11000011; // 3264 : 195 - 0xc3 -- Sprite 0xcc
      12'hCC1: dout <= 8'b01110000; // 3265 : 112 - 0x70
      12'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      12'hCC3: dout <= 8'b01100000; // 3267 :  96 - 0x60
      12'hCC4: dout <= 8'b11110000; // 3268 : 240 - 0xf0
      12'hCC5: dout <= 8'b11010000; // 3269 : 208 - 0xd0
      12'hCC6: dout <= 8'b10010000; // 3270 : 144 - 0x90
      12'hCC7: dout <= 8'b01100000; // 3271 :  96 - 0x60
      12'hCC8: dout <= 8'b00110000; // 3272 :  48 - 0x30 -- plane 1
      12'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      12'hCCA: dout <= 8'b00000000; // 3274 :   0 - 0x0
      12'hCCB: dout <= 8'b00000000; // 3275 :   0 - 0x0
      12'hCCC: dout <= 8'b00000000; // 3276 :   0 - 0x0
      12'hCCD: dout <= 8'b01100000; // 3277 :  96 - 0x60
      12'hCCE: dout <= 8'b01100000; // 3278 :  96 - 0x60
      12'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout <= 8'b11000000; // 3280 : 192 - 0xc0 -- Sprite 0xcd
      12'hCD1: dout <= 8'b00000000; // 3281 :   0 - 0x0
      12'hCD2: dout <= 8'b00000000; // 3282 :   0 - 0x0
      12'hCD3: dout <= 8'b00000110; // 3283 :   6 - 0x6
      12'hCD4: dout <= 8'b00001111; // 3284 :  15 - 0xf
      12'hCD5: dout <= 8'b00001101; // 3285 :  13 - 0xd
      12'hCD6: dout <= 8'b00001001; // 3286 :   9 - 0x9
      12'hCD7: dout <= 8'b00000110; // 3287 :   6 - 0x6
      12'hCD8: dout <= 8'b00000000; // 3288 :   0 - 0x0 -- plane 1
      12'hCD9: dout <= 8'b00000000; // 3289 :   0 - 0x0
      12'hCDA: dout <= 8'b00000000; // 3290 :   0 - 0x0
      12'hCDB: dout <= 8'b00000000; // 3291 :   0 - 0x0
      12'hCDC: dout <= 8'b00000000; // 3292 :   0 - 0x0
      12'hCDD: dout <= 8'b00000110; // 3293 :   6 - 0x6
      12'hCDE: dout <= 8'b00000110; // 3294 :   6 - 0x6
      12'hCDF: dout <= 8'b00000000; // 3295 :   0 - 0x0
      12'hCE0: dout <= 8'b11111100; // 3296 : 252 - 0xfc -- Sprite 0xce
      12'hCE1: dout <= 8'b11000000; // 3297 : 192 - 0xc0
      12'hCE2: dout <= 8'b11010001; // 3298 : 209 - 0xd1
      12'hCE3: dout <= 8'b11000010; // 3299 : 194 - 0xc2
      12'hCE4: dout <= 8'b10011110; // 3300 : 158 - 0x9e
      12'hCE5: dout <= 8'b10111111; // 3301 : 191 - 0xbf
      12'hCE6: dout <= 8'b10110000; // 3302 : 176 - 0xb0
      12'hCE7: dout <= 8'b10110011; // 3303 : 179 - 0xb3
      12'hCE8: dout <= 8'b00000000; // 3304 :   0 - 0x0 -- plane 1
      12'hCE9: dout <= 8'b00000001; // 3305 :   1 - 0x1
      12'hCEA: dout <= 8'b00011011; // 3306 :  27 - 0x1b
      12'hCEB: dout <= 8'b00010011; // 3307 :  19 - 0x13
      12'hCEC: dout <= 8'b00011111; // 3308 :  31 - 0x1f
      12'hCED: dout <= 8'b00111111; // 3309 :  63 - 0x3f
      12'hCEE: dout <= 8'b00111111; // 3310 :  63 - 0x3f
      12'hCEF: dout <= 8'b00111111; // 3311 :  63 - 0x3f
      12'hCF0: dout <= 8'b00000111; // 3312 :   7 - 0x7 -- Sprite 0xcf
      12'hCF1: dout <= 8'b11110011; // 3313 : 243 - 0xf3
      12'hCF2: dout <= 8'b00001011; // 3314 :  11 - 0xb
      12'hCF3: dout <= 8'b01111011; // 3315 : 123 - 0x7b
      12'hCF4: dout <= 8'b01111011; // 3316 : 123 - 0x7b
      12'hCF5: dout <= 8'b11111001; // 3317 : 249 - 0xf9
      12'hCF6: dout <= 8'b00001101; // 3318 :  13 - 0xd
      12'hCF7: dout <= 8'b11101101; // 3319 : 237 - 0xed
      12'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0 -- plane 1
      12'hCF9: dout <= 8'b11111000; // 3321 : 248 - 0xf8
      12'hCFA: dout <= 8'b00001000; // 3322 :   8 - 0x8
      12'hCFB: dout <= 8'b00001000; // 3323 :   8 - 0x8
      12'hCFC: dout <= 8'b00001000; // 3324 :   8 - 0x8
      12'hCFD: dout <= 8'b11111000; // 3325 : 248 - 0xf8
      12'hCFE: dout <= 8'b11110000; // 3326 : 240 - 0xf0
      12'hCFF: dout <= 8'b11010000; // 3327 : 208 - 0xd0
      12'hD00: dout <= 8'b11111111; // 3328 : 255 - 0xff -- Sprite 0xd0
      12'hD01: dout <= 8'b11111111; // 3329 : 255 - 0xff
      12'hD02: dout <= 8'b11111111; // 3330 : 255 - 0xff
      12'hD03: dout <= 8'b11111111; // 3331 : 255 - 0xff
      12'hD04: dout <= 8'b11101110; // 3332 : 238 - 0xee
      12'hD05: dout <= 8'b11101110; // 3333 : 238 - 0xee
      12'hD06: dout <= 8'b11101110; // 3334 : 238 - 0xee
      12'hD07: dout <= 8'b11101110; // 3335 : 238 - 0xee
      12'hD08: dout <= 8'b00000000; // 3336 :   0 - 0x0 -- plane 1
      12'hD09: dout <= 8'b00000000; // 3337 :   0 - 0x0
      12'hD0A: dout <= 8'b01111100; // 3338 : 124 - 0x7c
      12'hD0B: dout <= 8'b11111110; // 3339 : 254 - 0xfe
      12'hD0C: dout <= 8'b11101110; // 3340 : 238 - 0xee
      12'hD0D: dout <= 8'b11101110; // 3341 : 238 - 0xee
      12'hD0E: dout <= 8'b11101110; // 3342 : 238 - 0xee
      12'hD0F: dout <= 8'b11101110; // 3343 : 238 - 0xee
      12'hD10: dout <= 8'b11111111; // 3344 : 255 - 0xff -- Sprite 0xd1
      12'hD11: dout <= 8'b11111111; // 3345 : 255 - 0xff
      12'hD12: dout <= 8'b11111111; // 3346 : 255 - 0xff
      12'hD13: dout <= 8'b11111011; // 3347 : 251 - 0xfb
      12'hD14: dout <= 8'b11111011; // 3348 : 251 - 0xfb
      12'hD15: dout <= 8'b11111011; // 3349 : 251 - 0xfb
      12'hD16: dout <= 8'b11111011; // 3350 : 251 - 0xfb
      12'hD17: dout <= 8'b11111011; // 3351 : 251 - 0xfb
      12'hD18: dout <= 8'b00000000; // 3352 :   0 - 0x0 -- plane 1
      12'hD19: dout <= 8'b00000000; // 3353 :   0 - 0x0
      12'hD1A: dout <= 8'b00111000; // 3354 :  56 - 0x38
      12'hD1B: dout <= 8'b01111000; // 3355 : 120 - 0x78
      12'hD1C: dout <= 8'b01111000; // 3356 : 120 - 0x78
      12'hD1D: dout <= 8'b00111000; // 3357 :  56 - 0x38
      12'hD1E: dout <= 8'b00111000; // 3358 :  56 - 0x38
      12'hD1F: dout <= 8'b00111000; // 3359 :  56 - 0x38
      12'hD20: dout <= 8'b11111111; // 3360 : 255 - 0xff -- Sprite 0xd2
      12'hD21: dout <= 8'b11111111; // 3361 : 255 - 0xff
      12'hD22: dout <= 8'b11111111; // 3362 : 255 - 0xff
      12'hD23: dout <= 8'b11111111; // 3363 : 255 - 0xff
      12'hD24: dout <= 8'b11101110; // 3364 : 238 - 0xee
      12'hD25: dout <= 8'b10001110; // 3365 : 142 - 0x8e
      12'hD26: dout <= 8'b11111110; // 3366 : 254 - 0xfe
      12'hD27: dout <= 8'b11111110; // 3367 : 254 - 0xfe
      12'hD28: dout <= 8'b00000000; // 3368 :   0 - 0x0 -- plane 1
      12'hD29: dout <= 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout <= 8'b01111100; // 3370 : 124 - 0x7c
      12'hD2B: dout <= 8'b11111110; // 3371 : 254 - 0xfe
      12'hD2C: dout <= 8'b11101110; // 3372 : 238 - 0xee
      12'hD2D: dout <= 8'b00001110; // 3373 :  14 - 0xe
      12'hD2E: dout <= 8'b00001110; // 3374 :  14 - 0xe
      12'hD2F: dout <= 8'b01111110; // 3375 : 126 - 0x7e
      12'hD30: dout <= 8'b11111111; // 3376 : 255 - 0xff -- Sprite 0xd3
      12'hD31: dout <= 8'b11111111; // 3377 : 255 - 0xff
      12'hD32: dout <= 8'b11111111; // 3378 : 255 - 0xff
      12'hD33: dout <= 8'b11111111; // 3379 : 255 - 0xff
      12'hD34: dout <= 8'b11101110; // 3380 : 238 - 0xee
      12'hD35: dout <= 8'b10001110; // 3381 : 142 - 0x8e
      12'hD36: dout <= 8'b11111100; // 3382 : 252 - 0xfc
      12'hD37: dout <= 8'b11111101; // 3383 : 253 - 0xfd
      12'hD38: dout <= 8'b00000000; // 3384 :   0 - 0x0 -- plane 1
      12'hD39: dout <= 8'b00000000; // 3385 :   0 - 0x0
      12'hD3A: dout <= 8'b01111100; // 3386 : 124 - 0x7c
      12'hD3B: dout <= 8'b11111110; // 3387 : 254 - 0xfe
      12'hD3C: dout <= 8'b11101110; // 3388 : 238 - 0xee
      12'hD3D: dout <= 8'b00001110; // 3389 :  14 - 0xe
      12'hD3E: dout <= 8'b00111100; // 3390 :  60 - 0x3c
      12'hD3F: dout <= 8'b00111100; // 3391 :  60 - 0x3c
      12'hD40: dout <= 8'b11111111; // 3392 : 255 - 0xff -- Sprite 0xd4
      12'hD41: dout <= 8'b11111111; // 3393 : 255 - 0xff
      12'hD42: dout <= 8'b11111111; // 3394 : 255 - 0xff
      12'hD43: dout <= 8'b11111110; // 3395 : 254 - 0xfe
      12'hD44: dout <= 8'b11101110; // 3396 : 238 - 0xee
      12'hD45: dout <= 8'b11101110; // 3397 : 238 - 0xee
      12'hD46: dout <= 8'b11101110; // 3398 : 238 - 0xee
      12'hD47: dout <= 8'b11101110; // 3399 : 238 - 0xee
      12'hD48: dout <= 8'b00000000; // 3400 :   0 - 0x0 -- plane 1
      12'hD49: dout <= 8'b00000000; // 3401 :   0 - 0x0
      12'hD4A: dout <= 8'b00111110; // 3402 :  62 - 0x3e
      12'hD4B: dout <= 8'b01111110; // 3403 : 126 - 0x7e
      12'hD4C: dout <= 8'b11101110; // 3404 : 238 - 0xee
      12'hD4D: dout <= 8'b11101110; // 3405 : 238 - 0xee
      12'hD4E: dout <= 8'b11101110; // 3406 : 238 - 0xee
      12'hD4F: dout <= 8'b11101110; // 3407 : 238 - 0xee
      12'hD50: dout <= 8'b11111111; // 3408 : 255 - 0xff -- Sprite 0xd5
      12'hD51: dout <= 8'b11111111; // 3409 : 255 - 0xff
      12'hD52: dout <= 8'b11111111; // 3410 : 255 - 0xff
      12'hD53: dout <= 8'b11111101; // 3411 : 253 - 0xfd
      12'hD54: dout <= 8'b11100001; // 3412 : 225 - 0xe1
      12'hD55: dout <= 8'b11101111; // 3413 : 239 - 0xef
      12'hD56: dout <= 8'b11111111; // 3414 : 255 - 0xff
      12'hD57: dout <= 8'b11111111; // 3415 : 255 - 0xff
      12'hD58: dout <= 8'b00000000; // 3416 :   0 - 0x0 -- plane 1
      12'hD59: dout <= 8'b00000000; // 3417 :   0 - 0x0
      12'hD5A: dout <= 8'b11111100; // 3418 : 252 - 0xfc
      12'hD5B: dout <= 8'b11111100; // 3419 : 252 - 0xfc
      12'hD5C: dout <= 8'b11100000; // 3420 : 224 - 0xe0
      12'hD5D: dout <= 8'b11100000; // 3421 : 224 - 0xe0
      12'hD5E: dout <= 8'b11111100; // 3422 : 252 - 0xfc
      12'hD5F: dout <= 8'b11111110; // 3423 : 254 - 0xfe
      12'hD60: dout <= 8'b11111111; // 3424 : 255 - 0xff -- Sprite 0xd6
      12'hD61: dout <= 8'b11111111; // 3425 : 255 - 0xff
      12'hD62: dout <= 8'b11111111; // 3426 : 255 - 0xff
      12'hD63: dout <= 8'b11111101; // 3427 : 253 - 0xfd
      12'hD64: dout <= 8'b11100001; // 3428 : 225 - 0xe1
      12'hD65: dout <= 8'b11101111; // 3429 : 239 - 0xef
      12'hD66: dout <= 8'b11111111; // 3430 : 255 - 0xff
      12'hD67: dout <= 8'b11111111; // 3431 : 255 - 0xff
      12'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0 -- plane 1
      12'hD69: dout <= 8'b00000000; // 3433 :   0 - 0x0
      12'hD6A: dout <= 8'b01111100; // 3434 : 124 - 0x7c
      12'hD6B: dout <= 8'b11111100; // 3435 : 252 - 0xfc
      12'hD6C: dout <= 8'b11100000; // 3436 : 224 - 0xe0
      12'hD6D: dout <= 8'b11100000; // 3437 : 224 - 0xe0
      12'hD6E: dout <= 8'b11111100; // 3438 : 252 - 0xfc
      12'hD6F: dout <= 8'b11111110; // 3439 : 254 - 0xfe
      12'hD70: dout <= 8'b11111111; // 3440 : 255 - 0xff -- Sprite 0xd7
      12'hD71: dout <= 8'b11111111; // 3441 : 255 - 0xff
      12'hD72: dout <= 8'b11111111; // 3442 : 255 - 0xff
      12'hD73: dout <= 8'b11111110; // 3443 : 254 - 0xfe
      12'hD74: dout <= 8'b11101110; // 3444 : 238 - 0xee
      12'hD75: dout <= 8'b10001110; // 3445 : 142 - 0x8e
      12'hD76: dout <= 8'b11111110; // 3446 : 254 - 0xfe
      12'hD77: dout <= 8'b11111100; // 3447 : 252 - 0xfc
      12'hD78: dout <= 8'b00000000; // 3448 :   0 - 0x0 -- plane 1
      12'hD79: dout <= 8'b00000000; // 3449 :   0 - 0x0
      12'hD7A: dout <= 8'b11111110; // 3450 : 254 - 0xfe
      12'hD7B: dout <= 8'b11111110; // 3451 : 254 - 0xfe
      12'hD7C: dout <= 8'b11101110; // 3452 : 238 - 0xee
      12'hD7D: dout <= 8'b00001110; // 3453 :  14 - 0xe
      12'hD7E: dout <= 8'b00001110; // 3454 :  14 - 0xe
      12'hD7F: dout <= 8'b00011100; // 3455 :  28 - 0x1c
      12'hD80: dout <= 8'b11111111; // 3456 : 255 - 0xff -- Sprite 0xd8
      12'hD81: dout <= 8'b11111111; // 3457 : 255 - 0xff
      12'hD82: dout <= 8'b11111111; // 3458 : 255 - 0xff
      12'hD83: dout <= 8'b11111111; // 3459 : 255 - 0xff
      12'hD84: dout <= 8'b11101110; // 3460 : 238 - 0xee
      12'hD85: dout <= 8'b11101110; // 3461 : 238 - 0xee
      12'hD86: dout <= 8'b11111100; // 3462 : 252 - 0xfc
      12'hD87: dout <= 8'b11111111; // 3463 : 255 - 0xff
      12'hD88: dout <= 8'b00000000; // 3464 :   0 - 0x0 -- plane 1
      12'hD89: dout <= 8'b00000000; // 3465 :   0 - 0x0
      12'hD8A: dout <= 8'b01111100; // 3466 : 124 - 0x7c
      12'hD8B: dout <= 8'b11111110; // 3467 : 254 - 0xfe
      12'hD8C: dout <= 8'b11101110; // 3468 : 238 - 0xee
      12'hD8D: dout <= 8'b11101110; // 3469 : 238 - 0xee
      12'hD8E: dout <= 8'b01111100; // 3470 : 124 - 0x7c
      12'hD8F: dout <= 8'b11111110; // 3471 : 254 - 0xfe
      12'hD90: dout <= 8'b11111111; // 3472 : 255 - 0xff -- Sprite 0xd9
      12'hD91: dout <= 8'b11111111; // 3473 : 255 - 0xff
      12'hD92: dout <= 8'b11111111; // 3474 : 255 - 0xff
      12'hD93: dout <= 8'b11111111; // 3475 : 255 - 0xff
      12'hD94: dout <= 8'b11101110; // 3476 : 238 - 0xee
      12'hD95: dout <= 8'b11101110; // 3477 : 238 - 0xee
      12'hD96: dout <= 8'b11101110; // 3478 : 238 - 0xee
      12'hD97: dout <= 8'b11101110; // 3479 : 238 - 0xee
      12'hD98: dout <= 8'b00000000; // 3480 :   0 - 0x0 -- plane 1
      12'hD99: dout <= 8'b00000000; // 3481 :   0 - 0x0
      12'hD9A: dout <= 8'b01111100; // 3482 : 124 - 0x7c
      12'hD9B: dout <= 8'b11111110; // 3483 : 254 - 0xfe
      12'hD9C: dout <= 8'b11101110; // 3484 : 238 - 0xee
      12'hD9D: dout <= 8'b11101110; // 3485 : 238 - 0xee
      12'hD9E: dout <= 8'b11101110; // 3486 : 238 - 0xee
      12'hD9F: dout <= 8'b11101110; // 3487 : 238 - 0xee
      12'hDA0: dout <= 8'b00000000; // 3488 :   0 - 0x0 -- Sprite 0xda
      12'hDA1: dout <= 8'b00000000; // 3489 :   0 - 0x0
      12'hDA2: dout <= 8'b00000000; // 3490 :   0 - 0x0
      12'hDA3: dout <= 8'b10000000; // 3491 : 128 - 0x80
      12'hDA4: dout <= 8'b00000000; // 3492 :   0 - 0x0
      12'hDA5: dout <= 8'b00000000; // 3493 :   0 - 0x0
      12'hDA6: dout <= 8'b00000100; // 3494 :   4 - 0x4
      12'hDA7: dout <= 8'b00000000; // 3495 :   0 - 0x0
      12'hDA8: dout <= 8'b00000000; // 3496 :   0 - 0x0 -- plane 1
      12'hDA9: dout <= 8'b00100000; // 3497 :  32 - 0x20
      12'hDAA: dout <= 8'b00000000; // 3498 :   0 - 0x0
      12'hDAB: dout <= 8'b00000010; // 3499 :   2 - 0x2
      12'hDAC: dout <= 8'b00000000; // 3500 :   0 - 0x0
      12'hDAD: dout <= 8'b00100000; // 3501 :  32 - 0x20
      12'hDAE: dout <= 8'b00000000; // 3502 :   0 - 0x0
      12'hDAF: dout <= 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout <= 8'b00000000; // 3504 :   0 - 0x0 -- Sprite 0xdb
      12'hDB1: dout <= 8'b00000100; // 3505 :   4 - 0x4
      12'hDB2: dout <= 8'b00000000; // 3506 :   0 - 0x0
      12'hDB3: dout <= 8'b00010001; // 3507 :  17 - 0x11
      12'hDB4: dout <= 8'b00000000; // 3508 :   0 - 0x0
      12'hDB5: dout <= 8'b00000000; // 3509 :   0 - 0x0
      12'hDB6: dout <= 8'b00000000; // 3510 :   0 - 0x0
      12'hDB7: dout <= 8'b00100000; // 3511 :  32 - 0x20
      12'hDB8: dout <= 8'b00100000; // 3512 :  32 - 0x20 -- plane 1
      12'hDB9: dout <= 8'b00000000; // 3513 :   0 - 0x0
      12'hDBA: dout <= 8'b00000000; // 3514 :   0 - 0x0
      12'hDBB: dout <= 8'b00000000; // 3515 :   0 - 0x0
      12'hDBC: dout <= 8'b10000000; // 3516 : 128 - 0x80
      12'hDBD: dout <= 8'b00000000; // 3517 :   0 - 0x0
      12'hDBE: dout <= 8'b00000100; // 3518 :   4 - 0x4
      12'hDBF: dout <= 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout <= 8'b00000000; // 3520 :   0 - 0x0 -- Sprite 0xdc
      12'hDC1: dout <= 8'b00000000; // 3521 :   0 - 0x0
      12'hDC2: dout <= 8'b00000000; // 3522 :   0 - 0x0
      12'hDC3: dout <= 8'b00100000; // 3523 :  32 - 0x20
      12'hDC4: dout <= 8'b00000000; // 3524 :   0 - 0x0
      12'hDC5: dout <= 8'b00000000; // 3525 :   0 - 0x0
      12'hDC6: dout <= 8'b00000000; // 3526 :   0 - 0x0
      12'hDC7: dout <= 8'b00000100; // 3527 :   4 - 0x4
      12'hDC8: dout <= 8'b00000000; // 3528 :   0 - 0x0 -- plane 1
      12'hDC9: dout <= 8'b00001000; // 3529 :   8 - 0x8
      12'hDCA: dout <= 8'b00000000; // 3530 :   0 - 0x0
      12'hDCB: dout <= 8'b00000000; // 3531 :   0 - 0x0
      12'hDCC: dout <= 8'b00000010; // 3532 :   2 - 0x2
      12'hDCD: dout <= 8'b00000000; // 3533 :   0 - 0x0
      12'hDCE: dout <= 8'b01000000; // 3534 :  64 - 0x40
      12'hDCF: dout <= 8'b00000000; // 3535 :   0 - 0x0
      12'hDD0: dout <= 8'b00000000; // 3536 :   0 - 0x0 -- Sprite 0xdd
      12'hDD1: dout <= 8'b00000000; // 3537 :   0 - 0x0
      12'hDD2: dout <= 8'b00010001; // 3538 :  17 - 0x11
      12'hDD3: dout <= 8'b00000000; // 3539 :   0 - 0x0
      12'hDD4: dout <= 8'b00000000; // 3540 :   0 - 0x0
      12'hDD5: dout <= 8'b10000000; // 3541 : 128 - 0x80
      12'hDD6: dout <= 8'b00000000; // 3542 :   0 - 0x0
      12'hDD7: dout <= 8'b00000000; // 3543 :   0 - 0x0
      12'hDD8: dout <= 8'b00000000; // 3544 :   0 - 0x0 -- plane 1
      12'hDD9: dout <= 8'b01000000; // 3545 :  64 - 0x40
      12'hDDA: dout <= 8'b00000000; // 3546 :   0 - 0x0
      12'hDDB: dout <= 8'b00000000; // 3547 :   0 - 0x0
      12'hDDC: dout <= 8'b00000000; // 3548 :   0 - 0x0
      12'hDDD: dout <= 8'b00000000; // 3549 :   0 - 0x0
      12'hDDE: dout <= 8'b00000010; // 3550 :   2 - 0x2
      12'hDDF: dout <= 8'b00100000; // 3551 :  32 - 0x20
      12'hDE0: dout <= 8'b10110011; // 3552 : 179 - 0xb3 -- Sprite 0xde
      12'hDE1: dout <= 8'b10110011; // 3553 : 179 - 0xb3
      12'hDE2: dout <= 8'b10110011; // 3554 : 179 - 0xb3
      12'hDE3: dout <= 8'b10110011; // 3555 : 179 - 0xb3
      12'hDE4: dout <= 8'b10110000; // 3556 : 176 - 0xb0
      12'hDE5: dout <= 8'b10101111; // 3557 : 175 - 0xaf
      12'hDE6: dout <= 8'b10011111; // 3558 : 159 - 0x9f
      12'hDE7: dout <= 8'b11000000; // 3559 : 192 - 0xc0
      12'hDE8: dout <= 8'b00111110; // 3560 :  62 - 0x3e -- plane 1
      12'hDE9: dout <= 8'b00111111; // 3561 :  63 - 0x3f
      12'hDEA: dout <= 8'b00111110; // 3562 :  62 - 0x3e
      12'hDEB: dout <= 8'b00111100; // 3563 :  60 - 0x3c
      12'hDEC: dout <= 8'b00111111; // 3564 :  63 - 0x3f
      12'hDED: dout <= 8'b00110000; // 3565 :  48 - 0x30
      12'hDEE: dout <= 8'b00000000; // 3566 :   0 - 0x0
      12'hDEF: dout <= 8'b00000000; // 3567 :   0 - 0x0
      12'hDF0: dout <= 8'b11101101; // 3568 : 237 - 0xed -- Sprite 0xdf
      12'hDF1: dout <= 8'b11001101; // 3569 : 205 - 0xcd
      12'hDF2: dout <= 8'b11001101; // 3570 : 205 - 0xcd
      12'hDF3: dout <= 8'b00001101; // 3571 :  13 - 0xd
      12'hDF4: dout <= 8'b00001101; // 3572 :  13 - 0xd
      12'hDF5: dout <= 8'b11111101; // 3573 : 253 - 0xfd
      12'hDF6: dout <= 8'b11111101; // 3574 : 253 - 0xfd
      12'hDF7: dout <= 8'b00000011; // 3575 :   3 - 0x3
      12'hDF8: dout <= 8'b00010000; // 3576 :  16 - 0x10 -- plane 1
      12'hDF9: dout <= 8'b10110000; // 3577 : 176 - 0xb0
      12'hDFA: dout <= 8'b00110000; // 3578 :  48 - 0x30
      12'hDFB: dout <= 8'b11110000; // 3579 : 240 - 0xf0
      12'hDFC: dout <= 8'b11110000; // 3580 : 240 - 0xf0
      12'hDFD: dout <= 8'b00000000; // 3581 :   0 - 0x0
      12'hDFE: dout <= 8'b00000000; // 3582 :   0 - 0x0
      12'hDFF: dout <= 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout <= 8'b11101110; // 3584 : 238 - 0xee -- Sprite 0xe0
      12'hE01: dout <= 8'b11101110; // 3585 : 238 - 0xee
      12'hE02: dout <= 8'b11101110; // 3586 : 238 - 0xee
      12'hE03: dout <= 8'b11101110; // 3587 : 238 - 0xee
      12'hE04: dout <= 8'b11111110; // 3588 : 254 - 0xfe
      12'hE05: dout <= 8'b11111100; // 3589 : 252 - 0xfc
      12'hE06: dout <= 8'b11000001; // 3590 : 193 - 0xc1
      12'hE07: dout <= 8'b11111111; // 3591 : 255 - 0xff
      12'hE08: dout <= 8'b11101110; // 3592 : 238 - 0xee -- plane 1
      12'hE09: dout <= 8'b11101110; // 3593 : 238 - 0xee
      12'hE0A: dout <= 8'b11101110; // 3594 : 238 - 0xee
      12'hE0B: dout <= 8'b11101110; // 3595 : 238 - 0xee
      12'hE0C: dout <= 8'b11111110; // 3596 : 254 - 0xfe
      12'hE0D: dout <= 8'b01111100; // 3597 : 124 - 0x7c
      12'hE0E: dout <= 8'b00000000; // 3598 :   0 - 0x0
      12'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout <= 8'b11111011; // 3600 : 251 - 0xfb -- Sprite 0xe1
      12'hE11: dout <= 8'b11111011; // 3601 : 251 - 0xfb
      12'hE12: dout <= 8'b11111011; // 3602 : 251 - 0xfb
      12'hE13: dout <= 8'b11111011; // 3603 : 251 - 0xfb
      12'hE14: dout <= 8'b11111111; // 3604 : 255 - 0xff
      12'hE15: dout <= 8'b11111101; // 3605 : 253 - 0xfd
      12'hE16: dout <= 8'b11000001; // 3606 : 193 - 0xc1
      12'hE17: dout <= 8'b11111111; // 3607 : 255 - 0xff
      12'hE18: dout <= 8'b00111000; // 3608 :  56 - 0x38 -- plane 1
      12'hE19: dout <= 8'b00111000; // 3609 :  56 - 0x38
      12'hE1A: dout <= 8'b00111000; // 3610 :  56 - 0x38
      12'hE1B: dout <= 8'b00111000; // 3611 :  56 - 0x38
      12'hE1C: dout <= 8'b01111100; // 3612 : 124 - 0x7c
      12'hE1D: dout <= 8'b01111100; // 3613 : 124 - 0x7c
      12'hE1E: dout <= 8'b00000000; // 3614 :   0 - 0x0
      12'hE1F: dout <= 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout <= 8'b11111100; // 3616 : 252 - 0xfc -- Sprite 0xe2
      12'hE21: dout <= 8'b11100001; // 3617 : 225 - 0xe1
      12'hE22: dout <= 8'b11101111; // 3618 : 239 - 0xef
      12'hE23: dout <= 8'b11101111; // 3619 : 239 - 0xef
      12'hE24: dout <= 8'b11111111; // 3620 : 255 - 0xff
      12'hE25: dout <= 8'b11111110; // 3621 : 254 - 0xfe
      12'hE26: dout <= 8'b10000000; // 3622 : 128 - 0x80
      12'hE27: dout <= 8'b11111111; // 3623 : 255 - 0xff
      12'hE28: dout <= 8'b11111100; // 3624 : 252 - 0xfc -- plane 1
      12'hE29: dout <= 8'b11100000; // 3625 : 224 - 0xe0
      12'hE2A: dout <= 8'b11100000; // 3626 : 224 - 0xe0
      12'hE2B: dout <= 8'b11100000; // 3627 : 224 - 0xe0
      12'hE2C: dout <= 8'b11111110; // 3628 : 254 - 0xfe
      12'hE2D: dout <= 8'b11111110; // 3629 : 254 - 0xfe
      12'hE2E: dout <= 8'b00000000; // 3630 :   0 - 0x0
      12'hE2F: dout <= 8'b00000000; // 3631 :   0 - 0x0
      12'hE30: dout <= 8'b11101110; // 3632 : 238 - 0xee -- Sprite 0xe3
      12'hE31: dout <= 8'b11111110; // 3633 : 254 - 0xfe
      12'hE32: dout <= 8'b11111110; // 3634 : 254 - 0xfe
      12'hE33: dout <= 8'b11111110; // 3635 : 254 - 0xfe
      12'hE34: dout <= 8'b11111110; // 3636 : 254 - 0xfe
      12'hE35: dout <= 8'b11111100; // 3637 : 252 - 0xfc
      12'hE36: dout <= 8'b11000001; // 3638 : 193 - 0xc1
      12'hE37: dout <= 8'b11111111; // 3639 : 255 - 0xff
      12'hE38: dout <= 8'b00001110; // 3640 :  14 - 0xe -- plane 1
      12'hE39: dout <= 8'b00001110; // 3641 :  14 - 0xe
      12'hE3A: dout <= 8'b00001110; // 3642 :  14 - 0xe
      12'hE3B: dout <= 8'b11101110; // 3643 : 238 - 0xee
      12'hE3C: dout <= 8'b11111110; // 3644 : 254 - 0xfe
      12'hE3D: dout <= 8'b01111100; // 3645 : 124 - 0x7c
      12'hE3E: dout <= 8'b00000000; // 3646 :   0 - 0x0
      12'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout <= 8'b11101110; // 3648 : 238 - 0xee -- Sprite 0xe4
      12'hE41: dout <= 8'b11101110; // 3649 : 238 - 0xee
      12'hE42: dout <= 8'b11111110; // 3650 : 254 - 0xfe
      12'hE43: dout <= 8'b11111110; // 3651 : 254 - 0xfe
      12'hE44: dout <= 8'b10001110; // 3652 : 142 - 0x8e
      12'hE45: dout <= 8'b11111110; // 3653 : 254 - 0xfe
      12'hE46: dout <= 8'b11111000; // 3654 : 248 - 0xf8
      12'hE47: dout <= 8'b11111111; // 3655 : 255 - 0xff
      12'hE48: dout <= 8'b11101110; // 3656 : 238 - 0xee -- plane 1
      12'hE49: dout <= 8'b11101110; // 3657 : 238 - 0xee
      12'hE4A: dout <= 8'b11111110; // 3658 : 254 - 0xfe
      12'hE4B: dout <= 8'b11111110; // 3659 : 254 - 0xfe
      12'hE4C: dout <= 8'b00001110; // 3660 :  14 - 0xe
      12'hE4D: dout <= 8'b00001110; // 3661 :  14 - 0xe
      12'hE4E: dout <= 8'b00000000; // 3662 :   0 - 0x0
      12'hE4F: dout <= 8'b00000000; // 3663 :   0 - 0x0
      12'hE50: dout <= 8'b10001110; // 3664 : 142 - 0x8e -- Sprite 0xe5
      12'hE51: dout <= 8'b11111110; // 3665 : 254 - 0xfe
      12'hE52: dout <= 8'b11111110; // 3666 : 254 - 0xfe
      12'hE53: dout <= 8'b11111110; // 3667 : 254 - 0xfe
      12'hE54: dout <= 8'b11111110; // 3668 : 254 - 0xfe
      12'hE55: dout <= 8'b11111100; // 3669 : 252 - 0xfc
      12'hE56: dout <= 8'b11000001; // 3670 : 193 - 0xc1
      12'hE57: dout <= 8'b11111111; // 3671 : 255 - 0xff
      12'hE58: dout <= 8'b00001110; // 3672 :  14 - 0xe -- plane 1
      12'hE59: dout <= 8'b00001110; // 3673 :  14 - 0xe
      12'hE5A: dout <= 8'b00001110; // 3674 :  14 - 0xe
      12'hE5B: dout <= 8'b11101110; // 3675 : 238 - 0xee
      12'hE5C: dout <= 8'b11111110; // 3676 : 254 - 0xfe
      12'hE5D: dout <= 8'b01111100; // 3677 : 124 - 0x7c
      12'hE5E: dout <= 8'b00000000; // 3678 :   0 - 0x0
      12'hE5F: dout <= 8'b00000000; // 3679 :   0 - 0x0
      12'hE60: dout <= 8'b11101110; // 3680 : 238 - 0xee -- Sprite 0xe6
      12'hE61: dout <= 8'b11101110; // 3681 : 238 - 0xee
      12'hE62: dout <= 8'b11101110; // 3682 : 238 - 0xee
      12'hE63: dout <= 8'b11101110; // 3683 : 238 - 0xee
      12'hE64: dout <= 8'b11111110; // 3684 : 254 - 0xfe
      12'hE65: dout <= 8'b11111100; // 3685 : 252 - 0xfc
      12'hE66: dout <= 8'b11000001; // 3686 : 193 - 0xc1
      12'hE67: dout <= 8'b11111111; // 3687 : 255 - 0xff
      12'hE68: dout <= 8'b11101110; // 3688 : 238 - 0xee -- plane 1
      12'hE69: dout <= 8'b11101110; // 3689 : 238 - 0xee
      12'hE6A: dout <= 8'b11101110; // 3690 : 238 - 0xee
      12'hE6B: dout <= 8'b11101110; // 3691 : 238 - 0xee
      12'hE6C: dout <= 8'b11111110; // 3692 : 254 - 0xfe
      12'hE6D: dout <= 8'b01111100; // 3693 : 124 - 0x7c
      12'hE6E: dout <= 8'b00000000; // 3694 :   0 - 0x0
      12'hE6F: dout <= 8'b00000000; // 3695 :   0 - 0x0
      12'hE70: dout <= 8'b11111101; // 3696 : 253 - 0xfd -- Sprite 0xe7
      12'hE71: dout <= 8'b11111101; // 3697 : 253 - 0xfd
      12'hE72: dout <= 8'b11111001; // 3698 : 249 - 0xf9
      12'hE73: dout <= 8'b11111011; // 3699 : 251 - 0xfb
      12'hE74: dout <= 8'b11111011; // 3700 : 251 - 0xfb
      12'hE75: dout <= 8'b11111011; // 3701 : 251 - 0xfb
      12'hE76: dout <= 8'b11100011; // 3702 : 227 - 0xe3
      12'hE77: dout <= 8'b11111111; // 3703 : 255 - 0xff
      12'hE78: dout <= 8'b00011100; // 3704 :  28 - 0x1c -- plane 1
      12'hE79: dout <= 8'b00011100; // 3705 :  28 - 0x1c
      12'hE7A: dout <= 8'b00111000; // 3706 :  56 - 0x38
      12'hE7B: dout <= 8'b00111000; // 3707 :  56 - 0x38
      12'hE7C: dout <= 8'b00111000; // 3708 :  56 - 0x38
      12'hE7D: dout <= 8'b00111000; // 3709 :  56 - 0x38
      12'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout <= 8'b11101110; // 3712 : 238 - 0xee -- Sprite 0xe8
      12'hE81: dout <= 8'b11101110; // 3713 : 238 - 0xee
      12'hE82: dout <= 8'b11101110; // 3714 : 238 - 0xee
      12'hE83: dout <= 8'b11101110; // 3715 : 238 - 0xee
      12'hE84: dout <= 8'b11111110; // 3716 : 254 - 0xfe
      12'hE85: dout <= 8'b11111100; // 3717 : 252 - 0xfc
      12'hE86: dout <= 8'b11000001; // 3718 : 193 - 0xc1
      12'hE87: dout <= 8'b11111111; // 3719 : 255 - 0xff
      12'hE88: dout <= 8'b11101110; // 3720 : 238 - 0xee -- plane 1
      12'hE89: dout <= 8'b11101110; // 3721 : 238 - 0xee
      12'hE8A: dout <= 8'b11101110; // 3722 : 238 - 0xee
      12'hE8B: dout <= 8'b11101110; // 3723 : 238 - 0xee
      12'hE8C: dout <= 8'b11111110; // 3724 : 254 - 0xfe
      12'hE8D: dout <= 8'b01111100; // 3725 : 124 - 0x7c
      12'hE8E: dout <= 8'b00000000; // 3726 :   0 - 0x0
      12'hE8F: dout <= 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout <= 8'b11111110; // 3728 : 254 - 0xfe -- Sprite 0xe9
      12'hE91: dout <= 8'b11111110; // 3729 : 254 - 0xfe
      12'hE92: dout <= 8'b11001110; // 3730 : 206 - 0xce
      12'hE93: dout <= 8'b11111110; // 3731 : 254 - 0xfe
      12'hE94: dout <= 8'b11111110; // 3732 : 254 - 0xfe
      12'hE95: dout <= 8'b11111100; // 3733 : 252 - 0xfc
      12'hE96: dout <= 8'b11000001; // 3734 : 193 - 0xc1
      12'hE97: dout <= 8'b11111111; // 3735 : 255 - 0xff
      12'hE98: dout <= 8'b11111110; // 3736 : 254 - 0xfe -- plane 1
      12'hE99: dout <= 8'b01111110; // 3737 : 126 - 0x7e
      12'hE9A: dout <= 8'b00001110; // 3738 :  14 - 0xe
      12'hE9B: dout <= 8'b00001110; // 3739 :  14 - 0xe
      12'hE9C: dout <= 8'b01111110; // 3740 : 126 - 0x7e
      12'hE9D: dout <= 8'b01111100; // 3741 : 124 - 0x7c
      12'hE9E: dout <= 8'b00000000; // 3742 :   0 - 0x0
      12'hE9F: dout <= 8'b00000000; // 3743 :   0 - 0x0
      12'hEA0: dout <= 8'b00000000; // 3744 :   0 - 0x0 -- Sprite 0xea
      12'hEA1: dout <= 8'b01110000; // 3745 : 112 - 0x70
      12'hEA2: dout <= 8'b00111000; // 3746 :  56 - 0x38
      12'hEA3: dout <= 8'b00000000; // 3747 :   0 - 0x0
      12'hEA4: dout <= 8'b00000010; // 3748 :   2 - 0x2
      12'hEA5: dout <= 8'b00000111; // 3749 :   7 - 0x7
      12'hEA6: dout <= 8'b00000011; // 3750 :   3 - 0x3
      12'hEA7: dout <= 8'b00000000; // 3751 :   0 - 0x0
      12'hEA8: dout <= 8'b00000000; // 3752 :   0 - 0x0 -- plane 1
      12'hEA9: dout <= 8'b01110000; // 3753 : 112 - 0x70
      12'hEAA: dout <= 8'b00111000; // 3754 :  56 - 0x38
      12'hEAB: dout <= 8'b00000000; // 3755 :   0 - 0x0
      12'hEAC: dout <= 8'b00000010; // 3756 :   2 - 0x2
      12'hEAD: dout <= 8'b00000111; // 3757 :   7 - 0x7
      12'hEAE: dout <= 8'b00000011; // 3758 :   3 - 0x3
      12'hEAF: dout <= 8'b00000000; // 3759 :   0 - 0x0
      12'hEB0: dout <= 8'b00000000; // 3760 :   0 - 0x0 -- Sprite 0xeb
      12'hEB1: dout <= 8'b00001100; // 3761 :  12 - 0xc
      12'hEB2: dout <= 8'b00000110; // 3762 :   6 - 0x6
      12'hEB3: dout <= 8'b00000110; // 3763 :   6 - 0x6
      12'hEB4: dout <= 8'b01100000; // 3764 :  96 - 0x60
      12'hEB5: dout <= 8'b01110000; // 3765 : 112 - 0x70
      12'hEB6: dout <= 8'b00110000; // 3766 :  48 - 0x30
      12'hEB7: dout <= 8'b00000000; // 3767 :   0 - 0x0
      12'hEB8: dout <= 8'b00000000; // 3768 :   0 - 0x0 -- plane 1
      12'hEB9: dout <= 8'b00001100; // 3769 :  12 - 0xc
      12'hEBA: dout <= 8'b00000110; // 3770 :   6 - 0x6
      12'hEBB: dout <= 8'b00000110; // 3771 :   6 - 0x6
      12'hEBC: dout <= 8'b01100000; // 3772 :  96 - 0x60
      12'hEBD: dout <= 8'b01110000; // 3773 : 112 - 0x70
      12'hEBE: dout <= 8'b00110000; // 3774 :  48 - 0x30
      12'hEBF: dout <= 8'b00000000; // 3775 :   0 - 0x0
      12'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Sprite 0xec
      12'hEC1: dout <= 8'b11000000; // 3777 : 192 - 0xc0
      12'hEC2: dout <= 8'b11100000; // 3778 : 224 - 0xe0
      12'hEC3: dout <= 8'b01100000; // 3779 :  96 - 0x60
      12'hEC4: dout <= 8'b00000000; // 3780 :   0 - 0x0
      12'hEC5: dout <= 8'b00001100; // 3781 :  12 - 0xc
      12'hEC6: dout <= 8'b00001110; // 3782 :  14 - 0xe
      12'hEC7: dout <= 8'b00000110; // 3783 :   6 - 0x6
      12'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0 -- plane 1
      12'hEC9: dout <= 8'b11000000; // 3785 : 192 - 0xc0
      12'hECA: dout <= 8'b11100000; // 3786 : 224 - 0xe0
      12'hECB: dout <= 8'b01100000; // 3787 :  96 - 0x60
      12'hECC: dout <= 8'b00000000; // 3788 :   0 - 0x0
      12'hECD: dout <= 8'b00001100; // 3789 :  12 - 0xc
      12'hECE: dout <= 8'b00001110; // 3790 :  14 - 0xe
      12'hECF: dout <= 8'b00000110; // 3791 :   6 - 0x6
      12'hED0: dout <= 8'b01100000; // 3792 :  96 - 0x60 -- Sprite 0xed
      12'hED1: dout <= 8'b01110000; // 3793 : 112 - 0x70
      12'hED2: dout <= 8'b00110000; // 3794 :  48 - 0x30
      12'hED3: dout <= 8'b00000000; // 3795 :   0 - 0x0
      12'hED4: dout <= 8'b00000000; // 3796 :   0 - 0x0
      12'hED5: dout <= 8'b00001100; // 3797 :  12 - 0xc
      12'hED6: dout <= 8'b00001110; // 3798 :  14 - 0xe
      12'hED7: dout <= 8'b00000110; // 3799 :   6 - 0x6
      12'hED8: dout <= 8'b01100000; // 3800 :  96 - 0x60 -- plane 1
      12'hED9: dout <= 8'b01110000; // 3801 : 112 - 0x70
      12'hEDA: dout <= 8'b00110000; // 3802 :  48 - 0x30
      12'hEDB: dout <= 8'b00000000; // 3803 :   0 - 0x0
      12'hEDC: dout <= 8'b00000000; // 3804 :   0 - 0x0
      12'hEDD: dout <= 8'b00001100; // 3805 :  12 - 0xc
      12'hEDE: dout <= 8'b00001110; // 3806 :  14 - 0xe
      12'hEDF: dout <= 8'b00000110; // 3807 :   6 - 0x6
      12'hEE0: dout <= 8'b11111111; // 3808 : 255 - 0xff -- Sprite 0xee
      12'hEE1: dout <= 8'b11111111; // 3809 : 255 - 0xff
      12'hEE2: dout <= 8'b10111101; // 3810 : 189 - 0xbd
      12'hEE3: dout <= 8'b11111111; // 3811 : 255 - 0xff
      12'hEE4: dout <= 8'b11111111; // 3812 : 255 - 0xff
      12'hEE5: dout <= 8'b11111011; // 3813 : 251 - 0xfb
      12'hEE6: dout <= 8'b11111111; // 3814 : 255 - 0xff
      12'hEE7: dout <= 8'b11111111; // 3815 : 255 - 0xff
      12'hEE8: dout <= 8'b00000000; // 3816 :   0 - 0x0 -- plane 1
      12'hEE9: dout <= 8'b00000000; // 3817 :   0 - 0x0
      12'hEEA: dout <= 8'b01000010; // 3818 :  66 - 0x42
      12'hEEB: dout <= 8'b00000000; // 3819 :   0 - 0x0
      12'hEEC: dout <= 8'b00000000; // 3820 :   0 - 0x0
      12'hEED: dout <= 8'b00000100; // 3821 :   4 - 0x4
      12'hEEE: dout <= 8'b00000000; // 3822 :   0 - 0x0
      12'hEEF: dout <= 8'b00000000; // 3823 :   0 - 0x0
      12'hEF0: dout <= 8'b11111111; // 3824 : 255 - 0xff -- Sprite 0xef
      12'hEF1: dout <= 8'b11111111; // 3825 : 255 - 0xff
      12'hEF2: dout <= 8'b11111011; // 3826 : 251 - 0xfb
      12'hEF3: dout <= 8'b11111111; // 3827 : 255 - 0xff
      12'hEF4: dout <= 8'b11011111; // 3828 : 223 - 0xdf
      12'hEF5: dout <= 8'b11111111; // 3829 : 255 - 0xff
      12'hEF6: dout <= 8'b11111111; // 3830 : 255 - 0xff
      12'hEF7: dout <= 8'b11111111; // 3831 : 255 - 0xff
      12'hEF8: dout <= 8'b00000000; // 3832 :   0 - 0x0 -- plane 1
      12'hEF9: dout <= 8'b00000000; // 3833 :   0 - 0x0
      12'hEFA: dout <= 8'b00000100; // 3834 :   4 - 0x4
      12'hEFB: dout <= 8'b00000000; // 3835 :   0 - 0x0
      12'hEFC: dout <= 8'b00100000; // 3836 :  32 - 0x20
      12'hEFD: dout <= 8'b00000000; // 3837 :   0 - 0x0
      12'hEFE: dout <= 8'b00000000; // 3838 :   0 - 0x0
      12'hEFF: dout <= 8'b00000000; // 3839 :   0 - 0x0
      12'hF00: dout <= 8'b00000000; // 3840 :   0 - 0x0 -- Sprite 0xf0
      12'hF01: dout <= 8'b00000000; // 3841 :   0 - 0x0
      12'hF02: dout <= 8'b00000000; // 3842 :   0 - 0x0
      12'hF03: dout <= 8'b00000000; // 3843 :   0 - 0x0
      12'hF04: dout <= 8'b00000000; // 3844 :   0 - 0x0
      12'hF05: dout <= 8'b00000000; // 3845 :   0 - 0x0
      12'hF06: dout <= 8'b00000000; // 3846 :   0 - 0x0
      12'hF07: dout <= 8'b00000000; // 3847 :   0 - 0x0
      12'hF08: dout <= 8'b00000000; // 3848 :   0 - 0x0 -- plane 1
      12'hF09: dout <= 8'b00000000; // 3849 :   0 - 0x0
      12'hF0A: dout <= 8'b00000000; // 3850 :   0 - 0x0
      12'hF0B: dout <= 8'b00000000; // 3851 :   0 - 0x0
      12'hF0C: dout <= 8'b00000000; // 3852 :   0 - 0x0
      12'hF0D: dout <= 8'b00000000; // 3853 :   0 - 0x0
      12'hF0E: dout <= 8'b00000000; // 3854 :   0 - 0x0
      12'hF0F: dout <= 8'b00000000; // 3855 :   0 - 0x0
      12'hF10: dout <= 8'b00000000; // 3856 :   0 - 0x0 -- Sprite 0xf1
      12'hF11: dout <= 8'b10000000; // 3857 : 128 - 0x80
      12'hF12: dout <= 8'b00000000; // 3858 :   0 - 0x0
      12'hF13: dout <= 8'b00000000; // 3859 :   0 - 0x0
      12'hF14: dout <= 8'b00000000; // 3860 :   0 - 0x0
      12'hF15: dout <= 8'b00000000; // 3861 :   0 - 0x0
      12'hF16: dout <= 8'b00000000; // 3862 :   0 - 0x0
      12'hF17: dout <= 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout <= 8'b10000000; // 3864 : 128 - 0x80 -- plane 1
      12'hF19: dout <= 8'b10000000; // 3865 : 128 - 0x80
      12'hF1A: dout <= 8'b10000000; // 3866 : 128 - 0x80
      12'hF1B: dout <= 8'b10000000; // 3867 : 128 - 0x80
      12'hF1C: dout <= 8'b00000000; // 3868 :   0 - 0x0
      12'hF1D: dout <= 8'b00000000; // 3869 :   0 - 0x0
      12'hF1E: dout <= 8'b00000000; // 3870 :   0 - 0x0
      12'hF1F: dout <= 8'b00000000; // 3871 :   0 - 0x0
      12'hF20: dout <= 8'b00000000; // 3872 :   0 - 0x0 -- Sprite 0xf2
      12'hF21: dout <= 8'b11000000; // 3873 : 192 - 0xc0
      12'hF22: dout <= 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout <= 8'b00000000; // 3875 :   0 - 0x0
      12'hF24: dout <= 8'b00000000; // 3876 :   0 - 0x0
      12'hF25: dout <= 8'b00000000; // 3877 :   0 - 0x0
      12'hF26: dout <= 8'b00000000; // 3878 :   0 - 0x0
      12'hF27: dout <= 8'b00000000; // 3879 :   0 - 0x0
      12'hF28: dout <= 8'b11000000; // 3880 : 192 - 0xc0 -- plane 1
      12'hF29: dout <= 8'b11000000; // 3881 : 192 - 0xc0
      12'hF2A: dout <= 8'b11000000; // 3882 : 192 - 0xc0
      12'hF2B: dout <= 8'b11000000; // 3883 : 192 - 0xc0
      12'hF2C: dout <= 8'b00000000; // 3884 :   0 - 0x0
      12'hF2D: dout <= 8'b00000000; // 3885 :   0 - 0x0
      12'hF2E: dout <= 8'b00000000; // 3886 :   0 - 0x0
      12'hF2F: dout <= 8'b00000000; // 3887 :   0 - 0x0
      12'hF30: dout <= 8'b00000000; // 3888 :   0 - 0x0 -- Sprite 0xf3
      12'hF31: dout <= 8'b11100000; // 3889 : 224 - 0xe0
      12'hF32: dout <= 8'b00000000; // 3890 :   0 - 0x0
      12'hF33: dout <= 8'b00000000; // 3891 :   0 - 0x0
      12'hF34: dout <= 8'b00000000; // 3892 :   0 - 0x0
      12'hF35: dout <= 8'b00000000; // 3893 :   0 - 0x0
      12'hF36: dout <= 8'b00000000; // 3894 :   0 - 0x0
      12'hF37: dout <= 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout <= 8'b11100000; // 3896 : 224 - 0xe0 -- plane 1
      12'hF39: dout <= 8'b11100000; // 3897 : 224 - 0xe0
      12'hF3A: dout <= 8'b11100000; // 3898 : 224 - 0xe0
      12'hF3B: dout <= 8'b11100000; // 3899 : 224 - 0xe0
      12'hF3C: dout <= 8'b00000000; // 3900 :   0 - 0x0
      12'hF3D: dout <= 8'b00000000; // 3901 :   0 - 0x0
      12'hF3E: dout <= 8'b00000000; // 3902 :   0 - 0x0
      12'hF3F: dout <= 8'b00000000; // 3903 :   0 - 0x0
      12'hF40: dout <= 8'b00000000; // 3904 :   0 - 0x0 -- Sprite 0xf4
      12'hF41: dout <= 8'b11110000; // 3905 : 240 - 0xf0
      12'hF42: dout <= 8'b00000000; // 3906 :   0 - 0x0
      12'hF43: dout <= 8'b00000000; // 3907 :   0 - 0x0
      12'hF44: dout <= 8'b00000000; // 3908 :   0 - 0x0
      12'hF45: dout <= 8'b00000000; // 3909 :   0 - 0x0
      12'hF46: dout <= 8'b00000000; // 3910 :   0 - 0x0
      12'hF47: dout <= 8'b00000000; // 3911 :   0 - 0x0
      12'hF48: dout <= 8'b11110000; // 3912 : 240 - 0xf0 -- plane 1
      12'hF49: dout <= 8'b11110000; // 3913 : 240 - 0xf0
      12'hF4A: dout <= 8'b11110000; // 3914 : 240 - 0xf0
      12'hF4B: dout <= 8'b11110000; // 3915 : 240 - 0xf0
      12'hF4C: dout <= 8'b00000000; // 3916 :   0 - 0x0
      12'hF4D: dout <= 8'b00000000; // 3917 :   0 - 0x0
      12'hF4E: dout <= 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout <= 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout <= 8'b00000000; // 3920 :   0 - 0x0 -- Sprite 0xf5
      12'hF51: dout <= 8'b11111000; // 3921 : 248 - 0xf8
      12'hF52: dout <= 8'b00000000; // 3922 :   0 - 0x0
      12'hF53: dout <= 8'b00000000; // 3923 :   0 - 0x0
      12'hF54: dout <= 8'b00000000; // 3924 :   0 - 0x0
      12'hF55: dout <= 8'b00000000; // 3925 :   0 - 0x0
      12'hF56: dout <= 8'b00000000; // 3926 :   0 - 0x0
      12'hF57: dout <= 8'b00000000; // 3927 :   0 - 0x0
      12'hF58: dout <= 8'b11111000; // 3928 : 248 - 0xf8 -- plane 1
      12'hF59: dout <= 8'b11111000; // 3929 : 248 - 0xf8
      12'hF5A: dout <= 8'b11111000; // 3930 : 248 - 0xf8
      12'hF5B: dout <= 8'b11111000; // 3931 : 248 - 0xf8
      12'hF5C: dout <= 8'b00000000; // 3932 :   0 - 0x0
      12'hF5D: dout <= 8'b00000000; // 3933 :   0 - 0x0
      12'hF5E: dout <= 8'b00000000; // 3934 :   0 - 0x0
      12'hF5F: dout <= 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Sprite 0xf6
      12'hF61: dout <= 8'b11111100; // 3937 : 252 - 0xfc
      12'hF62: dout <= 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout <= 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout <= 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout <= 8'b00000000; // 3941 :   0 - 0x0
      12'hF66: dout <= 8'b00000000; // 3942 :   0 - 0x0
      12'hF67: dout <= 8'b00000000; // 3943 :   0 - 0x0
      12'hF68: dout <= 8'b11111100; // 3944 : 252 - 0xfc -- plane 1
      12'hF69: dout <= 8'b11111100; // 3945 : 252 - 0xfc
      12'hF6A: dout <= 8'b11111100; // 3946 : 252 - 0xfc
      12'hF6B: dout <= 8'b11111100; // 3947 : 252 - 0xfc
      12'hF6C: dout <= 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout <= 8'b00000000; // 3949 :   0 - 0x0
      12'hF6E: dout <= 8'b00000000; // 3950 :   0 - 0x0
      12'hF6F: dout <= 8'b00000000; // 3951 :   0 - 0x0
      12'hF70: dout <= 8'b00000000; // 3952 :   0 - 0x0 -- Sprite 0xf7
      12'hF71: dout <= 8'b11111110; // 3953 : 254 - 0xfe
      12'hF72: dout <= 8'b00000000; // 3954 :   0 - 0x0
      12'hF73: dout <= 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout <= 8'b00000000; // 3956 :   0 - 0x0
      12'hF75: dout <= 8'b00000000; // 3957 :   0 - 0x0
      12'hF76: dout <= 8'b00000000; // 3958 :   0 - 0x0
      12'hF77: dout <= 8'b00000000; // 3959 :   0 - 0x0
      12'hF78: dout <= 8'b11111110; // 3960 : 254 - 0xfe -- plane 1
      12'hF79: dout <= 8'b11111110; // 3961 : 254 - 0xfe
      12'hF7A: dout <= 8'b11111110; // 3962 : 254 - 0xfe
      12'hF7B: dout <= 8'b11111110; // 3963 : 254 - 0xfe
      12'hF7C: dout <= 8'b00000000; // 3964 :   0 - 0x0
      12'hF7D: dout <= 8'b00000000; // 3965 :   0 - 0x0
      12'hF7E: dout <= 8'b00000000; // 3966 :   0 - 0x0
      12'hF7F: dout <= 8'b00000000; // 3967 :   0 - 0x0
      12'hF80: dout <= 8'b00000000; // 3968 :   0 - 0x0 -- Sprite 0xf8
      12'hF81: dout <= 8'b11111111; // 3969 : 255 - 0xff
      12'hF82: dout <= 8'b00000000; // 3970 :   0 - 0x0
      12'hF83: dout <= 8'b00000000; // 3971 :   0 - 0x0
      12'hF84: dout <= 8'b00000000; // 3972 :   0 - 0x0
      12'hF85: dout <= 8'b00000000; // 3973 :   0 - 0x0
      12'hF86: dout <= 8'b00000000; // 3974 :   0 - 0x0
      12'hF87: dout <= 8'b00000000; // 3975 :   0 - 0x0
      12'hF88: dout <= 8'b11111111; // 3976 : 255 - 0xff -- plane 1
      12'hF89: dout <= 8'b11111111; // 3977 : 255 - 0xff
      12'hF8A: dout <= 8'b11111111; // 3978 : 255 - 0xff
      12'hF8B: dout <= 8'b11111111; // 3979 : 255 - 0xff
      12'hF8C: dout <= 8'b00000000; // 3980 :   0 - 0x0
      12'hF8D: dout <= 8'b00000000; // 3981 :   0 - 0x0
      12'hF8E: dout <= 8'b00000000; // 3982 :   0 - 0x0
      12'hF8F: dout <= 8'b00000000; // 3983 :   0 - 0x0
      12'hF90: dout <= 8'b11111111; // 3984 : 255 - 0xff -- Sprite 0xf9
      12'hF91: dout <= 8'b11111111; // 3985 : 255 - 0xff
      12'hF92: dout <= 8'b11111111; // 3986 : 255 - 0xff
      12'hF93: dout <= 8'b11111111; // 3987 : 255 - 0xff
      12'hF94: dout <= 8'b10000000; // 3988 : 128 - 0x80
      12'hF95: dout <= 8'b10000000; // 3989 : 128 - 0x80
      12'hF96: dout <= 8'b11000000; // 3990 : 192 - 0xc0
      12'hF97: dout <= 8'b11000000; // 3991 : 192 - 0xc0
      12'hF98: dout <= 8'b00000000; // 3992 :   0 - 0x0 -- plane 1
      12'hF99: dout <= 8'b00000000; // 3993 :   0 - 0x0
      12'hF9A: dout <= 8'b00000000; // 3994 :   0 - 0x0
      12'hF9B: dout <= 8'b00000000; // 3995 :   0 - 0x0
      12'hF9C: dout <= 8'b01111111; // 3996 : 127 - 0x7f
      12'hF9D: dout <= 8'b01000000; // 3997 :  64 - 0x40
      12'hF9E: dout <= 8'b01000000; // 3998 :  64 - 0x40
      12'hF9F: dout <= 8'b01000000; // 3999 :  64 - 0x40
      12'hFA0: dout <= 8'b11111111; // 4000 : 255 - 0xff -- Sprite 0xfa
      12'hFA1: dout <= 8'b11111111; // 4001 : 255 - 0xff
      12'hFA2: dout <= 8'b11111111; // 4002 : 255 - 0xff
      12'hFA3: dout <= 8'b11111111; // 4003 : 255 - 0xff
      12'hFA4: dout <= 8'b00000000; // 4004 :   0 - 0x0
      12'hFA5: dout <= 8'b00000000; // 4005 :   0 - 0x0
      12'hFA6: dout <= 8'b00000000; // 4006 :   0 - 0x0
      12'hFA7: dout <= 8'b00000000; // 4007 :   0 - 0x0
      12'hFA8: dout <= 8'b00000000; // 4008 :   0 - 0x0 -- plane 1
      12'hFA9: dout <= 8'b00000000; // 4009 :   0 - 0x0
      12'hFAA: dout <= 8'b00000000; // 4010 :   0 - 0x0
      12'hFAB: dout <= 8'b00000000; // 4011 :   0 - 0x0
      12'hFAC: dout <= 8'b11111111; // 4012 : 255 - 0xff
      12'hFAD: dout <= 8'b00000000; // 4013 :   0 - 0x0
      12'hFAE: dout <= 8'b00000000; // 4014 :   0 - 0x0
      12'hFAF: dout <= 8'b00000000; // 4015 :   0 - 0x0
      12'hFB0: dout <= 8'b11111111; // 4016 : 255 - 0xff -- Sprite 0xfb
      12'hFB1: dout <= 8'b11111111; // 4017 : 255 - 0xff
      12'hFB2: dout <= 8'b11111111; // 4018 : 255 - 0xff
      12'hFB3: dout <= 8'b11111111; // 4019 : 255 - 0xff
      12'hFB4: dout <= 8'b00000001; // 4020 :   1 - 0x1
      12'hFB5: dout <= 8'b00000000; // 4021 :   0 - 0x0
      12'hFB6: dout <= 8'b00000010; // 4022 :   2 - 0x2
      12'hFB7: dout <= 8'b00000010; // 4023 :   2 - 0x2
      12'hFB8: dout <= 8'b00000000; // 4024 :   0 - 0x0 -- plane 1
      12'hFB9: dout <= 8'b00000000; // 4025 :   0 - 0x0
      12'hFBA: dout <= 8'b00000000; // 4026 :   0 - 0x0
      12'hFBB: dout <= 8'b00000000; // 4027 :   0 - 0x0
      12'hFBC: dout <= 8'b11111110; // 4028 : 254 - 0xfe
      12'hFBD: dout <= 8'b00000010; // 4029 :   2 - 0x2
      12'hFBE: dout <= 8'b00000010; // 4030 :   2 - 0x2
      12'hFBF: dout <= 8'b00000010; // 4031 :   2 - 0x2
      12'hFC0: dout <= 8'b11000000; // 4032 : 192 - 0xc0 -- Sprite 0xfc
      12'hFC1: dout <= 8'b11000000; // 4033 : 192 - 0xc0
      12'hFC2: dout <= 8'b10000000; // 4034 : 128 - 0x80
      12'hFC3: dout <= 8'b10000000; // 4035 : 128 - 0x80
      12'hFC4: dout <= 8'b11000000; // 4036 : 192 - 0xc0
      12'hFC5: dout <= 8'b11111111; // 4037 : 255 - 0xff
      12'hFC6: dout <= 8'b11111111; // 4038 : 255 - 0xff
      12'hFC7: dout <= 8'b11111111; // 4039 : 255 - 0xff
      12'hFC8: dout <= 8'b01000000; // 4040 :  64 - 0x40 -- plane 1
      12'hFC9: dout <= 8'b01000000; // 4041 :  64 - 0x40
      12'hFCA: dout <= 8'b01000000; // 4042 :  64 - 0x40
      12'hFCB: dout <= 8'b01111111; // 4043 : 127 - 0x7f
      12'hFCC: dout <= 8'b00000000; // 4044 :   0 - 0x0
      12'hFCD: dout <= 8'b00000000; // 4045 :   0 - 0x0
      12'hFCE: dout <= 8'b00000000; // 4046 :   0 - 0x0
      12'hFCF: dout <= 8'b00000000; // 4047 :   0 - 0x0
      12'hFD0: dout <= 8'b00000000; // 4048 :   0 - 0x0 -- Sprite 0xfd
      12'hFD1: dout <= 8'b00000000; // 4049 :   0 - 0x0
      12'hFD2: dout <= 8'b00000000; // 4050 :   0 - 0x0
      12'hFD3: dout <= 8'b00000000; // 4051 :   0 - 0x0
      12'hFD4: dout <= 8'b00000000; // 4052 :   0 - 0x0
      12'hFD5: dout <= 8'b11111111; // 4053 : 255 - 0xff
      12'hFD6: dout <= 8'b11111111; // 4054 : 255 - 0xff
      12'hFD7: dout <= 8'b11111111; // 4055 : 255 - 0xff
      12'hFD8: dout <= 8'b00000000; // 4056 :   0 - 0x0 -- plane 1
      12'hFD9: dout <= 8'b00000000; // 4057 :   0 - 0x0
      12'hFDA: dout <= 8'b00000000; // 4058 :   0 - 0x0
      12'hFDB: dout <= 8'b11111111; // 4059 : 255 - 0xff
      12'hFDC: dout <= 8'b00000000; // 4060 :   0 - 0x0
      12'hFDD: dout <= 8'b00000000; // 4061 :   0 - 0x0
      12'hFDE: dout <= 8'b00000000; // 4062 :   0 - 0x0
      12'hFDF: dout <= 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout <= 8'b00000010; // 4064 :   2 - 0x2 -- Sprite 0xfe
      12'hFE1: dout <= 8'b00000010; // 4065 :   2 - 0x2
      12'hFE2: dout <= 8'b00000000; // 4066 :   0 - 0x0
      12'hFE3: dout <= 8'b00000000; // 4067 :   0 - 0x0
      12'hFE4: dout <= 8'b00000000; // 4068 :   0 - 0x0
      12'hFE5: dout <= 8'b11111111; // 4069 : 255 - 0xff
      12'hFE6: dout <= 8'b11111111; // 4070 : 255 - 0xff
      12'hFE7: dout <= 8'b11111111; // 4071 : 255 - 0xff
      12'hFE8: dout <= 8'b00000010; // 4072 :   2 - 0x2 -- plane 1
      12'hFE9: dout <= 8'b00000010; // 4073 :   2 - 0x2
      12'hFEA: dout <= 8'b00000010; // 4074 :   2 - 0x2
      12'hFEB: dout <= 8'b11111110; // 4075 : 254 - 0xfe
      12'hFEC: dout <= 8'b00000000; // 4076 :   0 - 0x0
      12'hFED: dout <= 8'b00000000; // 4077 :   0 - 0x0
      12'hFEE: dout <= 8'b00000000; // 4078 :   0 - 0x0
      12'hFEF: dout <= 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout <= 8'b11111111; // 4080 : 255 - 0xff -- Sprite 0xff
      12'hFF1: dout <= 8'b11111111; // 4081 : 255 - 0xff
      12'hFF2: dout <= 8'b11111111; // 4082 : 255 - 0xff
      12'hFF3: dout <= 8'b11111111; // 4083 : 255 - 0xff
      12'hFF4: dout <= 8'b11111111; // 4084 : 255 - 0xff
      12'hFF5: dout <= 8'b11111111; // 4085 : 255 - 0xff
      12'hFF6: dout <= 8'b11111111; // 4086 : 255 - 0xff
      12'hFF7: dout <= 8'b11111111; // 4087 : 255 - 0xff
      12'hFF8: dout <= 8'b00000000; // 4088 :   0 - 0x0 -- plane 1
      12'hFF9: dout <= 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout <= 8'b00000000; // 4090 :   0 - 0x0
      12'hFFB: dout <= 8'b00000000; // 4091 :   0 - 0x0
      12'hFFC: dout <= 8'b00000000; // 4092 :   0 - 0x0
      12'hFFD: dout <= 8'b00000000; // 4093 :   0 - 0x0
      12'hFFE: dout <= 8'b00000000; // 4094 :   0 - 0x0
      12'hFFF: dout <= 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
