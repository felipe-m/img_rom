//-   Sprites Pattern table COLOR PLANE 0
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: lawnmower_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_LAWN_SPR_PLN0
  (
     input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table COLOR PLANE 0
      11'h0: dout <= 8'b11111111; //    0 : 255 - 0xff -- Sprite 0x0
      11'h1: dout <= 8'b11111111; //    1 : 255 - 0xff
      11'h2: dout <= 8'b11111111; //    2 : 255 - 0xff
      11'h3: dout <= 8'b11111111; //    3 : 255 - 0xff
      11'h4: dout <= 8'b11111111; //    4 : 255 - 0xff
      11'h5: dout <= 8'b11111111; //    5 : 255 - 0xff
      11'h6: dout <= 8'b11111111; //    6 : 255 - 0xff
      11'h7: dout <= 8'b11111111; //    7 : 255 - 0xff
      11'h8: dout <= 8'b11111111; //    8 : 255 - 0xff -- Sprite 0x1
      11'h9: dout <= 8'b11111111; //    9 : 255 - 0xff
      11'hA: dout <= 8'b11111111; //   10 : 255 - 0xff
      11'hB: dout <= 8'b11111111; //   11 : 255 - 0xff
      11'hC: dout <= 8'b11111111; //   12 : 255 - 0xff
      11'hD: dout <= 8'b11111111; //   13 : 255 - 0xff
      11'hE: dout <= 8'b11111100; //   14 : 252 - 0xfc
      11'hF: dout <= 8'b11111100; //   15 : 252 - 0xfc
      11'h10: dout <= 8'b11111111; //   16 : 255 - 0xff -- Sprite 0x2
      11'h11: dout <= 8'b11111111; //   17 : 255 - 0xff
      11'h12: dout <= 8'b11111111; //   18 : 255 - 0xff
      11'h13: dout <= 8'b11111111; //   19 : 255 - 0xff
      11'h14: dout <= 8'b11111111; //   20 : 255 - 0xff
      11'h15: dout <= 8'b11111111; //   21 : 255 - 0xff
      11'h16: dout <= 8'b00000000; //   22 :   0 - 0x0
      11'h17: dout <= 8'b00000000; //   23 :   0 - 0x0
      11'h18: dout <= 8'b11111111; //   24 : 255 - 0xff -- Sprite 0x3
      11'h19: dout <= 8'b11111111; //   25 : 255 - 0xff
      11'h1A: dout <= 8'b11111111; //   26 : 255 - 0xff
      11'h1B: dout <= 8'b11111111; //   27 : 255 - 0xff
      11'h1C: dout <= 8'b11111111; //   28 : 255 - 0xff
      11'h1D: dout <= 8'b11111111; //   29 : 255 - 0xff
      11'h1E: dout <= 8'b00011111; //   30 :  31 - 0x1f
      11'h1F: dout <= 8'b01000111; //   31 :  71 - 0x47
      11'h20: dout <= 8'b11111111; //   32 : 255 - 0xff -- Sprite 0x4
      11'h21: dout <= 8'b11111111; //   33 : 255 - 0xff
      11'h22: dout <= 8'b11111111; //   34 : 255 - 0xff
      11'h23: dout <= 8'b11111111; //   35 : 255 - 0xff
      11'h24: dout <= 8'b11111111; //   36 : 255 - 0xff
      11'h25: dout <= 8'b11111111; //   37 : 255 - 0xff
      11'h26: dout <= 8'b11100000; //   38 : 224 - 0xe0
      11'h27: dout <= 8'b10000000; //   39 : 128 - 0x80
      11'h28: dout <= 8'b11111111; //   40 : 255 - 0xff -- Sprite 0x5
      11'h29: dout <= 8'b11111111; //   41 : 255 - 0xff
      11'h2A: dout <= 8'b11111111; //   42 : 255 - 0xff
      11'h2B: dout <= 8'b11111111; //   43 : 255 - 0xff
      11'h2C: dout <= 8'b11111111; //   44 : 255 - 0xff
      11'h2D: dout <= 8'b11110111; //   45 : 247 - 0xf7
      11'h2E: dout <= 8'b00000001; //   46 :   1 - 0x1
      11'h2F: dout <= 8'b00000100; //   47 :   4 - 0x4
      11'h30: dout <= 8'b11111111; //   48 : 255 - 0xff -- Sprite 0x6
      11'h31: dout <= 8'b11111111; //   49 : 255 - 0xff
      11'h32: dout <= 8'b11111111; //   50 : 255 - 0xff
      11'h33: dout <= 8'b11111111; //   51 : 255 - 0xff
      11'h34: dout <= 8'b11111111; //   52 : 255 - 0xff
      11'h35: dout <= 8'b11011111; //   53 : 223 - 0xdf
      11'h36: dout <= 8'b00011100; //   54 :  28 - 0x1c
      11'h37: dout <= 8'b01000100; //   55 :  68 - 0x44
      11'h38: dout <= 8'b11111111; //   56 : 255 - 0xff -- Sprite 0x7
      11'h39: dout <= 8'b11111111; //   57 : 255 - 0xff
      11'h3A: dout <= 8'b11111111; //   58 : 255 - 0xff
      11'h3B: dout <= 8'b11111111; //   59 : 255 - 0xff
      11'h3C: dout <= 8'b11111111; //   60 : 255 - 0xff
      11'h3D: dout <= 8'b10111111; //   61 : 191 - 0xbf
      11'h3E: dout <= 8'b00111100; //   62 :  60 - 0x3c
      11'h3F: dout <= 8'b01001100; //   63 :  76 - 0x4c
      11'h40: dout <= 8'b11111100; //   64 : 252 - 0xfc -- Sprite 0x8
      11'h41: dout <= 8'b11111100; //   65 : 252 - 0xfc
      11'h42: dout <= 8'b11111100; //   66 : 252 - 0xfc
      11'h43: dout <= 8'b11111100; //   67 : 252 - 0xfc
      11'h44: dout <= 8'b11111100; //   68 : 252 - 0xfc
      11'h45: dout <= 8'b11111100; //   69 : 252 - 0xfc
      11'h46: dout <= 8'b11111100; //   70 : 252 - 0xfc
      11'h47: dout <= 8'b11111100; //   71 : 252 - 0xfc
      11'h48: dout <= 8'b00010000; //   72 :  16 - 0x10 -- Sprite 0x9
      11'h49: dout <= 8'b00111000; //   73 :  56 - 0x38
      11'h4A: dout <= 8'b01111100; //   74 : 124 - 0x7c
      11'h4B: dout <= 8'b11111000; //   75 : 248 - 0xf8
      11'h4C: dout <= 8'b01110000; //   76 : 112 - 0x70
      11'h4D: dout <= 8'b00100010; //   77 :  34 - 0x22
      11'h4E: dout <= 8'b00000101; //   78 :   5 - 0x5
      11'h4F: dout <= 8'b00000010; //   79 :   2 - 0x2
      11'h50: dout <= 8'b01000111; //   80 :  71 - 0x47 -- Sprite 0xa
      11'h51: dout <= 8'b01000111; //   81 :  71 - 0x47
      11'h52: dout <= 8'b01000111; //   82 :  71 - 0x47
      11'h53: dout <= 8'b01000111; //   83 :  71 - 0x47
      11'h54: dout <= 8'b01000111; //   84 :  71 - 0x47
      11'h55: dout <= 8'b01000111; //   85 :  71 - 0x47
      11'h56: dout <= 8'b01000111; //   86 :  71 - 0x47
      11'h57: dout <= 8'b01000111; //   87 :  71 - 0x47
      11'h58: dout <= 8'b11111111; //   88 : 255 - 0xff -- Sprite 0xb
      11'h59: dout <= 8'b11111110; //   89 : 254 - 0xfe
      11'h5A: dout <= 8'b11111110; //   90 : 254 - 0xfe
      11'h5B: dout <= 8'b11111100; //   91 : 252 - 0xfc
      11'h5C: dout <= 8'b11111100; //   92 : 252 - 0xfc
      11'h5D: dout <= 8'b11111100; //   93 : 252 - 0xfc
      11'h5E: dout <= 8'b11111100; //   94 : 252 - 0xfc
      11'h5F: dout <= 8'b11111100; //   95 : 252 - 0xfc
      11'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0xc
      11'h61: dout <= 8'b00001000; //   97 :   8 - 0x8
      11'h62: dout <= 8'b00011100; //   98 :  28 - 0x1c
      11'h63: dout <= 8'b00111000; //   99 :  56 - 0x38
      11'h64: dout <= 8'b01110000; //  100 : 112 - 0x70
      11'h65: dout <= 8'b00100010; //  101 :  34 - 0x22
      11'h66: dout <= 8'b00000101; //  102 :   5 - 0x5
      11'h67: dout <= 8'b00000010; //  103 :   2 - 0x2
      11'h68: dout <= 8'b00000010; //  104 :   2 - 0x2 -- Sprite 0xd
      11'h69: dout <= 8'b00110001; //  105 :  49 - 0x31
      11'h6A: dout <= 8'b01111000; //  106 : 120 - 0x78
      11'h6B: dout <= 8'b11111000; //  107 : 248 - 0xf8
      11'h6C: dout <= 8'b01110000; //  108 : 112 - 0x70
      11'h6D: dout <= 8'b00100010; //  109 :  34 - 0x22
      11'h6E: dout <= 8'b00000101; //  110 :   5 - 0x5
      11'h6F: dout <= 8'b00000010; //  111 :   2 - 0x2
      11'h70: dout <= 8'b01111100; //  112 : 124 - 0x7c -- Sprite 0xe
      11'h71: dout <= 8'b00111100; //  113 :  60 - 0x3c
      11'h72: dout <= 8'b10011100; //  114 : 156 - 0x9c
      11'h73: dout <= 8'b10001100; //  115 : 140 - 0x8c
      11'h74: dout <= 8'b01001100; //  116 :  76 - 0x4c
      11'h75: dout <= 8'b01000100; //  117 :  68 - 0x44
      11'h76: dout <= 8'b01000100; //  118 :  68 - 0x44
      11'h77: dout <= 8'b01000100; //  119 :  68 - 0x44
      11'h78: dout <= 8'b01000100; //  120 :  68 - 0x44 -- Sprite 0xf
      11'h79: dout <= 8'b01000100; //  121 :  68 - 0x44
      11'h7A: dout <= 8'b01000100; //  122 :  68 - 0x44
      11'h7B: dout <= 8'b01000100; //  123 :  68 - 0x44
      11'h7C: dout <= 8'b01000100; //  124 :  68 - 0x44
      11'h7D: dout <= 8'b01000100; //  125 :  68 - 0x44
      11'h7E: dout <= 8'b01000100; //  126 :  68 - 0x44
      11'h7F: dout <= 8'b01000100; //  127 :  68 - 0x44
      11'h80: dout <= 8'b01001100; //  128 :  76 - 0x4c -- Sprite 0x10
      11'h81: dout <= 8'b00100100; //  129 :  36 - 0x24
      11'h82: dout <= 8'b00100100; //  130 :  36 - 0x24
      11'h83: dout <= 8'b10010100; //  131 : 148 - 0x94
      11'h84: dout <= 8'b00010000; //  132 :  16 - 0x10
      11'h85: dout <= 8'b00001000; //  133 :   8 - 0x8
      11'h86: dout <= 8'b00001000; //  134 :   8 - 0x8
      11'h87: dout <= 8'b00000100; //  135 :   4 - 0x4
      11'h88: dout <= 8'b00000000; //  136 :   0 - 0x0 -- Sprite 0x11
      11'h89: dout <= 8'b00111100; //  137 :  60 - 0x3c
      11'h8A: dout <= 8'b01000000; //  138 :  64 - 0x40
      11'h8B: dout <= 8'b01000100; //  139 :  68 - 0x44
      11'h8C: dout <= 8'b01000100; //  140 :  68 - 0x44
      11'h8D: dout <= 8'b01000100; //  141 :  68 - 0x44
      11'h8E: dout <= 8'b01000100; //  142 :  68 - 0x44
      11'h8F: dout <= 8'b01000100; //  143 :  68 - 0x44
      11'h90: dout <= 8'b00000100; //  144 :   4 - 0x4 -- Sprite 0x12
      11'h91: dout <= 8'b00010010; //  145 :  18 - 0x12
      11'h92: dout <= 8'b00110010; //  146 :  50 - 0x32
      11'h93: dout <= 8'b01111000; //  147 : 120 - 0x78
      11'h94: dout <= 8'b11111000; //  148 : 248 - 0xf8
      11'h95: dout <= 8'b01110000; //  149 : 112 - 0x70
      11'h96: dout <= 8'b00100100; //  150 :  36 - 0x24
      11'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      11'h98: dout <= 8'b01000100; //  152 :  68 - 0x44 -- Sprite 0x13
      11'h99: dout <= 8'b01000100; //  153 :  68 - 0x44
      11'h9A: dout <= 8'b01000100; //  154 :  68 - 0x44
      11'h9B: dout <= 8'b01000100; //  155 :  68 - 0x44
      11'h9C: dout <= 8'b01000100; //  156 :  68 - 0x44
      11'h9D: dout <= 8'b01000100; //  157 :  68 - 0x44
      11'h9E: dout <= 8'b01000100; //  158 :  68 - 0x44
      11'h9F: dout <= 8'b01011100; //  159 :  92 - 0x5c
      11'hA0: dout <= 8'b00010000; //  160 :  16 - 0x10 -- Sprite 0x14
      11'hA1: dout <= 8'b00111000; //  161 :  56 - 0x38
      11'hA2: dout <= 8'b00111100; //  162 :  60 - 0x3c
      11'hA3: dout <= 8'b00111000; //  163 :  56 - 0x38
      11'hA4: dout <= 8'b00010000; //  164 :  16 - 0x10
      11'hA5: dout <= 8'b00000010; //  165 :   2 - 0x2
      11'hA6: dout <= 8'b01000101; //  166 :  69 - 0x45
      11'hA7: dout <= 8'b01000010; //  167 :  66 - 0x42
      11'hA8: dout <= 8'b01000100; //  168 :  68 - 0x44 -- Sprite 0x15
      11'hA9: dout <= 8'b01000100; //  169 :  68 - 0x44
      11'hAA: dout <= 8'b01000100; //  170 :  68 - 0x44
      11'hAB: dout <= 8'b01000100; //  171 :  68 - 0x44
      11'hAC: dout <= 8'b01000100; //  172 :  68 - 0x44
      11'hAD: dout <= 8'b01011100; //  173 :  92 - 0x5c
      11'hAE: dout <= 8'b01000000; //  174 :  64 - 0x40
      11'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      11'hB0: dout <= 8'b01000000; //  176 :  64 - 0x40 -- Sprite 0x16
      11'hB1: dout <= 8'b01000000; //  177 :  64 - 0x40
      11'hB2: dout <= 8'b00000000; //  178 :   0 - 0x0
      11'hB3: dout <= 8'b00000000; //  179 :   0 - 0x0
      11'hB4: dout <= 8'b00011000; //  180 :  24 - 0x18
      11'hB5: dout <= 8'b00111000; //  181 :  56 - 0x38
      11'hB6: dout <= 8'b00010000; //  182 :  16 - 0x10
      11'hB7: dout <= 8'b00000000; //  183 :   0 - 0x0
      11'hB8: dout <= 8'b01000000; //  184 :  64 - 0x40 -- Sprite 0x17
      11'hB9: dout <= 8'b01000000; //  185 :  64 - 0x40
      11'hBA: dout <= 8'b01000000; //  186 :  64 - 0x40
      11'hBB: dout <= 8'b01000000; //  187 :  64 - 0x40
      11'hBC: dout <= 8'b01010000; //  188 :  80 - 0x50
      11'hBD: dout <= 8'b01010000; //  189 :  80 - 0x50
      11'hBE: dout <= 8'b01001000; //  190 :  72 - 0x48
      11'hBF: dout <= 8'b01001000; //  191 :  72 - 0x48
      11'hC0: dout <= 8'b01000111; //  192 :  71 - 0x47 -- Sprite 0x18
      11'hC1: dout <= 8'b01000111; //  193 :  71 - 0x47
      11'hC2: dout <= 8'b01000111; //  194 :  71 - 0x47
      11'hC3: dout <= 8'b01000111; //  195 :  71 - 0x47
      11'hC4: dout <= 8'b01000111; //  196 :  71 - 0x47
      11'hC5: dout <= 8'b01011111; //  197 :  95 - 0x5f
      11'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      11'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      11'hC8: dout <= 8'b11111100; //  200 : 252 - 0xfc -- Sprite 0x19
      11'hC9: dout <= 8'b11111100; //  201 : 252 - 0xfc
      11'hCA: dout <= 8'b11111100; //  202 : 252 - 0xfc
      11'hCB: dout <= 8'b11111100; //  203 : 252 - 0xfc
      11'hCC: dout <= 8'b11111100; //  204 : 252 - 0xfc
      11'hCD: dout <= 8'b11011100; //  205 : 220 - 0xdc
      11'hCE: dout <= 8'b00011100; //  206 :  28 - 0x1c
      11'hCF: dout <= 8'b01000100; //  207 :  68 - 0x44
      11'hD0: dout <= 8'b00010000; //  208 :  16 - 0x10 -- Sprite 0x1a
      11'hD1: dout <= 8'b00111000; //  209 :  56 - 0x38
      11'hD2: dout <= 8'b01111100; //  210 : 124 - 0x7c
      11'hD3: dout <= 8'b11100000; //  211 : 224 - 0xe0
      11'hD4: dout <= 8'b01000000; //  212 :  64 - 0x40
      11'hD5: dout <= 8'b00000000; //  213 :   0 - 0x0
      11'hD6: dout <= 8'b00010000; //  214 :  16 - 0x10
      11'hD7: dout <= 8'b00100000; //  215 :  32 - 0x20
      11'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x1b
      11'hD9: dout <= 8'b01111100; //  217 : 124 - 0x7c
      11'hDA: dout <= 8'b01000000; //  218 :  64 - 0x40
      11'hDB: dout <= 8'b01000100; //  219 :  68 - 0x44
      11'hDC: dout <= 8'b01000100; //  220 :  68 - 0x44
      11'hDD: dout <= 8'b01000100; //  221 :  68 - 0x44
      11'hDE: dout <= 8'b01000100; //  222 :  68 - 0x44
      11'hDF: dout <= 8'b01000100; //  223 :  68 - 0x44
      11'hE0: dout <= 8'b00010000; //  224 :  16 - 0x10 -- Sprite 0x1c
      11'hE1: dout <= 8'b00111000; //  225 :  56 - 0x38
      11'hE2: dout <= 8'b01110001; //  226 : 113 - 0x71
      11'hE3: dout <= 8'b11100010; //  227 : 226 - 0xe2
      11'hE4: dout <= 8'b01000100; //  228 :  68 - 0x44
      11'hE5: dout <= 8'b00001000; //  229 :   8 - 0x8
      11'hE6: dout <= 8'b00010000; //  230 :  16 - 0x10
      11'hE7: dout <= 8'b00100000; //  231 :  32 - 0x20
      11'hE8: dout <= 8'b01000000; //  232 :  64 - 0x40 -- Sprite 0x1d
      11'hE9: dout <= 8'b10000100; //  233 : 132 - 0x84
      11'hEA: dout <= 8'b00000010; //  234 :   2 - 0x2
      11'hEB: dout <= 8'b00000111; //  235 :   7 - 0x7
      11'hEC: dout <= 8'b00001111; //  236 :  15 - 0xf
      11'hED: dout <= 8'b00011111; //  237 :  31 - 0x1f
      11'hEE: dout <= 8'b00111111; //  238 :  63 - 0x3f
      11'hEF: dout <= 8'b01111111; //  239 : 127 - 0x7f
      11'hF0: dout <= 8'b00010000; //  240 :  16 - 0x10 -- Sprite 0x1e
      11'hF1: dout <= 8'b00011000; //  241 :  24 - 0x18
      11'hF2: dout <= 8'b00001100; //  242 :  12 - 0xc
      11'hF3: dout <= 8'b00000110; //  243 :   6 - 0x6
      11'hF4: dout <= 8'b10000000; //  244 : 128 - 0x80
      11'hF5: dout <= 8'b11000000; //  245 : 192 - 0xc0
      11'hF6: dout <= 8'b11100000; //  246 : 224 - 0xe0
      11'hF7: dout <= 8'b11110000; //  247 : 240 - 0xf0
      11'hF8: dout <= 8'b11111100; //  248 : 252 - 0xfc -- Sprite 0x1f
      11'hF9: dout <= 8'b11111101; //  249 : 253 - 0xfd
      11'hFA: dout <= 8'b11111100; //  250 : 252 - 0xfc
      11'hFB: dout <= 8'b11111110; //  251 : 254 - 0xfe
      11'hFC: dout <= 8'b11111110; //  252 : 254 - 0xfe
      11'hFD: dout <= 8'b11111111; //  253 : 255 - 0xff
      11'hFE: dout <= 8'b11111111; //  254 : 255 - 0xff
      11'hFF: dout <= 8'b11111111; //  255 : 255 - 0xff
      11'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      11'h101: dout <= 8'b11111111; //  257 : 255 - 0xff
      11'h102: dout <= 8'b00000000; //  258 :   0 - 0x0
      11'h103: dout <= 8'b00000000; //  259 :   0 - 0x0
      11'h104: dout <= 8'b00000000; //  260 :   0 - 0x0
      11'h105: dout <= 8'b11111111; //  261 : 255 - 0xff
      11'h106: dout <= 8'b11111111; //  262 : 255 - 0xff
      11'h107: dout <= 8'b11111111; //  263 : 255 - 0xff
      11'h108: dout <= 8'b01000100; //  264 :  68 - 0x44 -- Sprite 0x21
      11'h109: dout <= 8'b11000101; //  265 : 197 - 0xc5
      11'h10A: dout <= 8'b00000000; //  266 :   0 - 0x0
      11'h10B: dout <= 8'b00000110; //  267 :   6 - 0x6
      11'h10C: dout <= 8'b00000110; //  268 :   6 - 0x6
      11'h10D: dout <= 8'b11111111; //  269 : 255 - 0xff
      11'h10E: dout <= 8'b11111111; //  270 : 255 - 0xff
      11'h10F: dout <= 8'b11111111; //  271 : 255 - 0xff
      11'h110: dout <= 8'b01000000; //  272 :  64 - 0x40 -- Sprite 0x22
      11'h111: dout <= 8'b10000001; //  273 : 129 - 0x81
      11'h112: dout <= 8'b00000011; //  274 :   3 - 0x3
      11'h113: dout <= 8'b00000111; //  275 :   7 - 0x7
      11'h114: dout <= 8'b00001111; //  276 :  15 - 0xf
      11'h115: dout <= 8'b11111111; //  277 : 255 - 0xff
      11'h116: dout <= 8'b11111111; //  278 : 255 - 0xff
      11'h117: dout <= 8'b11111111; //  279 : 255 - 0xff
      11'h118: dout <= 8'b11111000; //  280 : 248 - 0xf8 -- Sprite 0x23
      11'h119: dout <= 8'b11111100; //  281 : 252 - 0xfc
      11'h11A: dout <= 8'b11111110; //  282 : 254 - 0xfe
      11'h11B: dout <= 8'b11111110; //  283 : 254 - 0xfe
      11'h11C: dout <= 8'b11111111; //  284 : 255 - 0xff
      11'h11D: dout <= 8'b11111111; //  285 : 255 - 0xff
      11'h11E: dout <= 8'b11111111; //  286 : 255 - 0xff
      11'h11F: dout <= 8'b11111111; //  287 : 255 - 0xff
      11'h120: dout <= 8'b01000111; //  288 :  71 - 0x47 -- Sprite 0x24
      11'h121: dout <= 8'b11000111; //  289 : 199 - 0xc7
      11'h122: dout <= 8'b00000111; //  290 :   7 - 0x7
      11'h123: dout <= 8'b00000111; //  291 :   7 - 0x7
      11'h124: dout <= 8'b00000111; //  292 :   7 - 0x7
      11'h125: dout <= 8'b11111111; //  293 : 255 - 0xff
      11'h126: dout <= 8'b11111111; //  294 : 255 - 0xff
      11'h127: dout <= 8'b11111111; //  295 : 255 - 0xff
      11'h128: dout <= 8'b11111111; //  296 : 255 - 0xff -- Sprite 0x25
      11'h129: dout <= 8'b11111111; //  297 : 255 - 0xff
      11'h12A: dout <= 8'b11111111; //  298 : 255 - 0xff
      11'h12B: dout <= 8'b11111111; //  299 : 255 - 0xff
      11'h12C: dout <= 8'b11111111; //  300 : 255 - 0xff
      11'h12D: dout <= 8'b11111111; //  301 : 255 - 0xff
      11'h12E: dout <= 8'b00011111; //  302 :  31 - 0x1f
      11'h12F: dout <= 8'b00001111; //  303 :  15 - 0xf
      11'h130: dout <= 8'b11111111; //  304 : 255 - 0xff -- Sprite 0x26
      11'h131: dout <= 8'b11111111; //  305 : 255 - 0xff
      11'h132: dout <= 8'b11111111; //  306 : 255 - 0xff
      11'h133: dout <= 8'b11111111; //  307 : 255 - 0xff
      11'h134: dout <= 8'b11111111; //  308 : 255 - 0xff
      11'h135: dout <= 8'b11111111; //  309 : 255 - 0xff
      11'h136: dout <= 8'b11111100; //  310 : 252 - 0xfc
      11'h137: dout <= 8'b11111000; //  311 : 248 - 0xf8
      11'h138: dout <= 8'b00100111; //  312 :  39 - 0x27 -- Sprite 0x27
      11'h139: dout <= 8'b00010011; //  313 :  19 - 0x13
      11'h13A: dout <= 8'b00001001; //  314 :   9 - 0x9
      11'h13B: dout <= 8'b11000100; //  315 : 196 - 0xc4
      11'h13C: dout <= 8'b01100010; //  316 :  98 - 0x62
      11'h13D: dout <= 8'b00100001; //  317 :  33 - 0x21
      11'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      11'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      11'h140: dout <= 8'b11111111; //  320 : 255 - 0xff -- Sprite 0x28
      11'h141: dout <= 8'b11111111; //  321 : 255 - 0xff
      11'h142: dout <= 8'b11111111; //  322 : 255 - 0xff
      11'h143: dout <= 8'b11111111; //  323 : 255 - 0xff
      11'h144: dout <= 8'b01111111; //  324 : 127 - 0x7f
      11'h145: dout <= 8'b00111110; //  325 :  62 - 0x3e
      11'h146: dout <= 8'b10011100; //  326 : 156 - 0x9c
      11'h147: dout <= 8'b01001000; //  327 :  72 - 0x48
      11'h148: dout <= 8'b11110000; //  328 : 240 - 0xf0 -- Sprite 0x29
      11'h149: dout <= 8'b11100000; //  329 : 224 - 0xe0
      11'h14A: dout <= 8'b11000000; //  330 : 192 - 0xc0
      11'h14B: dout <= 8'b10000000; //  331 : 128 - 0x80
      11'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      11'h14D: dout <= 8'b00000010; //  333 :   2 - 0x2
      11'h14E: dout <= 8'b00000101; //  334 :   5 - 0x5
      11'h14F: dout <= 8'b00000010; //  335 :   2 - 0x2
      11'h150: dout <= 8'b01000111; //  336 :  71 - 0x47 -- Sprite 0x2a
      11'h151: dout <= 8'b01000110; //  337 :  70 - 0x46
      11'h152: dout <= 8'b01000110; //  338 :  70 - 0x46
      11'h153: dout <= 8'b01000100; //  339 :  68 - 0x44
      11'h154: dout <= 8'b01000100; //  340 :  68 - 0x44
      11'h155: dout <= 8'b01000100; //  341 :  68 - 0x44
      11'h156: dout <= 8'b01000100; //  342 :  68 - 0x44
      11'h157: dout <= 8'b01000100; //  343 :  68 - 0x44
      11'h158: dout <= 8'b01111111; //  344 : 127 - 0x7f -- Sprite 0x2b
      11'h159: dout <= 8'b00111111; //  345 :  63 - 0x3f
      11'h15A: dout <= 8'b10011111; //  346 : 159 - 0x9f
      11'h15B: dout <= 8'b10001111; //  347 : 143 - 0x8f
      11'h15C: dout <= 8'b01001111; //  348 :  79 - 0x4f
      11'h15D: dout <= 8'b01000111; //  349 :  71 - 0x47
      11'h15E: dout <= 8'b01000111; //  350 :  71 - 0x47
      11'h15F: dout <= 8'b01000111; //  351 :  71 - 0x47
      11'h160: dout <= 8'b00100000; //  352 :  32 - 0x20 -- Sprite 0x2c
      11'h161: dout <= 8'b00010000; //  353 :  16 - 0x10
      11'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      11'h163: dout <= 8'b11000000; //  355 : 192 - 0xc0
      11'h164: dout <= 8'b01100000; //  356 :  96 - 0x60
      11'h165: dout <= 8'b00100010; //  357 :  34 - 0x22
      11'h166: dout <= 8'b00000101; //  358 :   5 - 0x5
      11'h167: dout <= 8'b00000010; //  359 :   2 - 0x2
      11'h168: dout <= 8'b00000000; //  360 :   0 - 0x0 -- Sprite 0x2d
      11'h169: dout <= 8'b01111111; //  361 : 127 - 0x7f
      11'h16A: dout <= 8'b01000000; //  362 :  64 - 0x40
      11'h16B: dout <= 8'b01000000; //  363 :  64 - 0x40
      11'h16C: dout <= 8'b01000000; //  364 :  64 - 0x40
      11'h16D: dout <= 8'b01000111; //  365 :  71 - 0x47
      11'h16E: dout <= 8'b01000111; //  366 :  71 - 0x47
      11'h16F: dout <= 8'b01000111; //  367 :  71 - 0x47
      11'h170: dout <= 8'b01000100; //  368 :  68 - 0x44 -- Sprite 0x2e
      11'h171: dout <= 8'b11000100; //  369 : 196 - 0xc4
      11'h172: dout <= 8'b00000100; //  370 :   4 - 0x4
      11'h173: dout <= 8'b00000100; //  371 :   4 - 0x4
      11'h174: dout <= 8'b00000100; //  372 :   4 - 0x4
      11'h175: dout <= 8'b11111100; //  373 : 252 - 0xfc
      11'h176: dout <= 8'b11111100; //  374 : 252 - 0xfc
      11'h177: dout <= 8'b11111100; //  375 : 252 - 0xfc
      11'h178: dout <= 8'b00000001; //  376 :   1 - 0x1 -- Sprite 0x2f
      11'h179: dout <= 8'b01111100; //  377 : 124 - 0x7c
      11'h17A: dout <= 8'b01000000; //  378 :  64 - 0x40
      11'h17B: dout <= 8'b01000100; //  379 :  68 - 0x44
      11'h17C: dout <= 8'b01000100; //  380 :  68 - 0x44
      11'h17D: dout <= 8'b01000100; //  381 :  68 - 0x44
      11'h17E: dout <= 8'b01000100; //  382 :  68 - 0x44
      11'h17F: dout <= 8'b01000100; //  383 :  68 - 0x44
      11'h180: dout <= 8'b00010000; //  384 :  16 - 0x10 -- Sprite 0x30
      11'h181: dout <= 8'b00111000; //  385 :  56 - 0x38
      11'h182: dout <= 8'b00111100; //  386 :  60 - 0x3c
      11'h183: dout <= 8'b00011000; //  387 :  24 - 0x18
      11'h184: dout <= 8'b00000000; //  388 :   0 - 0x0
      11'h185: dout <= 8'b01000010; //  389 :  66 - 0x42
      11'h186: dout <= 8'b01000100; //  390 :  68 - 0x44
      11'h187: dout <= 8'b01001000; //  391 :  72 - 0x48
      11'h188: dout <= 8'b01000111; //  392 :  71 - 0x47 -- Sprite 0x31
      11'h189: dout <= 8'b01011111; //  393 :  95 - 0x5f
      11'h18A: dout <= 8'b00000000; //  394 :   0 - 0x0
      11'h18B: dout <= 8'b00000000; //  395 :   0 - 0x0
      11'h18C: dout <= 8'b01110000; //  396 : 112 - 0x70
      11'h18D: dout <= 8'b00100010; //  397 :  34 - 0x22
      11'h18E: dout <= 8'b00000101; //  398 :   5 - 0x5
      11'h18F: dout <= 8'b00000010; //  399 :   2 - 0x2
      11'h190: dout <= 8'b11111111; //  400 : 255 - 0xff -- Sprite 0x32
      11'h191: dout <= 8'b11111111; //  401 : 255 - 0xff
      11'h192: dout <= 8'b00000000; //  402 :   0 - 0x0
      11'h193: dout <= 8'b00000000; //  403 :   0 - 0x0
      11'h194: dout <= 8'b01110000; //  404 : 112 - 0x70
      11'h195: dout <= 8'b00100010; //  405 :  34 - 0x22
      11'h196: dout <= 8'b00000101; //  406 :   5 - 0x5
      11'h197: dout <= 8'b00000010; //  407 :   2 - 0x2
      11'h198: dout <= 8'b11111111; //  408 : 255 - 0xff -- Sprite 0x33
      11'h199: dout <= 8'b11011111; //  409 : 223 - 0xdf
      11'h19A: dout <= 8'b00011111; //  410 :  31 - 0x1f
      11'h19B: dout <= 8'b01000111; //  411 :  71 - 0x47
      11'h19C: dout <= 8'b01000111; //  412 :  71 - 0x47
      11'h19D: dout <= 8'b01000111; //  413 :  71 - 0x47
      11'h19E: dout <= 8'b01000111; //  414 :  71 - 0x47
      11'h19F: dout <= 8'b01000111; //  415 :  71 - 0x47
      11'h1A0: dout <= 8'b01000100; //  416 :  68 - 0x44 -- Sprite 0x34
      11'h1A1: dout <= 8'b01000100; //  417 :  68 - 0x44
      11'h1A2: dout <= 8'b01000100; //  418 :  68 - 0x44
      11'h1A3: dout <= 8'b01000100; //  419 :  68 - 0x44
      11'h1A4: dout <= 8'b01000100; //  420 :  68 - 0x44
      11'h1A5: dout <= 8'b01000100; //  421 :  68 - 0x44
      11'h1A6: dout <= 8'b01000100; //  422 :  68 - 0x44
      11'h1A7: dout <= 8'b01000100; //  423 :  68 - 0x44
      11'h1A8: dout <= 8'b00010000; //  424 :  16 - 0x10 -- Sprite 0x35
      11'h1A9: dout <= 8'b00111000; //  425 :  56 - 0x38
      11'h1AA: dout <= 8'b01111100; //  426 : 124 - 0x7c
      11'h1AB: dout <= 8'b11111000; //  427 : 248 - 0xf8
      11'h1AC: dout <= 8'b00000000; //  428 :   0 - 0x0
      11'h1AD: dout <= 8'b01111111; //  429 : 127 - 0x7f
      11'h1AE: dout <= 8'b01000000; //  430 :  64 - 0x40
      11'h1AF: dout <= 8'b01000000; //  431 :  64 - 0x40
      11'h1B0: dout <= 8'b00010000; //  432 :  16 - 0x10 -- Sprite 0x36
      11'h1B1: dout <= 8'b00111000; //  433 :  56 - 0x38
      11'h1B2: dout <= 8'b01111100; //  434 : 124 - 0x7c
      11'h1B3: dout <= 8'b11111000; //  435 : 248 - 0xf8
      11'h1B4: dout <= 8'b00000000; //  436 :   0 - 0x0
      11'h1B5: dout <= 8'b11111111; //  437 : 255 - 0xff
      11'h1B6: dout <= 8'b00000000; //  438 :   0 - 0x0
      11'h1B7: dout <= 8'b00000000; //  439 :   0 - 0x0
      11'h1B8: dout <= 8'b01000111; //  440 :  71 - 0x47 -- Sprite 0x37
      11'h1B9: dout <= 8'b01000111; //  441 :  71 - 0x47
      11'h1BA: dout <= 8'b01000111; //  442 :  71 - 0x47
      11'h1BB: dout <= 8'b01000111; //  443 :  71 - 0x47
      11'h1BC: dout <= 8'b01000111; //  444 :  71 - 0x47
      11'h1BD: dout <= 8'b11000111; //  445 : 199 - 0xc7
      11'h1BE: dout <= 8'b00000111; //  446 :   7 - 0x7
      11'h1BF: dout <= 8'b00000111; //  447 :   7 - 0x7
      11'h1C0: dout <= 8'b01000100; //  448 :  68 - 0x44 -- Sprite 0x38
      11'h1C1: dout <= 8'b01000100; //  449 :  68 - 0x44
      11'h1C2: dout <= 8'b01000100; //  450 :  68 - 0x44
      11'h1C3: dout <= 8'b01000100; //  451 :  68 - 0x44
      11'h1C4: dout <= 8'b01000100; //  452 :  68 - 0x44
      11'h1C5: dout <= 8'b01011000; //  453 :  88 - 0x58
      11'h1C6: dout <= 8'b00000000; //  454 :   0 - 0x0
      11'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      11'h1C8: dout <= 8'b00010000; //  456 :  16 - 0x10 -- Sprite 0x39
      11'h1C9: dout <= 8'b00111000; //  457 :  56 - 0x38
      11'h1CA: dout <= 8'b01111100; //  458 : 124 - 0x7c
      11'h1CB: dout <= 8'b11111000; //  459 : 248 - 0xf8
      11'h1CC: dout <= 8'b01110000; //  460 : 112 - 0x70
      11'h1CD: dout <= 8'b00100010; //  461 :  34 - 0x22
      11'h1CE: dout <= 8'b00000100; //  462 :   4 - 0x4
      11'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout <= 8'b01000100; //  464 :  68 - 0x44 -- Sprite 0x3a
      11'h1D1: dout <= 8'b01000100; //  465 :  68 - 0x44
      11'h1D2: dout <= 8'b01000100; //  466 :  68 - 0x44
      11'h1D3: dout <= 8'b01000100; //  467 :  68 - 0x44
      11'h1D4: dout <= 8'b01000100; //  468 :  68 - 0x44
      11'h1D5: dout <= 8'b01011000; //  469 :  88 - 0x58
      11'h1D6: dout <= 8'b00000000; //  470 :   0 - 0x0
      11'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      11'h1D8: dout <= 8'b01000000; //  472 :  64 - 0x40 -- Sprite 0x3b
      11'h1D9: dout <= 8'b01000111; //  473 :  71 - 0x47
      11'h1DA: dout <= 8'b01000111; //  474 :  71 - 0x47
      11'h1DB: dout <= 8'b01000111; //  475 :  71 - 0x47
      11'h1DC: dout <= 8'b01000111; //  476 :  71 - 0x47
      11'h1DD: dout <= 8'b01011111; //  477 :  95 - 0x5f
      11'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      11'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      11'h1E1: dout <= 8'b11111111; //  481 : 255 - 0xff
      11'h1E2: dout <= 8'b11111111; //  482 : 255 - 0xff
      11'h1E3: dout <= 8'b11111111; //  483 : 255 - 0xff
      11'h1E4: dout <= 8'b11111111; //  484 : 255 - 0xff
      11'h1E5: dout <= 8'b11111111; //  485 : 255 - 0xff
      11'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      11'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout <= 8'b00000111; //  488 :   7 - 0x7 -- Sprite 0x3d
      11'h1E9: dout <= 8'b11111111; //  489 : 255 - 0xff
      11'h1EA: dout <= 8'b11111111; //  490 : 255 - 0xff
      11'h1EB: dout <= 8'b11111111; //  491 : 255 - 0xff
      11'h1EC: dout <= 8'b11111111; //  492 : 255 - 0xff
      11'h1ED: dout <= 8'b11111111; //  493 : 255 - 0xff
      11'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      11'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      11'h1F0: dout <= 8'b00010000; //  496 :  16 - 0x10 -- Sprite 0x3e
      11'h1F1: dout <= 8'b00111000; //  497 :  56 - 0x38
      11'h1F2: dout <= 8'b01110001; //  498 : 113 - 0x71
      11'h1F3: dout <= 8'b11100010; //  499 : 226 - 0xe2
      11'h1F4: dout <= 8'b01100010; //  500 :  98 - 0x62
      11'h1F5: dout <= 8'b00100001; //  501 :  33 - 0x21
      11'h1F6: dout <= 8'b00000000; //  502 :   0 - 0x0
      11'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      11'h1F8: dout <= 8'b10000111; //  504 : 135 - 0x87 -- Sprite 0x3f
      11'h1F9: dout <= 8'b10000111; //  505 : 135 - 0x87
      11'h1FA: dout <= 8'b00000111; //  506 :   7 - 0x7
      11'h1FB: dout <= 8'b00001111; //  507 :  15 - 0xf
      11'h1FC: dout <= 8'b00001111; //  508 :  15 - 0xf
      11'h1FD: dout <= 8'b00011111; //  509 :  31 - 0x1f
      11'h1FE: dout <= 8'b10011111; //  510 : 159 - 0x9f
      11'h1FF: dout <= 8'b10001111; //  511 : 143 - 0x8f
      11'h200: dout <= 8'b01000100; //  512 :  68 - 0x44 -- Sprite 0x40
      11'h201: dout <= 8'b01000100; //  513 :  68 - 0x44
      11'h202: dout <= 8'b01000100; //  514 :  68 - 0x44
      11'h203: dout <= 8'b01000100; //  515 :  68 - 0x44
      11'h204: dout <= 8'b01000100; //  516 :  68 - 0x44
      11'h205: dout <= 8'b01000110; //  517 :  70 - 0x46
      11'h206: dout <= 8'b01000110; //  518 :  70 - 0x46
      11'h207: dout <= 8'b01000111; //  519 :  71 - 0x47
      11'h208: dout <= 8'b00010000; //  520 :  16 - 0x10 -- Sprite 0x41
      11'h209: dout <= 8'b00111000; //  521 :  56 - 0x38
      11'h20A: dout <= 8'b01111100; //  522 : 124 - 0x7c
      11'h20B: dout <= 8'b01111000; //  523 : 120 - 0x78
      11'h20C: dout <= 8'b00110000; //  524 :  48 - 0x30
      11'h20D: dout <= 8'b00000010; //  525 :   2 - 0x2
      11'h20E: dout <= 8'b00000101; //  526 :   5 - 0x5
      11'h20F: dout <= 8'b00000010; //  527 :   2 - 0x2
      11'h210: dout <= 8'b00010000; //  528 :  16 - 0x10 -- Sprite 0x42
      11'h211: dout <= 8'b00111000; //  529 :  56 - 0x38
      11'h212: dout <= 8'b01111100; //  530 : 124 - 0x7c
      11'h213: dout <= 8'b11111000; //  531 : 248 - 0xf8
      11'h214: dout <= 8'b01110000; //  532 : 112 - 0x70
      11'h215: dout <= 8'b00100000; //  533 :  32 - 0x20
      11'h216: dout <= 8'b00000001; //  534 :   1 - 0x1
      11'h217: dout <= 8'b00000010; //  535 :   2 - 0x2
      11'h218: dout <= 8'b01000100; //  536 :  68 - 0x44 -- Sprite 0x43
      11'h219: dout <= 8'b01000100; //  537 :  68 - 0x44
      11'h21A: dout <= 8'b01000100; //  538 :  68 - 0x44
      11'h21B: dout <= 8'b01000100; //  539 :  68 - 0x44
      11'h21C: dout <= 8'b10000100; //  540 : 132 - 0x84
      11'h21D: dout <= 8'b10000100; //  541 : 132 - 0x84
      11'h21E: dout <= 8'b00000100; //  542 :   4 - 0x4
      11'h21F: dout <= 8'b00001100; //  543 :  12 - 0xc
      11'h220: dout <= 8'b00010000; //  544 :  16 - 0x10 -- Sprite 0x44
      11'h221: dout <= 8'b00111000; //  545 :  56 - 0x38
      11'h222: dout <= 8'b01111100; //  546 : 124 - 0x7c
      11'h223: dout <= 8'b11111000; //  547 : 248 - 0xf8
      11'h224: dout <= 8'b01110000; //  548 : 112 - 0x70
      11'h225: dout <= 8'b00100010; //  549 :  34 - 0x22
      11'h226: dout <= 8'b00000101; //  550 :   5 - 0x5
      11'h227: dout <= 8'b00000010; //  551 :   2 - 0x2
      11'h228: dout <= 8'b01001111; //  552 :  79 - 0x4f -- Sprite 0x45
      11'h229: dout <= 8'b01000111; //  553 :  71 - 0x47
      11'h22A: dout <= 8'b01000111; //  554 :  71 - 0x47
      11'h22B: dout <= 8'b01000111; //  555 :  71 - 0x47
      11'h22C: dout <= 8'b01000111; //  556 :  71 - 0x47
      11'h22D: dout <= 8'b01000111; //  557 :  71 - 0x47
      11'h22E: dout <= 8'b01000111; //  558 :  71 - 0x47
      11'h22F: dout <= 8'b01000111; //  559 :  71 - 0x47
      11'h230: dout <= 8'b10100000; //  560 : 160 - 0xa0 -- Sprite 0x46
      11'h231: dout <= 8'b10011111; //  561 : 159 - 0x9f
      11'h232: dout <= 8'b11000000; //  562 : 192 - 0xc0
      11'h233: dout <= 8'b11100000; //  563 : 224 - 0xe0
      11'h234: dout <= 8'b11111000; //  564 : 248 - 0xf8
      11'h235: dout <= 8'b11111111; //  565 : 255 - 0xff
      11'h236: dout <= 8'b11111111; //  566 : 255 - 0xff
      11'h237: dout <= 8'b11111111; //  567 : 255 - 0xff
      11'h238: dout <= 8'b00001100; //  568 :  12 - 0xc -- Sprite 0x47
      11'h239: dout <= 8'b11110000; //  569 : 240 - 0xf0
      11'h23A: dout <= 8'b00000000; //  570 :   0 - 0x0
      11'h23B: dout <= 8'b00000000; //  571 :   0 - 0x0
      11'h23C: dout <= 8'b00000001; //  572 :   1 - 0x1
      11'h23D: dout <= 8'b11111111; //  573 : 255 - 0xff
      11'h23E: dout <= 8'b11111111; //  574 : 255 - 0xff
      11'h23F: dout <= 8'b11111111; //  575 : 255 - 0xff
      11'h240: dout <= 8'b00001100; //  576 :  12 - 0xc -- Sprite 0x48
      11'h241: dout <= 8'b00011101; //  577 :  29 - 0x1d
      11'h242: dout <= 8'b00111000; //  578 :  56 - 0x38
      11'h243: dout <= 8'b01111110; //  579 : 126 - 0x7e
      11'h244: dout <= 8'b11111110; //  580 : 254 - 0xfe
      11'h245: dout <= 8'b11111111; //  581 : 255 - 0xff
      11'h246: dout <= 8'b11111111; //  582 : 255 - 0xff
      11'h247: dout <= 8'b11111111; //  583 : 255 - 0xff
      11'h248: dout <= 8'b11111111; //  584 : 255 - 0xff -- Sprite 0x49
      11'h249: dout <= 8'b11111111; //  585 : 255 - 0xff
      11'h24A: dout <= 8'b11111111; //  586 : 255 - 0xff
      11'h24B: dout <= 8'b11111111; //  587 : 255 - 0xff
      11'h24C: dout <= 8'b11111111; //  588 : 255 - 0xff
      11'h24D: dout <= 8'b11111111; //  589 : 255 - 0xff
      11'h24E: dout <= 8'b11111111; //  590 : 255 - 0xff
      11'h24F: dout <= 8'b11111111; //  591 : 255 - 0xff
      11'h250: dout <= 8'b11111111; //  592 : 255 - 0xff -- Sprite 0x4a
      11'h251: dout <= 8'b11101111; //  593 : 239 - 0xef
      11'h252: dout <= 8'b11111101; //  594 : 253 - 0xfd
      11'h253: dout <= 8'b11111111; //  595 : 255 - 0xff
      11'h254: dout <= 8'b11111111; //  596 : 255 - 0xff
      11'h255: dout <= 8'b11101111; //  597 : 239 - 0xef
      11'h256: dout <= 8'b11111110; //  598 : 254 - 0xfe
      11'h257: dout <= 8'b11111111; //  599 : 255 - 0xff
      11'h258: dout <= 8'b11111111; //  600 : 255 - 0xff -- Sprite 0x4b
      11'h259: dout <= 8'b11101010; //  601 : 234 - 0xea
      11'h25A: dout <= 8'b11111111; //  602 : 255 - 0xff
      11'h25B: dout <= 8'b10101111; //  603 : 175 - 0xaf
      11'h25C: dout <= 8'b11111111; //  604 : 255 - 0xff
      11'h25D: dout <= 8'b11111111; //  605 : 255 - 0xff
      11'h25E: dout <= 8'b11111010; //  606 : 250 - 0xfa
      11'h25F: dout <= 8'b11111111; //  607 : 255 - 0xff
      11'h260: dout <= 8'b11111111; //  608 : 255 - 0xff -- Sprite 0x4c
      11'h261: dout <= 8'b11111111; //  609 : 255 - 0xff
      11'h262: dout <= 8'b11111111; //  610 : 255 - 0xff
      11'h263: dout <= 8'b11111111; //  611 : 255 - 0xff
      11'h264: dout <= 8'b11111111; //  612 : 255 - 0xff
      11'h265: dout <= 8'b11111111; //  613 : 255 - 0xff
      11'h266: dout <= 8'b11111110; //  614 : 254 - 0xfe
      11'h267: dout <= 8'b11111111; //  615 : 255 - 0xff
      11'h268: dout <= 8'b11111111; //  616 : 255 - 0xff -- Sprite 0x4d
      11'h269: dout <= 8'b10111111; //  617 : 191 - 0xbf
      11'h26A: dout <= 8'b11111110; //  618 : 254 - 0xfe
      11'h26B: dout <= 8'b10101111; //  619 : 175 - 0xaf
      11'h26C: dout <= 8'b11111111; //  620 : 255 - 0xff
      11'h26D: dout <= 8'b11111111; //  621 : 255 - 0xff
      11'h26E: dout <= 8'b11101111; //  622 : 239 - 0xef
      11'h26F: dout <= 8'b11111111; //  623 : 255 - 0xff
      11'h270: dout <= 8'b11111111; //  624 : 255 - 0xff -- Sprite 0x4e
      11'h271: dout <= 8'b11111111; //  625 : 255 - 0xff
      11'h272: dout <= 8'b11111011; //  626 : 251 - 0xfb
      11'h273: dout <= 8'b11111111; //  627 : 255 - 0xff
      11'h274: dout <= 8'b11111111; //  628 : 255 - 0xff
      11'h275: dout <= 8'b11111111; //  629 : 255 - 0xff
      11'h276: dout <= 8'b11111110; //  630 : 254 - 0xfe
      11'h277: dout <= 8'b11111111; //  631 : 255 - 0xff
      11'h278: dout <= 8'b11111111; //  632 : 255 - 0xff -- Sprite 0x4f
      11'h279: dout <= 8'b11111111; //  633 : 255 - 0xff
      11'h27A: dout <= 8'b11110111; //  634 : 247 - 0xf7
      11'h27B: dout <= 8'b11111110; //  635 : 254 - 0xfe
      11'h27C: dout <= 8'b11111011; //  636 : 251 - 0xfb
      11'h27D: dout <= 8'b11111111; //  637 : 255 - 0xff
      11'h27E: dout <= 8'b11101111; //  638 : 239 - 0xef
      11'h27F: dout <= 8'b11111101; //  639 : 253 - 0xfd
      11'h280: dout <= 8'b11111111; //  640 : 255 - 0xff -- Sprite 0x50
      11'h281: dout <= 8'b11111111; //  641 : 255 - 0xff
      11'h282: dout <= 8'b00000011; //  642 :   3 - 0x3
      11'h283: dout <= 8'b00000001; //  643 :   1 - 0x1
      11'h284: dout <= 8'b11101110; //  644 : 238 - 0xee
      11'h285: dout <= 8'b00000000; //  645 :   0 - 0x0
      11'h286: dout <= 8'b11101110; //  646 : 238 - 0xee
      11'h287: dout <= 8'b11101110; //  647 : 238 - 0xee
      11'h288: dout <= 8'b11111111; //  648 : 255 - 0xff -- Sprite 0x51
      11'h289: dout <= 8'b11111111; //  649 : 255 - 0xff
      11'h28A: dout <= 8'b00000011; //  650 :   3 - 0x3
      11'h28B: dout <= 8'b00000001; //  651 :   1 - 0x1
      11'h28C: dout <= 8'b11101110; //  652 : 238 - 0xee
      11'h28D: dout <= 8'b00000000; //  653 :   0 - 0x0
      11'h28E: dout <= 8'b11101110; //  654 : 238 - 0xee
      11'h28F: dout <= 8'b11101110; //  655 : 238 - 0xee
      11'h290: dout <= 8'b11111111; //  656 : 255 - 0xff -- Sprite 0x52
      11'h291: dout <= 8'b11111111; //  657 : 255 - 0xff
      11'h292: dout <= 8'b00000001; //  658 :   1 - 0x1
      11'h293: dout <= 8'b00000000; //  659 :   0 - 0x0
      11'h294: dout <= 8'b11100000; //  660 : 224 - 0xe0
      11'h295: dout <= 8'b00001111; //  661 :  15 - 0xf
      11'h296: dout <= 8'b11111111; //  662 : 255 - 0xff
      11'h297: dout <= 8'b11111011; //  663 : 251 - 0xfb
      11'h298: dout <= 8'b11111111; //  664 : 255 - 0xff -- Sprite 0x53
      11'h299: dout <= 8'b11111111; //  665 : 255 - 0xff
      11'h29A: dout <= 8'b10000011; //  666 : 131 - 0x83
      11'h29B: dout <= 8'b00000001; //  667 :   1 - 0x1
      11'h29C: dout <= 8'b11101110; //  668 : 238 - 0xee
      11'h29D: dout <= 8'b00000000; //  669 :   0 - 0x0
      11'h29E: dout <= 8'b11111111; //  670 : 255 - 0xff
      11'h29F: dout <= 8'b11111111; //  671 : 255 - 0xff
      11'h2A0: dout <= 8'b11111111; //  672 : 255 - 0xff -- Sprite 0x54
      11'h2A1: dout <= 8'b11111111; //  673 : 255 - 0xff
      11'h2A2: dout <= 8'b00000001; //  674 :   1 - 0x1
      11'h2A3: dout <= 8'b00000000; //  675 :   0 - 0x0
      11'h2A4: dout <= 8'b10111000; //  676 : 184 - 0xb8
      11'h2A5: dout <= 8'b11000011; //  677 : 195 - 0xc3
      11'h2A6: dout <= 8'b11111011; //  678 : 251 - 0xfb
      11'h2A7: dout <= 8'b11111011; //  679 : 251 - 0xfb
      11'h2A8: dout <= 8'b11111111; //  680 : 255 - 0xff -- Sprite 0x55
      11'h2A9: dout <= 8'b11111111; //  681 : 255 - 0xff
      11'h2AA: dout <= 8'b10000011; //  682 : 131 - 0x83
      11'h2AB: dout <= 8'b00000001; //  683 :   1 - 0x1
      11'h2AC: dout <= 8'b11101110; //  684 : 238 - 0xee
      11'h2AD: dout <= 8'b00000000; //  685 :   0 - 0x0
      11'h2AE: dout <= 8'b11101110; //  686 : 238 - 0xee
      11'h2AF: dout <= 8'b11101110; //  687 : 238 - 0xee
      11'h2B0: dout <= 8'b11111111; //  688 : 255 - 0xff -- Sprite 0x56
      11'h2B1: dout <= 8'b11111111; //  689 : 255 - 0xff
      11'h2B2: dout <= 8'b00011111; //  690 :  31 - 0x1f
      11'h2B3: dout <= 8'b00001111; //  691 :  15 - 0xf
      11'h2B4: dout <= 8'b11101111; //  692 : 239 - 0xef
      11'h2B5: dout <= 8'b00001111; //  693 :  15 - 0xf
      11'h2B6: dout <= 8'b11101111; //  694 : 239 - 0xef
      11'h2B7: dout <= 8'b11101111; //  695 : 239 - 0xef
      11'h2B8: dout <= 8'b11111111; //  696 : 255 - 0xff -- Sprite 0x57
      11'h2B9: dout <= 8'b11111111; //  697 : 255 - 0xff
      11'h2BA: dout <= 8'b00010001; //  698 :  17 - 0x11
      11'h2BB: dout <= 8'b00000000; //  699 :   0 - 0x0
      11'h2BC: dout <= 8'b11101110; //  700 : 238 - 0xee
      11'h2BD: dout <= 8'b00000000; //  701 :   0 - 0x0
      11'h2BE: dout <= 8'b11101110; //  702 : 238 - 0xee
      11'h2BF: dout <= 8'b11101110; //  703 : 238 - 0xee
      11'h2C0: dout <= 8'b11111111; //  704 : 255 - 0xff -- Sprite 0x58
      11'h2C1: dout <= 8'b11111111; //  705 : 255 - 0xff
      11'h2C2: dout <= 8'b01110001; //  706 : 113 - 0x71
      11'h2C3: dout <= 8'b00110000; //  707 :  48 - 0x30
      11'h2C4: dout <= 8'b11111110; //  708 : 254 - 0xfe
      11'h2C5: dout <= 8'b00000000; //  709 :   0 - 0x0
      11'h2C6: dout <= 8'b11111110; //  710 : 254 - 0xfe
      11'h2C7: dout <= 8'b11101110; //  711 : 238 - 0xee
      11'h2C8: dout <= 8'b11111111; //  712 : 255 - 0xff -- Sprite 0x59
      11'h2C9: dout <= 8'b11111111; //  713 : 255 - 0xff
      11'h2CA: dout <= 8'b00000011; //  714 :   3 - 0x3
      11'h2CB: dout <= 8'b00000001; //  715 :   1 - 0x1
      11'h2CC: dout <= 8'b11101110; //  716 : 238 - 0xee
      11'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      11'h2CE: dout <= 8'b11101110; //  718 : 238 - 0xee
      11'h2CF: dout <= 8'b11101110; //  719 : 238 - 0xee
      11'h2D0: dout <= 8'b11111111; //  720 : 255 - 0xff -- Sprite 0x5a
      11'h2D1: dout <= 8'b11111111; //  721 : 255 - 0xff
      11'h2D2: dout <= 8'b10000011; //  722 : 131 - 0x83
      11'h2D3: dout <= 8'b00000001; //  723 :   1 - 0x1
      11'h2D4: dout <= 8'b11101110; //  724 : 238 - 0xee
      11'h2D5: dout <= 8'b00000000; //  725 :   0 - 0x0
      11'h2D6: dout <= 8'b11101110; //  726 : 238 - 0xee
      11'h2D7: dout <= 8'b11101110; //  727 : 238 - 0xee
      11'h2D8: dout <= 8'b11111111; //  728 : 255 - 0xff -- Sprite 0x5b
      11'h2D9: dout <= 8'b11111111; //  729 : 255 - 0xff
      11'h2DA: dout <= 8'b00000001; //  730 :   1 - 0x1
      11'h2DB: dout <= 8'b00000000; //  731 :   0 - 0x0
      11'h2DC: dout <= 8'b11100000; //  732 : 224 - 0xe0
      11'h2DD: dout <= 8'b00001111; //  733 :  15 - 0xf
      11'h2DE: dout <= 8'b11111111; //  734 : 255 - 0xff
      11'h2DF: dout <= 8'b11111011; //  735 : 251 - 0xfb
      11'h2E0: dout <= 8'b11111111; //  736 : 255 - 0xff -- Sprite 0x5c
      11'h2E1: dout <= 8'b11111111; //  737 : 255 - 0xff
      11'h2E2: dout <= 8'b11111111; //  738 : 255 - 0xff
      11'h2E3: dout <= 8'b11111111; //  739 : 255 - 0xff
      11'h2E4: dout <= 8'b11111111; //  740 : 255 - 0xff
      11'h2E5: dout <= 8'b11111111; //  741 : 255 - 0xff
      11'h2E6: dout <= 8'b11111111; //  742 : 255 - 0xff
      11'h2E7: dout <= 8'b11011101; //  743 : 221 - 0xdd
      11'h2E8: dout <= 8'b11111111; //  744 : 255 - 0xff -- Sprite 0x5d
      11'h2E9: dout <= 8'b11111111; //  745 : 255 - 0xff
      11'h2EA: dout <= 8'b00000001; //  746 :   1 - 0x1
      11'h2EB: dout <= 8'b00000000; //  747 :   0 - 0x0
      11'h2EC: dout <= 8'b11100000; //  748 : 224 - 0xe0
      11'h2ED: dout <= 8'b00001111; //  749 :  15 - 0xf
      11'h2EE: dout <= 8'b11111111; //  750 : 255 - 0xff
      11'h2EF: dout <= 8'b11111011; //  751 : 251 - 0xfb
      11'h2F0: dout <= 8'b11111111; //  752 : 255 - 0xff -- Sprite 0x5e
      11'h2F1: dout <= 8'b11111111; //  753 : 255 - 0xff
      11'h2F2: dout <= 8'b00010001; //  754 :  17 - 0x11
      11'h2F3: dout <= 8'b00000000; //  755 :   0 - 0x0
      11'h2F4: dout <= 8'b11101110; //  756 : 238 - 0xee
      11'h2F5: dout <= 8'b00000000; //  757 :   0 - 0x0
      11'h2F6: dout <= 8'b11101110; //  758 : 238 - 0xee
      11'h2F7: dout <= 8'b11101110; //  759 : 238 - 0xee
      11'h2F8: dout <= 8'b10111101; //  760 : 189 - 0xbd -- Sprite 0x5f
      11'h2F9: dout <= 8'b11111111; //  761 : 255 - 0xff
      11'h2FA: dout <= 8'b11111111; //  762 : 255 - 0xff
      11'h2FB: dout <= 8'b11111111; //  763 : 255 - 0xff
      11'h2FC: dout <= 8'b11111111; //  764 : 255 - 0xff
      11'h2FD: dout <= 8'b11111111; //  765 : 255 - 0xff
      11'h2FE: dout <= 8'b11111111; //  766 : 255 - 0xff
      11'h2FF: dout <= 8'b11111111; //  767 : 255 - 0xff
      11'h300: dout <= 8'b11101110; //  768 : 238 - 0xee -- Sprite 0x60
      11'h301: dout <= 8'b00000000; //  769 :   0 - 0x0
      11'h302: dout <= 8'b11111110; //  770 : 254 - 0xfe
      11'h303: dout <= 8'b00000000; //  771 :   0 - 0x0
      11'h304: dout <= 8'b00000001; //  772 :   1 - 0x1
      11'h305: dout <= 8'b00001111; //  773 :  15 - 0xf
      11'h306: dout <= 8'b10001111; //  774 : 143 - 0x8f
      11'h307: dout <= 8'b11111111; //  775 : 255 - 0xff
      11'h308: dout <= 8'b11101110; //  776 : 238 - 0xee -- Sprite 0x61
      11'h309: dout <= 8'b00000000; //  777 :   0 - 0x0
      11'h30A: dout <= 8'b11111100; //  778 : 252 - 0xfc
      11'h30B: dout <= 8'b00000001; //  779 :   1 - 0x1
      11'h30C: dout <= 8'b00000001; //  780 :   1 - 0x1
      11'h30D: dout <= 8'b00000000; //  781 :   0 - 0x0
      11'h30E: dout <= 8'b10001000; //  782 : 136 - 0x88
      11'h30F: dout <= 8'b11111111; //  783 : 255 - 0xff
      11'h310: dout <= 8'b11100011; //  784 : 227 - 0xe3 -- Sprite 0x62
      11'h311: dout <= 8'b00001111; //  785 :  15 - 0xf
      11'h312: dout <= 8'b11101111; //  786 : 239 - 0xef
      11'h313: dout <= 8'b00001111; //  787 :  15 - 0xf
      11'h314: dout <= 8'b00000001; //  788 :   1 - 0x1
      11'h315: dout <= 8'b00000000; //  789 :   0 - 0x0
      11'h316: dout <= 8'b10000000; //  790 : 128 - 0x80
      11'h317: dout <= 8'b11111111; //  791 : 255 - 0xff
      11'h318: dout <= 8'b11001110; //  792 : 206 - 0xce -- Sprite 0x63
      11'h319: dout <= 8'b11110000; //  793 : 240 - 0xf0
      11'h31A: dout <= 8'b11111110; //  794 : 254 - 0xfe
      11'h31B: dout <= 8'b00010000; //  795 :  16 - 0x10
      11'h31C: dout <= 8'b00000000; //  796 :   0 - 0x0
      11'h31D: dout <= 8'b10000000; //  797 : 128 - 0x80
      11'h31E: dout <= 8'b11000001; //  798 : 193 - 0xc1
      11'h31F: dout <= 8'b11111111; //  799 : 255 - 0xff
      11'h320: dout <= 8'b11111011; //  800 : 251 - 0xfb -- Sprite 0x64
      11'h321: dout <= 8'b11000011; //  801 : 195 - 0xc3
      11'h322: dout <= 8'b11111011; //  802 : 251 - 0xfb
      11'h323: dout <= 8'b11000011; //  803 : 195 - 0xc3
      11'h324: dout <= 8'b11000011; //  804 : 195 - 0xc3
      11'h325: dout <= 8'b11000011; //  805 : 195 - 0xc3
      11'h326: dout <= 8'b11100011; //  806 : 227 - 0xe3
      11'h327: dout <= 8'b11111111; //  807 : 255 - 0xff
      11'h328: dout <= 8'b11101110; //  808 : 238 - 0xee -- Sprite 0x65
      11'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      11'h32A: dout <= 8'b11111110; //  810 : 254 - 0xfe
      11'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      11'h32C: dout <= 8'b00000000; //  812 :   0 - 0x0
      11'h32D: dout <= 8'b00000000; //  813 :   0 - 0x0
      11'h32E: dout <= 8'b10001000; //  814 : 136 - 0x88
      11'h32F: dout <= 8'b11111111; //  815 : 255 - 0xff
      11'h330: dout <= 8'b11101111; //  816 : 239 - 0xef -- Sprite 0x66
      11'h331: dout <= 8'b00001111; //  817 :  15 - 0xf
      11'h332: dout <= 8'b11101111; //  818 : 239 - 0xef
      11'h333: dout <= 8'b00000001; //  819 :   1 - 0x1
      11'h334: dout <= 8'b00000000; //  820 :   0 - 0x0
      11'h335: dout <= 8'b00000000; //  821 :   0 - 0x0
      11'h336: dout <= 8'b10000000; //  822 : 128 - 0x80
      11'h337: dout <= 8'b11111111; //  823 : 255 - 0xff
      11'h338: dout <= 8'b11101110; //  824 : 238 - 0xee -- Sprite 0x67
      11'h339: dout <= 8'b00000000; //  825 :   0 - 0x0
      11'h33A: dout <= 8'b11111110; //  826 : 254 - 0xfe
      11'h33B: dout <= 8'b00000000; //  827 :   0 - 0x0
      11'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      11'h33D: dout <= 8'b00001000; //  829 :   8 - 0x8
      11'h33E: dout <= 8'b10011100; //  830 : 156 - 0x9c
      11'h33F: dout <= 8'b11111111; //  831 : 255 - 0xff
      11'h340: dout <= 8'b11101110; //  832 : 238 - 0xee -- Sprite 0x68
      11'h341: dout <= 8'b00000000; //  833 :   0 - 0x0
      11'h342: dout <= 8'b11101110; //  834 : 238 - 0xee
      11'h343: dout <= 8'b00000000; //  835 :   0 - 0x0
      11'h344: dout <= 8'b00000000; //  836 :   0 - 0x0
      11'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      11'h346: dout <= 8'b10001000; //  838 : 136 - 0x88
      11'h347: dout <= 8'b11111111; //  839 : 255 - 0xff
      11'h348: dout <= 8'b11101110; //  840 : 238 - 0xee -- Sprite 0x69
      11'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      11'h34A: dout <= 8'b11101110; //  842 : 238 - 0xee
      11'h34B: dout <= 8'b00000000; //  843 :   0 - 0x0
      11'h34C: dout <= 8'b00000000; //  844 :   0 - 0x0
      11'h34D: dout <= 8'b00000000; //  845 :   0 - 0x0
      11'h34E: dout <= 8'b10000001; //  846 : 129 - 0x81
      11'h34F: dout <= 8'b11111111; //  847 : 255 - 0xff
      11'h350: dout <= 8'b11101110; //  848 : 238 - 0xee -- Sprite 0x6a
      11'h351: dout <= 8'b00000000; //  849 :   0 - 0x0
      11'h352: dout <= 8'b11101110; //  850 : 238 - 0xee
      11'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      11'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      11'h355: dout <= 8'b10000000; //  853 : 128 - 0x80
      11'h356: dout <= 8'b11000001; //  854 : 193 - 0xc1
      11'h357: dout <= 8'b11111111; //  855 : 255 - 0xff
      11'h358: dout <= 8'b11100011; //  856 : 227 - 0xe3 -- Sprite 0x6b
      11'h359: dout <= 8'b00001111; //  857 :  15 - 0xf
      11'h35A: dout <= 8'b11101111; //  858 : 239 - 0xef
      11'h35B: dout <= 8'b00001111; //  859 :  15 - 0xf
      11'h35C: dout <= 8'b00000001; //  860 :   1 - 0x1
      11'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      11'h35E: dout <= 8'b10000000; //  862 : 128 - 0x80
      11'h35F: dout <= 8'b11111111; //  863 : 255 - 0xff
      11'h360: dout <= 8'b10011001; //  864 : 153 - 0x99 -- Sprite 0x6c
      11'h361: dout <= 8'b11100011; //  865 : 227 - 0xe3
      11'h362: dout <= 8'b11110011; //  866 : 243 - 0xf3
      11'h363: dout <= 8'b11000111; //  867 : 199 - 0xc7
      11'h364: dout <= 8'b10000001; //  868 : 129 - 0x81
      11'h365: dout <= 8'b10001000; //  869 : 136 - 0x88
      11'h366: dout <= 8'b11001100; //  870 : 204 - 0xcc
      11'h367: dout <= 8'b11111111; //  871 : 255 - 0xff
      11'h368: dout <= 8'b11100011; //  872 : 227 - 0xe3 -- Sprite 0x6d
      11'h369: dout <= 8'b00001111; //  873 :  15 - 0xf
      11'h36A: dout <= 8'b11101111; //  874 : 239 - 0xef
      11'h36B: dout <= 8'b00001111; //  875 :  15 - 0xf
      11'h36C: dout <= 8'b00001111; //  876 :  15 - 0xf
      11'h36D: dout <= 8'b00001111; //  877 :  15 - 0xf
      11'h36E: dout <= 8'b10001111; //  878 : 143 - 0x8f
      11'h36F: dout <= 8'b11111111; //  879 : 255 - 0xff
      11'h370: dout <= 8'b11101110; //  880 : 238 - 0xee -- Sprite 0x6e
      11'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout <= 8'b11101110; //  882 : 238 - 0xee
      11'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      11'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      11'h375: dout <= 8'b10000000; //  885 : 128 - 0x80
      11'h376: dout <= 8'b11000001; //  886 : 193 - 0xc1
      11'h377: dout <= 8'b11111111; //  887 : 255 - 0xff
      11'h378: dout <= 8'b11111111; //  888 : 255 - 0xff -- Sprite 0x6f
      11'h379: dout <= 8'b11111111; //  889 : 255 - 0xff
      11'h37A: dout <= 8'b11111111; //  890 : 255 - 0xff
      11'h37B: dout <= 8'b10111101; //  891 : 189 - 0xbd
      11'h37C: dout <= 8'b11111111; //  892 : 255 - 0xff
      11'h37D: dout <= 8'b11011011; //  893 : 219 - 0xdb
      11'h37E: dout <= 8'b11111111; //  894 : 255 - 0xff
      11'h37F: dout <= 8'b11111111; //  895 : 255 - 0xff
      11'h380: dout <= 8'b11111011; //  896 : 251 - 0xfb -- Sprite 0x70
      11'h381: dout <= 8'b11101111; //  897 : 239 - 0xef
      11'h382: dout <= 8'b11011111; //  898 : 223 - 0xdf
      11'h383: dout <= 8'b11111111; //  899 : 255 - 0xff
      11'h384: dout <= 8'b10111111; //  900 : 191 - 0xbf
      11'h385: dout <= 8'b10111111; //  901 : 191 - 0xbf
      11'h386: dout <= 8'b11111110; //  902 : 254 - 0xfe
      11'h387: dout <= 8'b11111111; //  903 : 255 - 0xff
      11'h388: dout <= 8'b11011111; //  904 : 223 - 0xdf -- Sprite 0x71
      11'h389: dout <= 8'b11110111; //  905 : 247 - 0xf7
      11'h38A: dout <= 8'b11111011; //  906 : 251 - 0xfb
      11'h38B: dout <= 8'b11111111; //  907 : 255 - 0xff
      11'h38C: dout <= 8'b11111101; //  908 : 253 - 0xfd
      11'h38D: dout <= 8'b11111101; //  909 : 253 - 0xfd
      11'h38E: dout <= 8'b01111111; //  910 : 127 - 0x7f
      11'h38F: dout <= 8'b11111111; //  911 : 255 - 0xff
      11'h390: dout <= 8'b11111111; //  912 : 255 - 0xff -- Sprite 0x72
      11'h391: dout <= 8'b11111111; //  913 : 255 - 0xff
      11'h392: dout <= 8'b11111111; //  914 : 255 - 0xff
      11'h393: dout <= 8'b11111111; //  915 : 255 - 0xff
      11'h394: dout <= 8'b11111111; //  916 : 255 - 0xff
      11'h395: dout <= 8'b11111111; //  917 : 255 - 0xff
      11'h396: dout <= 8'b11111111; //  918 : 255 - 0xff
      11'h397: dout <= 8'b11111111; //  919 : 255 - 0xff
      11'h398: dout <= 8'b11111111; //  920 : 255 - 0xff -- Sprite 0x73
      11'h399: dout <= 8'b11111110; //  921 : 254 - 0xfe
      11'h39A: dout <= 8'b10111111; //  922 : 191 - 0xbf
      11'h39B: dout <= 8'b10111111; //  923 : 191 - 0xbf
      11'h39C: dout <= 8'b11111111; //  924 : 255 - 0xff
      11'h39D: dout <= 8'b11011111; //  925 : 223 - 0xdf
      11'h39E: dout <= 8'b11101111; //  926 : 239 - 0xef
      11'h39F: dout <= 8'b11111011; //  927 : 251 - 0xfb
      11'h3A0: dout <= 8'b11111111; //  928 : 255 - 0xff -- Sprite 0x74
      11'h3A1: dout <= 8'b01111111; //  929 : 127 - 0x7f
      11'h3A2: dout <= 8'b11111101; //  930 : 253 - 0xfd
      11'h3A3: dout <= 8'b11111101; //  931 : 253 - 0xfd
      11'h3A4: dout <= 8'b11111111; //  932 : 255 - 0xff
      11'h3A5: dout <= 8'b11111011; //  933 : 251 - 0xfb
      11'h3A6: dout <= 8'b11110111; //  934 : 247 - 0xf7
      11'h3A7: dout <= 8'b11011111; //  935 : 223 - 0xdf
      11'h3A8: dout <= 8'b11111111; //  936 : 255 - 0xff -- Sprite 0x75
      11'h3A9: dout <= 8'b11111111; //  937 : 255 - 0xff
      11'h3AA: dout <= 8'b11111111; //  938 : 255 - 0xff
      11'h3AB: dout <= 8'b11111111; //  939 : 255 - 0xff
      11'h3AC: dout <= 8'b11111111; //  940 : 255 - 0xff
      11'h3AD: dout <= 8'b11111111; //  941 : 255 - 0xff
      11'h3AE: dout <= 8'b11111111; //  942 : 255 - 0xff
      11'h3AF: dout <= 8'b11111111; //  943 : 255 - 0xff
      11'h3B0: dout <= 8'b11111111; //  944 : 255 - 0xff -- Sprite 0x76
      11'h3B1: dout <= 8'b11111111; //  945 : 255 - 0xff
      11'h3B2: dout <= 8'b11111111; //  946 : 255 - 0xff
      11'h3B3: dout <= 8'b11111111; //  947 : 255 - 0xff
      11'h3B4: dout <= 8'b11111111; //  948 : 255 - 0xff
      11'h3B5: dout <= 8'b11111111; //  949 : 255 - 0xff
      11'h3B6: dout <= 8'b11111111; //  950 : 255 - 0xff
      11'h3B7: dout <= 8'b11111111; //  951 : 255 - 0xff
      11'h3B8: dout <= 8'b11111111; //  952 : 255 - 0xff -- Sprite 0x77
      11'h3B9: dout <= 8'b11111111; //  953 : 255 - 0xff
      11'h3BA: dout <= 8'b11111111; //  954 : 255 - 0xff
      11'h3BB: dout <= 8'b11111111; //  955 : 255 - 0xff
      11'h3BC: dout <= 8'b11111111; //  956 : 255 - 0xff
      11'h3BD: dout <= 8'b11111111; //  957 : 255 - 0xff
      11'h3BE: dout <= 8'b11111111; //  958 : 255 - 0xff
      11'h3BF: dout <= 8'b11111111; //  959 : 255 - 0xff
      11'h3C0: dout <= 8'b11111111; //  960 : 255 - 0xff -- Sprite 0x78
      11'h3C1: dout <= 8'b11111111; //  961 : 255 - 0xff
      11'h3C2: dout <= 8'b11111111; //  962 : 255 - 0xff
      11'h3C3: dout <= 8'b11111111; //  963 : 255 - 0xff
      11'h3C4: dout <= 8'b11111111; //  964 : 255 - 0xff
      11'h3C5: dout <= 8'b11111111; //  965 : 255 - 0xff
      11'h3C6: dout <= 8'b11111111; //  966 : 255 - 0xff
      11'h3C7: dout <= 8'b11111111; //  967 : 255 - 0xff
      11'h3C8: dout <= 8'b11111111; //  968 : 255 - 0xff -- Sprite 0x79
      11'h3C9: dout <= 8'b11111111; //  969 : 255 - 0xff
      11'h3CA: dout <= 8'b11111111; //  970 : 255 - 0xff
      11'h3CB: dout <= 8'b11111111; //  971 : 255 - 0xff
      11'h3CC: dout <= 8'b11111111; //  972 : 255 - 0xff
      11'h3CD: dout <= 8'b11111111; //  973 : 255 - 0xff
      11'h3CE: dout <= 8'b11111111; //  974 : 255 - 0xff
      11'h3CF: dout <= 8'b11111111; //  975 : 255 - 0xff
      11'h3D0: dout <= 8'b11111111; //  976 : 255 - 0xff -- Sprite 0x7a
      11'h3D1: dout <= 8'b11111111; //  977 : 255 - 0xff
      11'h3D2: dout <= 8'b11111111; //  978 : 255 - 0xff
      11'h3D3: dout <= 8'b11111111; //  979 : 255 - 0xff
      11'h3D4: dout <= 8'b11111111; //  980 : 255 - 0xff
      11'h3D5: dout <= 8'b11111111; //  981 : 255 - 0xff
      11'h3D6: dout <= 8'b11111111; //  982 : 255 - 0xff
      11'h3D7: dout <= 8'b11111111; //  983 : 255 - 0xff
      11'h3D8: dout <= 8'b11111111; //  984 : 255 - 0xff -- Sprite 0x7b
      11'h3D9: dout <= 8'b11111111; //  985 : 255 - 0xff
      11'h3DA: dout <= 8'b11111111; //  986 : 255 - 0xff
      11'h3DB: dout <= 8'b11111111; //  987 : 255 - 0xff
      11'h3DC: dout <= 8'b11111111; //  988 : 255 - 0xff
      11'h3DD: dout <= 8'b11111111; //  989 : 255 - 0xff
      11'h3DE: dout <= 8'b11111111; //  990 : 255 - 0xff
      11'h3DF: dout <= 8'b11111111; //  991 : 255 - 0xff
      11'h3E0: dout <= 8'b11111111; //  992 : 255 - 0xff -- Sprite 0x7c
      11'h3E1: dout <= 8'b11111111; //  993 : 255 - 0xff
      11'h3E2: dout <= 8'b11111111; //  994 : 255 - 0xff
      11'h3E3: dout <= 8'b11111111; //  995 : 255 - 0xff
      11'h3E4: dout <= 8'b11111111; //  996 : 255 - 0xff
      11'h3E5: dout <= 8'b11111111; //  997 : 255 - 0xff
      11'h3E6: dout <= 8'b11111111; //  998 : 255 - 0xff
      11'h3E7: dout <= 8'b11111111; //  999 : 255 - 0xff
      11'h3E8: dout <= 8'b11111111; // 1000 : 255 - 0xff -- Sprite 0x7d
      11'h3E9: dout <= 8'b11111111; // 1001 : 255 - 0xff
      11'h3EA: dout <= 8'b11111111; // 1002 : 255 - 0xff
      11'h3EB: dout <= 8'b11111111; // 1003 : 255 - 0xff
      11'h3EC: dout <= 8'b11111111; // 1004 : 255 - 0xff
      11'h3ED: dout <= 8'b11111111; // 1005 : 255 - 0xff
      11'h3EE: dout <= 8'b11111111; // 1006 : 255 - 0xff
      11'h3EF: dout <= 8'b11111111; // 1007 : 255 - 0xff
      11'h3F0: dout <= 8'b11111111; // 1008 : 255 - 0xff -- Sprite 0x7e
      11'h3F1: dout <= 8'b11111111; // 1009 : 255 - 0xff
      11'h3F2: dout <= 8'b11111111; // 1010 : 255 - 0xff
      11'h3F3: dout <= 8'b11111111; // 1011 : 255 - 0xff
      11'h3F4: dout <= 8'b11111111; // 1012 : 255 - 0xff
      11'h3F5: dout <= 8'b11111111; // 1013 : 255 - 0xff
      11'h3F6: dout <= 8'b11111111; // 1014 : 255 - 0xff
      11'h3F7: dout <= 8'b11111111; // 1015 : 255 - 0xff
      11'h3F8: dout <= 8'b11111111; // 1016 : 255 - 0xff -- Sprite 0x7f
      11'h3F9: dout <= 8'b11111111; // 1017 : 255 - 0xff
      11'h3FA: dout <= 8'b11111111; // 1018 : 255 - 0xff
      11'h3FB: dout <= 8'b11111111; // 1019 : 255 - 0xff
      11'h3FC: dout <= 8'b11111111; // 1020 : 255 - 0xff
      11'h3FD: dout <= 8'b11111111; // 1021 : 255 - 0xff
      11'h3FE: dout <= 8'b11111111; // 1022 : 255 - 0xff
      11'h3FF: dout <= 8'b11111111; // 1023 : 255 - 0xff
      11'h400: dout <= 8'b10111111; // 1024 : 191 - 0xbf -- Sprite 0x80
      11'h401: dout <= 8'b11110111; // 1025 : 247 - 0xf7
      11'h402: dout <= 8'b11111101; // 1026 : 253 - 0xfd
      11'h403: dout <= 8'b11011111; // 1027 : 223 - 0xdf
      11'h404: dout <= 8'b11111011; // 1028 : 251 - 0xfb
      11'h405: dout <= 8'b10111111; // 1029 : 191 - 0xbf
      11'h406: dout <= 8'b11111110; // 1030 : 254 - 0xfe
      11'h407: dout <= 8'b11101111; // 1031 : 239 - 0xef
      11'h408: dout <= 8'b11111111; // 1032 : 255 - 0xff -- Sprite 0x81
      11'h409: dout <= 8'b11101110; // 1033 : 238 - 0xee
      11'h40A: dout <= 8'b11111111; // 1034 : 255 - 0xff
      11'h40B: dout <= 8'b11011111; // 1035 : 223 - 0xdf
      11'h40C: dout <= 8'b01110111; // 1036 : 119 - 0x77
      11'h40D: dout <= 8'b11111101; // 1037 : 253 - 0xfd
      11'h40E: dout <= 8'b11011111; // 1038 : 223 - 0xdf
      11'h40F: dout <= 8'b10111111; // 1039 : 191 - 0xbf
      11'h410: dout <= 8'b11111110; // 1040 : 254 - 0xfe -- Sprite 0x82
      11'h411: dout <= 8'b11101111; // 1041 : 239 - 0xef
      11'h412: dout <= 8'b10111111; // 1042 : 191 - 0xbf
      11'h413: dout <= 8'b11110111; // 1043 : 247 - 0xf7
      11'h414: dout <= 8'b11111101; // 1044 : 253 - 0xfd
      11'h415: dout <= 8'b11011111; // 1045 : 223 - 0xdf
      11'h416: dout <= 8'b11111011; // 1046 : 251 - 0xfb
      11'h417: dout <= 8'b10111111; // 1047 : 191 - 0xbf
      11'h418: dout <= 8'b11101111; // 1048 : 239 - 0xef -- Sprite 0x83
      11'h419: dout <= 8'b11111111; // 1049 : 255 - 0xff
      11'h41A: dout <= 8'b10111011; // 1050 : 187 - 0xbb
      11'h41B: dout <= 8'b11111111; // 1051 : 255 - 0xff
      11'h41C: dout <= 8'b11110111; // 1052 : 247 - 0xf7
      11'h41D: dout <= 8'b11011101; // 1053 : 221 - 0xdd
      11'h41E: dout <= 8'b01111111; // 1054 : 127 - 0x7f
      11'h41F: dout <= 8'b11110111; // 1055 : 247 - 0xf7
      11'h420: dout <= 8'b11111111; // 1056 : 255 - 0xff -- Sprite 0x84
      11'h421: dout <= 8'b11101110; // 1057 : 238 - 0xee
      11'h422: dout <= 8'b11111011; // 1058 : 251 - 0xfb
      11'h423: dout <= 8'b10111111; // 1059 : 191 - 0xbf
      11'h424: dout <= 8'b01111111; // 1060 : 127 - 0x7f
      11'h425: dout <= 8'b11101101; // 1061 : 237 - 0xed
      11'h426: dout <= 8'b11111111; // 1062 : 255 - 0xff
      11'h427: dout <= 8'b10111111; // 1063 : 191 - 0xbf
      11'h428: dout <= 8'b11111111; // 1064 : 255 - 0xff -- Sprite 0x85
      11'h429: dout <= 8'b10111111; // 1065 : 191 - 0xbf
      11'h42A: dout <= 8'b01111101; // 1066 : 125 - 0x7d
      11'h42B: dout <= 8'b11110111; // 1067 : 247 - 0xf7
      11'h42C: dout <= 8'b11011011; // 1068 : 219 - 0xdb
      11'h42D: dout <= 8'b11111101; // 1069 : 253 - 0xfd
      11'h42E: dout <= 8'b01111110; // 1070 : 126 - 0x7e
      11'h42F: dout <= 8'b11111011; // 1071 : 251 - 0xfb
      11'h430: dout <= 8'b11111111; // 1072 : 255 - 0xff -- Sprite 0x86
      11'h431: dout <= 8'b11110111; // 1073 : 247 - 0xf7
      11'h432: dout <= 8'b11111111; // 1074 : 255 - 0xff
      11'h433: dout <= 8'b11011101; // 1075 : 221 - 0xdd
      11'h434: dout <= 8'b01111111; // 1076 : 127 - 0x7f
      11'h435: dout <= 8'b11110111; // 1077 : 247 - 0xf7
      11'h436: dout <= 8'b11101111; // 1078 : 239 - 0xef
      11'h437: dout <= 8'b10111101; // 1079 : 189 - 0xbd
      11'h438: dout <= 8'b01011111; // 1080 :  95 - 0x5f -- Sprite 0x87
      11'h439: dout <= 8'b11111101; // 1081 : 253 - 0xfd
      11'h43A: dout <= 8'b11110110; // 1082 : 246 - 0xf6
      11'h43B: dout <= 8'b01111111; // 1083 : 127 - 0x7f
      11'h43C: dout <= 8'b10011111; // 1084 : 159 - 0x9f
      11'h43D: dout <= 8'b11111110; // 1085 : 254 - 0xfe
      11'h43E: dout <= 8'b11111111; // 1086 : 255 - 0xff
      11'h43F: dout <= 8'b11101111; // 1087 : 239 - 0xef
      11'h440: dout <= 8'b11111111; // 1088 : 255 - 0xff -- Sprite 0x88
      11'h441: dout <= 8'b11111111; // 1089 : 255 - 0xff
      11'h442: dout <= 8'b10011111; // 1090 : 159 - 0x9f
      11'h443: dout <= 8'b10110011; // 1091 : 179 - 0xb3
      11'h444: dout <= 8'b11110011; // 1092 : 243 - 0xf3
      11'h445: dout <= 8'b11111111; // 1093 : 255 - 0xff
      11'h446: dout <= 8'b11111111; // 1094 : 255 - 0xff
      11'h447: dout <= 8'b11111111; // 1095 : 255 - 0xff
      11'h448: dout <= 8'b11111111; // 1096 : 255 - 0xff -- Sprite 0x89
      11'h449: dout <= 8'b11001111; // 1097 : 207 - 0xcf
      11'h44A: dout <= 8'b11011111; // 1098 : 223 - 0xdf
      11'h44B: dout <= 8'b11111111; // 1099 : 255 - 0xff
      11'h44C: dout <= 8'b11110011; // 1100 : 243 - 0xf3
      11'h44D: dout <= 8'b11110011; // 1101 : 243 - 0xf3
      11'h44E: dout <= 8'b11111111; // 1102 : 255 - 0xff
      11'h44F: dout <= 8'b11111111; // 1103 : 255 - 0xff
      11'h450: dout <= 8'b10111111; // 1104 : 191 - 0xbf -- Sprite 0x8a
      11'h451: dout <= 8'b11110111; // 1105 : 247 - 0xf7
      11'h452: dout <= 8'b11111101; // 1106 : 253 - 0xfd
      11'h453: dout <= 8'b11111111; // 1107 : 255 - 0xff
      11'h454: dout <= 8'b11111011; // 1108 : 251 - 0xfb
      11'h455: dout <= 8'b10111111; // 1109 : 191 - 0xbf
      11'h456: dout <= 8'b11111110; // 1110 : 254 - 0xfe
      11'h457: dout <= 8'b11101111; // 1111 : 239 - 0xef
      11'h458: dout <= 8'b10111111; // 1112 : 191 - 0xbf -- Sprite 0x8b
      11'h459: dout <= 8'b11111111; // 1113 : 255 - 0xff
      11'h45A: dout <= 8'b11101110; // 1114 : 238 - 0xee
      11'h45B: dout <= 8'b11111111; // 1115 : 255 - 0xff
      11'h45C: dout <= 8'b11011111; // 1116 : 223 - 0xdf
      11'h45D: dout <= 8'b01111101; // 1117 : 125 - 0x7d
      11'h45E: dout <= 8'b11111111; // 1118 : 255 - 0xff
      11'h45F: dout <= 8'b11011111; // 1119 : 223 - 0xdf
      11'h460: dout <= 8'b11111111; // 1120 : 255 - 0xff -- Sprite 0x8c
      11'h461: dout <= 8'b11111000; // 1121 : 248 - 0xf8
      11'h462: dout <= 8'b11100010; // 1122 : 226 - 0xe2
      11'h463: dout <= 8'b11010111; // 1123 : 215 - 0xd7
      11'h464: dout <= 8'b11001111; // 1124 : 207 - 0xcf
      11'h465: dout <= 8'b10011111; // 1125 : 159 - 0x9f
      11'h466: dout <= 8'b10111110; // 1126 : 190 - 0xbe
      11'h467: dout <= 8'b10011101; // 1127 : 157 - 0x9d
      11'h468: dout <= 8'b11111111; // 1128 : 255 - 0xff -- Sprite 0x8d
      11'h469: dout <= 8'b00011111; // 1129 :  31 - 0x1f
      11'h46A: dout <= 8'b10100111; // 1130 : 167 - 0xa7
      11'h46B: dout <= 8'b11000011; // 1131 : 195 - 0xc3
      11'h46C: dout <= 8'b11100011; // 1132 : 227 - 0xe3
      11'h46D: dout <= 8'b01000001; // 1133 :  65 - 0x41
      11'h46E: dout <= 8'b10100001; // 1134 : 161 - 0xa1
      11'h46F: dout <= 8'b00000001; // 1135 :   1 - 0x1
      11'h470: dout <= 8'b10111110; // 1136 : 190 - 0xbe -- Sprite 0x8e
      11'h471: dout <= 8'b11111111; // 1137 : 255 - 0xff
      11'h472: dout <= 8'b11011111; // 1138 : 223 - 0xdf
      11'h473: dout <= 8'b11111111; // 1139 : 255 - 0xff
      11'h474: dout <= 8'b11101111; // 1140 : 239 - 0xef
      11'h475: dout <= 8'b11111111; // 1141 : 255 - 0xff
      11'h476: dout <= 8'b11110111; // 1142 : 247 - 0xf7
      11'h477: dout <= 8'b11111111; // 1143 : 255 - 0xff
      11'h478: dout <= 8'b01111101; // 1144 : 125 - 0x7d -- Sprite 0x8f
      11'h479: dout <= 8'b11111111; // 1145 : 255 - 0xff
      11'h47A: dout <= 8'b11111011; // 1146 : 251 - 0xfb
      11'h47B: dout <= 8'b11111111; // 1147 : 255 - 0xff
      11'h47C: dout <= 8'b11110111; // 1148 : 247 - 0xf7
      11'h47D: dout <= 8'b11111111; // 1149 : 255 - 0xff
      11'h47E: dout <= 8'b11101111; // 1150 : 239 - 0xef
      11'h47F: dout <= 8'b11111111; // 1151 : 255 - 0xff
      11'h480: dout <= 8'b10111110; // 1152 : 190 - 0xbe -- Sprite 0x90
      11'h481: dout <= 8'b11110111; // 1153 : 247 - 0xf7
      11'h482: dout <= 8'b11111111; // 1154 : 255 - 0xff
      11'h483: dout <= 8'b11011111; // 1155 : 223 - 0xdf
      11'h484: dout <= 8'b11111011; // 1156 : 251 - 0xfb
      11'h485: dout <= 8'b11111110; // 1157 : 254 - 0xfe
      11'h486: dout <= 8'b10111111; // 1158 : 191 - 0xbf
      11'h487: dout <= 8'b11110111; // 1159 : 247 - 0xf7
      11'h488: dout <= 8'b11101110; // 1160 : 238 - 0xee -- Sprite 0x91
      11'h489: dout <= 8'b11111111; // 1161 : 255 - 0xff
      11'h48A: dout <= 8'b01111011; // 1162 : 123 - 0x7b
      11'h48B: dout <= 8'b11111101; // 1163 : 253 - 0xfd
      11'h48C: dout <= 8'b11101111; // 1164 : 239 - 0xef
      11'h48D: dout <= 8'b11111111; // 1165 : 255 - 0xff
      11'h48E: dout <= 8'b10111101; // 1166 : 189 - 0xbd
      11'h48F: dout <= 8'b11111111; // 1167 : 255 - 0xff
      11'h490: dout <= 8'b11111011; // 1168 : 251 - 0xfb -- Sprite 0x92
      11'h491: dout <= 8'b10111111; // 1169 : 191 - 0xbf
      11'h492: dout <= 8'b11101111; // 1170 : 239 - 0xef
      11'h493: dout <= 8'b11111101; // 1171 : 253 - 0xfd
      11'h494: dout <= 8'b11111111; // 1172 : 255 - 0xff
      11'h495: dout <= 8'b10111111; // 1173 : 191 - 0xbf
      11'h496: dout <= 8'b11111011; // 1174 : 251 - 0xfb
      11'h497: dout <= 8'b11011111; // 1175 : 223 - 0xdf
      11'h498: dout <= 8'b10111101; // 1176 : 189 - 0xbd -- Sprite 0x93
      11'h499: dout <= 8'b11111111; // 1177 : 255 - 0xff
      11'h49A: dout <= 8'b01110111; // 1178 : 119 - 0x77
      11'h49B: dout <= 8'b11111110; // 1179 : 254 - 0xfe
      11'h49C: dout <= 8'b11011111; // 1180 : 223 - 0xdf
      11'h49D: dout <= 8'b11111011; // 1181 : 251 - 0xfb
      11'h49E: dout <= 8'b11101111; // 1182 : 239 - 0xef
      11'h49F: dout <= 8'b01111111; // 1183 : 127 - 0x7f
      11'h4A0: dout <= 8'b01111111; // 1184 : 127 - 0x7f -- Sprite 0x94
      11'h4A1: dout <= 8'b11110111; // 1185 : 247 - 0xf7
      11'h4A2: dout <= 8'b11011101; // 1186 : 221 - 0xdd
      11'h4A3: dout <= 8'b01111011; // 1187 : 123 - 0x7b
      11'h4A4: dout <= 8'b11111111; // 1188 : 255 - 0xff
      11'h4A5: dout <= 8'b11101110; // 1189 : 238 - 0xee
      11'h4A6: dout <= 8'b10111011; // 1190 : 187 - 0xbb
      11'h4A7: dout <= 8'b11111101; // 1191 : 253 - 0xfd
      11'h4A8: dout <= 8'b11010111; // 1192 : 215 - 0xd7 -- Sprite 0x95
      11'h4A9: dout <= 8'b01111111; // 1193 : 127 - 0x7f
      11'h4AA: dout <= 8'b11111101; // 1194 : 253 - 0xfd
      11'h4AB: dout <= 8'b11101110; // 1195 : 238 - 0xee
      11'h4AC: dout <= 8'b11110111; // 1196 : 247 - 0xf7
      11'h4AD: dout <= 8'b10111011; // 1197 : 187 - 0xbb
      11'h4AE: dout <= 8'b11101111; // 1198 : 239 - 0xef
      11'h4AF: dout <= 8'b11110111; // 1199 : 247 - 0xf7
      11'h4B0: dout <= 8'b10111111; // 1200 : 191 - 0xbf -- Sprite 0x96
      11'h4B1: dout <= 8'b11101110; // 1201 : 238 - 0xee
      11'h4B2: dout <= 8'b11011011; // 1202 : 219 - 0xdb
      11'h4B3: dout <= 8'b11111111; // 1203 : 255 - 0xff
      11'h4B4: dout <= 8'b01110111; // 1204 : 119 - 0x77
      11'h4B5: dout <= 8'b11011101; // 1205 : 221 - 0xdd
      11'h4B6: dout <= 8'b11101111; // 1206 : 239 - 0xef
      11'h4B7: dout <= 8'b11111011; // 1207 : 251 - 0xfb
      11'h4B8: dout <= 8'b11111101; // 1208 : 253 - 0xfd -- Sprite 0x97
      11'h4B9: dout <= 8'b11101110; // 1209 : 238 - 0xee
      11'h4BA: dout <= 8'b11111011; // 1210 : 251 - 0xfb
      11'h4BB: dout <= 8'b11111101; // 1211 : 253 - 0xfd
      11'h4BC: dout <= 8'b11110101; // 1212 : 245 - 0xf5
      11'h4BD: dout <= 8'b11011111; // 1213 : 223 - 0xdf
      11'h4BE: dout <= 8'b01111111; // 1214 : 127 - 0x7f
      11'h4BF: dout <= 8'b10111011; // 1215 : 187 - 0xbb
      11'h4C0: dout <= 8'b11111111; // 1216 : 255 - 0xff -- Sprite 0x98
      11'h4C1: dout <= 8'b11001111; // 1217 : 207 - 0xcf
      11'h4C2: dout <= 8'b11011111; // 1218 : 223 - 0xdf
      11'h4C3: dout <= 8'b11111111; // 1219 : 255 - 0xff
      11'h4C4: dout <= 8'b11110011; // 1220 : 243 - 0xf3
      11'h4C5: dout <= 8'b11110011; // 1221 : 243 - 0xf3
      11'h4C6: dout <= 8'b11111111; // 1222 : 255 - 0xff
      11'h4C7: dout <= 8'b11111111; // 1223 : 255 - 0xff
      11'h4C8: dout <= 8'b11111111; // 1224 : 255 - 0xff -- Sprite 0x99
      11'h4C9: dout <= 8'b11111111; // 1225 : 255 - 0xff
      11'h4CA: dout <= 8'b10011111; // 1226 : 159 - 0x9f
      11'h4CB: dout <= 8'b10110011; // 1227 : 179 - 0xb3
      11'h4CC: dout <= 8'b11110011; // 1228 : 243 - 0xf3
      11'h4CD: dout <= 8'b11111111; // 1229 : 255 - 0xff
      11'h4CE: dout <= 8'b11111111; // 1230 : 255 - 0xff
      11'h4CF: dout <= 8'b11111111; // 1231 : 255 - 0xff
      11'h4D0: dout <= 8'b10111111; // 1232 : 191 - 0xbf -- Sprite 0x9a
      11'h4D1: dout <= 8'b11110111; // 1233 : 247 - 0xf7
      11'h4D2: dout <= 8'b11111111; // 1234 : 255 - 0xff
      11'h4D3: dout <= 8'b11011111; // 1235 : 223 - 0xdf
      11'h4D4: dout <= 8'b11111011; // 1236 : 251 - 0xfb
      11'h4D5: dout <= 8'b11111111; // 1237 : 255 - 0xff
      11'h4D6: dout <= 8'b10111111; // 1238 : 191 - 0xbf
      11'h4D7: dout <= 8'b11110111; // 1239 : 247 - 0xf7
      11'h4D8: dout <= 8'b11011111; // 1240 : 223 - 0xdf -- Sprite 0x9b
      11'h4D9: dout <= 8'b11111111; // 1241 : 255 - 0xff
      11'h4DA: dout <= 8'b01111011; // 1242 : 123 - 0x7b
      11'h4DB: dout <= 8'b11111111; // 1243 : 255 - 0xff
      11'h4DC: dout <= 8'b11101111; // 1244 : 239 - 0xef
      11'h4DD: dout <= 8'b11111101; // 1245 : 253 - 0xfd
      11'h4DE: dout <= 8'b10111111; // 1246 : 191 - 0xbf
      11'h4DF: dout <= 8'b11111111; // 1247 : 255 - 0xff
      11'h4E0: dout <= 8'b10111010; // 1248 : 186 - 0xba -- Sprite 0x9c
      11'h4E1: dout <= 8'b10011100; // 1249 : 156 - 0x9c
      11'h4E2: dout <= 8'b10101010; // 1250 : 170 - 0xaa
      11'h4E3: dout <= 8'b11000000; // 1251 : 192 - 0xc0
      11'h4E4: dout <= 8'b11000000; // 1252 : 192 - 0xc0
      11'h4E5: dout <= 8'b11100000; // 1253 : 224 - 0xe0
      11'h4E6: dout <= 8'b11111000; // 1254 : 248 - 0xf8
      11'h4E7: dout <= 8'b11111111; // 1255 : 255 - 0xff
      11'h4E8: dout <= 8'b00000001; // 1256 :   1 - 0x1 -- Sprite 0x9d
      11'h4E9: dout <= 8'b00000001; // 1257 :   1 - 0x1
      11'h4EA: dout <= 8'b00000001; // 1258 :   1 - 0x1
      11'h4EB: dout <= 8'b00000011; // 1259 :   3 - 0x3
      11'h4EC: dout <= 8'b00000011; // 1260 :   3 - 0x3
      11'h4ED: dout <= 8'b00000111; // 1261 :   7 - 0x7
      11'h4EE: dout <= 8'b00011111; // 1262 :  31 - 0x1f
      11'h4EF: dout <= 8'b11111111; // 1263 : 255 - 0xff
      11'h4F0: dout <= 8'b01111101; // 1264 : 125 - 0x7d -- Sprite 0x9e
      11'h4F1: dout <= 8'b11111111; // 1265 : 255 - 0xff
      11'h4F2: dout <= 8'b11111011; // 1266 : 251 - 0xfb
      11'h4F3: dout <= 8'b11111111; // 1267 : 255 - 0xff
      11'h4F4: dout <= 8'b11111111; // 1268 : 255 - 0xff
      11'h4F5: dout <= 8'b11111011; // 1269 : 251 - 0xfb
      11'h4F6: dout <= 8'b11111111; // 1270 : 255 - 0xff
      11'h4F7: dout <= 8'b01111101; // 1271 : 125 - 0x7d
      11'h4F8: dout <= 8'b11111111; // 1272 : 255 - 0xff -- Sprite 0x9f
      11'h4F9: dout <= 8'b11111111; // 1273 : 255 - 0xff
      11'h4FA: dout <= 8'b10111101; // 1274 : 189 - 0xbd
      11'h4FB: dout <= 8'b11111111; // 1275 : 255 - 0xff
      11'h4FC: dout <= 8'b11111111; // 1276 : 255 - 0xff
      11'h4FD: dout <= 8'b11111111; // 1277 : 255 - 0xff
      11'h4FE: dout <= 8'b11111111; // 1278 : 255 - 0xff
      11'h4FF: dout <= 8'b10111101; // 1279 : 189 - 0xbd
      11'h500: dout <= 8'b11101111; // 1280 : 239 - 0xef -- Sprite 0xa0
      11'h501: dout <= 8'b11000111; // 1281 : 199 - 0xc7
      11'h502: dout <= 8'b10000011; // 1282 : 131 - 0x83
      11'h503: dout <= 8'b00000111; // 1283 :   7 - 0x7
      11'h504: dout <= 8'b10001111; // 1284 : 143 - 0x8f
      11'h505: dout <= 8'b11011101; // 1285 : 221 - 0xdd
      11'h506: dout <= 8'b11111010; // 1286 : 250 - 0xfa
      11'h507: dout <= 8'b11111101; // 1287 : 253 - 0xfd
      11'h508: dout <= 8'b11101111; // 1288 : 239 - 0xef -- Sprite 0xa1
      11'h509: dout <= 8'b11000111; // 1289 : 199 - 0xc7
      11'h50A: dout <= 8'b10000011; // 1290 : 131 - 0x83
      11'h50B: dout <= 8'b00011111; // 1291 :  31 - 0x1f
      11'h50C: dout <= 8'b10010000; // 1292 : 144 - 0x90
      11'h50D: dout <= 8'b11010100; // 1293 : 212 - 0xd4
      11'h50E: dout <= 8'b11110011; // 1294 : 243 - 0xf3
      11'h50F: dout <= 8'b11110010; // 1295 : 242 - 0xf2
      11'h510: dout <= 8'b11101111; // 1296 : 239 - 0xef -- Sprite 0xa2
      11'h511: dout <= 8'b11000111; // 1297 : 199 - 0xc7
      11'h512: dout <= 8'b10000011; // 1298 : 131 - 0x83
      11'h513: dout <= 8'b11111111; // 1299 : 255 - 0xff
      11'h514: dout <= 8'b00000000; // 1300 :   0 - 0x0
      11'h515: dout <= 8'b00000000; // 1301 :   0 - 0x0
      11'h516: dout <= 8'b01010101; // 1302 :  85 - 0x55
      11'h517: dout <= 8'b00000000; // 1303 :   0 - 0x0
      11'h518: dout <= 8'b11110000; // 1304 : 240 - 0xf0 -- Sprite 0xa3
      11'h519: dout <= 8'b11010010; // 1305 : 210 - 0xd2
      11'h51A: dout <= 8'b10010000; // 1306 : 144 - 0x90
      11'h51B: dout <= 8'b00010010; // 1307 :  18 - 0x12
      11'h51C: dout <= 8'b10010000; // 1308 : 144 - 0x90
      11'h51D: dout <= 8'b11010010; // 1309 : 210 - 0xd2
      11'h51E: dout <= 8'b11110000; // 1310 : 240 - 0xf0
      11'h51F: dout <= 8'b11110010; // 1311 : 242 - 0xf2
      11'h520: dout <= 8'b11110000; // 1312 : 240 - 0xf0 -- Sprite 0xa4
      11'h521: dout <= 8'b11010011; // 1313 : 211 - 0xd3
      11'h522: dout <= 8'b10010100; // 1314 : 148 - 0x94
      11'h523: dout <= 8'b00011000; // 1315 :  24 - 0x18
      11'h524: dout <= 8'b10011111; // 1316 : 159 - 0x9f
      11'h525: dout <= 8'b11011101; // 1317 : 221 - 0xdd
      11'h526: dout <= 8'b11111010; // 1318 : 250 - 0xfa
      11'h527: dout <= 8'b11111101; // 1319 : 253 - 0xfd
      11'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0 -- Sprite 0xa5
      11'h529: dout <= 8'b11111111; // 1321 : 255 - 0xff
      11'h52A: dout <= 8'b00000000; // 1322 :   0 - 0x0
      11'h52B: dout <= 8'b00000000; // 1323 :   0 - 0x0
      11'h52C: dout <= 8'b11111111; // 1324 : 255 - 0xff
      11'h52D: dout <= 8'b11011101; // 1325 : 221 - 0xdd
      11'h52E: dout <= 8'b11111010; // 1326 : 250 - 0xfa
      11'h52F: dout <= 8'b11111101; // 1327 : 253 - 0xfd
      11'h530: dout <= 8'b11101111; // 1328 : 239 - 0xef -- Sprite 0xa6
      11'h531: dout <= 8'b11000111; // 1329 : 199 - 0xc7
      11'h532: dout <= 8'b10000011; // 1330 : 131 - 0x83
      11'h533: dout <= 8'b11111111; // 1331 : 255 - 0xff
      11'h534: dout <= 8'b00011111; // 1332 :  31 - 0x1f
      11'h535: dout <= 8'b00101101; // 1333 :  45 - 0x2d
      11'h536: dout <= 8'b01001010; // 1334 :  74 - 0x4a
      11'h537: dout <= 8'b01001101; // 1335 :  77 - 0x4d
      11'h538: dout <= 8'b01001111; // 1336 :  79 - 0x4f -- Sprite 0xa7
      11'h539: dout <= 8'b01001111; // 1337 :  79 - 0x4f
      11'h53A: dout <= 8'b01001011; // 1338 :  75 - 0x4b
      11'h53B: dout <= 8'b01001111; // 1339 :  79 - 0x4f
      11'h53C: dout <= 8'b01001111; // 1340 :  79 - 0x4f
      11'h53D: dout <= 8'b01001101; // 1341 :  77 - 0x4d
      11'h53E: dout <= 8'b01001010; // 1342 :  74 - 0x4a
      11'h53F: dout <= 8'b01001101; // 1343 :  77 - 0x4d
      11'h540: dout <= 8'b01001111; // 1344 :  79 - 0x4f -- Sprite 0xa8
      11'h541: dout <= 8'b11001111; // 1345 : 207 - 0xcf
      11'h542: dout <= 8'b00001011; // 1346 :  11 - 0xb
      11'h543: dout <= 8'b00001111; // 1347 :  15 - 0xf
      11'h544: dout <= 8'b11111111; // 1348 : 255 - 0xff
      11'h545: dout <= 8'b11011101; // 1349 : 221 - 0xdd
      11'h546: dout <= 8'b11111010; // 1350 : 250 - 0xfa
      11'h547: dout <= 8'b11111101; // 1351 : 253 - 0xfd
      11'h548: dout <= 8'b11111111; // 1352 : 255 - 0xff -- Sprite 0xa9
      11'h549: dout <= 8'b11111111; // 1353 : 255 - 0xff
      11'h54A: dout <= 8'b11111111; // 1354 : 255 - 0xff
      11'h54B: dout <= 8'b11111111; // 1355 : 255 - 0xff
      11'h54C: dout <= 8'b11111111; // 1356 : 255 - 0xff
      11'h54D: dout <= 8'b11111111; // 1357 : 255 - 0xff
      11'h54E: dout <= 8'b11111111; // 1358 : 255 - 0xff
      11'h54F: dout <= 8'b11111111; // 1359 : 255 - 0xff
      11'h550: dout <= 8'b11111111; // 1360 : 255 - 0xff -- Sprite 0xaa
      11'h551: dout <= 8'b11111111; // 1361 : 255 - 0xff
      11'h552: dout <= 8'b10101111; // 1362 : 175 - 0xaf
      11'h553: dout <= 8'b01010111; // 1363 :  87 - 0x57
      11'h554: dout <= 8'b10001111; // 1364 : 143 - 0x8f
      11'h555: dout <= 8'b11011101; // 1365 : 221 - 0xdd
      11'h556: dout <= 8'b11111010; // 1366 : 250 - 0xfa
      11'h557: dout <= 8'b11111101; // 1367 : 253 - 0xfd
      11'h558: dout <= 8'b11111111; // 1368 : 255 - 0xff -- Sprite 0xab
      11'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      11'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      11'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      11'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      11'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      11'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      11'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      11'h560: dout <= 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      11'h561: dout <= 8'b00000000; // 1377 :   0 - 0x0
      11'h562: dout <= 8'b00000000; // 1378 :   0 - 0x0
      11'h563: dout <= 8'b00000000; // 1379 :   0 - 0x0
      11'h564: dout <= 8'b00000000; // 1380 :   0 - 0x0
      11'h565: dout <= 8'b00000000; // 1381 :   0 - 0x0
      11'h566: dout <= 8'b00000000; // 1382 :   0 - 0x0
      11'h567: dout <= 8'b00000000; // 1383 :   0 - 0x0
      11'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0 -- Sprite 0xad
      11'h569: dout <= 8'b11111111; // 1385 : 255 - 0xff
      11'h56A: dout <= 8'b00000000; // 1386 :   0 - 0x0
      11'h56B: dout <= 8'b11111111; // 1387 : 255 - 0xff
      11'h56C: dout <= 8'b11111111; // 1388 : 255 - 0xff
      11'h56D: dout <= 8'b11111111; // 1389 : 255 - 0xff
      11'h56E: dout <= 8'b11111111; // 1390 : 255 - 0xff
      11'h56F: dout <= 8'b11111111; // 1391 : 255 - 0xff
      11'h570: dout <= 8'b11111111; // 1392 : 255 - 0xff -- Sprite 0xae
      11'h571: dout <= 8'b11111111; // 1393 : 255 - 0xff
      11'h572: dout <= 8'b11111111; // 1394 : 255 - 0xff
      11'h573: dout <= 8'b11111111; // 1395 : 255 - 0xff
      11'h574: dout <= 8'b11111111; // 1396 : 255 - 0xff
      11'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      11'h576: dout <= 8'b11111111; // 1398 : 255 - 0xff
      11'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      11'h578: dout <= 8'b11111111; // 1400 : 255 - 0xff -- Sprite 0xaf
      11'h579: dout <= 8'b11111111; // 1401 : 255 - 0xff
      11'h57A: dout <= 8'b11111111; // 1402 : 255 - 0xff
      11'h57B: dout <= 8'b11111111; // 1403 : 255 - 0xff
      11'h57C: dout <= 8'b11111111; // 1404 : 255 - 0xff
      11'h57D: dout <= 8'b11111111; // 1405 : 255 - 0xff
      11'h57E: dout <= 8'b11111111; // 1406 : 255 - 0xff
      11'h57F: dout <= 8'b11111111; // 1407 : 255 - 0xff
      11'h580: dout <= 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      11'h581: dout <= 8'b00011111; // 1409 :  31 - 0x1f
      11'h582: dout <= 8'b00010000; // 1410 :  16 - 0x10
      11'h583: dout <= 8'b00010000; // 1411 :  16 - 0x10
      11'h584: dout <= 8'b00010000; // 1412 :  16 - 0x10
      11'h585: dout <= 8'b00010000; // 1413 :  16 - 0x10
      11'h586: dout <= 8'b00010000; // 1414 :  16 - 0x10
      11'h587: dout <= 8'b00010000; // 1415 :  16 - 0x10
      11'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0 -- Sprite 0xb1
      11'h589: dout <= 8'b11111000; // 1417 : 248 - 0xf8
      11'h58A: dout <= 8'b00001000; // 1418 :   8 - 0x8
      11'h58B: dout <= 8'b00001000; // 1419 :   8 - 0x8
      11'h58C: dout <= 8'b00001000; // 1420 :   8 - 0x8
      11'h58D: dout <= 8'b00001000; // 1421 :   8 - 0x8
      11'h58E: dout <= 8'b00001000; // 1422 :   8 - 0x8
      11'h58F: dout <= 8'b00001000; // 1423 :   8 - 0x8
      11'h590: dout <= 8'b00010000; // 1424 :  16 - 0x10 -- Sprite 0xb2
      11'h591: dout <= 8'b00010000; // 1425 :  16 - 0x10
      11'h592: dout <= 8'b00010000; // 1426 :  16 - 0x10
      11'h593: dout <= 8'b00010000; // 1427 :  16 - 0x10
      11'h594: dout <= 8'b00011111; // 1428 :  31 - 0x1f
      11'h595: dout <= 8'b00011111; // 1429 :  31 - 0x1f
      11'h596: dout <= 8'b00001111; // 1430 :  15 - 0xf
      11'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      11'h598: dout <= 8'b00001000; // 1432 :   8 - 0x8 -- Sprite 0xb3
      11'h599: dout <= 8'b00001000; // 1433 :   8 - 0x8
      11'h59A: dout <= 8'b00001000; // 1434 :   8 - 0x8
      11'h59B: dout <= 8'b00001000; // 1435 :   8 - 0x8
      11'h59C: dout <= 8'b11111000; // 1436 : 248 - 0xf8
      11'h59D: dout <= 8'b11111000; // 1437 : 248 - 0xf8
      11'h59E: dout <= 8'b11110000; // 1438 : 240 - 0xf0
      11'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      11'h5A0: dout <= 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0xb4
      11'h5A1: dout <= 8'b00000000; // 1441 :   0 - 0x0
      11'h5A2: dout <= 8'b00111111; // 1442 :  63 - 0x3f
      11'h5A3: dout <= 8'b01100000; // 1443 :  96 - 0x60
      11'h5A4: dout <= 8'b01100000; // 1444 :  96 - 0x60
      11'h5A5: dout <= 8'b01100000; // 1445 :  96 - 0x60
      11'h5A6: dout <= 8'b01100000; // 1446 :  96 - 0x60
      11'h5A7: dout <= 8'b01100000; // 1447 :  96 - 0x60
      11'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0 -- Sprite 0xb5
      11'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      11'h5AA: dout <= 8'b11111100; // 1450 : 252 - 0xfc
      11'h5AB: dout <= 8'b00000110; // 1451 :   6 - 0x6
      11'h5AC: dout <= 8'b00000110; // 1452 :   6 - 0x6
      11'h5AD: dout <= 8'b00000110; // 1453 :   6 - 0x6
      11'h5AE: dout <= 8'b00000110; // 1454 :   6 - 0x6
      11'h5AF: dout <= 8'b00000110; // 1455 :   6 - 0x6
      11'h5B0: dout <= 8'b01100000; // 1456 :  96 - 0x60 -- Sprite 0xb6
      11'h5B1: dout <= 8'b01100000; // 1457 :  96 - 0x60
      11'h5B2: dout <= 8'b01100000; // 1458 :  96 - 0x60
      11'h5B3: dout <= 8'b01111111; // 1459 : 127 - 0x7f
      11'h5B4: dout <= 8'b01111111; // 1460 : 127 - 0x7f
      11'h5B5: dout <= 8'b00111111; // 1461 :  63 - 0x3f
      11'h5B6: dout <= 8'b00000000; // 1462 :   0 - 0x0
      11'h5B7: dout <= 8'b00000000; // 1463 :   0 - 0x0
      11'h5B8: dout <= 8'b00000110; // 1464 :   6 - 0x6 -- Sprite 0xb7
      11'h5B9: dout <= 8'b00000110; // 1465 :   6 - 0x6
      11'h5BA: dout <= 8'b00000110; // 1466 :   6 - 0x6
      11'h5BB: dout <= 8'b11111110; // 1467 : 254 - 0xfe
      11'h5BC: dout <= 8'b11111110; // 1468 : 254 - 0xfe
      11'h5BD: dout <= 8'b11111100; // 1469 : 252 - 0xfc
      11'h5BE: dout <= 8'b00000000; // 1470 :   0 - 0x0
      11'h5BF: dout <= 8'b00000000; // 1471 :   0 - 0x0
      11'h5C0: dout <= 8'b01100000; // 1472 :  96 - 0x60 -- Sprite 0xb8
      11'h5C1: dout <= 8'b11110011; // 1473 : 243 - 0xf3
      11'h5C2: dout <= 8'b11000111; // 1474 : 199 - 0xc7
      11'h5C3: dout <= 8'b10000110; // 1475 : 134 - 0x86
      11'h5C4: dout <= 8'b00000100; // 1476 :   4 - 0x4
      11'h5C5: dout <= 8'b00000100; // 1477 :   4 - 0x4
      11'h5C6: dout <= 8'b00000111; // 1478 :   7 - 0x7
      11'h5C7: dout <= 8'b00000111; // 1479 :   7 - 0x7
      11'h5C8: dout <= 8'b00000110; // 1480 :   6 - 0x6 -- Sprite 0xb9
      11'h5C9: dout <= 8'b10001111; // 1481 : 143 - 0x8f
      11'h5CA: dout <= 8'b11000101; // 1482 : 197 - 0xc5
      11'h5CB: dout <= 8'b00100011; // 1483 :  35 - 0x23
      11'h5CC: dout <= 8'b00101110; // 1484 :  46 - 0x2e
      11'h5CD: dout <= 8'b01100000; // 1485 :  96 - 0x60
      11'h5CE: dout <= 8'b11100001; // 1486 : 225 - 0xe1
      11'h5CF: dout <= 8'b11100001; // 1487 : 225 - 0xe1
      11'h5D0: dout <= 8'b11001000; // 1488 : 200 - 0xc8 -- Sprite 0xba
      11'h5D1: dout <= 8'b11111000; // 1489 : 248 - 0xf8
      11'h5D2: dout <= 8'b10110000; // 1490 : 176 - 0xb0
      11'h5D3: dout <= 8'b00010000; // 1491 :  16 - 0x10
      11'h5D4: dout <= 8'b00110000; // 1492 :  48 - 0x30
      11'h5D5: dout <= 8'b11001000; // 1493 : 200 - 0xc8
      11'h5D6: dout <= 8'b11111000; // 1494 : 248 - 0xf8
      11'h5D7: dout <= 8'b10000000; // 1495 : 128 - 0x80
      11'h5D8: dout <= 8'b00000011; // 1496 :   3 - 0x3 -- Sprite 0xbb
      11'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      11'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      11'h5DB: dout <= 8'b01100000; // 1499 :  96 - 0x60
      11'h5DC: dout <= 8'b11110000; // 1500 : 240 - 0xf0
      11'h5DD: dout <= 8'b11010000; // 1501 : 208 - 0xd0
      11'h5DE: dout <= 8'b10010000; // 1502 : 144 - 0x90
      11'h5DF: dout <= 8'b01100000; // 1503 :  96 - 0x60
      11'h5E0: dout <= 8'b11000011; // 1504 : 195 - 0xc3 -- Sprite 0xbc
      11'h5E1: dout <= 8'b00001110; // 1505 :  14 - 0xe
      11'h5E2: dout <= 8'b00000000; // 1506 :   0 - 0x0
      11'h5E3: dout <= 8'b00000110; // 1507 :   6 - 0x6
      11'h5E4: dout <= 8'b00001111; // 1508 :  15 - 0xf
      11'h5E5: dout <= 8'b00001101; // 1509 :  13 - 0xd
      11'h5E6: dout <= 8'b00001001; // 1510 :   9 - 0x9
      11'h5E7: dout <= 8'b00000110; // 1511 :   6 - 0x6
      11'h5E8: dout <= 8'b11100000; // 1512 : 224 - 0xe0 -- Sprite 0xbd
      11'h5E9: dout <= 8'b01100011; // 1513 :  99 - 0x63
      11'h5EA: dout <= 8'b11100111; // 1514 : 231 - 0xe7
      11'h5EB: dout <= 8'b11100110; // 1515 : 230 - 0xe6
      11'h5EC: dout <= 8'b00000100; // 1516 :   4 - 0x4
      11'h5ED: dout <= 8'b00000100; // 1517 :   4 - 0x4
      11'h5EE: dout <= 8'b00000111; // 1518 :   7 - 0x7
      11'h5EF: dout <= 8'b00000111; // 1519 :   7 - 0x7
      11'h5F0: dout <= 8'b00000111; // 1520 :   7 - 0x7 -- Sprite 0xbe
      11'h5F1: dout <= 8'b10000011; // 1521 : 131 - 0x83
      11'h5F2: dout <= 8'b11000111; // 1522 : 199 - 0xc7
      11'h5F3: dout <= 8'b00100111; // 1523 :  39 - 0x27
      11'h5F4: dout <= 8'b00100000; // 1524 :  32 - 0x20
      11'h5F5: dout <= 8'b01100000; // 1525 :  96 - 0x60
      11'h5F6: dout <= 8'b11100000; // 1526 : 224 - 0xe0
      11'h5F7: dout <= 8'b11100000; // 1527 : 224 - 0xe0
      11'h5F8: dout <= 8'b00000011; // 1528 :   3 - 0x3 -- Sprite 0xbf
      11'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      11'h5FA: dout <= 8'b00001100; // 1530 :  12 - 0xc
      11'h5FB: dout <= 8'b00001100; // 1531 :  12 - 0xc
      11'h5FC: dout <= 8'b11100100; // 1532 : 228 - 0xe4
      11'h5FD: dout <= 8'b01101100; // 1533 : 108 - 0x6c
      11'h5FE: dout <= 8'b11101101; // 1534 : 237 - 0xed
      11'h5FF: dout <= 8'b11100111; // 1535 : 231 - 0xe7
      11'h600: dout <= 8'b11000000; // 1536 : 192 - 0xc0 -- Sprite 0xc0
      11'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      11'h602: dout <= 8'b00110000; // 1538 :  48 - 0x30
      11'h603: dout <= 8'b00110000; // 1539 :  48 - 0x30
      11'h604: dout <= 8'b00010111; // 1540 :  23 - 0x17
      11'h605: dout <= 8'b00110011; // 1541 :  51 - 0x33
      11'h606: dout <= 8'b01110111; // 1542 : 119 - 0x77
      11'h607: dout <= 8'b11010111; // 1543 : 215 - 0xd7
      11'h608: dout <= 8'b00001100; // 1544 :  12 - 0xc -- Sprite 0xc1
      11'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      11'h60A: dout <= 8'b00000000; // 1546 :   0 - 0x0
      11'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      11'h60C: dout <= 8'b00000000; // 1548 :   0 - 0x0
      11'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      11'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      11'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout <= 8'b00110000; // 1552 :  48 - 0x30 -- Sprite 0xc2
      11'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      11'h612: dout <= 8'b00000000; // 1554 :   0 - 0x0
      11'h613: dout <= 8'b00000000; // 1555 :   0 - 0x0
      11'h614: dout <= 8'b00000000; // 1556 :   0 - 0x0
      11'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      11'h616: dout <= 8'b00000000; // 1558 :   0 - 0x0
      11'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      11'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0 -- Sprite 0xc3
      11'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      11'h61A: dout <= 8'b00000100; // 1562 :   4 - 0x4
      11'h61B: dout <= 8'b00001101; // 1563 :  13 - 0xd
      11'h61C: dout <= 8'b00001111; // 1564 :  15 - 0xf
      11'h61D: dout <= 8'b00001100; // 1565 :  12 - 0xc
      11'h61E: dout <= 8'b00001100; // 1566 :  12 - 0xc
      11'h61F: dout <= 8'b00000100; // 1567 :   4 - 0x4
      11'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      11'h621: dout <= 8'b00000000; // 1569 :   0 - 0x0
      11'h622: dout <= 8'b00010000; // 1570 :  16 - 0x10
      11'h623: dout <= 8'b01110000; // 1571 : 112 - 0x70
      11'h624: dout <= 8'b11110000; // 1572 : 240 - 0xf0
      11'h625: dout <= 8'b00110000; // 1573 :  48 - 0x30
      11'h626: dout <= 8'b00110000; // 1574 :  48 - 0x30
      11'h627: dout <= 8'b00010000; // 1575 :  16 - 0x10
      11'h628: dout <= 8'b11100100; // 1576 : 228 - 0xe4 -- Sprite 0xc5
      11'h629: dout <= 8'b00100100; // 1577 :  36 - 0x24
      11'h62A: dout <= 8'b11101111; // 1578 : 239 - 0xef
      11'h62B: dout <= 8'b11100111; // 1579 : 231 - 0xe7
      11'h62C: dout <= 8'b00000110; // 1580 :   6 - 0x6
      11'h62D: dout <= 8'b00000100; // 1581 :   4 - 0x4
      11'h62E: dout <= 8'b00000100; // 1582 :   4 - 0x4
      11'h62F: dout <= 8'b00000111; // 1583 :   7 - 0x7
      11'h630: dout <= 8'b00010111; // 1584 :  23 - 0x17 -- Sprite 0xc6
      11'h631: dout <= 8'b00010001; // 1585 :  17 - 0x11
      11'h632: dout <= 8'b10110111; // 1586 : 183 - 0xb7
      11'h633: dout <= 8'b11000111; // 1587 : 199 - 0xc7
      11'h634: dout <= 8'b00100000; // 1588 :  32 - 0x20
      11'h635: dout <= 8'b00100000; // 1589 :  32 - 0x20
      11'h636: dout <= 8'b01100000; // 1590 :  96 - 0x60
      11'h637: dout <= 8'b11100000; // 1591 : 224 - 0xe0
      11'h638: dout <= 8'b00000111; // 1592 :   7 - 0x7 -- Sprite 0xc7
      11'h639: dout <= 8'b00000011; // 1593 :   3 - 0x3
      11'h63A: dout <= 8'b00000000; // 1594 :   0 - 0x0
      11'h63B: dout <= 8'b00000000; // 1595 :   0 - 0x0
      11'h63C: dout <= 8'b11100000; // 1596 : 224 - 0xe0
      11'h63D: dout <= 8'b00100000; // 1597 :  32 - 0x20
      11'h63E: dout <= 8'b11100000; // 1598 : 224 - 0xe0
      11'h63F: dout <= 8'b11100000; // 1599 : 224 - 0xe0
      11'h640: dout <= 8'b11100000; // 1600 : 224 - 0xe0 -- Sprite 0xc8
      11'h641: dout <= 8'b11000000; // 1601 : 192 - 0xc0
      11'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      11'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      11'h644: dout <= 8'b00000111; // 1604 :   7 - 0x7
      11'h645: dout <= 8'b00000001; // 1605 :   1 - 0x1
      11'h646: dout <= 8'b00000111; // 1606 :   7 - 0x7
      11'h647: dout <= 8'b00000111; // 1607 :   7 - 0x7
      11'h648: dout <= 8'b00010011; // 1608 :  19 - 0x13 -- Sprite 0xc9
      11'h649: dout <= 8'b00011111; // 1609 :  31 - 0x1f
      11'h64A: dout <= 8'b00001101; // 1610 :  13 - 0xd
      11'h64B: dout <= 8'b00000100; // 1611 :   4 - 0x4
      11'h64C: dout <= 8'b00001100; // 1612 :  12 - 0xc
      11'h64D: dout <= 8'b00010011; // 1613 :  19 - 0x13
      11'h64E: dout <= 8'b00011111; // 1614 :  31 - 0x1f
      11'h64F: dout <= 8'b00000001; // 1615 :   1 - 0x1
      11'h650: dout <= 8'b01100000; // 1616 :  96 - 0x60 -- Sprite 0xca
      11'h651: dout <= 8'b11110011; // 1617 : 243 - 0xf3
      11'h652: dout <= 8'b10100111; // 1618 : 167 - 0xa7
      11'h653: dout <= 8'b11000110; // 1619 : 198 - 0xc6
      11'h654: dout <= 8'b01110100; // 1620 : 116 - 0x74
      11'h655: dout <= 8'b00000100; // 1621 :   4 - 0x4
      11'h656: dout <= 8'b10000111; // 1622 : 135 - 0x87
      11'h657: dout <= 8'b10000111; // 1623 : 135 - 0x87
      11'h658: dout <= 8'b00000110; // 1624 :   6 - 0x6 -- Sprite 0xcb
      11'h659: dout <= 8'b10001111; // 1625 : 143 - 0x8f
      11'h65A: dout <= 8'b11000011; // 1626 : 195 - 0xc3
      11'h65B: dout <= 8'b00100001; // 1627 :  33 - 0x21
      11'h65C: dout <= 8'b00100000; // 1628 :  32 - 0x20
      11'h65D: dout <= 8'b01100000; // 1629 :  96 - 0x60
      11'h65E: dout <= 8'b11100000; // 1630 : 224 - 0xe0
      11'h65F: dout <= 8'b11100000; // 1631 : 224 - 0xe0
      11'h660: dout <= 8'b11000011; // 1632 : 195 - 0xc3 -- Sprite 0xcc
      11'h661: dout <= 8'b01110000; // 1633 : 112 - 0x70
      11'h662: dout <= 8'b00000000; // 1634 :   0 - 0x0
      11'h663: dout <= 8'b01100000; // 1635 :  96 - 0x60
      11'h664: dout <= 8'b11110000; // 1636 : 240 - 0xf0
      11'h665: dout <= 8'b11010000; // 1637 : 208 - 0xd0
      11'h666: dout <= 8'b10010000; // 1638 : 144 - 0x90
      11'h667: dout <= 8'b01100000; // 1639 :  96 - 0x60
      11'h668: dout <= 8'b11000000; // 1640 : 192 - 0xc0 -- Sprite 0xcd
      11'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      11'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      11'h66B: dout <= 8'b00000110; // 1643 :   6 - 0x6
      11'h66C: dout <= 8'b00001111; // 1644 :  15 - 0xf
      11'h66D: dout <= 8'b00001101; // 1645 :  13 - 0xd
      11'h66E: dout <= 8'b00001001; // 1646 :   9 - 0x9
      11'h66F: dout <= 8'b00000110; // 1647 :   6 - 0x6
      11'h670: dout <= 8'b11111100; // 1648 : 252 - 0xfc -- Sprite 0xce
      11'h671: dout <= 8'b11000000; // 1649 : 192 - 0xc0
      11'h672: dout <= 8'b11010001; // 1650 : 209 - 0xd1
      11'h673: dout <= 8'b11000010; // 1651 : 194 - 0xc2
      11'h674: dout <= 8'b10011110; // 1652 : 158 - 0x9e
      11'h675: dout <= 8'b10111111; // 1653 : 191 - 0xbf
      11'h676: dout <= 8'b10110000; // 1654 : 176 - 0xb0
      11'h677: dout <= 8'b10110011; // 1655 : 179 - 0xb3
      11'h678: dout <= 8'b00000111; // 1656 :   7 - 0x7 -- Sprite 0xcf
      11'h679: dout <= 8'b11110011; // 1657 : 243 - 0xf3
      11'h67A: dout <= 8'b00001011; // 1658 :  11 - 0xb
      11'h67B: dout <= 8'b01111011; // 1659 : 123 - 0x7b
      11'h67C: dout <= 8'b01111011; // 1660 : 123 - 0x7b
      11'h67D: dout <= 8'b11111001; // 1661 : 249 - 0xf9
      11'h67E: dout <= 8'b00001101; // 1662 :  13 - 0xd
      11'h67F: dout <= 8'b11101101; // 1663 : 237 - 0xed
      11'h680: dout <= 8'b11111111; // 1664 : 255 - 0xff -- Sprite 0xd0
      11'h681: dout <= 8'b11111111; // 1665 : 255 - 0xff
      11'h682: dout <= 8'b11111111; // 1666 : 255 - 0xff
      11'h683: dout <= 8'b11111111; // 1667 : 255 - 0xff
      11'h684: dout <= 8'b11101110; // 1668 : 238 - 0xee
      11'h685: dout <= 8'b11101110; // 1669 : 238 - 0xee
      11'h686: dout <= 8'b11101110; // 1670 : 238 - 0xee
      11'h687: dout <= 8'b11101110; // 1671 : 238 - 0xee
      11'h688: dout <= 8'b11111111; // 1672 : 255 - 0xff -- Sprite 0xd1
      11'h689: dout <= 8'b11111111; // 1673 : 255 - 0xff
      11'h68A: dout <= 8'b11111111; // 1674 : 255 - 0xff
      11'h68B: dout <= 8'b11111011; // 1675 : 251 - 0xfb
      11'h68C: dout <= 8'b11111011; // 1676 : 251 - 0xfb
      11'h68D: dout <= 8'b11111011; // 1677 : 251 - 0xfb
      11'h68E: dout <= 8'b11111011; // 1678 : 251 - 0xfb
      11'h68F: dout <= 8'b11111011; // 1679 : 251 - 0xfb
      11'h690: dout <= 8'b11111111; // 1680 : 255 - 0xff -- Sprite 0xd2
      11'h691: dout <= 8'b11111111; // 1681 : 255 - 0xff
      11'h692: dout <= 8'b11111111; // 1682 : 255 - 0xff
      11'h693: dout <= 8'b11111111; // 1683 : 255 - 0xff
      11'h694: dout <= 8'b11101110; // 1684 : 238 - 0xee
      11'h695: dout <= 8'b10001110; // 1685 : 142 - 0x8e
      11'h696: dout <= 8'b11111110; // 1686 : 254 - 0xfe
      11'h697: dout <= 8'b11111110; // 1687 : 254 - 0xfe
      11'h698: dout <= 8'b11111111; // 1688 : 255 - 0xff -- Sprite 0xd3
      11'h699: dout <= 8'b11111111; // 1689 : 255 - 0xff
      11'h69A: dout <= 8'b11111111; // 1690 : 255 - 0xff
      11'h69B: dout <= 8'b11111111; // 1691 : 255 - 0xff
      11'h69C: dout <= 8'b11101110; // 1692 : 238 - 0xee
      11'h69D: dout <= 8'b10001110; // 1693 : 142 - 0x8e
      11'h69E: dout <= 8'b11111100; // 1694 : 252 - 0xfc
      11'h69F: dout <= 8'b11111101; // 1695 : 253 - 0xfd
      11'h6A0: dout <= 8'b11111111; // 1696 : 255 - 0xff -- Sprite 0xd4
      11'h6A1: dout <= 8'b11111111; // 1697 : 255 - 0xff
      11'h6A2: dout <= 8'b11111111; // 1698 : 255 - 0xff
      11'h6A3: dout <= 8'b11111110; // 1699 : 254 - 0xfe
      11'h6A4: dout <= 8'b11101110; // 1700 : 238 - 0xee
      11'h6A5: dout <= 8'b11101110; // 1701 : 238 - 0xee
      11'h6A6: dout <= 8'b11101110; // 1702 : 238 - 0xee
      11'h6A7: dout <= 8'b11101110; // 1703 : 238 - 0xee
      11'h6A8: dout <= 8'b11111111; // 1704 : 255 - 0xff -- Sprite 0xd5
      11'h6A9: dout <= 8'b11111111; // 1705 : 255 - 0xff
      11'h6AA: dout <= 8'b11111111; // 1706 : 255 - 0xff
      11'h6AB: dout <= 8'b11111101; // 1707 : 253 - 0xfd
      11'h6AC: dout <= 8'b11100001; // 1708 : 225 - 0xe1
      11'h6AD: dout <= 8'b11101111; // 1709 : 239 - 0xef
      11'h6AE: dout <= 8'b11111111; // 1710 : 255 - 0xff
      11'h6AF: dout <= 8'b11111111; // 1711 : 255 - 0xff
      11'h6B0: dout <= 8'b11111111; // 1712 : 255 - 0xff -- Sprite 0xd6
      11'h6B1: dout <= 8'b11111111; // 1713 : 255 - 0xff
      11'h6B2: dout <= 8'b11111111; // 1714 : 255 - 0xff
      11'h6B3: dout <= 8'b11111101; // 1715 : 253 - 0xfd
      11'h6B4: dout <= 8'b11100001; // 1716 : 225 - 0xe1
      11'h6B5: dout <= 8'b11101111; // 1717 : 239 - 0xef
      11'h6B6: dout <= 8'b11111111; // 1718 : 255 - 0xff
      11'h6B7: dout <= 8'b11111111; // 1719 : 255 - 0xff
      11'h6B8: dout <= 8'b11111111; // 1720 : 255 - 0xff -- Sprite 0xd7
      11'h6B9: dout <= 8'b11111111; // 1721 : 255 - 0xff
      11'h6BA: dout <= 8'b11111111; // 1722 : 255 - 0xff
      11'h6BB: dout <= 8'b11111110; // 1723 : 254 - 0xfe
      11'h6BC: dout <= 8'b11101110; // 1724 : 238 - 0xee
      11'h6BD: dout <= 8'b10001110; // 1725 : 142 - 0x8e
      11'h6BE: dout <= 8'b11111110; // 1726 : 254 - 0xfe
      11'h6BF: dout <= 8'b11111100; // 1727 : 252 - 0xfc
      11'h6C0: dout <= 8'b11111111; // 1728 : 255 - 0xff -- Sprite 0xd8
      11'h6C1: dout <= 8'b11111111; // 1729 : 255 - 0xff
      11'h6C2: dout <= 8'b11111111; // 1730 : 255 - 0xff
      11'h6C3: dout <= 8'b11111111; // 1731 : 255 - 0xff
      11'h6C4: dout <= 8'b11101110; // 1732 : 238 - 0xee
      11'h6C5: dout <= 8'b11101110; // 1733 : 238 - 0xee
      11'h6C6: dout <= 8'b11111100; // 1734 : 252 - 0xfc
      11'h6C7: dout <= 8'b11111111; // 1735 : 255 - 0xff
      11'h6C8: dout <= 8'b11111111; // 1736 : 255 - 0xff -- Sprite 0xd9
      11'h6C9: dout <= 8'b11111111; // 1737 : 255 - 0xff
      11'h6CA: dout <= 8'b11111111; // 1738 : 255 - 0xff
      11'h6CB: dout <= 8'b11111111; // 1739 : 255 - 0xff
      11'h6CC: dout <= 8'b11101110; // 1740 : 238 - 0xee
      11'h6CD: dout <= 8'b11101110; // 1741 : 238 - 0xee
      11'h6CE: dout <= 8'b11101110; // 1742 : 238 - 0xee
      11'h6CF: dout <= 8'b11101110; // 1743 : 238 - 0xee
      11'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0xda
      11'h6D1: dout <= 8'b00000000; // 1745 :   0 - 0x0
      11'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      11'h6D3: dout <= 8'b10000000; // 1747 : 128 - 0x80
      11'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      11'h6D5: dout <= 8'b00000000; // 1749 :   0 - 0x0
      11'h6D6: dout <= 8'b00000100; // 1750 :   4 - 0x4
      11'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      11'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0 -- Sprite 0xdb
      11'h6D9: dout <= 8'b00000100; // 1753 :   4 - 0x4
      11'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      11'h6DB: dout <= 8'b00010001; // 1755 :  17 - 0x11
      11'h6DC: dout <= 8'b00000000; // 1756 :   0 - 0x0
      11'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      11'h6DE: dout <= 8'b00000000; // 1758 :   0 - 0x0
      11'h6DF: dout <= 8'b00100000; // 1759 :  32 - 0x20
      11'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0xdc
      11'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      11'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      11'h6E3: dout <= 8'b00100000; // 1763 :  32 - 0x20
      11'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      11'h6E5: dout <= 8'b00000000; // 1765 :   0 - 0x0
      11'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      11'h6E7: dout <= 8'b00000100; // 1767 :   4 - 0x4
      11'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- Sprite 0xdd
      11'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      11'h6EA: dout <= 8'b00010001; // 1770 :  17 - 0x11
      11'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      11'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      11'h6ED: dout <= 8'b10000000; // 1773 : 128 - 0x80
      11'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      11'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      11'h6F0: dout <= 8'b10110011; // 1776 : 179 - 0xb3 -- Sprite 0xde
      11'h6F1: dout <= 8'b10110011; // 1777 : 179 - 0xb3
      11'h6F2: dout <= 8'b10110011; // 1778 : 179 - 0xb3
      11'h6F3: dout <= 8'b10110011; // 1779 : 179 - 0xb3
      11'h6F4: dout <= 8'b10110000; // 1780 : 176 - 0xb0
      11'h6F5: dout <= 8'b10101111; // 1781 : 175 - 0xaf
      11'h6F6: dout <= 8'b10011111; // 1782 : 159 - 0x9f
      11'h6F7: dout <= 8'b11000000; // 1783 : 192 - 0xc0
      11'h6F8: dout <= 8'b11101101; // 1784 : 237 - 0xed -- Sprite 0xdf
      11'h6F9: dout <= 8'b11001101; // 1785 : 205 - 0xcd
      11'h6FA: dout <= 8'b11001101; // 1786 : 205 - 0xcd
      11'h6FB: dout <= 8'b00001101; // 1787 :  13 - 0xd
      11'h6FC: dout <= 8'b00001101; // 1788 :  13 - 0xd
      11'h6FD: dout <= 8'b11111101; // 1789 : 253 - 0xfd
      11'h6FE: dout <= 8'b11111101; // 1790 : 253 - 0xfd
      11'h6FF: dout <= 8'b00000011; // 1791 :   3 - 0x3
      11'h700: dout <= 8'b11101110; // 1792 : 238 - 0xee -- Sprite 0xe0
      11'h701: dout <= 8'b11101110; // 1793 : 238 - 0xee
      11'h702: dout <= 8'b11101110; // 1794 : 238 - 0xee
      11'h703: dout <= 8'b11101110; // 1795 : 238 - 0xee
      11'h704: dout <= 8'b11111110; // 1796 : 254 - 0xfe
      11'h705: dout <= 8'b11111100; // 1797 : 252 - 0xfc
      11'h706: dout <= 8'b11000001; // 1798 : 193 - 0xc1
      11'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      11'h708: dout <= 8'b11111011; // 1800 : 251 - 0xfb -- Sprite 0xe1
      11'h709: dout <= 8'b11111011; // 1801 : 251 - 0xfb
      11'h70A: dout <= 8'b11111011; // 1802 : 251 - 0xfb
      11'h70B: dout <= 8'b11111011; // 1803 : 251 - 0xfb
      11'h70C: dout <= 8'b11111111; // 1804 : 255 - 0xff
      11'h70D: dout <= 8'b11111101; // 1805 : 253 - 0xfd
      11'h70E: dout <= 8'b11000001; // 1806 : 193 - 0xc1
      11'h70F: dout <= 8'b11111111; // 1807 : 255 - 0xff
      11'h710: dout <= 8'b11111100; // 1808 : 252 - 0xfc -- Sprite 0xe2
      11'h711: dout <= 8'b11100001; // 1809 : 225 - 0xe1
      11'h712: dout <= 8'b11101111; // 1810 : 239 - 0xef
      11'h713: dout <= 8'b11101111; // 1811 : 239 - 0xef
      11'h714: dout <= 8'b11111111; // 1812 : 255 - 0xff
      11'h715: dout <= 8'b11111110; // 1813 : 254 - 0xfe
      11'h716: dout <= 8'b10000000; // 1814 : 128 - 0x80
      11'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      11'h718: dout <= 8'b11101110; // 1816 : 238 - 0xee -- Sprite 0xe3
      11'h719: dout <= 8'b11111110; // 1817 : 254 - 0xfe
      11'h71A: dout <= 8'b11111110; // 1818 : 254 - 0xfe
      11'h71B: dout <= 8'b11111110; // 1819 : 254 - 0xfe
      11'h71C: dout <= 8'b11111110; // 1820 : 254 - 0xfe
      11'h71D: dout <= 8'b11111100; // 1821 : 252 - 0xfc
      11'h71E: dout <= 8'b11000001; // 1822 : 193 - 0xc1
      11'h71F: dout <= 8'b11111111; // 1823 : 255 - 0xff
      11'h720: dout <= 8'b11101110; // 1824 : 238 - 0xee -- Sprite 0xe4
      11'h721: dout <= 8'b11101110; // 1825 : 238 - 0xee
      11'h722: dout <= 8'b11111110; // 1826 : 254 - 0xfe
      11'h723: dout <= 8'b11111110; // 1827 : 254 - 0xfe
      11'h724: dout <= 8'b10001110; // 1828 : 142 - 0x8e
      11'h725: dout <= 8'b11111110; // 1829 : 254 - 0xfe
      11'h726: dout <= 8'b11111000; // 1830 : 248 - 0xf8
      11'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      11'h728: dout <= 8'b10001110; // 1832 : 142 - 0x8e -- Sprite 0xe5
      11'h729: dout <= 8'b11111110; // 1833 : 254 - 0xfe
      11'h72A: dout <= 8'b11111110; // 1834 : 254 - 0xfe
      11'h72B: dout <= 8'b11111110; // 1835 : 254 - 0xfe
      11'h72C: dout <= 8'b11111110; // 1836 : 254 - 0xfe
      11'h72D: dout <= 8'b11111100; // 1837 : 252 - 0xfc
      11'h72E: dout <= 8'b11000001; // 1838 : 193 - 0xc1
      11'h72F: dout <= 8'b11111111; // 1839 : 255 - 0xff
      11'h730: dout <= 8'b11101110; // 1840 : 238 - 0xee -- Sprite 0xe6
      11'h731: dout <= 8'b11101110; // 1841 : 238 - 0xee
      11'h732: dout <= 8'b11101110; // 1842 : 238 - 0xee
      11'h733: dout <= 8'b11101110; // 1843 : 238 - 0xee
      11'h734: dout <= 8'b11111110; // 1844 : 254 - 0xfe
      11'h735: dout <= 8'b11111100; // 1845 : 252 - 0xfc
      11'h736: dout <= 8'b11000001; // 1846 : 193 - 0xc1
      11'h737: dout <= 8'b11111111; // 1847 : 255 - 0xff
      11'h738: dout <= 8'b11111101; // 1848 : 253 - 0xfd -- Sprite 0xe7
      11'h739: dout <= 8'b11111101; // 1849 : 253 - 0xfd
      11'h73A: dout <= 8'b11111001; // 1850 : 249 - 0xf9
      11'h73B: dout <= 8'b11111011; // 1851 : 251 - 0xfb
      11'h73C: dout <= 8'b11111011; // 1852 : 251 - 0xfb
      11'h73D: dout <= 8'b11111011; // 1853 : 251 - 0xfb
      11'h73E: dout <= 8'b11100011; // 1854 : 227 - 0xe3
      11'h73F: dout <= 8'b11111111; // 1855 : 255 - 0xff
      11'h740: dout <= 8'b11101110; // 1856 : 238 - 0xee -- Sprite 0xe8
      11'h741: dout <= 8'b11101110; // 1857 : 238 - 0xee
      11'h742: dout <= 8'b11101110; // 1858 : 238 - 0xee
      11'h743: dout <= 8'b11101110; // 1859 : 238 - 0xee
      11'h744: dout <= 8'b11111110; // 1860 : 254 - 0xfe
      11'h745: dout <= 8'b11111100; // 1861 : 252 - 0xfc
      11'h746: dout <= 8'b11000001; // 1862 : 193 - 0xc1
      11'h747: dout <= 8'b11111111; // 1863 : 255 - 0xff
      11'h748: dout <= 8'b11111110; // 1864 : 254 - 0xfe -- Sprite 0xe9
      11'h749: dout <= 8'b11111110; // 1865 : 254 - 0xfe
      11'h74A: dout <= 8'b11001110; // 1866 : 206 - 0xce
      11'h74B: dout <= 8'b11111110; // 1867 : 254 - 0xfe
      11'h74C: dout <= 8'b11111110; // 1868 : 254 - 0xfe
      11'h74D: dout <= 8'b11111100; // 1869 : 252 - 0xfc
      11'h74E: dout <= 8'b11000001; // 1870 : 193 - 0xc1
      11'h74F: dout <= 8'b11111111; // 1871 : 255 - 0xff
      11'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0xea
      11'h751: dout <= 8'b01110000; // 1873 : 112 - 0x70
      11'h752: dout <= 8'b00111000; // 1874 :  56 - 0x38
      11'h753: dout <= 8'b00000000; // 1875 :   0 - 0x0
      11'h754: dout <= 8'b00000010; // 1876 :   2 - 0x2
      11'h755: dout <= 8'b00000111; // 1877 :   7 - 0x7
      11'h756: dout <= 8'b00000011; // 1878 :   3 - 0x3
      11'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      11'h758: dout <= 8'b00000000; // 1880 :   0 - 0x0 -- Sprite 0xeb
      11'h759: dout <= 8'b00001100; // 1881 :  12 - 0xc
      11'h75A: dout <= 8'b00000110; // 1882 :   6 - 0x6
      11'h75B: dout <= 8'b00000110; // 1883 :   6 - 0x6
      11'h75C: dout <= 8'b01100000; // 1884 :  96 - 0x60
      11'h75D: dout <= 8'b01110000; // 1885 : 112 - 0x70
      11'h75E: dout <= 8'b00110000; // 1886 :  48 - 0x30
      11'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      11'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      11'h761: dout <= 8'b11000000; // 1889 : 192 - 0xc0
      11'h762: dout <= 8'b11100000; // 1890 : 224 - 0xe0
      11'h763: dout <= 8'b01100000; // 1891 :  96 - 0x60
      11'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      11'h765: dout <= 8'b00001100; // 1893 :  12 - 0xc
      11'h766: dout <= 8'b00001110; // 1894 :  14 - 0xe
      11'h767: dout <= 8'b00000110; // 1895 :   6 - 0x6
      11'h768: dout <= 8'b01100000; // 1896 :  96 - 0x60 -- Sprite 0xed
      11'h769: dout <= 8'b01110000; // 1897 : 112 - 0x70
      11'h76A: dout <= 8'b00110000; // 1898 :  48 - 0x30
      11'h76B: dout <= 8'b00000000; // 1899 :   0 - 0x0
      11'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      11'h76D: dout <= 8'b00001100; // 1901 :  12 - 0xc
      11'h76E: dout <= 8'b00001110; // 1902 :  14 - 0xe
      11'h76F: dout <= 8'b00000110; // 1903 :   6 - 0x6
      11'h770: dout <= 8'b11111111; // 1904 : 255 - 0xff -- Sprite 0xee
      11'h771: dout <= 8'b11111111; // 1905 : 255 - 0xff
      11'h772: dout <= 8'b10111101; // 1906 : 189 - 0xbd
      11'h773: dout <= 8'b11111111; // 1907 : 255 - 0xff
      11'h774: dout <= 8'b11111111; // 1908 : 255 - 0xff
      11'h775: dout <= 8'b11111011; // 1909 : 251 - 0xfb
      11'h776: dout <= 8'b11111111; // 1910 : 255 - 0xff
      11'h777: dout <= 8'b11111111; // 1911 : 255 - 0xff
      11'h778: dout <= 8'b11111111; // 1912 : 255 - 0xff -- Sprite 0xef
      11'h779: dout <= 8'b11111111; // 1913 : 255 - 0xff
      11'h77A: dout <= 8'b11111011; // 1914 : 251 - 0xfb
      11'h77B: dout <= 8'b11111111; // 1915 : 255 - 0xff
      11'h77C: dout <= 8'b11011111; // 1916 : 223 - 0xdf
      11'h77D: dout <= 8'b11111111; // 1917 : 255 - 0xff
      11'h77E: dout <= 8'b11111111; // 1918 : 255 - 0xff
      11'h77F: dout <= 8'b11111111; // 1919 : 255 - 0xff
      11'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      11'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      11'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      11'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      11'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      11'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      11'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      11'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      11'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0 -- Sprite 0xf1
      11'h789: dout <= 8'b10000000; // 1929 : 128 - 0x80
      11'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      11'h78B: dout <= 8'b00000000; // 1931 :   0 - 0x0
      11'h78C: dout <= 8'b00000000; // 1932 :   0 - 0x0
      11'h78D: dout <= 8'b00000000; // 1933 :   0 - 0x0
      11'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      11'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      11'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0xf2
      11'h791: dout <= 8'b11000000; // 1937 : 192 - 0xc0
      11'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      11'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      11'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      11'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      11'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      11'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      11'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0 -- Sprite 0xf3
      11'h799: dout <= 8'b11100000; // 1945 : 224 - 0xe0
      11'h79A: dout <= 8'b00000000; // 1946 :   0 - 0x0
      11'h79B: dout <= 8'b00000000; // 1947 :   0 - 0x0
      11'h79C: dout <= 8'b00000000; // 1948 :   0 - 0x0
      11'h79D: dout <= 8'b00000000; // 1949 :   0 - 0x0
      11'h79E: dout <= 8'b00000000; // 1950 :   0 - 0x0
      11'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      11'h7A0: dout <= 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0xf4
      11'h7A1: dout <= 8'b11110000; // 1953 : 240 - 0xf0
      11'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      11'h7A3: dout <= 8'b00000000; // 1955 :   0 - 0x0
      11'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      11'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      11'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      11'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      11'h7A8: dout <= 8'b00000000; // 1960 :   0 - 0x0 -- Sprite 0xf5
      11'h7A9: dout <= 8'b11111000; // 1961 : 248 - 0xf8
      11'h7AA: dout <= 8'b00000000; // 1962 :   0 - 0x0
      11'h7AB: dout <= 8'b00000000; // 1963 :   0 - 0x0
      11'h7AC: dout <= 8'b00000000; // 1964 :   0 - 0x0
      11'h7AD: dout <= 8'b00000000; // 1965 :   0 - 0x0
      11'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      11'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      11'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      11'h7B1: dout <= 8'b11111100; // 1969 : 252 - 0xfc
      11'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      11'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      11'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      11'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      11'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      11'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      11'h7B8: dout <= 8'b00000000; // 1976 :   0 - 0x0 -- Sprite 0xf7
      11'h7B9: dout <= 8'b11111110; // 1977 : 254 - 0xfe
      11'h7BA: dout <= 8'b00000000; // 1978 :   0 - 0x0
      11'h7BB: dout <= 8'b00000000; // 1979 :   0 - 0x0
      11'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      11'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      11'h7BE: dout <= 8'b00000000; // 1982 :   0 - 0x0
      11'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      11'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0xf8
      11'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      11'h7C2: dout <= 8'b00000000; // 1986 :   0 - 0x0
      11'h7C3: dout <= 8'b00000000; // 1987 :   0 - 0x0
      11'h7C4: dout <= 8'b00000000; // 1988 :   0 - 0x0
      11'h7C5: dout <= 8'b00000000; // 1989 :   0 - 0x0
      11'h7C6: dout <= 8'b00000000; // 1990 :   0 - 0x0
      11'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout <= 8'b11111111; // 1992 : 255 - 0xff -- Sprite 0xf9
      11'h7C9: dout <= 8'b11111111; // 1993 : 255 - 0xff
      11'h7CA: dout <= 8'b11111111; // 1994 : 255 - 0xff
      11'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      11'h7CC: dout <= 8'b10000000; // 1996 : 128 - 0x80
      11'h7CD: dout <= 8'b10000000; // 1997 : 128 - 0x80
      11'h7CE: dout <= 8'b11000000; // 1998 : 192 - 0xc0
      11'h7CF: dout <= 8'b11000000; // 1999 : 192 - 0xc0
      11'h7D0: dout <= 8'b11111111; // 2000 : 255 - 0xff -- Sprite 0xfa
      11'h7D1: dout <= 8'b11111111; // 2001 : 255 - 0xff
      11'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      11'h7D3: dout <= 8'b11111111; // 2003 : 255 - 0xff
      11'h7D4: dout <= 8'b00000000; // 2004 :   0 - 0x0
      11'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      11'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout <= 8'b11111111; // 2008 : 255 - 0xff -- Sprite 0xfb
      11'h7D9: dout <= 8'b11111111; // 2009 : 255 - 0xff
      11'h7DA: dout <= 8'b11111111; // 2010 : 255 - 0xff
      11'h7DB: dout <= 8'b11111111; // 2011 : 255 - 0xff
      11'h7DC: dout <= 8'b00000001; // 2012 :   1 - 0x1
      11'h7DD: dout <= 8'b00000000; // 2013 :   0 - 0x0
      11'h7DE: dout <= 8'b00000010; // 2014 :   2 - 0x2
      11'h7DF: dout <= 8'b00000010; // 2015 :   2 - 0x2
      11'h7E0: dout <= 8'b11000000; // 2016 : 192 - 0xc0 -- Sprite 0xfc
      11'h7E1: dout <= 8'b11000000; // 2017 : 192 - 0xc0
      11'h7E2: dout <= 8'b10000000; // 2018 : 128 - 0x80
      11'h7E3: dout <= 8'b10000000; // 2019 : 128 - 0x80
      11'h7E4: dout <= 8'b11000000; // 2020 : 192 - 0xc0
      11'h7E5: dout <= 8'b11111111; // 2021 : 255 - 0xff
      11'h7E6: dout <= 8'b11111111; // 2022 : 255 - 0xff
      11'h7E7: dout <= 8'b11111111; // 2023 : 255 - 0xff
      11'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0 -- Sprite 0xfd
      11'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      11'h7EA: dout <= 8'b00000000; // 2026 :   0 - 0x0
      11'h7EB: dout <= 8'b00000000; // 2027 :   0 - 0x0
      11'h7EC: dout <= 8'b00000000; // 2028 :   0 - 0x0
      11'h7ED: dout <= 8'b11111111; // 2029 : 255 - 0xff
      11'h7EE: dout <= 8'b11111111; // 2030 : 255 - 0xff
      11'h7EF: dout <= 8'b11111111; // 2031 : 255 - 0xff
      11'h7F0: dout <= 8'b00000010; // 2032 :   2 - 0x2 -- Sprite 0xfe
      11'h7F1: dout <= 8'b00000010; // 2033 :   2 - 0x2
      11'h7F2: dout <= 8'b00000000; // 2034 :   0 - 0x0
      11'h7F3: dout <= 8'b00000000; // 2035 :   0 - 0x0
      11'h7F4: dout <= 8'b00000000; // 2036 :   0 - 0x0
      11'h7F5: dout <= 8'b11111111; // 2037 : 255 - 0xff
      11'h7F6: dout <= 8'b11111111; // 2038 : 255 - 0xff
      11'h7F7: dout <= 8'b11111111; // 2039 : 255 - 0xff
      11'h7F8: dout <= 8'b11111111; // 2040 : 255 - 0xff -- Sprite 0xff
      11'h7F9: dout <= 8'b11111111; // 2041 : 255 - 0xff
      11'h7FA: dout <= 8'b11111111; // 2042 : 255 - 0xff
      11'h7FB: dout <= 8'b11111111; // 2043 : 255 - 0xff
      11'h7FC: dout <= 8'b11111111; // 2044 : 255 - 0xff
      11'h7FD: dout <= 8'b11111111; // 2045 : 255 - 0xff
      11'h7FE: dout <= 8'b11111111; // 2046 : 255 - 0xff
      11'h7FF: dout <= 8'b11111111; // 2047 : 255 - 0xff
    endcase
  end

endmodule
