//-   Sprites Pattern table COLOR PLANE 1
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_NOVA_SPR_PLN1
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table COLOR PLANE 1
      11'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      11'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      11'h2: dout  = 8'b00000011; //    2 :   3 - 0x3
      11'h3: dout  = 8'b00000001; //    3 :   1 - 0x1
      11'h4: dout  = 8'b00000001; //    4 :   1 - 0x1
      11'h5: dout  = 8'b00000000; //    5 :   0 - 0x0
      11'h6: dout  = 8'b00000011; //    6 :   3 - 0x3
      11'h7: dout  = 8'b00000001; //    7 :   1 - 0x1
      11'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      11'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      11'hA: dout  = 8'b00111000; //   10 :  56 - 0x38
      11'hB: dout  = 8'b10110100; //   11 : 180 - 0xb4
      11'hC: dout  = 8'b10101000; //   12 : 168 - 0xa8
      11'hD: dout  = 8'b11010100; //   13 : 212 - 0xd4
      11'hE: dout  = 8'b01110100; //   14 : 116 - 0x74
      11'hF: dout  = 8'b01111110; //   15 : 126 - 0x7e
      11'h10: dout  = 8'b00111000; //   16 :  56 - 0x38 -- Sprite 0x2
      11'h11: dout  = 8'b01111000; //   17 : 120 - 0x78
      11'h12: dout  = 8'b01111100; //   18 : 124 - 0x7c
      11'h13: dout  = 8'b01111110; //   19 : 126 - 0x7e
      11'h14: dout  = 8'b01111110; //   20 : 126 - 0x7e
      11'h15: dout  = 8'b01111110; //   21 : 126 - 0x7e
      11'h16: dout  = 8'b00111110; //   22 :  62 - 0x3e
      11'h17: dout  = 8'b00011110; //   23 :  30 - 0x1e
      11'h18: dout  = 8'b11110110; //   24 : 246 - 0xf6 -- Sprite 0x3
      11'h19: dout  = 8'b11110000; //   25 : 240 - 0xf0
      11'h1A: dout  = 8'b00111000; //   26 :  56 - 0x38
      11'h1B: dout  = 8'b11010000; //   27 : 208 - 0xd0
      11'h1C: dout  = 8'b11100000; //   28 : 224 - 0xe0
      11'h1D: dout  = 8'b01110000; //   29 : 112 - 0x70
      11'h1E: dout  = 8'b10111000; //   30 : 184 - 0xb8
      11'h1F: dout  = 8'b01000000; //   31 :  64 - 0x40
      11'h20: dout  = 8'b00011100; //   32 :  28 - 0x1c -- Sprite 0x4
      11'h21: dout  = 8'b00011100; //   33 :  28 - 0x1c
      11'h22: dout  = 8'b00011110; //   34 :  30 - 0x1e
      11'h23: dout  = 8'b00011111; //   35 :  31 - 0x1f
      11'h24: dout  = 8'b00001100; //   36 :  12 - 0xc
      11'h25: dout  = 8'b00000000; //   37 :   0 - 0x0
      11'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      11'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      11'h28: dout  = 8'b10101000; //   40 : 168 - 0xa8 -- Sprite 0x5
      11'h29: dout  = 8'b01010000; //   41 :  80 - 0x50
      11'h2A: dout  = 8'b10101000; //   42 : 168 - 0xa8
      11'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      11'h2C: dout  = 8'b01100000; //   44 :  96 - 0x60
      11'h2D: dout  = 8'b01100000; //   45 :  96 - 0x60
      11'h2E: dout  = 8'b01110000; //   46 : 112 - 0x70
      11'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      11'h30: dout  = 8'b00011100; //   48 :  28 - 0x1c -- Sprite 0x6
      11'h31: dout  = 8'b00011100; //   49 :  28 - 0x1c
      11'h32: dout  = 8'b00011110; //   50 :  30 - 0x1e
      11'h33: dout  = 8'b00011111; //   51 :  31 - 0x1f
      11'h34: dout  = 8'b00001100; //   52 :  12 - 0xc
      11'h35: dout  = 8'b00000000; //   53 :   0 - 0x0
      11'h36: dout  = 8'b00000001; //   54 :   1 - 0x1
      11'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      11'h38: dout  = 8'b10101000; //   56 : 168 - 0xa8 -- Sprite 0x7
      11'h39: dout  = 8'b01010000; //   57 :  80 - 0x50
      11'h3A: dout  = 8'b10101000; //   58 : 168 - 0xa8
      11'h3B: dout  = 8'b00000000; //   59 :   0 - 0x0
      11'h3C: dout  = 8'b01011000; //   60 :  88 - 0x58
      11'h3D: dout  = 8'b11011000; //   61 : 216 - 0xd8
      11'h3E: dout  = 8'b10001100; //   62 : 140 - 0x8c
      11'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      11'h40: dout  = 8'b00011100; //   64 :  28 - 0x1c -- Sprite 0x8
      11'h41: dout  = 8'b00011100; //   65 :  28 - 0x1c
      11'h42: dout  = 8'b00011110; //   66 :  30 - 0x1e
      11'h43: dout  = 8'b00011111; //   67 :  31 - 0x1f
      11'h44: dout  = 8'b00001100; //   68 :  12 - 0xc
      11'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      11'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      11'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      11'h48: dout  = 8'b10101000; //   72 : 168 - 0xa8 -- Sprite 0x9
      11'h49: dout  = 8'b01010100; //   73 :  84 - 0x54
      11'h4A: dout  = 8'b10101000; //   74 : 168 - 0xa8
      11'h4B: dout  = 8'b00000000; //   75 :   0 - 0x0
      11'h4C: dout  = 8'b01101110; //   76 : 110 - 0x6e
      11'h4D: dout  = 8'b11000000; //   77 : 192 - 0xc0
      11'h4E: dout  = 8'b10000000; //   78 : 128 - 0x80
      11'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      11'h50: dout  = 8'b00011100; //   80 :  28 - 0x1c -- Sprite 0xa
      11'h51: dout  = 8'b00011100; //   81 :  28 - 0x1c
      11'h52: dout  = 8'b00011110; //   82 :  30 - 0x1e
      11'h53: dout  = 8'b00011111; //   83 :  31 - 0x1f
      11'h54: dout  = 8'b00001100; //   84 :  12 - 0xc
      11'h55: dout  = 8'b00000001; //   85 :   1 - 0x1
      11'h56: dout  = 8'b00000000; //   86 :   0 - 0x0
      11'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      11'h58: dout  = 8'b10101000; //   88 : 168 - 0xa8 -- Sprite 0xb
      11'h59: dout  = 8'b01010100; //   89 :  84 - 0x54
      11'h5A: dout  = 8'b10101000; //   90 : 168 - 0xa8
      11'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      11'h5C: dout  = 8'b11011000; //   92 : 216 - 0xd8
      11'h5D: dout  = 8'b11011100; //   93 : 220 - 0xdc
      11'h5E: dout  = 8'b00001100; //   94 :  12 - 0xc
      11'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      11'h60: dout  = 8'b11110110; //   96 : 246 - 0xf6 -- Sprite 0xc
      11'h61: dout  = 8'b11110000; //   97 : 240 - 0xf0
      11'h62: dout  = 8'b00000000; //   98 :   0 - 0x0
      11'h63: dout  = 8'b11111100; //   99 : 252 - 0xfc
      11'h64: dout  = 8'b11111000; //  100 : 248 - 0xf8
      11'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      11'h66: dout  = 8'b10101000; //  102 : 168 - 0xa8
      11'h67: dout  = 8'b01010100; //  103 :  84 - 0x54
      11'h68: dout  = 8'b00111000; //  104 :  56 - 0x38 -- Sprite 0xd
      11'h69: dout  = 8'b01111000; //  105 : 120 - 0x78
      11'h6A: dout  = 8'b01111100; //  106 : 124 - 0x7c
      11'h6B: dout  = 8'b01111101; //  107 : 125 - 0x7d
      11'h6C: dout  = 8'b01111101; //  108 : 125 - 0x7d
      11'h6D: dout  = 8'b01111011; //  109 : 123 - 0x7b
      11'h6E: dout  = 8'b00111011; //  110 :  59 - 0x3b
      11'h6F: dout  = 8'b00011011; //  111 :  27 - 0x1b
      11'h70: dout  = 8'b11110110; //  112 : 246 - 0xf6 -- Sprite 0xe
      11'h71: dout  = 8'b11110000; //  113 : 240 - 0xf0
      11'h72: dout  = 8'b01111000; //  114 : 120 - 0x78
      11'h73: dout  = 8'b01110000; //  115 : 112 - 0x70
      11'h74: dout  = 8'b10100000; //  116 : 160 - 0xa0
      11'h75: dout  = 8'b10010000; //  117 : 144 - 0x90
      11'h76: dout  = 8'b00101000; //  118 :  40 - 0x28
      11'h77: dout  = 8'b01010100; //  119 :  84 - 0x54
      11'h78: dout  = 8'b00000000; //  120 :   0 - 0x0 -- Sprite 0xf
      11'h79: dout  = 8'b00000000; //  121 :   0 - 0x0
      11'h7A: dout  = 8'b00000011; //  122 :   3 - 0x3
      11'h7B: dout  = 8'b00000001; //  123 :   1 - 0x1
      11'h7C: dout  = 8'b00000001; //  124 :   1 - 0x1
      11'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      11'h7E: dout  = 8'b00000011; //  126 :   3 - 0x3
      11'h7F: dout  = 8'b00000001; //  127 :   1 - 0x1
      11'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      11'h81: dout  = 8'b00000011; //  129 :   3 - 0x3
      11'h82: dout  = 8'b00001111; //  130 :  15 - 0xf
      11'h83: dout  = 8'b00001111; //  131 :  15 - 0xf
      11'h84: dout  = 8'b00001111; //  132 :  15 - 0xf
      11'h85: dout  = 8'b00011111; //  133 :  31 - 0x1f
      11'h86: dout  = 8'b00011111; //  134 :  31 - 0x1f
      11'h87: dout  = 8'b00011110; //  135 :  30 - 0x1e
      11'h88: dout  = 8'b00110110; //  136 :  54 - 0x36 -- Sprite 0x11
      11'h89: dout  = 8'b10110000; //  137 : 176 - 0xb0
      11'h8A: dout  = 8'b10111000; //  138 : 184 - 0xb8
      11'h8B: dout  = 8'b10010000; //  139 : 144 - 0x90
      11'h8C: dout  = 8'b10100000; //  140 : 160 - 0xa0
      11'h8D: dout  = 8'b01110000; //  141 : 112 - 0x70
      11'h8E: dout  = 8'b00111000; //  142 :  56 - 0x38
      11'h8F: dout  = 8'b01000000; //  143 :  64 - 0x40
      11'h90: dout  = 8'b00011100; //  144 :  28 - 0x1c -- Sprite 0x12
      11'h91: dout  = 8'b00011100; //  145 :  28 - 0x1c
      11'h92: dout  = 8'b00011110; //  146 :  30 - 0x1e
      11'h93: dout  = 8'b00011111; //  147 :  31 - 0x1f
      11'h94: dout  = 8'b00001100; //  148 :  12 - 0xc
      11'h95: dout  = 8'b00000000; //  149 :   0 - 0x0
      11'h96: dout  = 8'b00000000; //  150 :   0 - 0x0
      11'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      11'h98: dout  = 8'b00000000; //  152 :   0 - 0x0 -- Sprite 0x13
      11'h99: dout  = 8'b00000000; //  153 :   0 - 0x0
      11'h9A: dout  = 8'b00000000; //  154 :   0 - 0x0
      11'h9B: dout  = 8'b00000011; //  155 :   3 - 0x3
      11'h9C: dout  = 8'b00000111; //  156 :   7 - 0x7
      11'h9D: dout  = 8'b00001111; //  157 :  15 - 0xf
      11'h9E: dout  = 8'b00001111; //  158 :  15 - 0xf
      11'h9F: dout  = 8'b00011111; //  159 :  31 - 0x1f
      11'hA0: dout  = 8'b11110110; //  160 : 246 - 0xf6 -- Sprite 0x14
      11'hA1: dout  = 8'b00000000; //  161 :   0 - 0x0
      11'hA2: dout  = 8'b11111000; //  162 : 248 - 0xf8
      11'hA3: dout  = 8'b11111110; //  163 : 254 - 0xfe
      11'hA4: dout  = 8'b11111110; //  164 : 254 - 0xfe
      11'hA5: dout  = 8'b11111110; //  165 : 254 - 0xfe
      11'hA6: dout  = 8'b11111000; //  166 : 248 - 0xf8
      11'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      11'hA8: dout  = 8'b00000011; //  168 :   3 - 0x3 -- Sprite 0x15
      11'hA9: dout  = 8'b00000011; //  169 :   3 - 0x3
      11'hAA: dout  = 8'b00000000; //  170 :   0 - 0x0
      11'hAB: dout  = 8'b00000011; //  171 :   3 - 0x3
      11'hAC: dout  = 8'b00000011; //  172 :   3 - 0x3
      11'hAD: dout  = 8'b00000000; //  173 :   0 - 0x0
      11'hAE: dout  = 8'b00001111; //  174 :  15 - 0xf
      11'hAF: dout  = 8'b00111111; //  175 :  63 - 0x3f
      11'hB0: dout  = 8'b11011000; //  176 : 216 - 0xd8 -- Sprite 0x16
      11'hB1: dout  = 8'b11000000; //  177 : 192 - 0xc0
      11'hB2: dout  = 8'b11100000; //  178 : 224 - 0xe0
      11'hB3: dout  = 8'b01000000; //  179 :  64 - 0x40
      11'hB4: dout  = 8'b10000000; //  180 : 128 - 0x80
      11'hB5: dout  = 8'b00000000; //  181 :   0 - 0x0
      11'hB6: dout  = 8'b11100000; //  182 : 224 - 0xe0
      11'hB7: dout  = 8'b11111100; //  183 : 252 - 0xfc
      11'hB8: dout  = 8'b01111111; //  184 : 127 - 0x7f -- Sprite 0x17
      11'hB9: dout  = 8'b01111111; //  185 : 127 - 0x7f
      11'hBA: dout  = 8'b01111111; //  186 : 127 - 0x7f
      11'hBB: dout  = 8'b01111100; //  187 : 124 - 0x7c
      11'hBC: dout  = 8'b00110000; //  188 :  48 - 0x30
      11'hBD: dout  = 8'b00000001; //  189 :   1 - 0x1
      11'hBE: dout  = 8'b00000001; //  190 :   1 - 0x1
      11'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      11'hC0: dout  = 8'b11111100; //  192 : 252 - 0xfc -- Sprite 0x18
      11'hC1: dout  = 8'b11111110; //  193 : 254 - 0xfe
      11'hC2: dout  = 8'b11111100; //  194 : 252 - 0xfc
      11'hC3: dout  = 8'b00000000; //  195 :   0 - 0x0
      11'hC4: dout  = 8'b00000000; //  196 :   0 - 0x0
      11'hC5: dout  = 8'b10000000; //  197 : 128 - 0x80
      11'hC6: dout  = 8'b11000000; //  198 : 192 - 0xc0
      11'hC7: dout  = 8'b00000000; //  199 :   0 - 0x0
      11'hC8: dout  = 8'b00000111; //  200 :   7 - 0x7 -- Sprite 0x19
      11'hC9: dout  = 8'b00000111; //  201 :   7 - 0x7
      11'hCA: dout  = 8'b00000001; //  202 :   1 - 0x1
      11'hCB: dout  = 8'b00000110; //  203 :   6 - 0x6
      11'hCC: dout  = 8'b00000111; //  204 :   7 - 0x7
      11'hCD: dout  = 8'b00000110; //  205 :   6 - 0x6
      11'hCE: dout  = 8'b00000000; //  206 :   0 - 0x0
      11'hCF: dout  = 8'b00001111; //  207 :  15 - 0xf
      11'hD0: dout  = 8'b10110000; //  208 : 176 - 0xb0 -- Sprite 0x1a
      11'hD1: dout  = 8'b10000000; //  209 : 128 - 0x80
      11'hD2: dout  = 8'b11000000; //  210 : 192 - 0xc0
      11'hD3: dout  = 8'b10000000; //  211 : 128 - 0x80
      11'hD4: dout  = 8'b00000000; //  212 :   0 - 0x0
      11'hD5: dout  = 8'b00000000; //  213 :   0 - 0x0
      11'hD6: dout  = 8'b00000000; //  214 :   0 - 0x0
      11'hD7: dout  = 8'b11100000; //  215 : 224 - 0xe0
      11'hD8: dout  = 8'b00111111; //  216 :  63 - 0x3f -- Sprite 0x1b
      11'hD9: dout  = 8'b00111111; //  217 :  63 - 0x3f
      11'hDA: dout  = 8'b01111111; //  218 : 127 - 0x7f
      11'hDB: dout  = 8'b01111111; //  219 : 127 - 0x7f
      11'hDC: dout  = 8'b00111111; //  220 :  63 - 0x3f
      11'hDD: dout  = 8'b00000000; //  221 :   0 - 0x0
      11'hDE: dout  = 8'b00000011; //  222 :   3 - 0x3
      11'hDF: dout  = 8'b00000000; //  223 :   0 - 0x0
      11'hE0: dout  = 8'b11111111; //  224 : 255 - 0xff -- Sprite 0x1c
      11'hE1: dout  = 8'b11111111; //  225 : 255 - 0xff
      11'hE2: dout  = 8'b11111111; //  226 : 255 - 0xff
      11'hE3: dout  = 8'b11111111; //  227 : 255 - 0xff
      11'hE4: dout  = 8'b11111111; //  228 : 255 - 0xff
      11'hE5: dout  = 8'b00000000; //  229 :   0 - 0x0
      11'hE6: dout  = 8'b10000000; //  230 : 128 - 0x80
      11'hE7: dout  = 8'b00000000; //  231 :   0 - 0x0
      11'hE8: dout  = 8'b00000000; //  232 :   0 - 0x0 -- Sprite 0x1d
      11'hE9: dout  = 8'b11000000; //  233 : 192 - 0xc0
      11'hEA: dout  = 8'b11000000; //  234 : 192 - 0xc0
      11'hEB: dout  = 8'b11000000; //  235 : 192 - 0xc0
      11'hEC: dout  = 8'b10000000; //  236 : 128 - 0x80
      11'hED: dout  = 8'b00000000; //  237 :   0 - 0x0
      11'hEE: dout  = 8'b00000000; //  238 :   0 - 0x0
      11'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      11'hF0: dout  = 8'b11100000; //  240 : 224 - 0xe0 -- Sprite 0x1e
      11'hF1: dout  = 8'b10011100; //  241 : 156 - 0x9c
      11'hF2: dout  = 8'b00111000; //  242 :  56 - 0x38
      11'hF3: dout  = 8'b11100000; //  243 : 224 - 0xe0
      11'hF4: dout  = 8'b11001000; //  244 : 200 - 0xc8
      11'hF5: dout  = 8'b00010100; //  245 :  20 - 0x14
      11'hF6: dout  = 8'b10101000; //  246 : 168 - 0xa8
      11'hF7: dout  = 8'b01010100; //  247 :  84 - 0x54
      11'hF8: dout  = 8'b00000000; //  248 :   0 - 0x0 -- Sprite 0x1f
      11'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      11'hFA: dout  = 8'b00111000; //  250 :  56 - 0x38
      11'hFB: dout  = 8'b10110100; //  251 : 180 - 0xb4
      11'hFC: dout  = 8'b10101000; //  252 : 168 - 0xa8
      11'hFD: dout  = 8'b11010100; //  253 : 212 - 0xd4
      11'hFE: dout  = 8'b01110100; //  254 : 116 - 0x74
      11'hFF: dout  = 8'b00011110; //  255 :  30 - 0x1e
      11'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      11'h101: dout  = 8'b00000000; //  257 :   0 - 0x0
      11'h102: dout  = 8'b00001100; //  258 :  12 - 0xc
      11'h103: dout  = 8'b00000111; //  259 :   7 - 0x7
      11'h104: dout  = 8'b00001111; //  260 :  15 - 0xf
      11'h105: dout  = 8'b00000111; //  261 :   7 - 0x7
      11'h106: dout  = 8'b00001111; //  262 :  15 - 0xf
      11'h107: dout  = 8'b00001111; //  263 :  15 - 0xf
      11'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- Sprite 0x21
      11'h109: dout  = 8'b00000000; //  265 :   0 - 0x0
      11'h10A: dout  = 8'b00110000; //  266 :  48 - 0x30
      11'h10B: dout  = 8'b11100000; //  267 : 224 - 0xe0
      11'h10C: dout  = 8'b11110000; //  268 : 240 - 0xf0
      11'h10D: dout  = 8'b11100000; //  269 : 224 - 0xe0
      11'h10E: dout  = 8'b11110000; //  270 : 240 - 0xf0
      11'h10F: dout  = 8'b11110000; //  271 : 240 - 0xf0
      11'h110: dout  = 8'b00000111; //  272 :   7 - 0x7 -- Sprite 0x22
      11'h111: dout  = 8'b00000011; //  273 :   3 - 0x3
      11'h112: dout  = 8'b00011000; //  274 :  24 - 0x18
      11'h113: dout  = 8'b00010101; //  275 :  21 - 0x15
      11'h114: dout  = 8'b00000010; //  276 :   2 - 0x2
      11'h115: dout  = 8'b00000101; //  277 :   5 - 0x5
      11'h116: dout  = 8'b00000010; //  278 :   2 - 0x2
      11'h117: dout  = 8'b00000100; //  279 :   4 - 0x4
      11'h118: dout  = 8'b11100000; //  280 : 224 - 0xe0 -- Sprite 0x23
      11'h119: dout  = 8'b11000000; //  281 : 192 - 0xc0
      11'h11A: dout  = 8'b00111100; //  282 :  60 - 0x3c
      11'h11B: dout  = 8'b01111100; //  283 : 124 - 0x7c
      11'h11C: dout  = 8'b01111100; //  284 : 124 - 0x7c
      11'h11D: dout  = 8'b01111100; //  285 : 124 - 0x7c
      11'h11E: dout  = 8'b11101100; //  286 : 236 - 0xec
      11'h11F: dout  = 8'b11100000; //  287 : 224 - 0xe0
      11'h120: dout  = 8'b00000010; //  288 :   2 - 0x2 -- Sprite 0x24
      11'h121: dout  = 8'b00000101; //  289 :   5 - 0x5
      11'h122: dout  = 8'b00001011; //  290 :  11 - 0xb
      11'h123: dout  = 8'b00001011; //  291 :  11 - 0xb
      11'h124: dout  = 8'b00001101; //  292 :  13 - 0xd
      11'h125: dout  = 8'b00011000; //  293 :  24 - 0x18
      11'h126: dout  = 8'b00111000; //  294 :  56 - 0x38
      11'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      11'h128: dout  = 8'b11100000; //  296 : 224 - 0xe0 -- Sprite 0x25
      11'h129: dout  = 8'b11100000; //  297 : 224 - 0xe0
      11'h12A: dout  = 8'b11100000; //  298 : 224 - 0xe0
      11'h12B: dout  = 8'b11010000; //  299 : 208 - 0xd0
      11'h12C: dout  = 8'b10111000; //  300 : 184 - 0xb8
      11'h12D: dout  = 8'b00111000; //  301 :  56 - 0x38
      11'h12E: dout  = 8'b00000000; //  302 :   0 - 0x0
      11'h12F: dout  = 8'b00000000; //  303 :   0 - 0x0
      11'h130: dout  = 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      11'h131: dout  = 8'b00000000; //  305 :   0 - 0x0
      11'h132: dout  = 8'b00000000; //  306 :   0 - 0x0
      11'h133: dout  = 8'b00000000; //  307 :   0 - 0x0
      11'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      11'h135: dout  = 8'b00000000; //  309 :   0 - 0x0
      11'h136: dout  = 8'b00000000; //  310 :   0 - 0x0
      11'h137: dout  = 8'b00000000; //  311 :   0 - 0x0
      11'h138: dout  = 8'b00000000; //  312 :   0 - 0x0 -- Sprite 0x27
      11'h139: dout  = 8'b00000000; //  313 :   0 - 0x0
      11'h13A: dout  = 8'b00000000; //  314 :   0 - 0x0
      11'h13B: dout  = 8'b00000000; //  315 :   0 - 0x0
      11'h13C: dout  = 8'b00000000; //  316 :   0 - 0x0
      11'h13D: dout  = 8'b00000000; //  317 :   0 - 0x0
      11'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      11'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      11'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      11'h141: dout  = 8'b00000000; //  321 :   0 - 0x0
      11'h142: dout  = 8'b00000000; //  322 :   0 - 0x0
      11'h143: dout  = 8'b00000000; //  323 :   0 - 0x0
      11'h144: dout  = 8'b00000000; //  324 :   0 - 0x0
      11'h145: dout  = 8'b00000000; //  325 :   0 - 0x0
      11'h146: dout  = 8'b00000000; //  326 :   0 - 0x0
      11'h147: dout  = 8'b00000000; //  327 :   0 - 0x0
      11'h148: dout  = 8'b00011111; //  328 :  31 - 0x1f -- Sprite 0x29
      11'h149: dout  = 8'b00011111; //  329 :  31 - 0x1f
      11'h14A: dout  = 8'b00011111; //  330 :  31 - 0x1f
      11'h14B: dout  = 8'b00011111; //  331 :  31 - 0x1f
      11'h14C: dout  = 8'b00001100; //  332 :  12 - 0xc
      11'h14D: dout  = 8'b00000000; //  333 :   0 - 0x0
      11'h14E: dout  = 8'b00000001; //  334 :   1 - 0x1
      11'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      11'h150: dout  = 8'b00011111; //  336 :  31 - 0x1f -- Sprite 0x2a
      11'h151: dout  = 8'b00011111; //  337 :  31 - 0x1f
      11'h152: dout  = 8'b00011111; //  338 :  31 - 0x1f
      11'h153: dout  = 8'b00011111; //  339 :  31 - 0x1f
      11'h154: dout  = 8'b00001100; //  340 :  12 - 0xc
      11'h155: dout  = 8'b00000000; //  341 :   0 - 0x0
      11'h156: dout  = 8'b00000000; //  342 :   0 - 0x0
      11'h157: dout  = 8'b00000000; //  343 :   0 - 0x0
      11'h158: dout  = 8'b00000000; //  344 :   0 - 0x0 -- Sprite 0x2b
      11'h159: dout  = 8'b00000000; //  345 :   0 - 0x0
      11'h15A: dout  = 8'b00000000; //  346 :   0 - 0x0
      11'h15B: dout  = 8'b00000000; //  347 :   0 - 0x0
      11'h15C: dout  = 8'b00000000; //  348 :   0 - 0x0
      11'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      11'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      11'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      11'h160: dout  = 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x2c
      11'h161: dout  = 8'b00000000; //  353 :   0 - 0x0
      11'h162: dout  = 8'b00000000; //  354 :   0 - 0x0
      11'h163: dout  = 8'b00000000; //  355 :   0 - 0x0
      11'h164: dout  = 8'b00000000; //  356 :   0 - 0x0
      11'h165: dout  = 8'b00000000; //  357 :   0 - 0x0
      11'h166: dout  = 8'b00000000; //  358 :   0 - 0x0
      11'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      11'h168: dout  = 8'b00000000; //  360 :   0 - 0x0 -- Sprite 0x2d
      11'h169: dout  = 8'b01111110; //  361 : 126 - 0x7e
      11'h16A: dout  = 8'b01000010; //  362 :  66 - 0x42
      11'h16B: dout  = 8'b01000010; //  363 :  66 - 0x42
      11'h16C: dout  = 8'b01000010; //  364 :  66 - 0x42
      11'h16D: dout  = 8'b01000010; //  365 :  66 - 0x42
      11'h16E: dout  = 8'b01111110; //  366 : 126 - 0x7e
      11'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      11'h170: dout  = 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x2e
      11'h171: dout  = 8'b00000000; //  369 :   0 - 0x0
      11'h172: dout  = 8'b00000000; //  370 :   0 - 0x0
      11'h173: dout  = 8'b00000000; //  371 :   0 - 0x0
      11'h174: dout  = 8'b00000000; //  372 :   0 - 0x0
      11'h175: dout  = 8'b00000000; //  373 :   0 - 0x0
      11'h176: dout  = 8'b00000000; //  374 :   0 - 0x0
      11'h177: dout  = 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout  = 8'b01100110; //  376 : 102 - 0x66 -- Sprite 0x2f
      11'h179: dout  = 8'b01100000; //  377 :  96 - 0x60
      11'h17A: dout  = 8'b01101000; //  378 : 104 - 0x68
      11'h17B: dout  = 8'b11100000; //  379 : 224 - 0xe0
      11'h17C: dout  = 8'b11000000; //  380 : 192 - 0xc0
      11'h17D: dout  = 8'b00010000; //  381 :  16 - 0x10
      11'h17E: dout  = 8'b00101000; //  382 :  40 - 0x28
      11'h17F: dout  = 8'b01010000; //  383 :  80 - 0x50
      11'h180: dout  = 8'b11110110; //  384 : 246 - 0xf6 -- Sprite 0x30
      11'h181: dout  = 8'b11110000; //  385 : 240 - 0xf0
      11'h182: dout  = 8'b00111000; //  386 :  56 - 0x38
      11'h183: dout  = 8'b11010000; //  387 : 208 - 0xd0
      11'h184: dout  = 8'b11000000; //  388 : 192 - 0xc0
      11'h185: dout  = 8'b11111000; //  389 : 248 - 0xf8
      11'h186: dout  = 8'b01111000; //  390 : 120 - 0x78
      11'h187: dout  = 8'b00000000; //  391 :   0 - 0x0
      11'h188: dout  = 8'b11110110; //  392 : 246 - 0xf6 -- Sprite 0x31
      11'h189: dout  = 8'b11110000; //  393 : 240 - 0xf0
      11'h18A: dout  = 8'b00111000; //  394 :  56 - 0x38
      11'h18B: dout  = 8'b11010000; //  395 : 208 - 0xd0
      11'h18C: dout  = 8'b11000000; //  396 : 192 - 0xc0
      11'h18D: dout  = 8'b11100000; //  397 : 224 - 0xe0
      11'h18E: dout  = 8'b01111000; //  398 : 120 - 0x78
      11'h18F: dout  = 8'b00111000; //  399 :  56 - 0x38
      11'h190: dout  = 8'b11110110; //  400 : 246 - 0xf6 -- Sprite 0x32
      11'h191: dout  = 8'b11110000; //  401 : 240 - 0xf0
      11'h192: dout  = 8'b00111000; //  402 :  56 - 0x38
      11'h193: dout  = 8'b11000000; //  403 : 192 - 0xc0
      11'h194: dout  = 8'b11011000; //  404 : 216 - 0xd8
      11'h195: dout  = 8'b11111000; //  405 : 248 - 0xf8
      11'h196: dout  = 8'b01100000; //  406 :  96 - 0x60
      11'h197: dout  = 8'b00010000; //  407 :  16 - 0x10
      11'h198: dout  = 8'b00011100; //  408 :  28 - 0x1c -- Sprite 0x33
      11'h199: dout  = 8'b00011100; //  409 :  28 - 0x1c
      11'h19A: dout  = 8'b00011110; //  410 :  30 - 0x1e
      11'h19B: dout  = 8'b00011111; //  411 :  31 - 0x1f
      11'h19C: dout  = 8'b00001100; //  412 :  12 - 0xc
      11'h19D: dout  = 8'b00000000; //  413 :   0 - 0x0
      11'h19E: dout  = 8'b00000000; //  414 :   0 - 0x0
      11'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      11'h1A0: dout  = 8'b10000000; //  416 : 128 - 0x80 -- Sprite 0x34
      11'h1A1: dout  = 8'b01010000; //  417 :  80 - 0x50
      11'h1A2: dout  = 8'b10101000; //  418 : 168 - 0xa8
      11'h1A3: dout  = 8'b00000000; //  419 :   0 - 0x0
      11'h1A4: dout  = 8'b01011000; //  420 :  88 - 0x58
      11'h1A5: dout  = 8'b11011000; //  421 : 216 - 0xd8
      11'h1A6: dout  = 8'b11101100; //  422 : 236 - 0xec
      11'h1A7: dout  = 8'b00000000; //  423 :   0 - 0x0
      11'h1A8: dout  = 8'b00011100; //  424 :  28 - 0x1c -- Sprite 0x35
      11'h1A9: dout  = 8'b00011100; //  425 :  28 - 0x1c
      11'h1AA: dout  = 8'b00011110; //  426 :  30 - 0x1e
      11'h1AB: dout  = 8'b00011111; //  427 :  31 - 0x1f
      11'h1AC: dout  = 8'b00001100; //  428 :  12 - 0xc
      11'h1AD: dout  = 8'b00000001; //  429 :   1 - 0x1
      11'h1AE: dout  = 8'b00000001; //  430 :   1 - 0x1
      11'h1AF: dout  = 8'b00000000; //  431 :   0 - 0x0
      11'h1B0: dout  = 8'b10101000; //  432 : 168 - 0xa8 -- Sprite 0x36
      11'h1B1: dout  = 8'b01010000; //  433 :  80 - 0x50
      11'h1B2: dout  = 8'b10101000; //  434 : 168 - 0xa8
      11'h1B3: dout  = 8'b00000000; //  435 :   0 - 0x0
      11'h1B4: dout  = 8'b01011000; //  436 :  88 - 0x58
      11'h1B5: dout  = 8'b11001110; //  437 : 206 - 0xce
      11'h1B6: dout  = 8'b10000110; //  438 : 134 - 0x86
      11'h1B7: dout  = 8'b00000000; //  439 :   0 - 0x0
      11'h1B8: dout  = 8'b10101000; //  440 : 168 - 0xa8 -- Sprite 0x37
      11'h1B9: dout  = 8'b01010000; //  441 :  80 - 0x50
      11'h1BA: dout  = 8'b10101000; //  442 : 168 - 0xa8
      11'h1BB: dout  = 8'b00000000; //  443 :   0 - 0x0
      11'h1BC: dout  = 8'b01011000; //  444 :  88 - 0x58
      11'h1BD: dout  = 8'b11011000; //  445 : 216 - 0xd8
      11'h1BE: dout  = 8'b11101100; //  446 : 236 - 0xec
      11'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      11'h1C0: dout  = 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      11'h1C1: dout  = 8'b00000000; //  449 :   0 - 0x0
      11'h1C2: dout  = 8'b00000000; //  450 :   0 - 0x0
      11'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      11'h1C4: dout  = 8'b00000000; //  452 :   0 - 0x0
      11'h1C5: dout  = 8'b00000000; //  453 :   0 - 0x0
      11'h1C6: dout  = 8'b00000000; //  454 :   0 - 0x0
      11'h1C7: dout  = 8'b00000000; //  455 :   0 - 0x0
      11'h1C8: dout  = 8'b00000000; //  456 :   0 - 0x0 -- Sprite 0x39
      11'h1C9: dout  = 8'b00000000; //  457 :   0 - 0x0
      11'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      11'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      11'h1CC: dout  = 8'b00000000; //  460 :   0 - 0x0
      11'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      11'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      11'h1D2: dout  = 8'b00000000; //  466 :   0 - 0x0
      11'h1D3: dout  = 8'b00000000; //  467 :   0 - 0x0
      11'h1D4: dout  = 8'b00000000; //  468 :   0 - 0x0
      11'h1D5: dout  = 8'b00000000; //  469 :   0 - 0x0
      11'h1D6: dout  = 8'b00000000; //  470 :   0 - 0x0
      11'h1D7: dout  = 8'b00000000; //  471 :   0 - 0x0
      11'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0 -- Sprite 0x3b
      11'h1D9: dout  = 8'b00000000; //  473 :   0 - 0x0
      11'h1DA: dout  = 8'b00000000; //  474 :   0 - 0x0
      11'h1DB: dout  = 8'b00000000; //  475 :   0 - 0x0
      11'h1DC: dout  = 8'b00000000; //  476 :   0 - 0x0
      11'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      11'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      11'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      11'h1E1: dout  = 8'b00000000; //  481 :   0 - 0x0
      11'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      11'h1E3: dout  = 8'b00000000; //  483 :   0 - 0x0
      11'h1E4: dout  = 8'b00000000; //  484 :   0 - 0x0
      11'h1E5: dout  = 8'b00000000; //  485 :   0 - 0x0
      11'h1E6: dout  = 8'b00000000; //  486 :   0 - 0x0
      11'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      11'h1E9: dout  = 8'b00000000; //  489 :   0 - 0x0
      11'h1EA: dout  = 8'b00000000; //  490 :   0 - 0x0
      11'h1EB: dout  = 8'b00000000; //  491 :   0 - 0x0
      11'h1EC: dout  = 8'b00000000; //  492 :   0 - 0x0
      11'h1ED: dout  = 8'b00000000; //  493 :   0 - 0x0
      11'h1EE: dout  = 8'b00000000; //  494 :   0 - 0x0
      11'h1EF: dout  = 8'b00000000; //  495 :   0 - 0x0
      11'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      11'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      11'h1F2: dout  = 8'b00000000; //  498 :   0 - 0x0
      11'h1F3: dout  = 8'b00000000; //  499 :   0 - 0x0
      11'h1F4: dout  = 8'b00000000; //  500 :   0 - 0x0
      11'h1F5: dout  = 8'b00000000; //  501 :   0 - 0x0
      11'h1F6: dout  = 8'b00000000; //  502 :   0 - 0x0
      11'h1F7: dout  = 8'b00000000; //  503 :   0 - 0x0
      11'h1F8: dout  = 8'b00000000; //  504 :   0 - 0x0 -- Sprite 0x3f
      11'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      11'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      11'h1FB: dout  = 8'b00000000; //  507 :   0 - 0x0
      11'h1FC: dout  = 8'b00000000; //  508 :   0 - 0x0
      11'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      11'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      11'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      11'h200: dout  = 8'b00111100; //  512 :  60 - 0x3c -- Sprite 0x40
      11'h201: dout  = 8'b01111100; //  513 : 124 - 0x7c
      11'h202: dout  = 8'b11100110; //  514 : 230 - 0xe6
      11'h203: dout  = 8'b11101110; //  515 : 238 - 0xee
      11'h204: dout  = 8'b11110110; //  516 : 246 - 0xf6
      11'h205: dout  = 8'b11100110; //  517 : 230 - 0xe6
      11'h206: dout  = 8'b00111100; //  518 :  60 - 0x3c
      11'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      11'h208: dout  = 8'b00111000; //  520 :  56 - 0x38 -- Sprite 0x41
      11'h209: dout  = 8'b01111000; //  521 : 120 - 0x78
      11'h20A: dout  = 8'b00111000; //  522 :  56 - 0x38
      11'h20B: dout  = 8'b00111000; //  523 :  56 - 0x38
      11'h20C: dout  = 8'b00111000; //  524 :  56 - 0x38
      11'h20D: dout  = 8'b00111000; //  525 :  56 - 0x38
      11'h20E: dout  = 8'b00111000; //  526 :  56 - 0x38
      11'h20F: dout  = 8'b00000000; //  527 :   0 - 0x0
      11'h210: dout  = 8'b01111100; //  528 : 124 - 0x7c -- Sprite 0x42
      11'h211: dout  = 8'b11111110; //  529 : 254 - 0xfe
      11'h212: dout  = 8'b11100110; //  530 : 230 - 0xe6
      11'h213: dout  = 8'b00011110; //  531 :  30 - 0x1e
      11'h214: dout  = 8'b01111100; //  532 : 124 - 0x7c
      11'h215: dout  = 8'b11100000; //  533 : 224 - 0xe0
      11'h216: dout  = 8'b11111110; //  534 : 254 - 0xfe
      11'h217: dout  = 8'b00000000; //  535 :   0 - 0x0
      11'h218: dout  = 8'b01111100; //  536 : 124 - 0x7c -- Sprite 0x43
      11'h219: dout  = 8'b11111100; //  537 : 252 - 0xfc
      11'h21A: dout  = 8'b11100110; //  538 : 230 - 0xe6
      11'h21B: dout  = 8'b00011100; //  539 :  28 - 0x1c
      11'h21C: dout  = 8'b01100110; //  540 : 102 - 0x66
      11'h21D: dout  = 8'b11101110; //  541 : 238 - 0xee
      11'h21E: dout  = 8'b11111100; //  542 : 252 - 0xfc
      11'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      11'h220: dout  = 8'b00001100; //  544 :  12 - 0xc -- Sprite 0x44
      11'h221: dout  = 8'b00011100; //  545 :  28 - 0x1c
      11'h222: dout  = 8'b00111100; //  546 :  60 - 0x3c
      11'h223: dout  = 8'b01111100; //  547 : 124 - 0x7c
      11'h224: dout  = 8'b11101100; //  548 : 236 - 0xec
      11'h225: dout  = 8'b11111110; //  549 : 254 - 0xfe
      11'h226: dout  = 8'b00001100; //  550 :  12 - 0xc
      11'h227: dout  = 8'b00000000; //  551 :   0 - 0x0
      11'h228: dout  = 8'b11111110; //  552 : 254 - 0xfe -- Sprite 0x45
      11'h229: dout  = 8'b11111110; //  553 : 254 - 0xfe
      11'h22A: dout  = 8'b11100000; //  554 : 224 - 0xe0
      11'h22B: dout  = 8'b11111110; //  555 : 254 - 0xfe
      11'h22C: dout  = 8'b00000110; //  556 :   6 - 0x6
      11'h22D: dout  = 8'b11101110; //  557 : 238 - 0xee
      11'h22E: dout  = 8'b11111100; //  558 : 252 - 0xfc
      11'h22F: dout  = 8'b00000000; //  559 :   0 - 0x0
      11'h230: dout  = 8'b00111100; //  560 :  60 - 0x3c -- Sprite 0x46
      11'h231: dout  = 8'b01111100; //  561 : 124 - 0x7c
      11'h232: dout  = 8'b11100000; //  562 : 224 - 0xe0
      11'h233: dout  = 8'b11111110; //  563 : 254 - 0xfe
      11'h234: dout  = 8'b11100110; //  564 : 230 - 0xe6
      11'h235: dout  = 8'b11101110; //  565 : 238 - 0xee
      11'h236: dout  = 8'b00111100; //  566 :  60 - 0x3c
      11'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      11'h238: dout  = 8'b11111110; //  568 : 254 - 0xfe -- Sprite 0x47
      11'h239: dout  = 8'b11111100; //  569 : 252 - 0xfc
      11'h23A: dout  = 8'b00001100; //  570 :  12 - 0xc
      11'h23B: dout  = 8'b00111000; //  571 :  56 - 0x38
      11'h23C: dout  = 8'b00111000; //  572 :  56 - 0x38
      11'h23D: dout  = 8'b01110000; //  573 : 112 - 0x70
      11'h23E: dout  = 8'b01110000; //  574 : 112 - 0x70
      11'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout  = 8'b00111110; //  576 :  62 - 0x3e -- Sprite 0x48
      11'h241: dout  = 8'b01111100; //  577 : 124 - 0x7c
      11'h242: dout  = 8'b11100110; //  578 : 230 - 0xe6
      11'h243: dout  = 8'b10111100; //  579 : 188 - 0xbc
      11'h244: dout  = 8'b11100110; //  580 : 230 - 0xe6
      11'h245: dout  = 8'b11101110; //  581 : 238 - 0xee
      11'h246: dout  = 8'b00111100; //  582 :  60 - 0x3c
      11'h247: dout  = 8'b00000000; //  583 :   0 - 0x0
      11'h248: dout  = 8'b00111100; //  584 :  60 - 0x3c -- Sprite 0x49
      11'h249: dout  = 8'b01111100; //  585 : 124 - 0x7c
      11'h24A: dout  = 8'b11100110; //  586 : 230 - 0xe6
      11'h24B: dout  = 8'b11101110; //  587 : 238 - 0xee
      11'h24C: dout  = 8'b11111110; //  588 : 254 - 0xfe
      11'h24D: dout  = 8'b10000110; //  589 : 134 - 0x86
      11'h24E: dout  = 8'b01111100; //  590 : 124 - 0x7c
      11'h24F: dout  = 8'b01000000; //  591 :  64 - 0x40
      11'h250: dout  = 8'b11101110; //  592 : 238 - 0xee -- Sprite 0x4a
      11'h251: dout  = 8'b11101110; //  593 : 238 - 0xee
      11'h252: dout  = 8'b11101110; //  594 : 238 - 0xee
      11'h253: dout  = 8'b11101110; //  595 : 238 - 0xee
      11'h254: dout  = 8'b11101110; //  596 : 238 - 0xee
      11'h255: dout  = 8'b11101110; //  597 : 238 - 0xee
      11'h256: dout  = 8'b11101110; //  598 : 238 - 0xee
      11'h257: dout  = 8'b10001000; //  599 : 136 - 0x88
      11'h258: dout  = 8'b11100000; //  600 : 224 - 0xe0 -- Sprite 0x4b
      11'h259: dout  = 8'b11100000; //  601 : 224 - 0xe0
      11'h25A: dout  = 8'b11100000; //  602 : 224 - 0xe0
      11'h25B: dout  = 8'b11100000; //  603 : 224 - 0xe0
      11'h25C: dout  = 8'b11100000; //  604 : 224 - 0xe0
      11'h25D: dout  = 8'b11100000; //  605 : 224 - 0xe0
      11'h25E: dout  = 8'b11100000; //  606 : 224 - 0xe0
      11'h25F: dout  = 8'b10000000; //  607 : 128 - 0x80
      11'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x4c
      11'h261: dout  = 8'b01111111; //  609 : 127 - 0x7f
      11'h262: dout  = 8'b01111111; //  610 : 127 - 0x7f
      11'h263: dout  = 8'b01111111; //  611 : 127 - 0x7f
      11'h264: dout  = 8'b01111111; //  612 : 127 - 0x7f
      11'h265: dout  = 8'b01111111; //  613 : 127 - 0x7f
      11'h266: dout  = 8'b01111111; //  614 : 127 - 0x7f
      11'h267: dout  = 8'b01111111; //  615 : 127 - 0x7f
      11'h268: dout  = 8'b01111111; //  616 : 127 - 0x7f -- Sprite 0x4d
      11'h269: dout  = 8'b01111111; //  617 : 127 - 0x7f
      11'h26A: dout  = 8'b01111111; //  618 : 127 - 0x7f
      11'h26B: dout  = 8'b01111111; //  619 : 127 - 0x7f
      11'h26C: dout  = 8'b01111111; //  620 : 127 - 0x7f
      11'h26D: dout  = 8'b01111111; //  621 : 127 - 0x7f
      11'h26E: dout  = 8'b01111111; //  622 : 127 - 0x7f
      11'h26F: dout  = 8'b00000000; //  623 :   0 - 0x0
      11'h270: dout  = 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x4e
      11'h271: dout  = 8'b11111110; //  625 : 254 - 0xfe
      11'h272: dout  = 8'b11111110; //  626 : 254 - 0xfe
      11'h273: dout  = 8'b11111110; //  627 : 254 - 0xfe
      11'h274: dout  = 8'b11111110; //  628 : 254 - 0xfe
      11'h275: dout  = 8'b11111110; //  629 : 254 - 0xfe
      11'h276: dout  = 8'b11111110; //  630 : 254 - 0xfe
      11'h277: dout  = 8'b11111110; //  631 : 254 - 0xfe
      11'h278: dout  = 8'b11111110; //  632 : 254 - 0xfe -- Sprite 0x4f
      11'h279: dout  = 8'b11111110; //  633 : 254 - 0xfe
      11'h27A: dout  = 8'b11111110; //  634 : 254 - 0xfe
      11'h27B: dout  = 8'b11111110; //  635 : 254 - 0xfe
      11'h27C: dout  = 8'b11111110; //  636 : 254 - 0xfe
      11'h27D: dout  = 8'b11111110; //  637 : 254 - 0xfe
      11'h27E: dout  = 8'b11111110; //  638 : 254 - 0xfe
      11'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      11'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x50
      11'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      11'h282: dout  = 8'b00000000; //  642 :   0 - 0x0
      11'h283: dout  = 8'b00000000; //  643 :   0 - 0x0
      11'h284: dout  = 8'b00000000; //  644 :   0 - 0x0
      11'h285: dout  = 8'b00000000; //  645 :   0 - 0x0
      11'h286: dout  = 8'b00000000; //  646 :   0 - 0x0
      11'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      11'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- Sprite 0x51
      11'h289: dout  = 8'b00010000; //  649 :  16 - 0x10
      11'h28A: dout  = 8'b00010000; //  650 :  16 - 0x10
      11'h28B: dout  = 8'b01111100; //  651 : 124 - 0x7c
      11'h28C: dout  = 8'b00111000; //  652 :  56 - 0x38
      11'h28D: dout  = 8'b00111000; //  653 :  56 - 0x38
      11'h28E: dout  = 8'b01101100; //  654 : 108 - 0x6c
      11'h28F: dout  = 8'b00000000; //  655 :   0 - 0x0
      11'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      11'h291: dout  = 8'b00010000; //  657 :  16 - 0x10
      11'h292: dout  = 8'b00010000; //  658 :  16 - 0x10
      11'h293: dout  = 8'b01111100; //  659 : 124 - 0x7c
      11'h294: dout  = 8'b00111000; //  660 :  56 - 0x38
      11'h295: dout  = 8'b00111000; //  661 :  56 - 0x38
      11'h296: dout  = 8'b01101100; //  662 : 108 - 0x6c
      11'h297: dout  = 8'b00000000; //  663 :   0 - 0x0
      11'h298: dout  = 8'b00000000; //  664 :   0 - 0x0 -- Sprite 0x53
      11'h299: dout  = 8'b00000000; //  665 :   0 - 0x0
      11'h29A: dout  = 8'b00000000; //  666 :   0 - 0x0
      11'h29B: dout  = 8'b00000000; //  667 :   0 - 0x0
      11'h29C: dout  = 8'b00000000; //  668 :   0 - 0x0
      11'h29D: dout  = 8'b00000000; //  669 :   0 - 0x0
      11'h29E: dout  = 8'b00000000; //  670 :   0 - 0x0
      11'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      11'h2A0: dout  = 8'b11111111; //  672 : 255 - 0xff -- Sprite 0x54
      11'h2A1: dout  = 8'b11111111; //  673 : 255 - 0xff
      11'h2A2: dout  = 8'b11111111; //  674 : 255 - 0xff
      11'h2A3: dout  = 8'b11111111; //  675 : 255 - 0xff
      11'h2A4: dout  = 8'b11111111; //  676 : 255 - 0xff
      11'h2A5: dout  = 8'b11111111; //  677 : 255 - 0xff
      11'h2A6: dout  = 8'b11111111; //  678 : 255 - 0xff
      11'h2A7: dout  = 8'b11111111; //  679 : 255 - 0xff
      11'h2A8: dout  = 8'b11111111; //  680 : 255 - 0xff -- Sprite 0x55
      11'h2A9: dout  = 8'b11111111; //  681 : 255 - 0xff
      11'h2AA: dout  = 8'b11111111; //  682 : 255 - 0xff
      11'h2AB: dout  = 8'b11111111; //  683 : 255 - 0xff
      11'h2AC: dout  = 8'b11111111; //  684 : 255 - 0xff
      11'h2AD: dout  = 8'b11111111; //  685 : 255 - 0xff
      11'h2AE: dout  = 8'b11111111; //  686 : 255 - 0xff
      11'h2AF: dout  = 8'b11111111; //  687 : 255 - 0xff
      11'h2B0: dout  = 8'b00000010; //  688 :   2 - 0x2 -- Sprite 0x56
      11'h2B1: dout  = 8'b00000101; //  689 :   5 - 0x5
      11'h2B2: dout  = 8'b10101010; //  690 : 170 - 0xaa
      11'h2B3: dout  = 8'b01010001; //  691 :  81 - 0x51
      11'h2B4: dout  = 8'b10101010; //  692 : 170 - 0xaa
      11'h2B5: dout  = 8'b01010001; //  693 :  81 - 0x51
      11'h2B6: dout  = 8'b10100010; //  694 : 162 - 0xa2
      11'h2B7: dout  = 8'b00000100; //  695 :   4 - 0x4
      11'h2B8: dout  = 8'b00001000; //  696 :   8 - 0x8 -- Sprite 0x57
      11'h2B9: dout  = 8'b01010101; //  697 :  85 - 0x55
      11'h2BA: dout  = 8'b00101010; //  698 :  42 - 0x2a
      11'h2BB: dout  = 8'b01010101; //  699 :  85 - 0x55
      11'h2BC: dout  = 8'b00101010; //  700 :  42 - 0x2a
      11'h2BD: dout  = 8'b01000101; //  701 :  69 - 0x45
      11'h2BE: dout  = 8'b00001010; //  702 :  10 - 0xa
      11'h2BF: dout  = 8'b00010000; //  703 :  16 - 0x10
      11'h2C0: dout  = 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x58
      11'h2C1: dout  = 8'b00111111; //  705 :  63 - 0x3f
      11'h2C2: dout  = 8'b01011111; //  706 :  95 - 0x5f
      11'h2C3: dout  = 8'b01101111; //  707 : 111 - 0x6f
      11'h2C4: dout  = 8'b01110000; //  708 : 112 - 0x70
      11'h2C5: dout  = 8'b01110111; //  709 : 119 - 0x77
      11'h2C6: dout  = 8'b01110111; //  710 : 119 - 0x77
      11'h2C7: dout  = 8'b01110111; //  711 : 119 - 0x77
      11'h2C8: dout  = 8'b01110111; //  712 : 119 - 0x77 -- Sprite 0x59
      11'h2C9: dout  = 8'b01110111; //  713 : 119 - 0x77
      11'h2CA: dout  = 8'b01110111; //  714 : 119 - 0x77
      11'h2CB: dout  = 8'b01110000; //  715 : 112 - 0x70
      11'h2CC: dout  = 8'b01101111; //  716 : 111 - 0x6f
      11'h2CD: dout  = 8'b01011111; //  717 :  95 - 0x5f
      11'h2CE: dout  = 8'b00010101; //  718 :  21 - 0x15
      11'h2CF: dout  = 8'b00000000; //  719 :   0 - 0x0
      11'h2D0: dout  = 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x5a
      11'h2D1: dout  = 8'b11111100; //  721 : 252 - 0xfc
      11'h2D2: dout  = 8'b11111000; //  722 : 248 - 0xf8
      11'h2D3: dout  = 8'b11110110; //  723 : 246 - 0xf6
      11'h2D4: dout  = 8'b00001100; //  724 :  12 - 0xc
      11'h2D5: dout  = 8'b11101110; //  725 : 238 - 0xee
      11'h2D6: dout  = 8'b11101100; //  726 : 236 - 0xec
      11'h2D7: dout  = 8'b11101110; //  727 : 238 - 0xee
      11'h2D8: dout  = 8'b11101100; //  728 : 236 - 0xec -- Sprite 0x5b
      11'h2D9: dout  = 8'b11101110; //  729 : 238 - 0xee
      11'h2DA: dout  = 8'b11101100; //  730 : 236 - 0xec
      11'h2DB: dout  = 8'b00001110; //  731 :  14 - 0xe
      11'h2DC: dout  = 8'b11110100; //  732 : 244 - 0xf4
      11'h2DD: dout  = 8'b11111010; //  733 : 250 - 0xfa
      11'h2DE: dout  = 8'b01010100; //  734 :  84 - 0x54
      11'h2DF: dout  = 8'b00000000; //  735 :   0 - 0x0
      11'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x5c
      11'h2E1: dout  = 8'b00011100; //  737 :  28 - 0x1c
      11'h2E2: dout  = 8'b00111110; //  738 :  62 - 0x3e
      11'h2E3: dout  = 8'b00111110; //  739 :  62 - 0x3e
      11'h2E4: dout  = 8'b00111110; //  740 :  62 - 0x3e
      11'h2E5: dout  = 8'b00011100; //  741 :  28 - 0x1c
      11'h2E6: dout  = 8'b00011100; //  742 :  28 - 0x1c
      11'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      11'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0 -- Sprite 0x5d
      11'h2E9: dout  = 8'b00000000; //  745 :   0 - 0x0
      11'h2EA: dout  = 8'b00000000; //  746 :   0 - 0x0
      11'h2EB: dout  = 8'b00000000; //  747 :   0 - 0x0
      11'h2EC: dout  = 8'b00000000; //  748 :   0 - 0x0
      11'h2ED: dout  = 8'b00000000; //  749 :   0 - 0x0
      11'h2EE: dout  = 8'b00000000; //  750 :   0 - 0x0
      11'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      11'h2F0: dout  = 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x5e
      11'h2F1: dout  = 8'b00010100; //  753 :  20 - 0x14
      11'h2F2: dout  = 8'b00110110; //  754 :  54 - 0x36
      11'h2F3: dout  = 8'b00111110; //  755 :  62 - 0x3e
      11'h2F4: dout  = 8'b00111110; //  756 :  62 - 0x3e
      11'h2F5: dout  = 8'b00011100; //  757 :  28 - 0x1c
      11'h2F6: dout  = 8'b00001000; //  758 :   8 - 0x8
      11'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      11'h2F8: dout  = 8'b00000000; //  760 :   0 - 0x0 -- Sprite 0x5f
      11'h2F9: dout  = 8'b00010100; //  761 :  20 - 0x14
      11'h2FA: dout  = 8'b00011100; //  762 :  28 - 0x1c
      11'h2FB: dout  = 8'b00011100; //  763 :  28 - 0x1c
      11'h2FC: dout  = 8'b00011100; //  764 :  28 - 0x1c
      11'h2FD: dout  = 8'b00011100; //  765 :  28 - 0x1c
      11'h2FE: dout  = 8'b00011100; //  766 :  28 - 0x1c
      11'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      11'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      11'h301: dout  = 8'b01111111; //  769 : 127 - 0x7f
      11'h302: dout  = 8'b01111111; //  770 : 127 - 0x7f
      11'h303: dout  = 8'b01111111; //  771 : 127 - 0x7f
      11'h304: dout  = 8'b01111111; //  772 : 127 - 0x7f
      11'h305: dout  = 8'b01111111; //  773 : 127 - 0x7f
      11'h306: dout  = 8'b00101010; //  774 :  42 - 0x2a
      11'h307: dout  = 8'b00000000; //  775 :   0 - 0x0
      11'h308: dout  = 8'b00000000; //  776 :   0 - 0x0 -- Sprite 0x61
      11'h309: dout  = 8'b11111111; //  777 : 255 - 0xff
      11'h30A: dout  = 8'b11111111; //  778 : 255 - 0xff
      11'h30B: dout  = 8'b11111111; //  779 : 255 - 0xff
      11'h30C: dout  = 8'b11111111; //  780 : 255 - 0xff
      11'h30D: dout  = 8'b11111111; //  781 : 255 - 0xff
      11'h30E: dout  = 8'b10101010; //  782 : 170 - 0xaa
      11'h30F: dout  = 8'b00000000; //  783 :   0 - 0x0
      11'h310: dout  = 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x62
      11'h311: dout  = 8'b11111110; //  785 : 254 - 0xfe
      11'h312: dout  = 8'b11111110; //  786 : 254 - 0xfe
      11'h313: dout  = 8'b11111110; //  787 : 254 - 0xfe
      11'h314: dout  = 8'b11111110; //  788 : 254 - 0xfe
      11'h315: dout  = 8'b11111110; //  789 : 254 - 0xfe
      11'h316: dout  = 8'b10101010; //  790 : 170 - 0xaa
      11'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      11'h318: dout  = 8'b00000000; //  792 :   0 - 0x0 -- Sprite 0x63
      11'h319: dout  = 8'b00000000; //  793 :   0 - 0x0
      11'h31A: dout  = 8'b00000000; //  794 :   0 - 0x0
      11'h31B: dout  = 8'b00000000; //  795 :   0 - 0x0
      11'h31C: dout  = 8'b00000000; //  796 :   0 - 0x0
      11'h31D: dout  = 8'b00000000; //  797 :   0 - 0x0
      11'h31E: dout  = 8'b00000000; //  798 :   0 - 0x0
      11'h31F: dout  = 8'b00000000; //  799 :   0 - 0x0
      11'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x64
      11'h321: dout  = 8'b00000000; //  801 :   0 - 0x0
      11'h322: dout  = 8'b00000001; //  802 :   1 - 0x1
      11'h323: dout  = 8'b00000001; //  803 :   1 - 0x1
      11'h324: dout  = 8'b00000011; //  804 :   3 - 0x3
      11'h325: dout  = 8'b00000011; //  805 :   3 - 0x3
      11'h326: dout  = 8'b00000111; //  806 :   7 - 0x7
      11'h327: dout  = 8'b00000111; //  807 :   7 - 0x7
      11'h328: dout  = 8'b00001111; //  808 :  15 - 0xf -- Sprite 0x65
      11'h329: dout  = 8'b00001111; //  809 :  15 - 0xf
      11'h32A: dout  = 8'b00011111; //  810 :  31 - 0x1f
      11'h32B: dout  = 8'b00011111; //  811 :  31 - 0x1f
      11'h32C: dout  = 8'b00111111; //  812 :  63 - 0x3f
      11'h32D: dout  = 8'b00111111; //  813 :  63 - 0x3f
      11'h32E: dout  = 8'b01010101; //  814 :  85 - 0x55
      11'h32F: dout  = 8'b00000000; //  815 :   0 - 0x0
      11'h330: dout  = 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x66
      11'h331: dout  = 8'b00000000; //  817 :   0 - 0x0
      11'h332: dout  = 8'b00000000; //  818 :   0 - 0x0
      11'h333: dout  = 8'b10000000; //  819 : 128 - 0x80
      11'h334: dout  = 8'b01000000; //  820 :  64 - 0x40
      11'h335: dout  = 8'b10000000; //  821 : 128 - 0x80
      11'h336: dout  = 8'b11000000; //  822 : 192 - 0xc0
      11'h337: dout  = 8'b11100000; //  823 : 224 - 0xe0
      11'h338: dout  = 8'b11010000; //  824 : 208 - 0xd0 -- Sprite 0x67
      11'h339: dout  = 8'b11100000; //  825 : 224 - 0xe0
      11'h33A: dout  = 8'b11110000; //  826 : 240 - 0xf0
      11'h33B: dout  = 8'b11101000; //  827 : 232 - 0xe8
      11'h33C: dout  = 8'b11110100; //  828 : 244 - 0xf4
      11'h33D: dout  = 8'b11111000; //  829 : 248 - 0xf8
      11'h33E: dout  = 8'b01010100; //  830 :  84 - 0x54
      11'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      11'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      11'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      11'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      11'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      11'h344: dout  = 8'b00000000; //  836 :   0 - 0x0
      11'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      11'h346: dout  = 8'b00000000; //  838 :   0 - 0x0
      11'h347: dout  = 8'b00000000; //  839 :   0 - 0x0
      11'h348: dout  = 8'b00000000; //  840 :   0 - 0x0 -- Sprite 0x69
      11'h349: dout  = 8'b00000000; //  841 :   0 - 0x0
      11'h34A: dout  = 8'b00000000; //  842 :   0 - 0x0
      11'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      11'h34C: dout  = 8'b00000000; //  844 :   0 - 0x0
      11'h34D: dout  = 8'b00000000; //  845 :   0 - 0x0
      11'h34E: dout  = 8'b00000000; //  846 :   0 - 0x0
      11'h34F: dout  = 8'b00000000; //  847 :   0 - 0x0
      11'h350: dout  = 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      11'h351: dout  = 8'b00000000; //  849 :   0 - 0x0
      11'h352: dout  = 8'b00000000; //  850 :   0 - 0x0
      11'h353: dout  = 8'b00000000; //  851 :   0 - 0x0
      11'h354: dout  = 8'b00000000; //  852 :   0 - 0x0
      11'h355: dout  = 8'b00000000; //  853 :   0 - 0x0
      11'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      11'h357: dout  = 8'b00000000; //  855 :   0 - 0x0
      11'h358: dout  = 8'b00000000; //  856 :   0 - 0x0 -- Sprite 0x6b
      11'h359: dout  = 8'b00000000; //  857 :   0 - 0x0
      11'h35A: dout  = 8'b00000000; //  858 :   0 - 0x0
      11'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      11'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      11'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      11'h35E: dout  = 8'b00000000; //  862 :   0 - 0x0
      11'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      11'h360: dout  = 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x6c
      11'h361: dout  = 8'b00000000; //  865 :   0 - 0x0
      11'h362: dout  = 8'b00000000; //  866 :   0 - 0x0
      11'h363: dout  = 8'b00000000; //  867 :   0 - 0x0
      11'h364: dout  = 8'b00000000; //  868 :   0 - 0x0
      11'h365: dout  = 8'b00000000; //  869 :   0 - 0x0
      11'h366: dout  = 8'b00000000; //  870 :   0 - 0x0
      11'h367: dout  = 8'b00000000; //  871 :   0 - 0x0
      11'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      11'h369: dout  = 8'b00000000; //  873 :   0 - 0x0
      11'h36A: dout  = 8'b00000000; //  874 :   0 - 0x0
      11'h36B: dout  = 8'b00000000; //  875 :   0 - 0x0
      11'h36C: dout  = 8'b00000000; //  876 :   0 - 0x0
      11'h36D: dout  = 8'b00000000; //  877 :   0 - 0x0
      11'h36E: dout  = 8'b00000000; //  878 :   0 - 0x0
      11'h36F: dout  = 8'b00000000; //  879 :   0 - 0x0
      11'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      11'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout  = 8'b00000000; //  882 :   0 - 0x0
      11'h373: dout  = 8'b00000000; //  883 :   0 - 0x0
      11'h374: dout  = 8'b00000000; //  884 :   0 - 0x0
      11'h375: dout  = 8'b00000000; //  885 :   0 - 0x0
      11'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      11'h377: dout  = 8'b00000000; //  887 :   0 - 0x0
      11'h378: dout  = 8'b00000000; //  888 :   0 - 0x0 -- Sprite 0x6f
      11'h379: dout  = 8'b00000000; //  889 :   0 - 0x0
      11'h37A: dout  = 8'b00000000; //  890 :   0 - 0x0
      11'h37B: dout  = 8'b00000000; //  891 :   0 - 0x0
      11'h37C: dout  = 8'b00000000; //  892 :   0 - 0x0
      11'h37D: dout  = 8'b00000000; //  893 :   0 - 0x0
      11'h37E: dout  = 8'b00000000; //  894 :   0 - 0x0
      11'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      11'h380: dout  = 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x70
      11'h381: dout  = 8'b00000000; //  897 :   0 - 0x0
      11'h382: dout  = 8'b00000000; //  898 :   0 - 0x0
      11'h383: dout  = 8'b00000000; //  899 :   0 - 0x0
      11'h384: dout  = 8'b00000000; //  900 :   0 - 0x0
      11'h385: dout  = 8'b00000000; //  901 :   0 - 0x0
      11'h386: dout  = 8'b00000000; //  902 :   0 - 0x0
      11'h387: dout  = 8'b00000000; //  903 :   0 - 0x0
      11'h388: dout  = 8'b00000000; //  904 :   0 - 0x0 -- Sprite 0x71
      11'h389: dout  = 8'b00000000; //  905 :   0 - 0x0
      11'h38A: dout  = 8'b00000000; //  906 :   0 - 0x0
      11'h38B: dout  = 8'b00000000; //  907 :   0 - 0x0
      11'h38C: dout  = 8'b00000000; //  908 :   0 - 0x0
      11'h38D: dout  = 8'b00000000; //  909 :   0 - 0x0
      11'h38E: dout  = 8'b00000000; //  910 :   0 - 0x0
      11'h38F: dout  = 8'b00000000; //  911 :   0 - 0x0
      11'h390: dout  = 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x72
      11'h391: dout  = 8'b00000000; //  913 :   0 - 0x0
      11'h392: dout  = 8'b00000000; //  914 :   0 - 0x0
      11'h393: dout  = 8'b00000000; //  915 :   0 - 0x0
      11'h394: dout  = 8'b00000000; //  916 :   0 - 0x0
      11'h395: dout  = 8'b00000000; //  917 :   0 - 0x0
      11'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      11'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      11'h398: dout  = 8'b00000000; //  920 :   0 - 0x0 -- Sprite 0x73
      11'h399: dout  = 8'b00000000; //  921 :   0 - 0x0
      11'h39A: dout  = 8'b00000000; //  922 :   0 - 0x0
      11'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      11'h39C: dout  = 8'b00000000; //  924 :   0 - 0x0
      11'h39D: dout  = 8'b00000000; //  925 :   0 - 0x0
      11'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      11'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      11'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x74
      11'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      11'h3A2: dout  = 8'b00000000; //  930 :   0 - 0x0
      11'h3A3: dout  = 8'b00000000; //  931 :   0 - 0x0
      11'h3A4: dout  = 8'b00000000; //  932 :   0 - 0x0
      11'h3A5: dout  = 8'b00000000; //  933 :   0 - 0x0
      11'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      11'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      11'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0 -- Sprite 0x75
      11'h3A9: dout  = 8'b00000000; //  937 :   0 - 0x0
      11'h3AA: dout  = 8'b00000000; //  938 :   0 - 0x0
      11'h3AB: dout  = 8'b00000000; //  939 :   0 - 0x0
      11'h3AC: dout  = 8'b00000000; //  940 :   0 - 0x0
      11'h3AD: dout  = 8'b00000000; //  941 :   0 - 0x0
      11'h3AE: dout  = 8'b00000000; //  942 :   0 - 0x0
      11'h3AF: dout  = 8'b00000000; //  943 :   0 - 0x0
      11'h3B0: dout  = 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x76
      11'h3B1: dout  = 8'b00000000; //  945 :   0 - 0x0
      11'h3B2: dout  = 8'b00000000; //  946 :   0 - 0x0
      11'h3B3: dout  = 8'b00000000; //  947 :   0 - 0x0
      11'h3B4: dout  = 8'b00000000; //  948 :   0 - 0x0
      11'h3B5: dout  = 8'b00000000; //  949 :   0 - 0x0
      11'h3B6: dout  = 8'b00000000; //  950 :   0 - 0x0
      11'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      11'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0 -- Sprite 0x77
      11'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      11'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      11'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      11'h3BC: dout  = 8'b00000000; //  956 :   0 - 0x0
      11'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      11'h3BE: dout  = 8'b00000000; //  958 :   0 - 0x0
      11'h3BF: dout  = 8'b00000000; //  959 :   0 - 0x0
      11'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x78
      11'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      11'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      11'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      11'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      11'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      11'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      11'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      11'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0 -- Sprite 0x79
      11'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      11'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      11'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      11'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      11'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      11'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      11'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      11'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x7a
      11'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      11'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      11'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      11'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      11'h3D5: dout  = 8'b00000000; //  981 :   0 - 0x0
      11'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      11'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      11'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0 -- Sprite 0x7b
      11'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      11'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      11'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      11'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      11'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      11'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      11'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      11'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      11'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      11'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      11'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      11'h3E4: dout  = 8'b00000000; //  996 :   0 - 0x0
      11'h3E5: dout  = 8'b00000000; //  997 :   0 - 0x0
      11'h3E6: dout  = 8'b00000000; //  998 :   0 - 0x0
      11'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      11'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- Sprite 0x7d
      11'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      11'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      11'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      11'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      11'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      11'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      11'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      11'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x7e
      11'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      11'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      11'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      11'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      11'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      11'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      11'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      11'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0 -- Sprite 0x7f
      11'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      11'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      11'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      11'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      11'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      11'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      11'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      11'h400: dout  = 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x80
      11'h401: dout  = 8'b00000011; // 1025 :   3 - 0x3
      11'h402: dout  = 8'b00001111; // 1026 :  15 - 0xf
      11'h403: dout  = 8'b00011111; // 1027 :  31 - 0x1f
      11'h404: dout  = 8'b00011111; // 1028 :  31 - 0x1f
      11'h405: dout  = 8'b00111111; // 1029 :  63 - 0x3f
      11'h406: dout  = 8'b00111111; // 1030 :  63 - 0x3f
      11'h407: dout  = 8'b00000000; // 1031 :   0 - 0x0
      11'h408: dout  = 8'b00000000; // 1032 :   0 - 0x0 -- Sprite 0x81
      11'h409: dout  = 8'b00000000; // 1033 :   0 - 0x0
      11'h40A: dout  = 8'b00000000; // 1034 :   0 - 0x0
      11'h40B: dout  = 8'b00000000; // 1035 :   0 - 0x0
      11'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      11'h40D: dout  = 8'b00000000; // 1037 :   0 - 0x0
      11'h40E: dout  = 8'b00000000; // 1038 :   0 - 0x0
      11'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      11'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x82
      11'h411: dout  = 8'b11000000; // 1041 : 192 - 0xc0
      11'h412: dout  = 8'b11110000; // 1042 : 240 - 0xf0
      11'h413: dout  = 8'b11110000; // 1043 : 240 - 0xf0
      11'h414: dout  = 8'b11101100; // 1044 : 236 - 0xec
      11'h415: dout  = 8'b11100000; // 1045 : 224 - 0xe0
      11'h416: dout  = 8'b11111100; // 1046 : 252 - 0xfc
      11'h417: dout  = 8'b00000000; // 1047 :   0 - 0x0
      11'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0 -- Sprite 0x83
      11'h419: dout  = 8'b00000000; // 1049 :   0 - 0x0
      11'h41A: dout  = 8'b00000000; // 1050 :   0 - 0x0
      11'h41B: dout  = 8'b00000000; // 1051 :   0 - 0x0
      11'h41C: dout  = 8'b00000000; // 1052 :   0 - 0x0
      11'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      11'h41E: dout  = 8'b11100000; // 1054 : 224 - 0xe0
      11'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      11'h420: dout  = 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x84
      11'h421: dout  = 8'b00000011; // 1057 :   3 - 0x3
      11'h422: dout  = 8'b00001111; // 1058 :  15 - 0xf
      11'h423: dout  = 8'b00011111; // 1059 :  31 - 0x1f
      11'h424: dout  = 8'b00011111; // 1060 :  31 - 0x1f
      11'h425: dout  = 8'b00111111; // 1061 :  63 - 0x3f
      11'h426: dout  = 8'b00111111; // 1062 :  63 - 0x3f
      11'h427: dout  = 8'b00000000; // 1063 :   0 - 0x0
      11'h428: dout  = 8'b00000000; // 1064 :   0 - 0x0 -- Sprite 0x85
      11'h429: dout  = 8'b00000000; // 1065 :   0 - 0x0
      11'h42A: dout  = 8'b00000000; // 1066 :   0 - 0x0
      11'h42B: dout  = 8'b00000000; // 1067 :   0 - 0x0
      11'h42C: dout  = 8'b00000000; // 1068 :   0 - 0x0
      11'h42D: dout  = 8'b00001000; // 1069 :   8 - 0x8
      11'h42E: dout  = 8'b00001110; // 1070 :  14 - 0xe
      11'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      11'h430: dout  = 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x86
      11'h431: dout  = 8'b11000000; // 1073 : 192 - 0xc0
      11'h432: dout  = 8'b11110000; // 1074 : 240 - 0xf0
      11'h433: dout  = 8'b11110000; // 1075 : 240 - 0xf0
      11'h434: dout  = 8'b11101100; // 1076 : 236 - 0xec
      11'h435: dout  = 8'b11100000; // 1077 : 224 - 0xe0
      11'h436: dout  = 8'b11111100; // 1078 : 252 - 0xfc
      11'h437: dout  = 8'b00000000; // 1079 :   0 - 0x0
      11'h438: dout  = 8'b00000000; // 1080 :   0 - 0x0 -- Sprite 0x87
      11'h439: dout  = 8'b00000000; // 1081 :   0 - 0x0
      11'h43A: dout  = 8'b00000000; // 1082 :   0 - 0x0
      11'h43B: dout  = 8'b00000000; // 1083 :   0 - 0x0
      11'h43C: dout  = 8'b00000000; // 1084 :   0 - 0x0
      11'h43D: dout  = 8'b00000110; // 1085 :   6 - 0x6
      11'h43E: dout  = 8'b00001100; // 1086 :  12 - 0xc
      11'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      11'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x88
      11'h441: dout  = 8'b00000011; // 1089 :   3 - 0x3
      11'h442: dout  = 8'b00000011; // 1090 :   3 - 0x3
      11'h443: dout  = 8'b00000100; // 1091 :   4 - 0x4
      11'h444: dout  = 8'b00001111; // 1092 :  15 - 0xf
      11'h445: dout  = 8'b00011111; // 1093 :  31 - 0x1f
      11'h446: dout  = 8'b01101111; // 1094 : 111 - 0x6f
      11'h447: dout  = 8'b01101111; // 1095 : 111 - 0x6f
      11'h448: dout  = 8'b01101111; // 1096 : 111 - 0x6f -- Sprite 0x89
      11'h449: dout  = 8'b01101111; // 1097 : 111 - 0x6f
      11'h44A: dout  = 8'b00011111; // 1098 :  31 - 0x1f
      11'h44B: dout  = 8'b00001111; // 1099 :  15 - 0xf
      11'h44C: dout  = 8'b00000100; // 1100 :   4 - 0x4
      11'h44D: dout  = 8'b00000011; // 1101 :   3 - 0x3
      11'h44E: dout  = 8'b00000011; // 1102 :   3 - 0x3
      11'h44F: dout  = 8'b00000000; // 1103 :   0 - 0x0
      11'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x8a
      11'h451: dout  = 8'b00000000; // 1105 :   0 - 0x0
      11'h452: dout  = 8'b00011000; // 1106 :  24 - 0x18
      11'h453: dout  = 8'b00110111; // 1107 :  55 - 0x37
      11'h454: dout  = 8'b00101111; // 1108 :  47 - 0x2f
      11'h455: dout  = 8'b00011111; // 1109 :  31 - 0x1f
      11'h456: dout  = 8'b00011111; // 1110 :  31 - 0x1f
      11'h457: dout  = 8'b00011111; // 1111 :  31 - 0x1f
      11'h458: dout  = 8'b00011111; // 1112 :  31 - 0x1f -- Sprite 0x8b
      11'h459: dout  = 8'b00011111; // 1113 :  31 - 0x1f
      11'h45A: dout  = 8'b00011111; // 1114 :  31 - 0x1f
      11'h45B: dout  = 8'b00101111; // 1115 :  47 - 0x2f
      11'h45C: dout  = 8'b00110111; // 1116 :  55 - 0x37
      11'h45D: dout  = 8'b00011000; // 1117 :  24 - 0x18
      11'h45E: dout  = 8'b00000000; // 1118 :   0 - 0x0
      11'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      11'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x8c
      11'h461: dout  = 8'b00000011; // 1121 :   3 - 0x3
      11'h462: dout  = 8'b00000001; // 1122 :   1 - 0x1
      11'h463: dout  = 8'b00011001; // 1123 :  25 - 0x19
      11'h464: dout  = 8'b00111001; // 1124 :  57 - 0x39
      11'h465: dout  = 8'b00011011; // 1125 :  27 - 0x1b
      11'h466: dout  = 8'b00001111; // 1126 :  15 - 0xf
      11'h467: dout  = 8'b00001111; // 1127 :  15 - 0xf
      11'h468: dout  = 8'b01111111; // 1128 : 127 - 0x7f -- Sprite 0x8d
      11'h469: dout  = 8'b01111111; // 1129 : 127 - 0x7f
      11'h46A: dout  = 8'b00111111; // 1130 :  63 - 0x3f
      11'h46B: dout  = 8'b00010111; // 1131 :  23 - 0x17
      11'h46C: dout  = 8'b00000110; // 1132 :   6 - 0x6
      11'h46D: dout  = 8'b00000100; // 1133 :   4 - 0x4
      11'h46E: dout  = 8'b00000111; // 1134 :   7 - 0x7
      11'h46F: dout  = 8'b00000000; // 1135 :   0 - 0x0
      11'h470: dout  = 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x8e
      11'h471: dout  = 8'b11000000; // 1137 : 192 - 0xc0
      11'h472: dout  = 8'b11110000; // 1138 : 240 - 0xf0
      11'h473: dout  = 8'b10111000; // 1139 : 184 - 0xb8
      11'h474: dout  = 8'b10011100; // 1140 : 156 - 0x9c
      11'h475: dout  = 8'b11111100; // 1141 : 252 - 0xfc
      11'h476: dout  = 8'b11111110; // 1142 : 254 - 0xfe
      11'h477: dout  = 8'b11000000; // 1143 : 192 - 0xc0
      11'h478: dout  = 8'b11111110; // 1144 : 254 - 0xfe -- Sprite 0x8f
      11'h479: dout  = 8'b11111110; // 1145 : 254 - 0xfe
      11'h47A: dout  = 8'b11111000; // 1146 : 248 - 0xf8
      11'h47B: dout  = 8'b11110000; // 1147 : 240 - 0xf0
      11'h47C: dout  = 8'b11000000; // 1148 : 192 - 0xc0
      11'h47D: dout  = 8'b00000000; // 1149 :   0 - 0x0
      11'h47E: dout  = 8'b00000000; // 1150 :   0 - 0x0
      11'h47F: dout  = 8'b10000000; // 1151 : 128 - 0x80
      11'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      11'h481: dout  = 8'b00000001; // 1153 :   1 - 0x1
      11'h482: dout  = 8'b00001001; // 1154 :   9 - 0x9
      11'h483: dout  = 8'b00011001; // 1155 :  25 - 0x19
      11'h484: dout  = 8'b00011100; // 1156 :  28 - 0x1c
      11'h485: dout  = 8'b00001101; // 1157 :  13 - 0xd
      11'h486: dout  = 8'b00001111; // 1158 :  15 - 0xf
      11'h487: dout  = 8'b00101111; // 1159 :  47 - 0x2f
      11'h488: dout  = 8'b01111111; // 1160 : 127 - 0x7f -- Sprite 0x91
      11'h489: dout  = 8'b01111111; // 1161 : 127 - 0x7f
      11'h48A: dout  = 8'b00111111; // 1162 :  63 - 0x3f
      11'h48B: dout  = 8'b00011011; // 1163 :  27 - 0x1b
      11'h48C: dout  = 8'b00000011; // 1164 :   3 - 0x3
      11'h48D: dout  = 8'b00000011; // 1165 :   3 - 0x3
      11'h48E: dout  = 8'b00000001; // 1166 :   1 - 0x1
      11'h48F: dout  = 8'b00000000; // 1167 :   0 - 0x0
      11'h490: dout  = 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x92
      11'h491: dout  = 8'b11000000; // 1169 : 192 - 0xc0
      11'h492: dout  = 8'b11110000; // 1170 : 240 - 0xf0
      11'h493: dout  = 8'b11011000; // 1171 : 216 - 0xd8
      11'h494: dout  = 8'b11001100; // 1172 : 204 - 0xcc
      11'h495: dout  = 8'b11111100; // 1173 : 252 - 0xfc
      11'h496: dout  = 8'b11111110; // 1174 : 254 - 0xfe
      11'h497: dout  = 8'b11100000; // 1175 : 224 - 0xe0
      11'h498: dout  = 8'b11111110; // 1176 : 254 - 0xfe -- Sprite 0x93
      11'h499: dout  = 8'b11111110; // 1177 : 254 - 0xfe
      11'h49A: dout  = 8'b11111000; // 1178 : 248 - 0xf8
      11'h49B: dout  = 8'b01110000; // 1179 : 112 - 0x70
      11'h49C: dout  = 8'b01000000; // 1180 :  64 - 0x40
      11'h49D: dout  = 8'b00000000; // 1181 :   0 - 0x0
      11'h49E: dout  = 8'b11000000; // 1182 : 192 - 0xc0
      11'h49F: dout  = 8'b00100000; // 1183 :  32 - 0x20
      11'h4A0: dout  = 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x94
      11'h4A1: dout  = 8'b00000000; // 1185 :   0 - 0x0
      11'h4A2: dout  = 8'b00001100; // 1186 :  12 - 0xc
      11'h4A3: dout  = 8'b00001110; // 1187 :  14 - 0xe
      11'h4A4: dout  = 8'b00000110; // 1188 :   6 - 0x6
      11'h4A5: dout  = 8'b00100110; // 1189 :  38 - 0x26
      11'h4A6: dout  = 8'b00110111; // 1190 :  55 - 0x37
      11'h4A7: dout  = 8'b00110011; // 1191 :  51 - 0x33
      11'h4A8: dout  = 8'b01111111; // 1192 : 127 - 0x7f -- Sprite 0x95
      11'h4A9: dout  = 8'b01111111; // 1193 : 127 - 0x7f
      11'h4AA: dout  = 8'b00111111; // 1194 :  63 - 0x3f
      11'h4AB: dout  = 8'b00011111; // 1195 :  31 - 0x1f
      11'h4AC: dout  = 8'b00001110; // 1196 :  14 - 0xe
      11'h4AD: dout  = 8'b00000000; // 1197 :   0 - 0x0
      11'h4AE: dout  = 8'b00000000; // 1198 :   0 - 0x0
      11'h4AF: dout  = 8'b00000000; // 1199 :   0 - 0x0
      11'h4B0: dout  = 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x96
      11'h4B1: dout  = 8'b11000000; // 1201 : 192 - 0xc0
      11'h4B2: dout  = 8'b11110000; // 1202 : 240 - 0xf0
      11'h4B3: dout  = 8'b01101000; // 1203 : 104 - 0x68
      11'h4B4: dout  = 8'b01100100; // 1204 : 100 - 0x64
      11'h4B5: dout  = 8'b11111100; // 1205 : 252 - 0xfc
      11'h4B6: dout  = 8'b11111110; // 1206 : 254 - 0xfe
      11'h4B7: dout  = 8'b11110000; // 1207 : 240 - 0xf0
      11'h4B8: dout  = 8'b11111111; // 1208 : 255 - 0xff -- Sprite 0x97
      11'h4B9: dout  = 8'b11111110; // 1209 : 254 - 0xfe
      11'h4BA: dout  = 8'b11111100; // 1210 : 252 - 0xfc
      11'h4BB: dout  = 8'b10110000; // 1211 : 176 - 0xb0
      11'h4BC: dout  = 8'b11000000; // 1212 : 192 - 0xc0
      11'h4BD: dout  = 8'b11000000; // 1213 : 192 - 0xc0
      11'h4BE: dout  = 8'b01110000; // 1214 : 112 - 0x70
      11'h4BF: dout  = 8'b00001000; // 1215 :   8 - 0x8
      11'h4C0: dout  = 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x98
      11'h4C1: dout  = 8'b00000001; // 1217 :   1 - 0x1
      11'h4C2: dout  = 8'b00000000; // 1218 :   0 - 0x0
      11'h4C3: dout  = 8'b00000000; // 1219 :   0 - 0x0
      11'h4C4: dout  = 8'b00000000; // 1220 :   0 - 0x0
      11'h4C5: dout  = 8'b00000000; // 1221 :   0 - 0x0
      11'h4C6: dout  = 8'b00000001; // 1222 :   1 - 0x1
      11'h4C7: dout  = 8'b00000011; // 1223 :   3 - 0x3
      11'h4C8: dout  = 8'b00000111; // 1224 :   7 - 0x7 -- Sprite 0x99
      11'h4C9: dout  = 8'b00010111; // 1225 :  23 - 0x17
      11'h4CA: dout  = 8'b00101111; // 1226 :  47 - 0x2f
      11'h4CB: dout  = 8'b00011110; // 1227 :  30 - 0x1e
      11'h4CC: dout  = 8'b00010001; // 1228 :  17 - 0x11
      11'h4CD: dout  = 8'b00000000; // 1229 :   0 - 0x0
      11'h4CE: dout  = 8'b00000001; // 1230 :   1 - 0x1
      11'h4CF: dout  = 8'b00000000; // 1231 :   0 - 0x0
      11'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      11'h4D1: dout  = 8'b00010000; // 1233 :  16 - 0x10
      11'h4D2: dout  = 8'b01111000; // 1234 : 120 - 0x78
      11'h4D3: dout  = 8'b01110100; // 1235 : 116 - 0x74
      11'h4D4: dout  = 8'b11111110; // 1236 : 254 - 0xfe
      11'h4D5: dout  = 8'b11111000; // 1237 : 248 - 0xf8
      11'h4D6: dout  = 8'b11111100; // 1238 : 252 - 0xfc
      11'h4D7: dout  = 8'b11111000; // 1239 : 248 - 0xf8
      11'h4D8: dout  = 8'b11111000; // 1240 : 248 - 0xf8 -- Sprite 0x9b
      11'h4D9: dout  = 8'b11010000; // 1241 : 208 - 0xd0
      11'h4DA: dout  = 8'b00110000; // 1242 :  48 - 0x30
      11'h4DB: dout  = 8'b01100000; // 1243 :  96 - 0x60
      11'h4DC: dout  = 8'b10000000; // 1244 : 128 - 0x80
      11'h4DD: dout  = 8'b00000000; // 1245 :   0 - 0x0
      11'h4DE: dout  = 8'b00000000; // 1246 :   0 - 0x0
      11'h4DF: dout  = 8'b00000000; // 1247 :   0 - 0x0
      11'h4E0: dout  = 8'b00000000; // 1248 :   0 - 0x0 -- Sprite 0x9c
      11'h4E1: dout  = 8'b00000001; // 1249 :   1 - 0x1
      11'h4E2: dout  = 8'b00000000; // 1250 :   0 - 0x0
      11'h4E3: dout  = 8'b00000000; // 1251 :   0 - 0x0
      11'h4E4: dout  = 8'b00000000; // 1252 :   0 - 0x0
      11'h4E5: dout  = 8'b00000000; // 1253 :   0 - 0x0
      11'h4E6: dout  = 8'b00000001; // 1254 :   1 - 0x1
      11'h4E7: dout  = 8'b00000011; // 1255 :   3 - 0x3
      11'h4E8: dout  = 8'b00000111; // 1256 :   7 - 0x7 -- Sprite 0x9d
      11'h4E9: dout  = 8'b00010111; // 1257 :  23 - 0x17
      11'h4EA: dout  = 8'b00101111; // 1258 :  47 - 0x2f
      11'h4EB: dout  = 8'b00011110; // 1259 :  30 - 0x1e
      11'h4EC: dout  = 8'b00010000; // 1260 :  16 - 0x10
      11'h4ED: dout  = 8'b00000100; // 1261 :   4 - 0x4
      11'h4EE: dout  = 8'b00000000; // 1262 :   0 - 0x0
      11'h4EF: dout  = 8'b00000000; // 1263 :   0 - 0x0
      11'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Sprite 0x9e
      11'h4F1: dout  = 8'b00010000; // 1265 :  16 - 0x10
      11'h4F2: dout  = 8'b01111000; // 1266 : 120 - 0x78
      11'h4F3: dout  = 8'b01110100; // 1267 : 116 - 0x74
      11'h4F4: dout  = 8'b11111110; // 1268 : 254 - 0xfe
      11'h4F5: dout  = 8'b11111000; // 1269 : 248 - 0xf8
      11'h4F6: dout  = 8'b11111100; // 1270 : 252 - 0xfc
      11'h4F7: dout  = 8'b11111000; // 1271 : 248 - 0xf8
      11'h4F8: dout  = 8'b11111000; // 1272 : 248 - 0xf8 -- Sprite 0x9f
      11'h4F9: dout  = 8'b11010000; // 1273 : 208 - 0xd0
      11'h4FA: dout  = 8'b00110000; // 1274 :  48 - 0x30
      11'h4FB: dout  = 8'b11000000; // 1275 : 192 - 0xc0
      11'h4FC: dout  = 8'b00000000; // 1276 :   0 - 0x0
      11'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      11'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      11'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0xa0
      11'h501: dout  = 8'b00000011; // 1281 :   3 - 0x3
      11'h502: dout  = 8'b00001111; // 1282 :  15 - 0xf
      11'h503: dout  = 8'b00011111; // 1283 :  31 - 0x1f
      11'h504: dout  = 8'b00111111; // 1284 :  63 - 0x3f
      11'h505: dout  = 8'b00111111; // 1285 :  63 - 0x3f
      11'h506: dout  = 8'b01111111; // 1286 : 127 - 0x7f
      11'h507: dout  = 8'b01111111; // 1287 : 127 - 0x7f
      11'h508: dout  = 8'b01111111; // 1288 : 127 - 0x7f -- Sprite 0xa1
      11'h509: dout  = 8'b01111111; // 1289 : 127 - 0x7f
      11'h50A: dout  = 8'b00111111; // 1290 :  63 - 0x3f
      11'h50B: dout  = 8'b00111111; // 1291 :  63 - 0x3f
      11'h50C: dout  = 8'b00011111; // 1292 :  31 - 0x1f
      11'h50D: dout  = 8'b00000101; // 1293 :   5 - 0x5
      11'h50E: dout  = 8'b00000010; // 1294 :   2 - 0x2
      11'h50F: dout  = 8'b00000000; // 1295 :   0 - 0x0
      11'h510: dout  = 8'b00000000; // 1296 :   0 - 0x0 -- Sprite 0xa2
      11'h511: dout  = 8'b11000000; // 1297 : 192 - 0xc0
      11'h512: dout  = 8'b11110000; // 1298 : 240 - 0xf0
      11'h513: dout  = 8'b11111000; // 1299 : 248 - 0xf8
      11'h514: dout  = 8'b11111000; // 1300 : 248 - 0xf8
      11'h515: dout  = 8'b11111100; // 1301 : 252 - 0xfc
      11'h516: dout  = 8'b11111010; // 1302 : 250 - 0xfa
      11'h517: dout  = 8'b11111100; // 1303 : 252 - 0xfc
      11'h518: dout  = 8'b11111010; // 1304 : 250 - 0xfa -- Sprite 0xa3
      11'h519: dout  = 8'b11110100; // 1305 : 244 - 0xf4
      11'h51A: dout  = 8'b11101000; // 1306 : 232 - 0xe8
      11'h51B: dout  = 8'b11010100; // 1307 : 212 - 0xd4
      11'h51C: dout  = 8'b10101000; // 1308 : 168 - 0xa8
      11'h51D: dout  = 8'b01010000; // 1309 :  80 - 0x50
      11'h51E: dout  = 8'b10000000; // 1310 : 128 - 0x80
      11'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      11'h520: dout  = 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0xa4
      11'h521: dout  = 8'b00000000; // 1313 :   0 - 0x0
      11'h522: dout  = 8'b00000000; // 1314 :   0 - 0x0
      11'h523: dout  = 8'b00001110; // 1315 :  14 - 0xe
      11'h524: dout  = 8'b00000000; // 1316 :   0 - 0x0
      11'h525: dout  = 8'b00001010; // 1317 :  10 - 0xa
      11'h526: dout  = 8'b01001010; // 1318 :  74 - 0x4a
      11'h527: dout  = 8'b01100000; // 1319 :  96 - 0x60
      11'h528: dout  = 8'b01111111; // 1320 : 127 - 0x7f -- Sprite 0xa5
      11'h529: dout  = 8'b01111000; // 1321 : 120 - 0x78
      11'h52A: dout  = 8'b00110111; // 1322 :  55 - 0x37
      11'h52B: dout  = 8'b00111011; // 1323 :  59 - 0x3b
      11'h52C: dout  = 8'b00111100; // 1324 :  60 - 0x3c
      11'h52D: dout  = 8'b00011111; // 1325 :  31 - 0x1f
      11'h52E: dout  = 8'b00000111; // 1326 :   7 - 0x7
      11'h52F: dout  = 8'b00000000; // 1327 :   0 - 0x0
      11'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0xa6
      11'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      11'h532: dout  = 8'b00000000; // 1330 :   0 - 0x0
      11'h533: dout  = 8'b01110000; // 1331 : 112 - 0x70
      11'h534: dout  = 8'b00000000; // 1332 :   0 - 0x0
      11'h535: dout  = 8'b01010000; // 1333 :  80 - 0x50
      11'h536: dout  = 8'b01010010; // 1334 :  82 - 0x52
      11'h537: dout  = 8'b00000110; // 1335 :   6 - 0x6
      11'h538: dout  = 8'b11111100; // 1336 : 252 - 0xfc -- Sprite 0xa7
      11'h539: dout  = 8'b00011010; // 1337 :  26 - 0x1a
      11'h53A: dout  = 8'b11101100; // 1338 : 236 - 0xec
      11'h53B: dout  = 8'b11011000; // 1339 : 216 - 0xd8
      11'h53C: dout  = 8'b00110100; // 1340 :  52 - 0x34
      11'h53D: dout  = 8'b11101000; // 1341 : 232 - 0xe8
      11'h53E: dout  = 8'b11000000; // 1342 : 192 - 0xc0
      11'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      11'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0xa8
      11'h541: dout  = 8'b00000000; // 1345 :   0 - 0x0
      11'h542: dout  = 8'b00000000; // 1346 :   0 - 0x0
      11'h543: dout  = 8'b00001110; // 1347 :  14 - 0xe
      11'h544: dout  = 8'b00000000; // 1348 :   0 - 0x0
      11'h545: dout  = 8'b00001110; // 1349 :  14 - 0xe
      11'h546: dout  = 8'b01001010; // 1350 :  74 - 0x4a
      11'h547: dout  = 8'b01100000; // 1351 :  96 - 0x60
      11'h548: dout  = 8'b01111111; // 1352 : 127 - 0x7f -- Sprite 0xa9
      11'h549: dout  = 8'b01111100; // 1353 : 124 - 0x7c
      11'h54A: dout  = 8'b01111011; // 1354 : 123 - 0x7b
      11'h54B: dout  = 8'b01110111; // 1355 : 119 - 0x77
      11'h54C: dout  = 8'b01111000; // 1356 : 120 - 0x78
      11'h54D: dout  = 8'b01111111; // 1357 : 127 - 0x7f
      11'h54E: dout  = 8'b01111111; // 1358 : 127 - 0x7f
      11'h54F: dout  = 8'b00000000; // 1359 :   0 - 0x0
      11'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      11'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      11'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      11'h553: dout  = 8'b01110000; // 1363 : 112 - 0x70
      11'h554: dout  = 8'b00000000; // 1364 :   0 - 0x0
      11'h555: dout  = 8'b01110000; // 1365 : 112 - 0x70
      11'h556: dout  = 8'b01010010; // 1366 :  82 - 0x52
      11'h557: dout  = 8'b00000110; // 1367 :   6 - 0x6
      11'h558: dout  = 8'b11111100; // 1368 : 252 - 0xfc -- Sprite 0xab
      11'h559: dout  = 8'b00111010; // 1369 :  58 - 0x3a
      11'h55A: dout  = 8'b11011100; // 1370 : 220 - 0xdc
      11'h55B: dout  = 8'b11101010; // 1371 : 234 - 0xea
      11'h55C: dout  = 8'b00011100; // 1372 :  28 - 0x1c
      11'h55D: dout  = 8'b11111010; // 1373 : 250 - 0xfa
      11'h55E: dout  = 8'b11110100; // 1374 : 244 - 0xf4
      11'h55F: dout  = 8'b00000000; // 1375 :   0 - 0x0
      11'h560: dout  = 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      11'h561: dout  = 8'b00000011; // 1377 :   3 - 0x3
      11'h562: dout  = 8'b00001111; // 1378 :  15 - 0xf
      11'h563: dout  = 8'b00001111; // 1379 :  15 - 0xf
      11'h564: dout  = 8'b00011111; // 1380 :  31 - 0x1f
      11'h565: dout  = 8'b01011111; // 1381 :  95 - 0x5f
      11'h566: dout  = 8'b01010000; // 1382 :  80 - 0x50
      11'h567: dout  = 8'b00010000; // 1383 :  16 - 0x10
      11'h568: dout  = 8'b00000000; // 1384 :   0 - 0x0 -- Sprite 0xad
      11'h569: dout  = 8'b11111010; // 1385 : 250 - 0xfa
      11'h56A: dout  = 8'b11111010; // 1386 : 250 - 0xfa
      11'h56B: dout  = 8'b11111010; // 1387 : 250 - 0xfa
      11'h56C: dout  = 8'b10111010; // 1388 : 186 - 0xba
      11'h56D: dout  = 8'b10011010; // 1389 : 154 - 0x9a
      11'h56E: dout  = 8'b00001010; // 1390 :  10 - 0xa
      11'h56F: dout  = 8'b00000010; // 1391 :   2 - 0x2
      11'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      11'h571: dout  = 8'b00000011; // 1393 :   3 - 0x3
      11'h572: dout  = 8'b00001111; // 1394 :  15 - 0xf
      11'h573: dout  = 8'b00001111; // 1395 :  15 - 0xf
      11'h574: dout  = 8'b00011111; // 1396 :  31 - 0x1f
      11'h575: dout  = 8'b01011111; // 1397 :  95 - 0x5f
      11'h576: dout  = 8'b01010000; // 1398 :  80 - 0x50
      11'h577: dout  = 8'b00010111; // 1399 :  23 - 0x17
      11'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Sprite 0xaf
      11'h579: dout  = 8'b11111010; // 1401 : 250 - 0xfa
      11'h57A: dout  = 8'b11111010; // 1402 : 250 - 0xfa
      11'h57B: dout  = 8'b11111010; // 1403 : 250 - 0xfa
      11'h57C: dout  = 8'b00111010; // 1404 :  58 - 0x3a
      11'h57D: dout  = 8'b01011010; // 1405 :  90 - 0x5a
      11'h57E: dout  = 8'b01101010; // 1406 : 106 - 0x6a
      11'h57F: dout  = 8'b11110010; // 1407 : 242 - 0xf2
      11'h580: dout  = 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      11'h581: dout  = 8'b00000000; // 1409 :   0 - 0x0
      11'h582: dout  = 8'b00000011; // 1410 :   3 - 0x3
      11'h583: dout  = 8'b00001111; // 1411 :  15 - 0xf
      11'h584: dout  = 8'b00111011; // 1412 :  59 - 0x3b
      11'h585: dout  = 8'b00111111; // 1413 :  63 - 0x3f
      11'h586: dout  = 8'b01101111; // 1414 : 111 - 0x6f
      11'h587: dout  = 8'b01111101; // 1415 : 125 - 0x7d
      11'h588: dout  = 8'b00001111; // 1416 :  15 - 0xf -- Sprite 0xb1
      11'h589: dout  = 8'b01110000; // 1417 : 112 - 0x70
      11'h58A: dout  = 8'b01111111; // 1418 : 127 - 0x7f
      11'h58B: dout  = 8'b00001111; // 1419 :  15 - 0xf
      11'h58C: dout  = 8'b01110000; // 1420 : 112 - 0x70
      11'h58D: dout  = 8'b01111111; // 1421 : 127 - 0x7f
      11'h58E: dout  = 8'b00001111; // 1422 :  15 - 0xf
      11'h58F: dout  = 8'b00000000; // 1423 :   0 - 0x0
      11'h590: dout  = 8'b00000000; // 1424 :   0 - 0x0 -- Sprite 0xb2
      11'h591: dout  = 8'b00000000; // 1425 :   0 - 0x0
      11'h592: dout  = 8'b11000000; // 1426 : 192 - 0xc0
      11'h593: dout  = 8'b11110000; // 1427 : 240 - 0xf0
      11'h594: dout  = 8'b10111100; // 1428 : 188 - 0xbc
      11'h595: dout  = 8'b11110100; // 1429 : 244 - 0xf4
      11'h596: dout  = 8'b11111110; // 1430 : 254 - 0xfe
      11'h597: dout  = 8'b11011110; // 1431 : 222 - 0xde
      11'h598: dout  = 8'b11110000; // 1432 : 240 - 0xf0 -- Sprite 0xb3
      11'h599: dout  = 8'b00001110; // 1433 :  14 - 0xe
      11'h59A: dout  = 8'b11111110; // 1434 : 254 - 0xfe
      11'h59B: dout  = 8'b11110000; // 1435 : 240 - 0xf0
      11'h59C: dout  = 8'b00001110; // 1436 :  14 - 0xe
      11'h59D: dout  = 8'b11111110; // 1437 : 254 - 0xfe
      11'h59E: dout  = 8'b11110000; // 1438 : 240 - 0xf0
      11'h59F: dout  = 8'b00000000; // 1439 :   0 - 0x0
      11'h5A0: dout  = 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0xb4
      11'h5A1: dout  = 8'b00000000; // 1441 :   0 - 0x0
      11'h5A2: dout  = 8'b00000011; // 1442 :   3 - 0x3
      11'h5A3: dout  = 8'b00001111; // 1443 :  15 - 0xf
      11'h5A4: dout  = 8'b00111011; // 1444 :  59 - 0x3b
      11'h5A5: dout  = 8'b00111111; // 1445 :  63 - 0x3f
      11'h5A6: dout  = 8'b01101111; // 1446 : 111 - 0x6f
      11'h5A7: dout  = 8'b01111101; // 1447 : 125 - 0x7d
      11'h5A8: dout  = 8'b00001111; // 1448 :  15 - 0xf -- Sprite 0xb5
      11'h5A9: dout  = 8'b01110000; // 1449 : 112 - 0x70
      11'h5AA: dout  = 8'b01111111; // 1450 : 127 - 0x7f
      11'h5AB: dout  = 8'b00001111; // 1451 :  15 - 0xf
      11'h5AC: dout  = 8'b01110000; // 1452 : 112 - 0x70
      11'h5AD: dout  = 8'b01111111; // 1453 : 127 - 0x7f
      11'h5AE: dout  = 8'b00001111; // 1454 :  15 - 0xf
      11'h5AF: dout  = 8'b00000000; // 1455 :   0 - 0x0
      11'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0xb6
      11'h5B1: dout  = 8'b00000000; // 1457 :   0 - 0x0
      11'h5B2: dout  = 8'b11000000; // 1458 : 192 - 0xc0
      11'h5B3: dout  = 8'b11110000; // 1459 : 240 - 0xf0
      11'h5B4: dout  = 8'b10111100; // 1460 : 188 - 0xbc
      11'h5B5: dout  = 8'b11110100; // 1461 : 244 - 0xf4
      11'h5B6: dout  = 8'b11111110; // 1462 : 254 - 0xfe
      11'h5B7: dout  = 8'b11011110; // 1463 : 222 - 0xde
      11'h5B8: dout  = 8'b11110000; // 1464 : 240 - 0xf0 -- Sprite 0xb7
      11'h5B9: dout  = 8'b00001110; // 1465 :  14 - 0xe
      11'h5BA: dout  = 8'b11111110; // 1466 : 254 - 0xfe
      11'h5BB: dout  = 8'b11110000; // 1467 : 240 - 0xf0
      11'h5BC: dout  = 8'b00001110; // 1468 :  14 - 0xe
      11'h5BD: dout  = 8'b11111110; // 1469 : 254 - 0xfe
      11'h5BE: dout  = 8'b11110000; // 1470 : 240 - 0xf0
      11'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      11'h5C0: dout  = 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0xb8
      11'h5C1: dout  = 8'b00000000; // 1473 :   0 - 0x0
      11'h5C2: dout  = 8'b00000011; // 1474 :   3 - 0x3
      11'h5C3: dout  = 8'b00001111; // 1475 :  15 - 0xf
      11'h5C4: dout  = 8'b00111011; // 1476 :  59 - 0x3b
      11'h5C5: dout  = 8'b00111111; // 1477 :  63 - 0x3f
      11'h5C6: dout  = 8'b01101111; // 1478 : 111 - 0x6f
      11'h5C7: dout  = 8'b01111101; // 1479 : 125 - 0x7d
      11'h5C8: dout  = 8'b00001111; // 1480 :  15 - 0xf -- Sprite 0xb9
      11'h5C9: dout  = 8'b00100000; // 1481 :  32 - 0x20
      11'h5CA: dout  = 8'b01010101; // 1482 :  85 - 0x55
      11'h5CB: dout  = 8'b00001010; // 1483 :  10 - 0xa
      11'h5CC: dout  = 8'b01110000; // 1484 : 112 - 0x70
      11'h5CD: dout  = 8'b01111111; // 1485 : 127 - 0x7f
      11'h5CE: dout  = 8'b00001111; // 1486 :  15 - 0xf
      11'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      11'h5D0: dout  = 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0xba
      11'h5D1: dout  = 8'b00000000; // 1489 :   0 - 0x0
      11'h5D2: dout  = 8'b11000000; // 1490 : 192 - 0xc0
      11'h5D3: dout  = 8'b11110000; // 1491 : 240 - 0xf0
      11'h5D4: dout  = 8'b10111100; // 1492 : 188 - 0xbc
      11'h5D5: dout  = 8'b11110100; // 1493 : 244 - 0xf4
      11'h5D6: dout  = 8'b11111110; // 1494 : 254 - 0xfe
      11'h5D7: dout  = 8'b11011110; // 1495 : 222 - 0xde
      11'h5D8: dout  = 8'b11110000; // 1496 : 240 - 0xf0 -- Sprite 0xbb
      11'h5D9: dout  = 8'b00001010; // 1497 :  10 - 0xa
      11'h5DA: dout  = 8'b01010100; // 1498 :  84 - 0x54
      11'h5DB: dout  = 8'b10100000; // 1499 : 160 - 0xa0
      11'h5DC: dout  = 8'b00001110; // 1500 :  14 - 0xe
      11'h5DD: dout  = 8'b11111110; // 1501 : 254 - 0xfe
      11'h5DE: dout  = 8'b11110000; // 1502 : 240 - 0xf0
      11'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      11'h5E0: dout  = 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0xbc
      11'h5E1: dout  = 8'b01110011; // 1505 : 115 - 0x73
      11'h5E2: dout  = 8'b01111011; // 1506 : 123 - 0x7b
      11'h5E3: dout  = 8'b01111111; // 1507 : 127 - 0x7f
      11'h5E4: dout  = 8'b00111111; // 1508 :  63 - 0x3f
      11'h5E5: dout  = 8'b00011100; // 1509 :  28 - 0x1c
      11'h5E6: dout  = 8'b01111011; // 1510 : 123 - 0x7b
      11'h5E7: dout  = 8'b01111011; // 1511 : 123 - 0x7b
      11'h5E8: dout  = 8'b01111011; // 1512 : 123 - 0x7b -- Sprite 0xbd
      11'h5E9: dout  = 8'b01111011; // 1513 : 123 - 0x7b
      11'h5EA: dout  = 8'b00011100; // 1514 :  28 - 0x1c
      11'h5EB: dout  = 8'b00111111; // 1515 :  63 - 0x3f
      11'h5EC: dout  = 8'b01111111; // 1516 : 127 - 0x7f
      11'h5ED: dout  = 8'b01111011; // 1517 : 123 - 0x7b
      11'h5EE: dout  = 8'b01110011; // 1518 : 115 - 0x73
      11'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      11'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      11'h5F1: dout  = 8'b11001110; // 1521 : 206 - 0xce
      11'h5F2: dout  = 8'b11011110; // 1522 : 222 - 0xde
      11'h5F3: dout  = 8'b11111110; // 1523 : 254 - 0xfe
      11'h5F4: dout  = 8'b11111100; // 1524 : 252 - 0xfc
      11'h5F5: dout  = 8'b00111000; // 1525 :  56 - 0x38
      11'h5F6: dout  = 8'b11011110; // 1526 : 222 - 0xde
      11'h5F7: dout  = 8'b11011110; // 1527 : 222 - 0xde
      11'h5F8: dout  = 8'b11011110; // 1528 : 222 - 0xde -- Sprite 0xbf
      11'h5F9: dout  = 8'b11011110; // 1529 : 222 - 0xde
      11'h5FA: dout  = 8'b00111000; // 1530 :  56 - 0x38
      11'h5FB: dout  = 8'b11111100; // 1531 : 252 - 0xfc
      11'h5FC: dout  = 8'b11111110; // 1532 : 254 - 0xfe
      11'h5FD: dout  = 8'b11011110; // 1533 : 222 - 0xde
      11'h5FE: dout  = 8'b11001110; // 1534 : 206 - 0xce
      11'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      11'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      11'h601: dout  = 8'b00000000; // 1537 :   0 - 0x0
      11'h602: dout  = 8'b01000000; // 1538 :  64 - 0x40
      11'h603: dout  = 8'b01100000; // 1539 :  96 - 0x60
      11'h604: dout  = 8'b01100001; // 1540 :  97 - 0x61
      11'h605: dout  = 8'b00000010; // 1541 :   2 - 0x2
      11'h606: dout  = 8'b00000010; // 1542 :   2 - 0x2
      11'h607: dout  = 8'b00000111; // 1543 :   7 - 0x7
      11'h608: dout  = 8'b00000111; // 1544 :   7 - 0x7 -- Sprite 0xc1
      11'h609: dout  = 8'b00000100; // 1545 :   4 - 0x4
      11'h60A: dout  = 8'b00000111; // 1546 :   7 - 0x7
      11'h60B: dout  = 8'b00000001; // 1547 :   1 - 0x1
      11'h60C: dout  = 8'b00000000; // 1548 :   0 - 0x0
      11'h60D: dout  = 8'b00010000; // 1549 :  16 - 0x10
      11'h60E: dout  = 8'b00101000; // 1550 :  40 - 0x28
      11'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      11'h611: dout  = 8'b00000000; // 1553 :   0 - 0x0
      11'h612: dout  = 8'b00000010; // 1554 :   2 - 0x2
      11'h613: dout  = 8'b00000110; // 1555 :   6 - 0x6
      11'h614: dout  = 8'b11100110; // 1556 : 230 - 0xe6
      11'h615: dout  = 8'b10100000; // 1557 : 160 - 0xa0
      11'h616: dout  = 8'b10100000; // 1558 : 160 - 0xa0
      11'h617: dout  = 8'b11110000; // 1559 : 240 - 0xf0
      11'h618: dout  = 8'b11110000; // 1560 : 240 - 0xf0 -- Sprite 0xc3
      11'h619: dout  = 8'b00110000; // 1561 :  48 - 0x30
      11'h61A: dout  = 8'b11000000; // 1562 : 192 - 0xc0
      11'h61B: dout  = 8'b10000000; // 1563 : 128 - 0x80
      11'h61C: dout  = 8'b00000000; // 1564 :   0 - 0x0
      11'h61D: dout  = 8'b00001000; // 1565 :   8 - 0x8
      11'h61E: dout  = 8'b00010100; // 1566 :  20 - 0x14
      11'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      11'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      11'h621: dout  = 8'b00000101; // 1569 :   5 - 0x5
      11'h622: dout  = 8'b00000111; // 1570 :   7 - 0x7
      11'h623: dout  = 8'b00000000; // 1571 :   0 - 0x0
      11'h624: dout  = 8'b00000000; // 1572 :   0 - 0x0
      11'h625: dout  = 8'b00000000; // 1573 :   0 - 0x0
      11'h626: dout  = 8'b00000000; // 1574 :   0 - 0x0
      11'h627: dout  = 8'b00000001; // 1575 :   1 - 0x1
      11'h628: dout  = 8'b00000010; // 1576 :   2 - 0x2 -- Sprite 0xc5
      11'h629: dout  = 8'b00000111; // 1577 :   7 - 0x7
      11'h62A: dout  = 8'b00100111; // 1578 :  39 - 0x27
      11'h62B: dout  = 8'b01010011; // 1579 :  83 - 0x53
      11'h62C: dout  = 8'b00000000; // 1580 :   0 - 0x0
      11'h62D: dout  = 8'b00000010; // 1581 :   2 - 0x2
      11'h62E: dout  = 8'b00000101; // 1582 :   5 - 0x5
      11'h62F: dout  = 8'b00000000; // 1583 :   0 - 0x0
      11'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0xc6
      11'h631: dout  = 8'b00000000; // 1585 :   0 - 0x0
      11'h632: dout  = 8'b00000000; // 1586 :   0 - 0x0
      11'h633: dout  = 8'b00000000; // 1587 :   0 - 0x0
      11'h634: dout  = 8'b00000000; // 1588 :   0 - 0x0
      11'h635: dout  = 8'b01100000; // 1589 :  96 - 0x60
      11'h636: dout  = 8'b11011000; // 1590 : 216 - 0xd8
      11'h637: dout  = 8'b10110000; // 1591 : 176 - 0xb0
      11'h638: dout  = 8'b11101000; // 1592 : 232 - 0xe8 -- Sprite 0xc7
      11'h639: dout  = 8'b01111000; // 1593 : 120 - 0x78
      11'h63A: dout  = 8'b10110110; // 1594 : 182 - 0xb6
      11'h63B: dout  = 8'b11100100; // 1595 : 228 - 0xe4
      11'h63C: dout  = 8'b00000110; // 1596 :   6 - 0x6
      11'h63D: dout  = 8'b00000000; // 1597 :   0 - 0x0
      11'h63E: dout  = 8'b00000000; // 1598 :   0 - 0x0
      11'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      11'h640: dout  = 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      11'h641: dout  = 8'b00000000; // 1601 :   0 - 0x0
      11'h642: dout  = 8'b01000000; // 1602 :  64 - 0x40
      11'h643: dout  = 8'b00100000; // 1603 :  32 - 0x20
      11'h644: dout  = 8'b01000000; // 1604 :  64 - 0x40
      11'h645: dout  = 8'b00000111; // 1605 :   7 - 0x7
      11'h646: dout  = 8'b00000101; // 1606 :   5 - 0x5
      11'h647: dout  = 8'b00001101; // 1607 :  13 - 0xd
      11'h648: dout  = 8'b00001101; // 1608 :  13 - 0xd -- Sprite 0xc9
      11'h649: dout  = 8'b00000101; // 1609 :   5 - 0x5
      11'h64A: dout  = 8'b00000011; // 1610 :   3 - 0x3
      11'h64B: dout  = 8'b01000011; // 1611 :  67 - 0x43
      11'h64C: dout  = 8'b00100000; // 1612 :  32 - 0x20
      11'h64D: dout  = 8'b01000000; // 1613 :  64 - 0x40
      11'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      11'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      11'h650: dout  = 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      11'h651: dout  = 8'b00011100; // 1617 :  28 - 0x1c
      11'h652: dout  = 8'b00011000; // 1618 :  24 - 0x18
      11'h653: dout  = 8'b00000000; // 1619 :   0 - 0x0
      11'h654: dout  = 8'b00000000; // 1620 :   0 - 0x0
      11'h655: dout  = 8'b10000000; // 1621 : 128 - 0x80
      11'h656: dout  = 8'b11100000; // 1622 : 224 - 0xe0
      11'h657: dout  = 8'b10010000; // 1623 : 144 - 0x90
      11'h658: dout  = 8'b11110000; // 1624 : 240 - 0xf0 -- Sprite 0xcb
      11'h659: dout  = 8'b10010000; // 1625 : 144 - 0x90
      11'h65A: dout  = 8'b11110000; // 1626 : 240 - 0xf0
      11'h65B: dout  = 8'b10000000; // 1627 : 128 - 0x80
      11'h65C: dout  = 8'b00000000; // 1628 :   0 - 0x0
      11'h65D: dout  = 8'b00011000; // 1629 :  24 - 0x18
      11'h65E: dout  = 8'b00011100; // 1630 :  28 - 0x1c
      11'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      11'h660: dout  = 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0xcc
      11'h661: dout  = 8'b00001000; // 1633 :   8 - 0x8
      11'h662: dout  = 8'b00000100; // 1634 :   4 - 0x4
      11'h663: dout  = 8'b00001000; // 1635 :   8 - 0x8
      11'h664: dout  = 8'b00000000; // 1636 :   0 - 0x0
      11'h665: dout  = 8'b01000110; // 1637 :  70 - 0x46
      11'h666: dout  = 8'b00101111; // 1638 :  47 - 0x2f
      11'h667: dout  = 8'b01001110; // 1639 :  78 - 0x4e
      11'h668: dout  = 8'b00001101; // 1640 :  13 - 0xd -- Sprite 0xcd
      11'h669: dout  = 8'b00001011; // 1641 :  11 - 0xb
      11'h66A: dout  = 8'b00001111; // 1642 :  15 - 0xf
      11'h66B: dout  = 8'b00000110; // 1643 :   6 - 0x6
      11'h66C: dout  = 8'b00000011; // 1644 :   3 - 0x3
      11'h66D: dout  = 8'b00011100; // 1645 :  28 - 0x1c
      11'h66E: dout  = 8'b00010100; // 1646 :  20 - 0x14
      11'h66F: dout  = 8'b00000000; // 1647 :   0 - 0x0
      11'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      11'h671: dout  = 8'b00000000; // 1649 :   0 - 0x0
      11'h672: dout  = 8'b00000000; // 1650 :   0 - 0x0
      11'h673: dout  = 8'b00000000; // 1651 :   0 - 0x0
      11'h674: dout  = 8'b00000000; // 1652 :   0 - 0x0
      11'h675: dout  = 8'b00000110; // 1653 :   6 - 0x6
      11'h676: dout  = 8'b00000100; // 1654 :   4 - 0x4
      11'h677: dout  = 8'b10000110; // 1655 : 134 - 0x86
      11'h678: dout  = 8'b11000000; // 1656 : 192 - 0xc0 -- Sprite 0xcf
      11'h679: dout  = 8'b01100000; // 1657 :  96 - 0x60
      11'h67A: dout  = 8'b10100000; // 1658 : 160 - 0xa0
      11'h67B: dout  = 8'b11000000; // 1659 : 192 - 0xc0
      11'h67C: dout  = 8'b01000000; // 1660 :  64 - 0x40
      11'h67D: dout  = 8'b00000000; // 1661 :   0 - 0x0
      11'h67E: dout  = 8'b00000000; // 1662 :   0 - 0x0
      11'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      11'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      11'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      11'h682: dout  = 8'b00000000; // 1666 :   0 - 0x0
      11'h683: dout  = 8'b00000000; // 1667 :   0 - 0x0
      11'h684: dout  = 8'b00000100; // 1668 :   4 - 0x4
      11'h685: dout  = 8'b00001110; // 1669 :  14 - 0xe
      11'h686: dout  = 8'b00111111; // 1670 :  63 - 0x3f
      11'h687: dout  = 8'b00111001; // 1671 :  57 - 0x39
      11'h688: dout  = 8'b01110000; // 1672 : 112 - 0x70 -- Sprite 0xd1
      11'h689: dout  = 8'b01111000; // 1673 : 120 - 0x78
      11'h68A: dout  = 8'b00111111; // 1674 :  63 - 0x3f
      11'h68B: dout  = 8'b00111111; // 1675 :  63 - 0x3f
      11'h68C: dout  = 8'b00000011; // 1676 :   3 - 0x3
      11'h68D: dout  = 8'b00001100; // 1677 :  12 - 0xc
      11'h68E: dout  = 8'b00001110; // 1678 :  14 - 0xe
      11'h68F: dout  = 8'b00000000; // 1679 :   0 - 0x0
      11'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0xd2
      11'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      11'h692: dout  = 8'b00000000; // 1682 :   0 - 0x0
      11'h693: dout  = 8'b00001000; // 1683 :   8 - 0x8
      11'h694: dout  = 8'b11011000; // 1684 : 216 - 0xd8
      11'h695: dout  = 8'b11111100; // 1685 : 252 - 0xfc
      11'h696: dout  = 8'b11111100; // 1686 : 252 - 0xfc
      11'h697: dout  = 8'b10011100; // 1687 : 156 - 0x9c
      11'h698: dout  = 8'b00001100; // 1688 :  12 - 0xc -- Sprite 0xd3
      11'h699: dout  = 8'b10011100; // 1689 : 156 - 0x9c
      11'h69A: dout  = 8'b11111000; // 1690 : 248 - 0xf8
      11'h69B: dout  = 8'b01111000; // 1691 : 120 - 0x78
      11'h69C: dout  = 8'b10001000; // 1692 : 136 - 0x88
      11'h69D: dout  = 8'b00110000; // 1693 :  48 - 0x30
      11'h69E: dout  = 8'b00111000; // 1694 :  56 - 0x38
      11'h69F: dout  = 8'b00000000; // 1695 :   0 - 0x0
      11'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      11'h6A1: dout  = 8'b00000000; // 1697 :   0 - 0x0
      11'h6A2: dout  = 8'b00000000; // 1698 :   0 - 0x0
      11'h6A3: dout  = 8'b00000000; // 1699 :   0 - 0x0
      11'h6A4: dout  = 8'b00000001; // 1700 :   1 - 0x1
      11'h6A5: dout  = 8'b00001011; // 1701 :  11 - 0xb
      11'h6A6: dout  = 8'b00011111; // 1702 :  31 - 0x1f
      11'h6A7: dout  = 8'b00111001; // 1703 :  57 - 0x39
      11'h6A8: dout  = 8'b01110000; // 1704 : 112 - 0x70 -- Sprite 0xd5
      11'h6A9: dout  = 8'b01111000; // 1705 : 120 - 0x78
      11'h6AA: dout  = 8'b00111111; // 1706 :  63 - 0x3f
      11'h6AB: dout  = 8'b00111111; // 1707 :  63 - 0x3f
      11'h6AC: dout  = 8'b00000011; // 1708 :   3 - 0x3
      11'h6AD: dout  = 8'b00111000; // 1709 :  56 - 0x38
      11'h6AE: dout  = 8'b00011100; // 1710 :  28 - 0x1c
      11'h6AF: dout  = 8'b00000000; // 1711 :   0 - 0x0
      11'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      11'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      11'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      11'h6B3: dout  = 8'b11000000; // 1715 : 192 - 0xc0
      11'h6B4: dout  = 8'b11001000; // 1716 : 200 - 0xc8
      11'h6B5: dout  = 8'b11111000; // 1717 : 248 - 0xf8
      11'h6B6: dout  = 8'b11111100; // 1718 : 252 - 0xfc
      11'h6B7: dout  = 8'b10011100; // 1719 : 156 - 0x9c
      11'h6B8: dout  = 8'b00001100; // 1720 :  12 - 0xc -- Sprite 0xd7
      11'h6B9: dout  = 8'b10011100; // 1721 : 156 - 0x9c
      11'h6BA: dout  = 8'b11111000; // 1722 : 248 - 0xf8
      11'h6BB: dout  = 8'b01111000; // 1723 : 120 - 0x78
      11'h6BC: dout  = 8'b11100010; // 1724 : 226 - 0xe2
      11'h6BD: dout  = 8'b00011110; // 1725 :  30 - 0x1e
      11'h6BE: dout  = 8'b00001100; // 1726 :  12 - 0xc
      11'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      11'h6C0: dout  = 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0xd8
      11'h6C1: dout  = 8'b00110000; // 1729 :  48 - 0x30
      11'h6C2: dout  = 8'b00111100; // 1730 :  60 - 0x3c
      11'h6C3: dout  = 8'b01111100; // 1731 : 124 - 0x7c
      11'h6C4: dout  = 8'b01111100; // 1732 : 124 - 0x7c
      11'h6C5: dout  = 8'b00111110; // 1733 :  62 - 0x3e
      11'h6C6: dout  = 8'b00011100; // 1734 :  28 - 0x1c
      11'h6C7: dout  = 8'b00000000; // 1735 :   0 - 0x0
      11'h6C8: dout  = 8'b00000000; // 1736 :   0 - 0x0 -- Sprite 0xd9
      11'h6C9: dout  = 8'b00001110; // 1737 :  14 - 0xe
      11'h6CA: dout  = 8'b00111110; // 1738 :  62 - 0x3e
      11'h6CB: dout  = 8'b01111110; // 1739 : 126 - 0x7e
      11'h6CC: dout  = 8'b01111110; // 1740 : 126 - 0x7e
      11'h6CD: dout  = 8'b00111100; // 1741 :  60 - 0x3c
      11'h6CE: dout  = 8'b00001100; // 1742 :  12 - 0xc
      11'h6CF: dout  = 8'b00000000; // 1743 :   0 - 0x0
      11'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0xda
      11'h6D1: dout  = 8'b00100000; // 1745 :  32 - 0x20
      11'h6D2: dout  = 8'b01111110; // 1746 : 126 - 0x7e
      11'h6D3: dout  = 8'b01111110; // 1747 : 126 - 0x7e
      11'h6D4: dout  = 8'b01111110; // 1748 : 126 - 0x7e
      11'h6D5: dout  = 8'b00111100; // 1749 :  60 - 0x3c
      11'h6D6: dout  = 8'b00111000; // 1750 :  56 - 0x38
      11'h6D7: dout  = 8'b00000000; // 1751 :   0 - 0x0
      11'h6D8: dout  = 8'b00000000; // 1752 :   0 - 0x0 -- Sprite 0xdb
      11'h6D9: dout  = 8'b00011100; // 1753 :  28 - 0x1c
      11'h6DA: dout  = 8'b00111110; // 1754 :  62 - 0x3e
      11'h6DB: dout  = 8'b01111110; // 1755 : 126 - 0x7e
      11'h6DC: dout  = 8'b01111110; // 1756 : 126 - 0x7e
      11'h6DD: dout  = 8'b00111100; // 1757 :  60 - 0x3c
      11'h6DE: dout  = 8'b00010000; // 1758 :  16 - 0x10
      11'h6DF: dout  = 8'b00000000; // 1759 :   0 - 0x0
      11'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0xdc
      11'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      11'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      11'h6E3: dout  = 8'b00000001; // 1763 :   1 - 0x1
      11'h6E4: dout  = 8'b00000011; // 1764 :   3 - 0x3
      11'h6E5: dout  = 8'b00000001; // 1765 :   1 - 0x1
      11'h6E6: dout  = 8'b00000001; // 1766 :   1 - 0x1
      11'h6E7: dout  = 8'b00001111; // 1767 :  15 - 0xf
      11'h6E8: dout  = 8'b00000111; // 1768 :   7 - 0x7 -- Sprite 0xdd
      11'h6E9: dout  = 8'b00000111; // 1769 :   7 - 0x7
      11'h6EA: dout  = 8'b00000111; // 1770 :   7 - 0x7
      11'h6EB: dout  = 8'b00011111; // 1771 :  31 - 0x1f
      11'h6EC: dout  = 8'b00001111; // 1772 :  15 - 0xf
      11'h6ED: dout  = 8'b00000111; // 1773 :   7 - 0x7
      11'h6EE: dout  = 8'b00000011; // 1774 :   3 - 0x3
      11'h6EF: dout  = 8'b00000000; // 1775 :   0 - 0x0
      11'h6F0: dout  = 8'b00000000; // 1776 :   0 - 0x0 -- Sprite 0xde
      11'h6F1: dout  = 8'b00000000; // 1777 :   0 - 0x0
      11'h6F2: dout  = 8'b00000000; // 1778 :   0 - 0x0
      11'h6F3: dout  = 8'b00000000; // 1779 :   0 - 0x0
      11'h6F4: dout  = 8'b10000000; // 1780 : 128 - 0x80
      11'h6F5: dout  = 8'b10000000; // 1781 : 128 - 0x80
      11'h6F6: dout  = 8'b10010000; // 1782 : 144 - 0x90
      11'h6F7: dout  = 8'b11110000; // 1783 : 240 - 0xf0
      11'h6F8: dout  = 8'b11100000; // 1784 : 224 - 0xe0 -- Sprite 0xdf
      11'h6F9: dout  = 8'b11100000; // 1785 : 224 - 0xe0
      11'h6FA: dout  = 8'b11110000; // 1786 : 240 - 0xf0
      11'h6FB: dout  = 8'b11110000; // 1787 : 240 - 0xf0
      11'h6FC: dout  = 8'b11100000; // 1788 : 224 - 0xe0
      11'h6FD: dout  = 8'b11000000; // 1789 : 192 - 0xc0
      11'h6FE: dout  = 8'b11000000; // 1790 : 192 - 0xc0
      11'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      11'h700: dout  = 8'b00001111; // 1792 :  15 - 0xf -- Sprite 0xe0
      11'h701: dout  = 8'b00011111; // 1793 :  31 - 0x1f
      11'h702: dout  = 8'b00011111; // 1794 :  31 - 0x1f
      11'h703: dout  = 8'b00111111; // 1795 :  63 - 0x3f
      11'h704: dout  = 8'b01111111; // 1796 : 127 - 0x7f
      11'h705: dout  = 8'b11111111; // 1797 : 255 - 0xff
      11'h706: dout  = 8'b11111111; // 1798 : 255 - 0xff
      11'h707: dout  = 8'b11111111; // 1799 : 255 - 0xff
      11'h708: dout  = 8'b11111111; // 1800 : 255 - 0xff -- Sprite 0xe1
      11'h709: dout  = 8'b11111111; // 1801 : 255 - 0xff
      11'h70A: dout  = 8'b01111111; // 1802 : 127 - 0x7f
      11'h70B: dout  = 8'b00111111; // 1803 :  63 - 0x3f
      11'h70C: dout  = 8'b00111111; // 1804 :  63 - 0x3f
      11'h70D: dout  = 8'b00011111; // 1805 :  31 - 0x1f
      11'h70E: dout  = 8'b00001111; // 1806 :  15 - 0xf
      11'h70F: dout  = 8'b00000111; // 1807 :   7 - 0x7
      11'h710: dout  = 8'b11111110; // 1808 : 254 - 0xfe -- Sprite 0xe2
      11'h711: dout  = 8'b11111111; // 1809 : 255 - 0xff
      11'h712: dout  = 8'b11111111; // 1810 : 255 - 0xff
      11'h713: dout  = 8'b00001111; // 1811 :  15 - 0xf
      11'h714: dout  = 8'b10111111; // 1812 : 191 - 0xbf
      11'h715: dout  = 8'b10100011; // 1813 : 163 - 0xa3
      11'h716: dout  = 8'b11110111; // 1814 : 247 - 0xf7
      11'h717: dout  = 8'b11110111; // 1815 : 247 - 0xf7
      11'h718: dout  = 8'b11111111; // 1816 : 255 - 0xff -- Sprite 0xe3
      11'h719: dout  = 8'b11111111; // 1817 : 255 - 0xff
      11'h71A: dout  = 8'b00111111; // 1818 :  63 - 0x3f
      11'h71B: dout  = 8'b00011111; // 1819 :  31 - 0x1f
      11'h71C: dout  = 8'b11111110; // 1820 : 254 - 0xfe
      11'h71D: dout  = 8'b11111100; // 1821 : 252 - 0xfc
      11'h71E: dout  = 8'b11111000; // 1822 : 248 - 0xf8
      11'h71F: dout  = 8'b11110000; // 1823 : 240 - 0xf0
      11'h720: dout  = 8'b00001111; // 1824 :  15 - 0xf -- Sprite 0xe4
      11'h721: dout  = 8'b00011111; // 1825 :  31 - 0x1f
      11'h722: dout  = 8'b00011111; // 1826 :  31 - 0x1f
      11'h723: dout  = 8'b00111111; // 1827 :  63 - 0x3f
      11'h724: dout  = 8'b01111111; // 1828 : 127 - 0x7f
      11'h725: dout  = 8'b11111111; // 1829 : 255 - 0xff
      11'h726: dout  = 8'b11111111; // 1830 : 255 - 0xff
      11'h727: dout  = 8'b11111111; // 1831 : 255 - 0xff
      11'h728: dout  = 8'b11111111; // 1832 : 255 - 0xff -- Sprite 0xe5
      11'h729: dout  = 8'b11111111; // 1833 : 255 - 0xff
      11'h72A: dout  = 8'b01111110; // 1834 : 126 - 0x7e
      11'h72B: dout  = 8'b00111111; // 1835 :  63 - 0x3f
      11'h72C: dout  = 8'b00111111; // 1836 :  63 - 0x3f
      11'h72D: dout  = 8'b00011111; // 1837 :  31 - 0x1f
      11'h72E: dout  = 8'b00001111; // 1838 :  15 - 0xf
      11'h72F: dout  = 8'b00000111; // 1839 :   7 - 0x7
      11'h730: dout  = 8'b11111110; // 1840 : 254 - 0xfe -- Sprite 0xe6
      11'h731: dout  = 8'b11111111; // 1841 : 255 - 0xff
      11'h732: dout  = 8'b11111111; // 1842 : 255 - 0xff
      11'h733: dout  = 8'b11100011; // 1843 : 227 - 0xe3
      11'h734: dout  = 8'b00010111; // 1844 :  23 - 0x17
      11'h735: dout  = 8'b10110111; // 1845 : 183 - 0xb7
      11'h736: dout  = 8'b10111111; // 1846 : 191 - 0xbf
      11'h737: dout  = 8'b11111111; // 1847 : 255 - 0xff
      11'h738: dout  = 8'b11111111; // 1848 : 255 - 0xff -- Sprite 0xe7
      11'h739: dout  = 8'b11111111; // 1849 : 255 - 0xff
      11'h73A: dout  = 8'b00111111; // 1850 :  63 - 0x3f
      11'h73B: dout  = 8'b00001111; // 1851 :  15 - 0xf
      11'h73C: dout  = 8'b00001110; // 1852 :  14 - 0xe
      11'h73D: dout  = 8'b11111100; // 1853 : 252 - 0xfc
      11'h73E: dout  = 8'b11111000; // 1854 : 248 - 0xf8
      11'h73F: dout  = 8'b11110000; // 1855 : 240 - 0xf0
      11'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0xe8
      11'h741: dout  = 8'b00000101; // 1857 :   5 - 0x5
      11'h742: dout  = 8'b00000111; // 1858 :   7 - 0x7
      11'h743: dout  = 8'b00000011; // 1859 :   3 - 0x3
      11'h744: dout  = 8'b00000000; // 1860 :   0 - 0x0
      11'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      11'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      11'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      11'h748: dout  = 8'b00000000; // 1864 :   0 - 0x0 -- Sprite 0xe9
      11'h749: dout  = 8'b00000000; // 1865 :   0 - 0x0
      11'h74A: dout  = 8'b00000000; // 1866 :   0 - 0x0
      11'h74B: dout  = 8'b00000000; // 1867 :   0 - 0x0
      11'h74C: dout  = 8'b00000000; // 1868 :   0 - 0x0
      11'h74D: dout  = 8'b00000000; // 1869 :   0 - 0x0
      11'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      11'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      11'h750: dout  = 8'b00000011; // 1872 :   3 - 0x3 -- Sprite 0xea
      11'h751: dout  = 8'b10011110; // 1873 : 158 - 0x9e
      11'h752: dout  = 8'b00001110; // 1874 :  14 - 0xe
      11'h753: dout  = 8'b00000000; // 1875 :   0 - 0x0
      11'h754: dout  = 8'b00000000; // 1876 :   0 - 0x0
      11'h755: dout  = 8'b00000000; // 1877 :   0 - 0x0
      11'h756: dout  = 8'b00000000; // 1878 :   0 - 0x0
      11'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      11'h758: dout  = 8'b00000000; // 1880 :   0 - 0x0 -- Sprite 0xeb
      11'h759: dout  = 8'b00000000; // 1881 :   0 - 0x0
      11'h75A: dout  = 8'b00000000; // 1882 :   0 - 0x0
      11'h75B: dout  = 8'b00000000; // 1883 :   0 - 0x0
      11'h75C: dout  = 8'b00000000; // 1884 :   0 - 0x0
      11'h75D: dout  = 8'b00000000; // 1885 :   0 - 0x0
      11'h75E: dout  = 8'b00000000; // 1886 :   0 - 0x0
      11'h75F: dout  = 8'b00000000; // 1887 :   0 - 0x0
      11'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      11'h761: dout  = 8'b00000000; // 1889 :   0 - 0x0
      11'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      11'h763: dout  = 8'b00000000; // 1891 :   0 - 0x0
      11'h764: dout  = 8'b00000100; // 1892 :   4 - 0x4
      11'h765: dout  = 8'b00001110; // 1893 :  14 - 0xe
      11'h766: dout  = 8'b00001111; // 1894 :  15 - 0xf
      11'h767: dout  = 8'b00001011; // 1895 :  11 - 0xb
      11'h768: dout  = 8'b00001111; // 1896 :  15 - 0xf -- Sprite 0xed
      11'h769: dout  = 8'b00001100; // 1897 :  12 - 0xc
      11'h76A: dout  = 8'b00001111; // 1898 :  15 - 0xf
      11'h76B: dout  = 8'b00001111; // 1899 :  15 - 0xf
      11'h76C: dout  = 8'b00000000; // 1900 :   0 - 0x0
      11'h76D: dout  = 8'b01111111; // 1901 : 127 - 0x7f
      11'h76E: dout  = 8'b11010101; // 1902 : 213 - 0xd5
      11'h76F: dout  = 8'b01111111; // 1903 : 127 - 0x7f
      11'h770: dout  = 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0xee
      11'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      11'h772: dout  = 8'b00000000; // 1906 :   0 - 0x0
      11'h773: dout  = 8'b00000000; // 1907 :   0 - 0x0
      11'h774: dout  = 8'b00100000; // 1908 :  32 - 0x20
      11'h775: dout  = 8'b01110000; // 1909 : 112 - 0x70
      11'h776: dout  = 8'b11110000; // 1910 : 240 - 0xf0
      11'h777: dout  = 8'b11100000; // 1911 : 224 - 0xe0
      11'h778: dout  = 8'b11110000; // 1912 : 240 - 0xf0 -- Sprite 0xef
      11'h779: dout  = 8'b00110000; // 1913 :  48 - 0x30
      11'h77A: dout  = 8'b11110000; // 1914 : 240 - 0xf0
      11'h77B: dout  = 8'b11110000; // 1915 : 240 - 0xf0
      11'h77C: dout  = 8'b00000000; // 1916 :   0 - 0x0
      11'h77D: dout  = 8'b11111110; // 1917 : 254 - 0xfe
      11'h77E: dout  = 8'b01010101; // 1918 :  85 - 0x55
      11'h77F: dout  = 8'b11111110; // 1919 : 254 - 0xfe
      11'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      11'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      11'h782: dout  = 8'b00000000; // 1922 :   0 - 0x0
      11'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      11'h784: dout  = 8'b00000100; // 1924 :   4 - 0x4
      11'h785: dout  = 8'b00001110; // 1925 :  14 - 0xe
      11'h786: dout  = 8'b00001111; // 1926 :  15 - 0xf
      11'h787: dout  = 8'b00001011; // 1927 :  11 - 0xb
      11'h788: dout  = 8'b00001111; // 1928 :  15 - 0xf -- Sprite 0xf1
      11'h789: dout  = 8'b00001100; // 1929 :  12 - 0xc
      11'h78A: dout  = 8'b00001111; // 1930 :  15 - 0xf
      11'h78B: dout  = 8'b00001111; // 1931 :  15 - 0xf
      11'h78C: dout  = 8'b00000000; // 1932 :   0 - 0x0
      11'h78D: dout  = 8'b01111111; // 1933 : 127 - 0x7f
      11'h78E: dout  = 8'b10101010; // 1934 : 170 - 0xaa
      11'h78F: dout  = 8'b01111111; // 1935 : 127 - 0x7f
      11'h790: dout  = 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0xf2
      11'h791: dout  = 8'b00000000; // 1937 :   0 - 0x0
      11'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      11'h793: dout  = 8'b00000000; // 1939 :   0 - 0x0
      11'h794: dout  = 8'b00100000; // 1940 :  32 - 0x20
      11'h795: dout  = 8'b01110000; // 1941 : 112 - 0x70
      11'h796: dout  = 8'b11110000; // 1942 : 240 - 0xf0
      11'h797: dout  = 8'b11100000; // 1943 : 224 - 0xe0
      11'h798: dout  = 8'b11110000; // 1944 : 240 - 0xf0 -- Sprite 0xf3
      11'h799: dout  = 8'b00110000; // 1945 :  48 - 0x30
      11'h79A: dout  = 8'b11110000; // 1946 : 240 - 0xf0
      11'h79B: dout  = 8'b11110000; // 1947 : 240 - 0xf0
      11'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      11'h79D: dout  = 8'b11111110; // 1949 : 254 - 0xfe
      11'h79E: dout  = 8'b10101011; // 1950 : 171 - 0xab
      11'h79F: dout  = 8'b11111110; // 1951 : 254 - 0xfe
      11'h7A0: dout  = 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0xf4
      11'h7A1: dout  = 8'b00010101; // 1953 :  21 - 0x15
      11'h7A2: dout  = 8'b00001010; // 1954 :  10 - 0xa
      11'h7A3: dout  = 8'b00000101; // 1955 :   5 - 0x5
      11'h7A4: dout  = 8'b00000010; // 1956 :   2 - 0x2
      11'h7A5: dout  = 8'b00000101; // 1957 :   5 - 0x5
      11'h7A6: dout  = 8'b00000111; // 1958 :   7 - 0x7
      11'h7A7: dout  = 8'b00000111; // 1959 :   7 - 0x7
      11'h7A8: dout  = 8'b00111100; // 1960 :  60 - 0x3c -- Sprite 0xf5
      11'h7A9: dout  = 8'b01111011; // 1961 : 123 - 0x7b
      11'h7AA: dout  = 8'b01111011; // 1962 : 123 - 0x7b
      11'h7AB: dout  = 8'b01111111; // 1963 : 127 - 0x7f
      11'h7AC: dout  = 8'b01111110; // 1964 : 126 - 0x7e
      11'h7AD: dout  = 8'b01111111; // 1965 : 127 - 0x7f
      11'h7AE: dout  = 8'b00111110; // 1966 :  62 - 0x3e
      11'h7AF: dout  = 8'b00000000; // 1967 :   0 - 0x0
      11'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      11'h7B1: dout  = 8'b01010000; // 1969 :  80 - 0x50
      11'h7B2: dout  = 8'b10100000; // 1970 : 160 - 0xa0
      11'h7B3: dout  = 8'b01000000; // 1971 :  64 - 0x40
      11'h7B4: dout  = 8'b10100000; // 1972 : 160 - 0xa0
      11'h7B5: dout  = 8'b01000000; // 1973 :  64 - 0x40
      11'h7B6: dout  = 8'b11100000; // 1974 : 224 - 0xe0
      11'h7B7: dout  = 8'b11100000; // 1975 : 224 - 0xe0
      11'h7B8: dout  = 8'b01111000; // 1976 : 120 - 0x78 -- Sprite 0xf7
      11'h7B9: dout  = 8'b10111100; // 1977 : 188 - 0xbc
      11'h7BA: dout  = 8'b10111000; // 1978 : 184 - 0xb8
      11'h7BB: dout  = 8'b10111110; // 1979 : 190 - 0xbe
      11'h7BC: dout  = 8'b01111100; // 1980 : 124 - 0x7c
      11'h7BD: dout  = 8'b11111110; // 1981 : 254 - 0xfe
      11'h7BE: dout  = 8'b01111000; // 1982 : 120 - 0x78
      11'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      11'h7C0: dout  = 8'b00000011; // 1984 :   3 - 0x3 -- Sprite 0xf8
      11'h7C1: dout  = 8'b00000011; // 1985 :   3 - 0x3
      11'h7C2: dout  = 8'b00000000; // 1986 :   0 - 0x0
      11'h7C3: dout  = 8'b00000011; // 1987 :   3 - 0x3
      11'h7C4: dout  = 8'b00000111; // 1988 :   7 - 0x7
      11'h7C5: dout  = 8'b00000110; // 1989 :   6 - 0x6
      11'h7C6: dout  = 8'b00000111; // 1990 :   7 - 0x7
      11'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0 -- Sprite 0xf9
      11'h7C9: dout  = 8'b00011111; // 1993 :  31 - 0x1f
      11'h7CA: dout  = 8'b00011111; // 1994 :  31 - 0x1f
      11'h7CB: dout  = 8'b00001111; // 1995 :  15 - 0xf
      11'h7CC: dout  = 8'b00000011; // 1996 :   3 - 0x3
      11'h7CD: dout  = 8'b00000000; // 1997 :   0 - 0x0
      11'h7CE: dout  = 8'b00000000; // 1998 :   0 - 0x0
      11'h7CF: dout  = 8'b00000000; // 1999 :   0 - 0x0
      11'h7D0: dout  = 8'b11100000; // 2000 : 224 - 0xe0 -- Sprite 0xfa
      11'h7D1: dout  = 8'b11100000; // 2001 : 224 - 0xe0
      11'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      11'h7D3: dout  = 8'b00110000; // 2003 :  48 - 0x30
      11'h7D4: dout  = 8'b01110000; // 2004 : 112 - 0x70
      11'h7D5: dout  = 8'b01100000; // 2005 :  96 - 0x60
      11'h7D6: dout  = 8'b01110000; // 2006 : 112 - 0x70
      11'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0 -- Sprite 0xfb
      11'h7D9: dout  = 8'b11111000; // 2009 : 248 - 0xf8
      11'h7DA: dout  = 8'b11111000; // 2010 : 248 - 0xf8
      11'h7DB: dout  = 8'b11110000; // 2011 : 240 - 0xf0
      11'h7DC: dout  = 8'b11000000; // 2012 : 192 - 0xc0
      11'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      11'h7DE: dout  = 8'b00000000; // 2014 :   0 - 0x0
      11'h7DF: dout  = 8'b00000000; // 2015 :   0 - 0x0
      11'h7E0: dout  = 8'b00111000; // 2016 :  56 - 0x38 -- Sprite 0xfc
      11'h7E1: dout  = 8'b00111000; // 2017 :  56 - 0x38
      11'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      11'h7E3: dout  = 8'b01111100; // 2019 : 124 - 0x7c
      11'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      11'h7E5: dout  = 8'b00111000; // 2021 :  56 - 0x38
      11'h7E6: dout  = 8'b00111000; // 2022 :  56 - 0x38
      11'h7E7: dout  = 8'b01111100; // 2023 : 124 - 0x7c
      11'h7E8: dout  = 8'b01111100; // 2024 : 124 - 0x7c -- Sprite 0xfd
      11'h7E9: dout  = 8'b01111100; // 2025 : 124 - 0x7c
      11'h7EA: dout  = 8'b01111100; // 2026 : 124 - 0x7c
      11'h7EB: dout  = 8'b00111000; // 2027 :  56 - 0x38
      11'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      11'h7ED: dout  = 8'b01111100; // 2029 : 124 - 0x7c
      11'h7EE: dout  = 8'b01111100; // 2030 : 124 - 0x7c
      11'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0xfe
      11'h7F1: dout  = 8'b00000000; // 2033 :   0 - 0x0
      11'h7F2: dout  = 8'b00010001; // 2034 :  17 - 0x11
      11'h7F3: dout  = 8'b11010111; // 2035 : 215 - 0xd7
      11'h7F4: dout  = 8'b11010111; // 2036 : 215 - 0xd7
      11'h7F5: dout  = 8'b11010111; // 2037 : 215 - 0xd7
      11'h7F6: dout  = 8'b00010001; // 2038 :  17 - 0x11
      11'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      11'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      11'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      11'h7FA: dout  = 8'b11100110; // 2042 : 230 - 0xe6
      11'h7FB: dout  = 8'b11110110; // 2043 : 246 - 0xf6
      11'h7FC: dout  = 8'b11110110; // 2044 : 246 - 0xf6
      11'h7FD: dout  = 8'b11110110; // 2045 : 246 - 0xf6
      11'h7FE: dout  = 8'b11100110; // 2046 : 230 - 0xe6
      11'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
    endcase
  end

endmodule
