---   Sprites Pattern table COLOR PLANE 0
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: nova_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_NOVA_SPR_PLN0 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_NOVA_SPR_PLN0;

architecture BEHAVIORAL of ROM_PTABLE_NOVA_SPR_PLN0 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table COLOR PLANE 0
    "11111111", --    0 -  0x0  :  255 - 0xff -- Sprite 0x0
    "11111111", --    1 -  0x1  :  255 - 0xff
    "11000000", --    2 -  0x2  :  192 - 0xc0
    "11000000", --    3 -  0x3  :  192 - 0xc0
    "11000000", --    4 -  0x4  :  192 - 0xc0
    "11000000", --    5 -  0x5  :  192 - 0xc0
    "11010101", --    6 -  0x6  :  213 - 0xd5
    "11111111", --    7 -  0x7  :  255 - 0xff
    "11111111", --    8 -  0x8  :  255 - 0xff -- Sprite 0x1
    "11111111", --    9 -  0x9  :  255 - 0xff
    "11001110", --   10 -  0xa  :  206 - 0xce
    "11000110", --   11 -  0xb  :  198 - 0xc6
    "11001110", --   12 -  0xc  :  206 - 0xce
    "11000110", --   13 -  0xd  :  198 - 0xc6
    "11101110", --   14 -  0xe  :  238 - 0xee
    "11111111", --   15 -  0xf  :  255 - 0xff
    "11111111", --   16 - 0x10  :  255 - 0xff -- Sprite 0x2
    "11111111", --   17 - 0x11  :  255 - 0xff
    "01110001", --   18 - 0x12  :  113 - 0x71
    "00110011", --   19 - 0x13  :   51 - 0x33
    "01110001", --   20 - 0x14  :  113 - 0x71
    "00110011", --   21 - 0x15  :   51 - 0x33
    "01110101", --   22 - 0x16  :  117 - 0x75
    "11111111", --   23 - 0x17  :  255 - 0xff
    "11111111", --   24 - 0x18  :  255 - 0xff -- Sprite 0x3
    "11111111", --   25 - 0x19  :  255 - 0xff
    "00000011", --   26 - 0x1a  :    3 - 0x3
    "00000001", --   27 - 0x1b  :    1 - 0x1
    "00000011", --   28 - 0x1c  :    3 - 0x3
    "00000001", --   29 - 0x1d  :    1 - 0x1
    "10101011", --   30 - 0x1e  :  171 - 0xab
    "11111111", --   31 - 0x1f  :  255 - 0xff
    "11111111", --   32 - 0x20  :  255 - 0xff -- Sprite 0x4
    "11111111", --   33 - 0x21  :  255 - 0xff
    "11100000", --   34 - 0x22  :  224 - 0xe0
    "11000110", --   35 - 0x23  :  198 - 0xc6
    "11000110", --   36 - 0x24  :  198 - 0xc6
    "11110110", --   37 - 0x25  :  246 - 0xf6
    "11110000", --   38 - 0x26  :  240 - 0xf0
    "11110001", --   39 - 0x27  :  241 - 0xf1
    "11000111", --   40 - 0x28  :  199 - 0xc7 -- Sprite 0x5
    "11001111", --   41 - 0x29  :  207 - 0xcf
    "11011111", --   42 - 0x2a  :  223 - 0xdf
    "11011111", --   43 - 0x2b  :  223 - 0xdf
    "11001110", --   44 - 0x2c  :  206 - 0xce
    "11100000", --   45 - 0x2d  :  224 - 0xe0
    "11111111", --   46 - 0x2e  :  255 - 0xff
    "11111111", --   47 - 0x2f  :  255 - 0xff
    "11111111", --   48 - 0x30  :  255 - 0xff -- Sprite 0x6
    "11111111", --   49 - 0x31  :  255 - 0xff
    "00000111", --   50 - 0x32  :    7 - 0x7
    "01100011", --   51 - 0x33  :   99 - 0x63
    "01100011", --   52 - 0x34  :   99 - 0x63
    "01101111", --   53 - 0x35  :  111 - 0x6f
    "00001111", --   54 - 0x36  :   15 - 0xf
    "10001111", --   55 - 0x37  :  143 - 0x8f
    "11100011", --   56 - 0x38  :  227 - 0xe3 -- Sprite 0x7
    "11110011", --   57 - 0x39  :  243 - 0xf3
    "11111011", --   58 - 0x3a  :  251 - 0xfb
    "11111011", --   59 - 0x3b  :  251 - 0xfb
    "01110011", --   60 - 0x3c  :  115 - 0x73
    "00000111", --   61 - 0x3d  :    7 - 0x7
    "11111111", --   62 - 0x3e  :  255 - 0xff
    "11111111", --   63 - 0x3f  :  255 - 0xff
    "11111111", --   64 - 0x40  :  255 - 0xff -- Sprite 0x8
    "11010101", --   65 - 0x41  :  213 - 0xd5
    "10101010", --   66 - 0x42  :  170 - 0xaa
    "11010101", --   67 - 0x43  :  213 - 0xd5
    "10101010", --   68 - 0x44  :  170 - 0xaa
    "11010101", --   69 - 0x45  :  213 - 0xd5
    "10101010", --   70 - 0x46  :  170 - 0xaa
    "11010101", --   71 - 0x47  :  213 - 0xd5
    "10101010", --   72 - 0x48  :  170 - 0xaa -- Sprite 0x9
    "11010101", --   73 - 0x49  :  213 - 0xd5
    "10101010", --   74 - 0x4a  :  170 - 0xaa
    "11010101", --   75 - 0x4b  :  213 - 0xd5
    "10101010", --   76 - 0x4c  :  170 - 0xaa
    "11110101", --   77 - 0x4d  :  245 - 0xf5
    "10101010", --   78 - 0x4e  :  170 - 0xaa
    "11111111", --   79 - 0x4f  :  255 - 0xff
    "11111111", --   80 - 0x50  :  255 - 0xff -- Sprite 0xa
    "01010101", --   81 - 0x51  :   85 - 0x55
    "10101111", --   82 - 0x52  :  175 - 0xaf
    "01010101", --   83 - 0x53  :   85 - 0x55
    "10101011", --   84 - 0x54  :  171 - 0xab
    "01010101", --   85 - 0x55  :   85 - 0x55
    "10101011", --   86 - 0x56  :  171 - 0xab
    "01010101", --   87 - 0x57  :   85 - 0x55
    "10101011", --   88 - 0x58  :  171 - 0xab -- Sprite 0xb
    "01010101", --   89 - 0x59  :   85 - 0x55
    "10101011", --   90 - 0x5a  :  171 - 0xab
    "01010101", --   91 - 0x5b  :   85 - 0x55
    "10101011", --   92 - 0x5c  :  171 - 0xab
    "01010101", --   93 - 0x5d  :   85 - 0x55
    "10101011", --   94 - 0x5e  :  171 - 0xab
    "11111111", --   95 - 0x5f  :  255 - 0xff
    "11111111", --   96 - 0x60  :  255 - 0xff -- Sprite 0xc
    "11010101", --   97 - 0x61  :  213 - 0xd5
    "10100000", --   98 - 0x62  :  160 - 0xa0
    "11010000", --   99 - 0x63  :  208 - 0xd0
    "10001111", --  100 - 0x64  :  143 - 0x8f
    "11001000", --  101 - 0x65  :  200 - 0xc8
    "10001000", --  102 - 0x66  :  136 - 0x88
    "11001000", --  103 - 0x67  :  200 - 0xc8
    "10001000", --  104 - 0x68  :  136 - 0x88 -- Sprite 0xd
    "11001000", --  105 - 0x69  :  200 - 0xc8
    "10001000", --  106 - 0x6a  :  136 - 0x88
    "11001111", --  107 - 0x6b  :  207 - 0xcf
    "10010000", --  108 - 0x6c  :  144 - 0x90
    "11100000", --  109 - 0x6d  :  224 - 0xe0
    "11101010", --  110 - 0x6e  :  234 - 0xea
    "11111111", --  111 - 0x6f  :  255 - 0xff
    "11111111", --  112 - 0x70  :  255 - 0xff -- Sprite 0xe
    "01011011", --  113 - 0x71  :   91 - 0x5b
    "00000111", --  114 - 0x72  :    7 - 0x7
    "00001001", --  115 - 0x73  :    9 - 0x9
    "11110011", --  116 - 0x74  :  243 - 0xf3
    "00010001", --  117 - 0x75  :   17 - 0x11
    "00010011", --  118 - 0x76  :   19 - 0x13
    "00010001", --  119 - 0x77  :   17 - 0x11
    "00010011", --  120 - 0x78  :   19 - 0x13 -- Sprite 0xf
    "00010001", --  121 - 0x79  :   17 - 0x11
    "00010011", --  122 - 0x7a  :   19 - 0x13
    "11110001", --  123 - 0x7b  :  241 - 0xf1
    "00001011", --  124 - 0x7c  :   11 - 0xb
    "00000101", --  125 - 0x7d  :    5 - 0x5
    "10101011", --  126 - 0x7e  :  171 - 0xab
    "11111111", --  127 - 0x7f  :  255 - 0xff
    "11010000", --  128 - 0x80  :  208 - 0xd0 -- Sprite 0x10
    "10010000", --  129 - 0x81  :  144 - 0x90
    "11011111", --  130 - 0x82  :  223 - 0xdf
    "10011010", --  131 - 0x83  :  154 - 0x9a
    "11010101", --  132 - 0x84  :  213 - 0xd5
    "10011111", --  133 - 0x85  :  159 - 0x9f
    "11010000", --  134 - 0x86  :  208 - 0xd0
    "10010000", --  135 - 0x87  :  144 - 0x90
    "00001001", --  136 - 0x88  :    9 - 0x9 -- Sprite 0x11
    "00001011", --  137 - 0x89  :   11 - 0xb
    "11111001", --  138 - 0x8a  :  249 - 0xf9
    "10101011", --  139 - 0x8b  :  171 - 0xab
    "01011001", --  140 - 0x8c  :   89 - 0x59
    "11111011", --  141 - 0x8d  :  251 - 0xfb
    "00001001", --  142 - 0x8e  :    9 - 0x9
    "00001011", --  143 - 0x8f  :   11 - 0xb
    "00011000", --  144 - 0x90  :   24 - 0x18 -- Sprite 0x12
    "00010100", --  145 - 0x91  :   20 - 0x14
    "00010100", --  146 - 0x92  :   20 - 0x14
    "00111010", --  147 - 0x93  :   58 - 0x3a
    "00111010", --  148 - 0x94  :   58 - 0x3a
    "01111010", --  149 - 0x95  :  122 - 0x7a
    "01111010", --  150 - 0x96  :  122 - 0x7a
    "01111010", --  151 - 0x97  :  122 - 0x7a
    "11111011", --  152 - 0x98  :  251 - 0xfb -- Sprite 0x13
    "11111101", --  153 - 0x99  :  253 - 0xfd
    "11111101", --  154 - 0x9a  :  253 - 0xfd
    "11111101", --  155 - 0x9b  :  253 - 0xfd
    "11111101", --  156 - 0x9c  :  253 - 0xfd
    "11111101", --  157 - 0x9d  :  253 - 0xfd
    "10000001", --  158 - 0x9e  :  129 - 0x81
    "11111111", --  159 - 0x9f  :  255 - 0xff
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Sprite 0x14
    "00000111", --  161 - 0xa1  :    7 - 0x7
    "00000010", --  162 - 0xa2  :    2 - 0x2
    "00000100", --  163 - 0xa3  :    4 - 0x4
    "00000011", --  164 - 0xa4  :    3 - 0x3
    "00000011", --  165 - 0xa5  :    3 - 0x3
    "00001101", --  166 - 0xa6  :   13 - 0xd
    "00010111", --  167 - 0xa7  :   23 - 0x17
    "00101111", --  168 - 0xa8  :   47 - 0x2f -- Sprite 0x15
    "01001111", --  169 - 0xa9  :   79 - 0x4f
    "01001111", --  170 - 0xaa  :   79 - 0x4f
    "01001111", --  171 - 0xab  :   79 - 0x4f
    "01001111", --  172 - 0xac  :   79 - 0x4f
    "00100111", --  173 - 0xad  :   39 - 0x27
    "00010000", --  174 - 0xae  :   16 - 0x10
    "00001111", --  175 - 0xaf  :   15 - 0xf
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0x16
    "11100000", --  177 - 0xb1  :  224 - 0xe0
    "10100000", --  178 - 0xb2  :  160 - 0xa0
    "00100000", --  179 - 0xb3  :   32 - 0x20
    "11000000", --  180 - 0xb4  :  192 - 0xc0
    "01000000", --  181 - 0xb5  :   64 - 0x40
    "00110000", --  182 - 0xb6  :   48 - 0x30
    "11101000", --  183 - 0xb7  :  232 - 0xe8
    "11110100", --  184 - 0xb8  :  244 - 0xf4 -- Sprite 0x17
    "11110010", --  185 - 0xb9  :  242 - 0xf2
    "11110010", --  186 - 0xba  :  242 - 0xf2
    "11110010", --  187 - 0xbb  :  242 - 0xf2
    "11110010", --  188 - 0xbc  :  242 - 0xf2
    "11100100", --  189 - 0xbd  :  228 - 0xe4
    "00001000", --  190 - 0xbe  :    8 - 0x8
    "11110000", --  191 - 0xbf  :  240 - 0xf0
    "00111111", --  192 - 0xc0  :   63 - 0x3f -- Sprite 0x18
    "01000000", --  193 - 0xc1  :   64 - 0x40
    "01000000", --  194 - 0xc2  :   64 - 0x40
    "10000000", --  195 - 0xc3  :  128 - 0x80
    "10000000", --  196 - 0xc4  :  128 - 0x80
    "01111111", --  197 - 0xc5  :  127 - 0x7f
    "00000001", --  198 - 0xc6  :    1 - 0x1
    "01111111", --  199 - 0xc7  :  127 - 0x7f
    "11111100", --  200 - 0xc8  :  252 - 0xfc -- Sprite 0x19
    "00000010", --  201 - 0xc9  :    2 - 0x2
    "00000010", --  202 - 0xca  :    2 - 0x2
    "00000001", --  203 - 0xcb  :    1 - 0x1
    "00000001", --  204 - 0xcc  :    1 - 0x1
    "11111110", --  205 - 0xcd  :  254 - 0xfe
    "10000000", --  206 - 0xce  :  128 - 0x80
    "11111110", --  207 - 0xcf  :  254 - 0xfe
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Sprite 0x1a
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00111111", --  210 - 0xd2  :   63 - 0x3f
    "01000000", --  211 - 0xd3  :   64 - 0x40
    "01000000", --  212 - 0xd4  :   64 - 0x40
    "10000000", --  213 - 0xd5  :  128 - 0x80
    "10000000", --  214 - 0xd6  :  128 - 0x80
    "01111111", --  215 - 0xd7  :  127 - 0x7f
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Sprite 0x1b
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "11111100", --  218 - 0xda  :  252 - 0xfc
    "00000010", --  219 - 0xdb  :    2 - 0x2
    "00000010", --  220 - 0xdc  :    2 - 0x2
    "00000001", --  221 - 0xdd  :    1 - 0x1
    "00000001", --  222 - 0xde  :    1 - 0x1
    "11111110", --  223 - 0xdf  :  254 - 0xfe
    "01111111", --  224 - 0xe0  :  127 - 0x7f -- Sprite 0x1c
    "10000000", --  225 - 0xe1  :  128 - 0x80
    "10000000", --  226 - 0xe2  :  128 - 0x80
    "10000000", --  227 - 0xe3  :  128 - 0x80
    "10011011", --  228 - 0xe4  :  155 - 0x9b
    "10100100", --  229 - 0xe5  :  164 - 0xa4
    "10100110", --  230 - 0xe6  :  166 - 0xa6
    "10000000", --  231 - 0xe7  :  128 - 0x80
    "10000000", --  232 - 0xe8  :  128 - 0x80 -- Sprite 0x1d
    "01111111", --  233 - 0xe9  :  127 - 0x7f
    "00000010", --  234 - 0xea  :    2 - 0x2
    "00000010", --  235 - 0xeb  :    2 - 0x2
    "00000010", --  236 - 0xec  :    2 - 0x2
    "00000010", --  237 - 0xed  :    2 - 0x2
    "00000010", --  238 - 0xee  :    2 - 0x2
    "00001111", --  239 - 0xef  :   15 - 0xf
    "11111110", --  240 - 0xf0  :  254 - 0xfe -- Sprite 0x1e
    "00000001", --  241 - 0xf1  :    1 - 0x1
    "00000001", --  242 - 0xf2  :    1 - 0x1
    "00000001", --  243 - 0xf3  :    1 - 0x1
    "01000001", --  244 - 0xf4  :   65 - 0x41
    "11110101", --  245 - 0xf5  :  245 - 0xf5
    "00011101", --  246 - 0xf6  :   29 - 0x1d
    "00000001", --  247 - 0xf7  :    1 - 0x1
    "00000001", --  248 - 0xf8  :    1 - 0x1 -- Sprite 0x1f
    "11111110", --  249 - 0xf9  :  254 - 0xfe
    "01000000", --  250 - 0xfa  :   64 - 0x40
    "01000000", --  251 - 0xfb  :   64 - 0x40
    "01000000", --  252 - 0xfc  :   64 - 0x40
    "01000000", --  253 - 0xfd  :   64 - 0x40
    "01000000", --  254 - 0xfe  :   64 - 0x40
    "11110000", --  255 - 0xff  :  240 - 0xf0
    "00000111", --  256 - 0x100  :    7 - 0x7 -- Sprite 0x20
    "00011111", --  257 - 0x101  :   31 - 0x1f
    "00111111", --  258 - 0x102  :   63 - 0x3f
    "01111111", --  259 - 0x103  :  127 - 0x7f
    "01111111", --  260 - 0x104  :  127 - 0x7f
    "11111111", --  261 - 0x105  :  255 - 0xff
    "11111111", --  262 - 0x106  :  255 - 0xff
    "11111111", --  263 - 0x107  :  255 - 0xff
    "11100000", --  264 - 0x108  :  224 - 0xe0 -- Sprite 0x21
    "11111000", --  265 - 0x109  :  248 - 0xf8
    "11111100", --  266 - 0x10a  :  252 - 0xfc
    "11111110", --  267 - 0x10b  :  254 - 0xfe
    "11111110", --  268 - 0x10c  :  254 - 0xfe
    "11111111", --  269 - 0x10d  :  255 - 0xff
    "11111111", --  270 - 0x10e  :  255 - 0xff
    "11111111", --  271 - 0x10f  :  255 - 0xff
    "00000111", --  272 - 0x110  :    7 - 0x7 -- Sprite 0x22
    "00011111", --  273 - 0x111  :   31 - 0x1f
    "00111111", --  274 - 0x112  :   63 - 0x3f
    "01111111", --  275 - 0x113  :  127 - 0x7f
    "01111111", --  276 - 0x114  :  127 - 0x7f
    "11111111", --  277 - 0x115  :  255 - 0xff
    "11111111", --  278 - 0x116  :  255 - 0xff
    "11111111", --  279 - 0x117  :  255 - 0xff
    "11100000", --  280 - 0x118  :  224 - 0xe0 -- Sprite 0x23
    "11111000", --  281 - 0x119  :  248 - 0xf8
    "11111100", --  282 - 0x11a  :  252 - 0xfc
    "11111110", --  283 - 0x11b  :  254 - 0xfe
    "11111110", --  284 - 0x11c  :  254 - 0xfe
    "11111111", --  285 - 0x11d  :  255 - 0xff
    "11111111", --  286 - 0x11e  :  255 - 0xff
    "11111111", --  287 - 0x11f  :  255 - 0xff
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Sprite 0x24
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00101111", --  296 - 0x128  :   47 - 0x2f -- Sprite 0x25
    "01001111", --  297 - 0x129  :   79 - 0x4f
    "01001111", --  298 - 0x12a  :   79 - 0x4f
    "01001111", --  299 - 0x12b  :   79 - 0x4f
    "01001111", --  300 - 0x12c  :   79 - 0x4f
    "00100111", --  301 - 0x12d  :   39 - 0x27
    "00010000", --  302 - 0x12e  :   16 - 0x10
    "00001111", --  303 - 0x12f  :   15 - 0xf
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x26
    "11100000", --  305 - 0x131  :  224 - 0xe0
    "10100000", --  306 - 0x132  :  160 - 0xa0
    "00100000", --  307 - 0x133  :   32 - 0x20
    "11000000", --  308 - 0x134  :  192 - 0xc0
    "01000000", --  309 - 0x135  :   64 - 0x40
    "00110000", --  310 - 0x136  :   48 - 0x30
    "11101000", --  311 - 0x137  :  232 - 0xe8
    "11110100", --  312 - 0x138  :  244 - 0xf4 -- Sprite 0x27
    "11110010", --  313 - 0x139  :  242 - 0xf2
    "11110010", --  314 - 0x13a  :  242 - 0xf2
    "11110010", --  315 - 0x13b  :  242 - 0xf2
    "11110010", --  316 - 0x13c  :  242 - 0xf2
    "11100100", --  317 - 0x13d  :  228 - 0xe4
    "00001000", --  318 - 0x13e  :    8 - 0x8
    "11110000", --  319 - 0x13f  :  240 - 0xf0
    "11111111", --  320 - 0x140  :  255 - 0xff -- Sprite 0x28
    "11010101", --  321 - 0x141  :  213 - 0xd5
    "10100011", --  322 - 0x142  :  163 - 0xa3
    "11010111", --  323 - 0x143  :  215 - 0xd7
    "10001111", --  324 - 0x144  :  143 - 0x8f
    "11001111", --  325 - 0x145  :  207 - 0xcf
    "10001011", --  326 - 0x146  :  139 - 0x8b
    "11001011", --  327 - 0x147  :  203 - 0xcb
    "10001111", --  328 - 0x148  :  143 - 0x8f -- Sprite 0x29
    "11001111", --  329 - 0x149  :  207 - 0xcf
    "10001111", --  330 - 0x14a  :  143 - 0x8f
    "11001111", --  331 - 0x14b  :  207 - 0xcf
    "10010000", --  332 - 0x14c  :  144 - 0x90
    "11100000", --  333 - 0x14d  :  224 - 0xe0
    "11101010", --  334 - 0x14e  :  234 - 0xea
    "11111111", --  335 - 0x14f  :  255 - 0xff
    "11111111", --  336 - 0x150  :  255 - 0xff -- Sprite 0x2a
    "11011011", --  337 - 0x151  :  219 - 0xdb
    "11000111", --  338 - 0x152  :  199 - 0xc7
    "11101001", --  339 - 0x153  :  233 - 0xe9
    "11110011", --  340 - 0x154  :  243 - 0xf3
    "11110001", --  341 - 0x155  :  241 - 0xf1
    "11010011", --  342 - 0x156  :  211 - 0xd3
    "11010001", --  343 - 0x157  :  209 - 0xd1
    "11110011", --  344 - 0x158  :  243 - 0xf3 -- Sprite 0x2b
    "11110001", --  345 - 0x159  :  241 - 0xf1
    "11110011", --  346 - 0x15a  :  243 - 0xf3
    "11110001", --  347 - 0x15b  :  241 - 0xf1
    "00001011", --  348 - 0x15c  :   11 - 0xb
    "00000101", --  349 - 0x15d  :    5 - 0x5
    "10101011", --  350 - 0x15e  :  171 - 0xab
    "11111111", --  351 - 0x15f  :  255 - 0xff
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00101111", --  360 - 0x168  :   47 - 0x2f -- Sprite 0x2d
    "01001111", --  361 - 0x169  :   79 - 0x4f
    "01001111", --  362 - 0x16a  :   79 - 0x4f
    "01001111", --  363 - 0x16b  :   79 - 0x4f
    "01001111", --  364 - 0x16c  :   79 - 0x4f
    "00100111", --  365 - 0x16d  :   39 - 0x27
    "00010000", --  366 - 0x16e  :   16 - 0x10
    "00001111", --  367 - 0x16f  :   15 - 0xf
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "11110100", --  376 - 0x178  :  244 - 0xf4 -- Sprite 0x2f
    "11110010", --  377 - 0x179  :  242 - 0xf2
    "11110010", --  378 - 0x17a  :  242 - 0xf2
    "11110010", --  379 - 0x17b  :  242 - 0xf2
    "11110010", --  380 - 0x17c  :  242 - 0xf2
    "11100100", --  381 - 0x17d  :  228 - 0xe4
    "00001000", --  382 - 0x17e  :    8 - 0x8
    "11110000", --  383 - 0x17f  :  240 - 0xf0
    "00011000", --  384 - 0x180  :   24 - 0x18 -- Sprite 0x30
    "00100100", --  385 - 0x181  :   36 - 0x24
    "01000010", --  386 - 0x182  :   66 - 0x42
    "10100101", --  387 - 0x183  :  165 - 0xa5
    "11100111", --  388 - 0x184  :  231 - 0xe7
    "00100100", --  389 - 0x185  :   36 - 0x24
    "00100100", --  390 - 0x186  :   36 - 0x24
    "00111100", --  391 - 0x187  :   60 - 0x3c
    "00111100", --  392 - 0x188  :   60 - 0x3c -- Sprite 0x31
    "00100100", --  393 - 0x189  :   36 - 0x24
    "00100100", --  394 - 0x18a  :   36 - 0x24
    "01100110", --  395 - 0x18b  :  102 - 0x66
    "10100101", --  396 - 0x18c  :  165 - 0xa5
    "01000010", --  397 - 0x18d  :   66 - 0x42
    "00100100", --  398 - 0x18e  :   36 - 0x24
    "00011000", --  399 - 0x18f  :   24 - 0x18
    "00000010", --  400 - 0x190  :    2 - 0x2 -- Sprite 0x32
    "00000010", --  401 - 0x191  :    2 - 0x2
    "00000011", --  402 - 0x192  :    3 - 0x3
    "00000010", --  403 - 0x193  :    2 - 0x2
    "00000010", --  404 - 0x194  :    2 - 0x2
    "00000010", --  405 - 0x195  :    2 - 0x2
    "00000011", --  406 - 0x196  :    3 - 0x3
    "00000010", --  407 - 0x197  :    2 - 0x2
    "01000000", --  408 - 0x198  :   64 - 0x40 -- Sprite 0x33
    "11000000", --  409 - 0x199  :  192 - 0xc0
    "01000000", --  410 - 0x19a  :   64 - 0x40
    "01000000", --  411 - 0x19b  :   64 - 0x40
    "01000000", --  412 - 0x19c  :   64 - 0x40
    "11000000", --  413 - 0x19d  :  192 - 0xc0
    "01000000", --  414 - 0x19e  :   64 - 0x40
    "01000000", --  415 - 0x19f  :   64 - 0x40
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- Sprite 0x34
    "00011000", --  417 - 0x1a1  :   24 - 0x18
    "00111100", --  418 - 0x1a2  :   60 - 0x3c
    "01100010", --  419 - 0x1a3  :   98 - 0x62
    "01100001", --  420 - 0x1a4  :   97 - 0x61
    "11000000", --  421 - 0x1a5  :  192 - 0xc0
    "11000000", --  422 - 0x1a6  :  192 - 0xc0
    "11000000", --  423 - 0x1a7  :  192 - 0xc0
    "01100000", --  424 - 0x1a8  :   96 - 0x60 -- Sprite 0x35
    "01100000", --  425 - 0x1a9  :   96 - 0x60
    "00110000", --  426 - 0x1aa  :   48 - 0x30
    "00011000", --  427 - 0x1ab  :   24 - 0x18
    "00001100", --  428 - 0x1ac  :   12 - 0xc
    "00000110", --  429 - 0x1ad  :    6 - 0x6
    "00000010", --  430 - 0x1ae  :    2 - 0x2
    "00000001", --  431 - 0x1af  :    1 - 0x1
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x36
    "00011000", --  433 - 0x1b1  :   24 - 0x18
    "00100100", --  434 - 0x1b2  :   36 - 0x24
    "01000010", --  435 - 0x1b3  :   66 - 0x42
    "10000010", --  436 - 0x1b4  :  130 - 0x82
    "00000001", --  437 - 0x1b5  :    1 - 0x1
    "00000001", --  438 - 0x1b6  :    1 - 0x1
    "00000001", --  439 - 0x1b7  :    1 - 0x1
    "00000010", --  440 - 0x1b8  :    2 - 0x2 -- Sprite 0x37
    "00000010", --  441 - 0x1b9  :    2 - 0x2
    "00000100", --  442 - 0x1ba  :    4 - 0x4
    "00001000", --  443 - 0x1bb  :    8 - 0x8
    "00010000", --  444 - 0x1bc  :   16 - 0x10
    "00100000", --  445 - 0x1bd  :   32 - 0x20
    "01000000", --  446 - 0x1be  :   64 - 0x40
    "10000000", --  447 - 0x1bf  :  128 - 0x80
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Sprite 0x38
    "00000110", --  449 - 0x1c1  :    6 - 0x6
    "00001101", --  450 - 0x1c2  :   13 - 0xd
    "00001100", --  451 - 0x1c3  :   12 - 0xc
    "00001100", --  452 - 0x1c4  :   12 - 0xc
    "00000110", --  453 - 0x1c5  :    6 - 0x6
    "00000010", --  454 - 0x1c6  :    2 - 0x2
    "00000001", --  455 - 0x1c7  :    1 - 0x1
    "11111111", --  456 - 0x1c8  :  255 - 0xff -- Sprite 0x39
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x3a
    "01100000", --  465 - 0x1d1  :   96 - 0x60
    "10010000", --  466 - 0x1d2  :  144 - 0x90
    "00010000", --  467 - 0x1d3  :   16 - 0x10
    "00010000", --  468 - 0x1d4  :   16 - 0x10
    "00100000", --  469 - 0x1d5  :   32 - 0x20
    "01000000", --  470 - 0x1d6  :   64 - 0x40
    "10000000", --  471 - 0x1d7  :  128 - 0x80
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Sprite 0x3b
    "01010100", --  473 - 0x1d9  :   84 - 0x54
    "00000010", --  474 - 0x1da  :    2 - 0x2
    "01000000", --  475 - 0x1db  :   64 - 0x40
    "00000010", --  476 - 0x1dc  :    2 - 0x2
    "01000000", --  477 - 0x1dd  :   64 - 0x40
    "00101010", --  478 - 0x1de  :   42 - 0x2a
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "11111111", --  480 - 0x1e0  :  255 - 0xff -- Sprite 0x3c
    "11111111", --  481 - 0x1e1  :  255 - 0xff
    "11111111", --  482 - 0x1e2  :  255 - 0xff
    "11111111", --  483 - 0x1e3  :  255 - 0xff
    "11111111", --  484 - 0x1e4  :  255 - 0xff
    "11111111", --  485 - 0x1e5  :  255 - 0xff
    "11111111", --  486 - 0x1e6  :  255 - 0xff
    "11111111", --  487 - 0x1e7  :  255 - 0xff
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Sprite 0x3d
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "11111111", --  496 - 0x1f0  :  255 - 0xff -- Sprite 0x3e
    "11111111", --  497 - 0x1f1  :  255 - 0xff
    "11111111", --  498 - 0x1f2  :  255 - 0xff
    "11111111", --  499 - 0x1f3  :  255 - 0xff
    "11111111", --  500 - 0x1f4  :  255 - 0xff
    "11111111", --  501 - 0x1f5  :  255 - 0xff
    "11111111", --  502 - 0x1f6  :  255 - 0xff
    "11111111", --  503 - 0x1f7  :  255 - 0xff
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- Sprite 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00111100", --  512 - 0x200  :   60 - 0x3c -- Sprite 0x40
    "01000010", --  513 - 0x201  :   66 - 0x42
    "10011001", --  514 - 0x202  :  153 - 0x99
    "10100101", --  515 - 0x203  :  165 - 0xa5
    "10100101", --  516 - 0x204  :  165 - 0xa5
    "10011010", --  517 - 0x205  :  154 - 0x9a
    "01000000", --  518 - 0x206  :   64 - 0x40
    "00111100", --  519 - 0x207  :   60 - 0x3c
    "00001100", --  520 - 0x208  :   12 - 0xc -- Sprite 0x41
    "00010010", --  521 - 0x209  :   18 - 0x12
    "00100010", --  522 - 0x20a  :   34 - 0x22
    "00100010", --  523 - 0x20b  :   34 - 0x22
    "01111110", --  524 - 0x20c  :  126 - 0x7e
    "00100010", --  525 - 0x20d  :   34 - 0x22
    "00100100", --  526 - 0x20e  :   36 - 0x24
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00111100", --  528 - 0x210  :   60 - 0x3c -- Sprite 0x42
    "01000010", --  529 - 0x211  :   66 - 0x42
    "01010010", --  530 - 0x212  :   82 - 0x52
    "00011100", --  531 - 0x213  :   28 - 0x1c
    "00010010", --  532 - 0x214  :   18 - 0x12
    "00110010", --  533 - 0x215  :   50 - 0x32
    "00011100", --  534 - 0x216  :   28 - 0x1c
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00011000", --  536 - 0x218  :   24 - 0x18 -- Sprite 0x43
    "00100100", --  537 - 0x219  :   36 - 0x24
    "01010100", --  538 - 0x21a  :   84 - 0x54
    "01001000", --  539 - 0x21b  :   72 - 0x48
    "01000010", --  540 - 0x21c  :   66 - 0x42
    "00100100", --  541 - 0x21d  :   36 - 0x24
    "00011000", --  542 - 0x21e  :   24 - 0x18
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "01011000", --  544 - 0x220  :   88 - 0x58 -- Sprite 0x44
    "11100100", --  545 - 0x221  :  228 - 0xe4
    "01000010", --  546 - 0x222  :   66 - 0x42
    "01000010", --  547 - 0x223  :   66 - 0x42
    "00100010", --  548 - 0x224  :   34 - 0x22
    "01100100", --  549 - 0x225  :  100 - 0x64
    "00111000", --  550 - 0x226  :   56 - 0x38
    "00000000", --  551 - 0x227  :    0 - 0x0
    "00011100", --  552 - 0x228  :   28 - 0x1c -- Sprite 0x45
    "00100000", --  553 - 0x229  :   32 - 0x20
    "00100000", --  554 - 0x22a  :   32 - 0x20
    "00101100", --  555 - 0x22b  :   44 - 0x2c
    "01110000", --  556 - 0x22c  :  112 - 0x70
    "00100010", --  557 - 0x22d  :   34 - 0x22
    "00011100", --  558 - 0x22e  :   28 - 0x1c
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00011100", --  560 - 0x230  :   28 - 0x1c -- Sprite 0x46
    "00100000", --  561 - 0x231  :   32 - 0x20
    "00100000", --  562 - 0x232  :   32 - 0x20
    "00101100", --  563 - 0x233  :   44 - 0x2c
    "01110000", --  564 - 0x234  :  112 - 0x70
    "00010000", --  565 - 0x235  :   16 - 0x10
    "00010000", --  566 - 0x236  :   16 - 0x10
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00011000", --  568 - 0x238  :   24 - 0x18 -- Sprite 0x47
    "00100100", --  569 - 0x239  :   36 - 0x24
    "01000000", --  570 - 0x23a  :   64 - 0x40
    "01001110", --  571 - 0x23b  :   78 - 0x4e
    "01000010", --  572 - 0x23c  :   66 - 0x42
    "00100100", --  573 - 0x23d  :   36 - 0x24
    "00011000", --  574 - 0x23e  :   24 - 0x18
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00100000", --  576 - 0x240  :   32 - 0x20 -- Sprite 0x48
    "01000100", --  577 - 0x241  :   68 - 0x44
    "01000100", --  578 - 0x242  :   68 - 0x44
    "01000100", --  579 - 0x243  :   68 - 0x44
    "11111100", --  580 - 0x244  :  252 - 0xfc
    "01000100", --  581 - 0x245  :   68 - 0x44
    "01001000", --  582 - 0x246  :   72 - 0x48
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00010000", --  584 - 0x248  :   16 - 0x10 -- Sprite 0x49
    "00010000", --  585 - 0x249  :   16 - 0x10
    "00010000", --  586 - 0x24a  :   16 - 0x10
    "00010000", --  587 - 0x24b  :   16 - 0x10
    "00010000", --  588 - 0x24c  :   16 - 0x10
    "00001000", --  589 - 0x24d  :    8 - 0x8
    "00001000", --  590 - 0x24e  :    8 - 0x8
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00001000", --  592 - 0x250  :    8 - 0x8 -- Sprite 0x4a
    "00001000", --  593 - 0x251  :    8 - 0x8
    "00000100", --  594 - 0x252  :    4 - 0x4
    "00000100", --  595 - 0x253  :    4 - 0x4
    "01000100", --  596 - 0x254  :   68 - 0x44
    "01001000", --  597 - 0x255  :   72 - 0x48
    "00110000", --  598 - 0x256  :   48 - 0x30
    "00000000", --  599 - 0x257  :    0 - 0x0
    "01000100", --  600 - 0x258  :   68 - 0x44 -- Sprite 0x4b
    "01000100", --  601 - 0x259  :   68 - 0x44
    "01001000", --  602 - 0x25a  :   72 - 0x48
    "01110000", --  603 - 0x25b  :  112 - 0x70
    "01001000", --  604 - 0x25c  :   72 - 0x48
    "00100100", --  605 - 0x25d  :   36 - 0x24
    "00100010", --  606 - 0x25e  :   34 - 0x22
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00010000", --  608 - 0x260  :   16 - 0x10 -- Sprite 0x4c
    "00100000", --  609 - 0x261  :   32 - 0x20
    "00100000", --  610 - 0x262  :   32 - 0x20
    "00100000", --  611 - 0x263  :   32 - 0x20
    "01000000", --  612 - 0x264  :   64 - 0x40
    "01000000", --  613 - 0x265  :   64 - 0x40
    "01000110", --  614 - 0x266  :   70 - 0x46
    "00111000", --  615 - 0x267  :   56 - 0x38
    "00100100", --  616 - 0x268  :   36 - 0x24 -- Sprite 0x4d
    "01011010", --  617 - 0x269  :   90 - 0x5a
    "01011010", --  618 - 0x26a  :   90 - 0x5a
    "01011010", --  619 - 0x26b  :   90 - 0x5a
    "01000010", --  620 - 0x26c  :   66 - 0x42
    "01000010", --  621 - 0x26d  :   66 - 0x42
    "00100010", --  622 - 0x26e  :   34 - 0x22
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00100100", --  624 - 0x270  :   36 - 0x24 -- Sprite 0x4e
    "01010010", --  625 - 0x271  :   82 - 0x52
    "01010010", --  626 - 0x272  :   82 - 0x52
    "01010010", --  627 - 0x273  :   82 - 0x52
    "01010010", --  628 - 0x274  :   82 - 0x52
    "01010010", --  629 - 0x275  :   82 - 0x52
    "01001100", --  630 - 0x276  :   76 - 0x4c
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00111000", --  632 - 0x278  :   56 - 0x38 -- Sprite 0x4f
    "01000100", --  633 - 0x279  :   68 - 0x44
    "10000010", --  634 - 0x27a  :  130 - 0x82
    "10000010", --  635 - 0x27b  :  130 - 0x82
    "10000010", --  636 - 0x27c  :  130 - 0x82
    "01000100", --  637 - 0x27d  :   68 - 0x44
    "00111000", --  638 - 0x27e  :   56 - 0x38
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "01111111", --  640 - 0x280  :  127 - 0x7f -- Sprite 0x50
    "11000000", --  641 - 0x281  :  192 - 0xc0
    "10000000", --  642 - 0x282  :  128 - 0x80
    "10000000", --  643 - 0x283  :  128 - 0x80
    "10000000", --  644 - 0x284  :  128 - 0x80
    "11000011", --  645 - 0x285  :  195 - 0xc3
    "11111111", --  646 - 0x286  :  255 - 0xff
    "11111111", --  647 - 0x287  :  255 - 0xff
    "11111110", --  648 - 0x288  :  254 - 0xfe -- Sprite 0x51
    "00000011", --  649 - 0x289  :    3 - 0x3
    "00000001", --  650 - 0x28a  :    1 - 0x1
    "00000001", --  651 - 0x28b  :    1 - 0x1
    "00000001", --  652 - 0x28c  :    1 - 0x1
    "11000011", --  653 - 0x28d  :  195 - 0xc3
    "11111111", --  654 - 0x28e  :  255 - 0xff
    "11111111", --  655 - 0x28f  :  255 - 0xff
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Sprite 0x52
    "00000111", --  657 - 0x291  :    7 - 0x7
    "00001100", --  658 - 0x292  :   12 - 0xc
    "00011000", --  659 - 0x293  :   24 - 0x18
    "00110000", --  660 - 0x294  :   48 - 0x30
    "01100000", --  661 - 0x295  :   96 - 0x60
    "01000000", --  662 - 0x296  :   64 - 0x40
    "01001111", --  663 - 0x297  :   79 - 0x4f
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Sprite 0x53
    "11110000", --  665 - 0x299  :  240 - 0xf0
    "01010000", --  666 - 0x29a  :   80 - 0x50
    "01001000", --  667 - 0x29b  :   72 - 0x48
    "01001100", --  668 - 0x29c  :   76 - 0x4c
    "01000100", --  669 - 0x29d  :   68 - 0x44
    "10000010", --  670 - 0x29e  :  130 - 0x82
    "10000011", --  671 - 0x29f  :  131 - 0x83
    "01111111", --  672 - 0x2a0  :  127 - 0x7f -- Sprite 0x54
    "11011110", --  673 - 0x2a1  :  222 - 0xde
    "10001110", --  674 - 0x2a2  :  142 - 0x8e
    "11000101", --  675 - 0x2a3  :  197 - 0xc5
    "10010010", --  676 - 0x2a4  :  146 - 0x92
    "11000111", --  677 - 0x2a5  :  199 - 0xc7
    "11100010", --  678 - 0x2a6  :  226 - 0xe2
    "11010000", --  679 - 0x2a7  :  208 - 0xd0
    "11111111", --  680 - 0x2a8  :  255 - 0xff -- Sprite 0x55
    "11011110", --  681 - 0x2a9  :  222 - 0xde
    "10001110", --  682 - 0x2aa  :  142 - 0x8e
    "11000101", --  683 - 0x2ab  :  197 - 0xc5
    "10010010", --  684 - 0x2ac  :  146 - 0x92
    "01000111", --  685 - 0x2ad  :   71 - 0x47
    "11100010", --  686 - 0x2ae  :  226 - 0xe2
    "01010000", --  687 - 0x2af  :   80 - 0x50
    "11111110", --  688 - 0x2b0  :  254 - 0xfe -- Sprite 0x56
    "11011111", --  689 - 0x2b1  :  223 - 0xdf
    "10001111", --  690 - 0x2b2  :  143 - 0x8f
    "11000101", --  691 - 0x2b3  :  197 - 0xc5
    "10010011", --  692 - 0x2b4  :  147 - 0x93
    "01000111", --  693 - 0x2b5  :   71 - 0x47
    "11100011", --  694 - 0x2b6  :  227 - 0xe3
    "01010001", --  695 - 0x2b7  :   81 - 0x51
    "01111111", --  696 - 0x2b8  :  127 - 0x7f -- Sprite 0x57
    "10000000", --  697 - 0x2b9  :  128 - 0x80
    "10110011", --  698 - 0x2ba  :  179 - 0xb3
    "01001100", --  699 - 0x2bb  :   76 - 0x4c
    "00111111", --  700 - 0x2bc  :   63 - 0x3f
    "00000011", --  701 - 0x2bd  :    3 - 0x3
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "11111111", --  704 - 0x2c0  :  255 - 0xff -- Sprite 0x58
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00110011", --  706 - 0x2c2  :   51 - 0x33
    "11001100", --  707 - 0x2c3  :  204 - 0xcc
    "00110011", --  708 - 0x2c4  :   51 - 0x33
    "11111111", --  709 - 0x2c5  :  255 - 0xff
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "11111110", --  712 - 0x2c8  :  254 - 0xfe -- Sprite 0x59
    "00000001", --  713 - 0x2c9  :    1 - 0x1
    "00110011", --  714 - 0x2ca  :   51 - 0x33
    "11001110", --  715 - 0x2cb  :  206 - 0xce
    "00111100", --  716 - 0x2cc  :   60 - 0x3c
    "11000000", --  717 - 0x2cd  :  192 - 0xc0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x5a
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Sprite 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000001", --  731 - 0x2db  :    1 - 0x1
    "00000011", --  732 - 0x2dc  :    3 - 0x3
    "00000011", --  733 - 0x2dd  :    3 - 0x3
    "00000111", --  734 - 0x2de  :    7 - 0x7
    "00111111", --  735 - 0x2df  :   63 - 0x3f
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Sprite 0x5c
    "00000001", --  737 - 0x2e1  :    1 - 0x1
    "01111111", --  738 - 0x2e2  :  127 - 0x7f
    "11111111", --  739 - 0x2e3  :  255 - 0xff
    "11111111", --  740 - 0x2e4  :  255 - 0xff
    "11111111", --  741 - 0x2e5  :  255 - 0xff
    "11111111", --  742 - 0x2e6  :  255 - 0xff
    "11111111", --  743 - 0x2e7  :  255 - 0xff
    "11111111", --  744 - 0x2e8  :  255 - 0xff -- Sprite 0x5d
    "11111111", --  745 - 0x2e9  :  255 - 0xff
    "11111111", --  746 - 0x2ea  :  255 - 0xff
    "11111111", --  747 - 0x2eb  :  255 - 0xff
    "11111111", --  748 - 0x2ec  :  255 - 0xff
    "11111111", --  749 - 0x2ed  :  255 - 0xff
    "11111111", --  750 - 0x2ee  :  255 - 0xff
    "11111111", --  751 - 0x2ef  :  255 - 0xff
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x5e
    "10000000", --  753 - 0x2f1  :  128 - 0x80
    "11111110", --  754 - 0x2f2  :  254 - 0xfe
    "11111111", --  755 - 0x2f3  :  255 - 0xff
    "11111111", --  756 - 0x2f4  :  255 - 0xff
    "11111111", --  757 - 0x2f5  :  255 - 0xff
    "11111111", --  758 - 0x2f6  :  255 - 0xff
    "11111111", --  759 - 0x2f7  :  255 - 0xff
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- Sprite 0x5f
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "10000000", --  763 - 0x2fb  :  128 - 0x80
    "11000000", --  764 - 0x2fc  :  192 - 0xc0
    "11000000", --  765 - 0x2fd  :  192 - 0xc0
    "11100000", --  766 - 0x2fe  :  224 - 0xe0
    "11111000", --  767 - 0x2ff  :  248 - 0xf8
    "11111111", --  768 - 0x300  :  255 - 0xff -- Sprite 0x60
    "11111111", --  769 - 0x301  :  255 - 0xff
    "11111111", --  770 - 0x302  :  255 - 0xff
    "11111111", --  771 - 0x303  :  255 - 0xff
    "11111111", --  772 - 0x304  :  255 - 0xff
    "11111111", --  773 - 0x305  :  255 - 0xff
    "11111111", --  774 - 0x306  :  255 - 0xff
    "11111111", --  775 - 0x307  :  255 - 0xff
    "11111111", --  776 - 0x308  :  255 - 0xff -- Sprite 0x61
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11111111", --  778 - 0x30a  :  255 - 0xff
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "11111111", --  780 - 0x30c  :  255 - 0xff
    "11111111", --  781 - 0x30d  :  255 - 0xff
    "11111111", --  782 - 0x30e  :  255 - 0xff
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "01111000", --  784 - 0x310  :  120 - 0x78 -- Sprite 0x62
    "01100000", --  785 - 0x311  :   96 - 0x60
    "01000000", --  786 - 0x312  :   64 - 0x40
    "01000000", --  787 - 0x313  :   64 - 0x40
    "01000000", --  788 - 0x314  :   64 - 0x40
    "01100000", --  789 - 0x315  :   96 - 0x60
    "00110000", --  790 - 0x316  :   48 - 0x30
    "00011111", --  791 - 0x317  :   31 - 0x1f
    "10000001", --  792 - 0x318  :  129 - 0x81 -- Sprite 0x63
    "10000011", --  793 - 0x319  :  131 - 0x83
    "11000001", --  794 - 0x31a  :  193 - 0xc1
    "01000011", --  795 - 0x31b  :   67 - 0x43
    "01000001", --  796 - 0x31c  :   65 - 0x41
    "01100011", --  797 - 0x31d  :   99 - 0x63
    "00100110", --  798 - 0x31e  :   38 - 0x26
    "11111000", --  799 - 0x31f  :  248 - 0xf8
    "10111001", --  800 - 0x320  :  185 - 0xb9 -- Sprite 0x64
    "10010100", --  801 - 0x321  :  148 - 0x94
    "10001110", --  802 - 0x322  :  142 - 0x8e
    "11000101", --  803 - 0x323  :  197 - 0xc5
    "10010010", --  804 - 0x324  :  146 - 0x92
    "11000111", --  805 - 0x325  :  199 - 0xc7
    "11100010", --  806 - 0x326  :  226 - 0xe2
    "11010000", --  807 - 0x327  :  208 - 0xd0
    "10111001", --  808 - 0x328  :  185 - 0xb9 -- Sprite 0x65
    "00010100", --  809 - 0x329  :   20 - 0x14
    "10001110", --  810 - 0x32a  :  142 - 0x8e
    "11000101", --  811 - 0x32b  :  197 - 0xc5
    "10010010", --  812 - 0x32c  :  146 - 0x92
    "01000111", --  813 - 0x32d  :   71 - 0x47
    "11100010", --  814 - 0x32e  :  226 - 0xe2
    "01010000", --  815 - 0x32f  :   80 - 0x50
    "10111001", --  816 - 0x330  :  185 - 0xb9 -- Sprite 0x66
    "00010101", --  817 - 0x331  :   21 - 0x15
    "10001111", --  818 - 0x332  :  143 - 0x8f
    "11000101", --  819 - 0x333  :  197 - 0xc5
    "10010011", --  820 - 0x334  :  147 - 0x93
    "01000111", --  821 - 0x335  :   71 - 0x47
    "11100011", --  822 - 0x336  :  227 - 0xe3
    "01010001", --  823 - 0x337  :   81 - 0x51
    "01111111", --  824 - 0x338  :  127 - 0x7f -- Sprite 0x67
    "10000000", --  825 - 0x339  :  128 - 0x80
    "11001100", --  826 - 0x33a  :  204 - 0xcc
    "01111111", --  827 - 0x33b  :  127 - 0x7f
    "00111111", --  828 - 0x33c  :   63 - 0x3f
    "00000011", --  829 - 0x33d  :    3 - 0x3
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "11111111", --  832 - 0x340  :  255 - 0xff -- Sprite 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "11001100", --  834 - 0x342  :  204 - 0xcc
    "00110011", --  835 - 0x343  :   51 - 0x33
    "11111111", --  836 - 0x344  :  255 - 0xff
    "11111111", --  837 - 0x345  :  255 - 0xff
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "11111110", --  840 - 0x348  :  254 - 0xfe -- Sprite 0x69
    "00000001", --  841 - 0x349  :    1 - 0x1
    "11001101", --  842 - 0x34a  :  205 - 0xcd
    "00111110", --  843 - 0x34b  :   62 - 0x3e
    "11111100", --  844 - 0x34c  :  252 - 0xfc
    "11000000", --  845 - 0x34d  :  192 - 0xc0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Sprite 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "01111111", --  856 - 0x358  :  127 - 0x7f -- Sprite 0x6b
    "11111111", --  857 - 0x359  :  255 - 0xff
    "11111111", --  858 - 0x35a  :  255 - 0xff
    "11111111", --  859 - 0x35b  :  255 - 0xff
    "01111111", --  860 - 0x35c  :  127 - 0x7f
    "00110000", --  861 - 0x35d  :   48 - 0x30
    "00001111", --  862 - 0x35e  :   15 - 0xf
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "11111111", --  864 - 0x360  :  255 - 0xff -- Sprite 0x6c
    "11111111", --  865 - 0x361  :  255 - 0xff
    "11111111", --  866 - 0x362  :  255 - 0xff
    "11111111", --  867 - 0x363  :  255 - 0xff
    "11111111", --  868 - 0x364  :  255 - 0xff
    "11111110", --  869 - 0x365  :  254 - 0xfe
    "00000001", --  870 - 0x366  :    1 - 0x1
    "11111110", --  871 - 0x367  :  254 - 0xfe
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Sprite 0x6d
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "11111100", --  888 - 0x378  :  252 - 0xfc -- Sprite 0x6f
    "11111110", --  889 - 0x379  :  254 - 0xfe
    "11111111", --  890 - 0x37a  :  255 - 0xff
    "11111111", --  891 - 0x37b  :  255 - 0xff
    "11110010", --  892 - 0x37c  :  242 - 0xf2
    "00001100", --  893 - 0x37d  :   12 - 0xc
    "11110000", --  894 - 0x37e  :  240 - 0xf0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "01111111", --  896 - 0x380  :  127 - 0x7f -- Sprite 0x70
    "11000000", --  897 - 0x381  :  192 - 0xc0
    "10000000", --  898 - 0x382  :  128 - 0x80
    "10000000", --  899 - 0x383  :  128 - 0x80
    "11100011", --  900 - 0x384  :  227 - 0xe3
    "11111111", --  901 - 0x385  :  255 - 0xff
    "11111111", --  902 - 0x386  :  255 - 0xff
    "11111111", --  903 - 0x387  :  255 - 0xff
    "11111111", --  904 - 0x388  :  255 - 0xff -- Sprite 0x71
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "11000011", --  909 - 0x38d  :  195 - 0xc3
    "11111111", --  910 - 0x38e  :  255 - 0xff
    "11111111", --  911 - 0x38f  :  255 - 0xff
    "11111110", --  912 - 0x390  :  254 - 0xfe -- Sprite 0x72
    "00000011", --  913 - 0x391  :    3 - 0x3
    "00000001", --  914 - 0x392  :    1 - 0x1
    "00000001", --  915 - 0x393  :    1 - 0x1
    "11000111", --  916 - 0x394  :  199 - 0xc7
    "11111111", --  917 - 0x395  :  255 - 0xff
    "11111111", --  918 - 0x396  :  255 - 0xff
    "11111111", --  919 - 0x397  :  255 - 0xff
    "11111111", --  920 - 0x398  :  255 - 0xff -- Sprite 0x73
    "11111111", --  921 - 0x399  :  255 - 0xff
    "11111111", --  922 - 0x39a  :  255 - 0xff
    "11111111", --  923 - 0x39b  :  255 - 0xff
    "11111111", --  924 - 0x39c  :  255 - 0xff
    "11111111", --  925 - 0x39d  :  255 - 0xff
    "11111111", --  926 - 0x39e  :  255 - 0xff
    "11111111", --  927 - 0x39f  :  255 - 0xff
    "10111001", --  928 - 0x3a0  :  185 - 0xb9 -- Sprite 0x74
    "10010100", --  929 - 0x3a1  :  148 - 0x94
    "10001110", --  930 - 0x3a2  :  142 - 0x8e
    "11000101", --  931 - 0x3a3  :  197 - 0xc5
    "10010010", --  932 - 0x3a4  :  146 - 0x92
    "11000111", --  933 - 0x3a5  :  199 - 0xc7
    "11100010", --  934 - 0x3a6  :  226 - 0xe2
    "01111111", --  935 - 0x3a7  :  127 - 0x7f
    "10111001", --  936 - 0x3a8  :  185 - 0xb9 -- Sprite 0x75
    "00010100", --  937 - 0x3a9  :   20 - 0x14
    "10001110", --  938 - 0x3aa  :  142 - 0x8e
    "11000101", --  939 - 0x3ab  :  197 - 0xc5
    "10010010", --  940 - 0x3ac  :  146 - 0x92
    "01000111", --  941 - 0x3ad  :   71 - 0x47
    "11100010", --  942 - 0x3ae  :  226 - 0xe2
    "11111111", --  943 - 0x3af  :  255 - 0xff
    "10111001", --  944 - 0x3b0  :  185 - 0xb9 -- Sprite 0x76
    "00010101", --  945 - 0x3b1  :   21 - 0x15
    "10001111", --  946 - 0x3b2  :  143 - 0x8f
    "11000101", --  947 - 0x3b3  :  197 - 0xc5
    "10010011", --  948 - 0x3b4  :  147 - 0x93
    "01000111", --  949 - 0x3b5  :   71 - 0x47
    "11100011", --  950 - 0x3b6  :  227 - 0xe3
    "11111110", --  951 - 0x3b7  :  254 - 0xfe
    "11111111", --  952 - 0x3b8  :  255 - 0xff -- Sprite 0x77
    "11111111", --  953 - 0x3b9  :  255 - 0xff
    "11111111", --  954 - 0x3ba  :  255 - 0xff
    "11111111", --  955 - 0x3bb  :  255 - 0xff
    "11111111", --  956 - 0x3bc  :  255 - 0xff
    "11111111", --  957 - 0x3bd  :  255 - 0xff
    "11111111", --  958 - 0x3be  :  255 - 0xff
    "11111111", --  959 - 0x3bf  :  255 - 0xff
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Sprite 0x79
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Sprite 0x7a
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Sprite 0x7b
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00100010", --  992 - 0x3e0  :   34 - 0x22 -- Sprite 0x7c
    "01010101", --  993 - 0x3e1  :   85 - 0x55
    "10101010", --  994 - 0x3e2  :  170 - 0xaa
    "00000101", --  995 - 0x3e3  :    5 - 0x5
    "00000100", --  996 - 0x3e4  :    4 - 0x4
    "00001010", --  997 - 0x3e5  :   10 - 0xa
    "01010000", --  998 - 0x3e6  :   80 - 0x50
    "00000010", --  999 - 0x3e7  :    2 - 0x2
    "01110011", -- 1000 - 0x3e8  :  115 - 0x73 -- Sprite 0x7d
    "11111111", -- 1001 - 0x3e9  :  255 - 0xff
    "11111111", -- 1002 - 0x3ea  :  255 - 0xff
    "10111101", -- 1003 - 0x3eb  :  189 - 0xbd
    "01101110", -- 1004 - 0x3ec  :  110 - 0x6e
    "00001010", -- 1005 - 0x3ed  :   10 - 0xa
    "01010000", -- 1006 - 0x3ee  :   80 - 0x50
    "00000010", -- 1007 - 0x3ef  :    2 - 0x2
    "00100000", -- 1008 - 0x3f0  :   32 - 0x20 -- Sprite 0x7e
    "01010000", -- 1009 - 0x3f1  :   80 - 0x50
    "10000100", -- 1010 - 0x3f2  :  132 - 0x84
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00100100", -- 1012 - 0x3f4  :   36 - 0x24
    "01011010", -- 1013 - 0x3f5  :   90 - 0x5a
    "00010000", -- 1014 - 0x3f6  :   16 - 0x10
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "11111111", -- 1016 - 0x3f8  :  255 - 0xff -- Sprite 0x7f
    "01010000", -- 1017 - 0x3f9  :   80 - 0x50
    "10000100", -- 1018 - 0x3fa  :  132 - 0x84
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00100100", -- 1020 - 0x3fc  :   36 - 0x24
    "01011010", -- 1021 - 0x3fd  :   90 - 0x5a
    "00010000", -- 1022 - 0x3fe  :   16 - 0x10
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "11111111", -- 1024 - 0x400  :  255 - 0xff -- Sprite 0x80
    "10000000", -- 1025 - 0x401  :  128 - 0x80
    "11001111", -- 1026 - 0x402  :  207 - 0xcf
    "01001000", -- 1027 - 0x403  :   72 - 0x48
    "11001111", -- 1028 - 0x404  :  207 - 0xcf
    "10000000", -- 1029 - 0x405  :  128 - 0x80
    "11001111", -- 1030 - 0x406  :  207 - 0xcf
    "01001000", -- 1031 - 0x407  :   72 - 0x48
    "11111111", -- 1032 - 0x408  :  255 - 0xff -- Sprite 0x81
    "10000000", -- 1033 - 0x409  :  128 - 0x80
    "11111111", -- 1034 - 0x40a  :  255 - 0xff
    "10000000", -- 1035 - 0x40b  :  128 - 0x80
    "10000000", -- 1036 - 0x40c  :  128 - 0x80
    "11011111", -- 1037 - 0x40d  :  223 - 0xdf
    "10110000", -- 1038 - 0x40e  :  176 - 0xb0
    "11000000", -- 1039 - 0x40f  :  192 - 0xc0
    "11111111", -- 1040 - 0x410  :  255 - 0xff -- Sprite 0x82
    "00000001", -- 1041 - 0x411  :    1 - 0x1
    "11110011", -- 1042 - 0x412  :  243 - 0xf3
    "00010010", -- 1043 - 0x413  :   18 - 0x12
    "11110011", -- 1044 - 0x414  :  243 - 0xf3
    "00000001", -- 1045 - 0x415  :    1 - 0x1
    "11110011", -- 1046 - 0x416  :  243 - 0xf3
    "00010010", -- 1047 - 0x417  :   18 - 0x12
    "11111111", -- 1048 - 0x418  :  255 - 0xff -- Sprite 0x83
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "11111111", -- 1050 - 0x41a  :  255 - 0xff
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "11111111", -- 1053 - 0x41d  :  255 - 0xff
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "11111111", -- 1056 - 0x420  :  255 - 0xff -- Sprite 0x84
    "10000010", -- 1057 - 0x421  :  130 - 0x82
    "00010000", -- 1058 - 0x422  :   16 - 0x10
    "00000000", -- 1059 - 0x423  :    0 - 0x0
    "00000000", -- 1060 - 0x424  :    0 - 0x0
    "00010000", -- 1061 - 0x425  :   16 - 0x10
    "01000100", -- 1062 - 0x426  :   68 - 0x44
    "11111111", -- 1063 - 0x427  :  255 - 0xff
    "11111111", -- 1064 - 0x428  :  255 - 0xff -- Sprite 0x85
    "00000001", -- 1065 - 0x429  :    1 - 0x1
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "00000001", -- 1067 - 0x42b  :    1 - 0x1
    "00000001", -- 1068 - 0x42c  :    1 - 0x1
    "11110011", -- 1069 - 0x42d  :  243 - 0xf3
    "00001101", -- 1070 - 0x42e  :   13 - 0xd
    "00000011", -- 1071 - 0x42f  :    3 - 0x3
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Sprite 0x86
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- Sprite 0x87
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000111", -- 1088 - 0x440  :    7 - 0x7 -- Sprite 0x88
    "00011110", -- 1089 - 0x441  :   30 - 0x1e
    "00101111", -- 1090 - 0x442  :   47 - 0x2f
    "01010011", -- 1091 - 0x443  :   83 - 0x53
    "01101110", -- 1092 - 0x444  :  110 - 0x6e
    "11011011", -- 1093 - 0x445  :  219 - 0xdb
    "11111010", -- 1094 - 0x446  :  250 - 0xfa
    "11010101", -- 1095 - 0x447  :  213 - 0xd5
    "10111011", -- 1096 - 0x448  :  187 - 0xbb -- Sprite 0x89
    "11110010", -- 1097 - 0x449  :  242 - 0xf2
    "11011101", -- 1098 - 0x44a  :  221 - 0xdd
    "01001111", -- 1099 - 0x44b  :   79 - 0x4f
    "01111011", -- 1100 - 0x44c  :  123 - 0x7b
    "00110010", -- 1101 - 0x44d  :   50 - 0x32
    "00011111", -- 1102 - 0x44e  :   31 - 0x1f
    "00000111", -- 1103 - 0x44f  :    7 - 0x7
    "11100000", -- 1104 - 0x450  :  224 - 0xe0 -- Sprite 0x8a
    "11011000", -- 1105 - 0x451  :  216 - 0xd8
    "01010100", -- 1106 - 0x452  :   84 - 0x54
    "11101010", -- 1107 - 0x453  :  234 - 0xea
    "10111010", -- 1108 - 0x454  :  186 - 0xba
    "10010011", -- 1109 - 0x455  :  147 - 0x93
    "11011111", -- 1110 - 0x456  :  223 - 0xdf
    "10111101", -- 1111 - 0x457  :  189 - 0xbd
    "01101011", -- 1112 - 0x458  :  107 - 0x6b -- Sprite 0x8b
    "10011111", -- 1113 - 0x459  :  159 - 0x9f
    "01011101", -- 1114 - 0x45a  :   93 - 0x5d
    "10110110", -- 1115 - 0x45b  :  182 - 0xb6
    "11101010", -- 1116 - 0x45c  :  234 - 0xea
    "11001100", -- 1117 - 0x45d  :  204 - 0xcc
    "01111000", -- 1118 - 0x45e  :  120 - 0x78
    "11100000", -- 1119 - 0x45f  :  224 - 0xe0
    "00000111", -- 1120 - 0x460  :    7 - 0x7 -- Sprite 0x8c
    "00011000", -- 1121 - 0x461  :   24 - 0x18
    "00100011", -- 1122 - 0x462  :   35 - 0x23
    "01001100", -- 1123 - 0x463  :   76 - 0x4c
    "01110000", -- 1124 - 0x464  :  112 - 0x70
    "10100001", -- 1125 - 0x465  :  161 - 0xa1
    "10100110", -- 1126 - 0x466  :  166 - 0xa6
    "10101000", -- 1127 - 0x467  :  168 - 0xa8
    "10100101", -- 1128 - 0x468  :  165 - 0xa5 -- Sprite 0x8d
    "10100010", -- 1129 - 0x469  :  162 - 0xa2
    "10010000", -- 1130 - 0x46a  :  144 - 0x90
    "01001000", -- 1131 - 0x46b  :   72 - 0x48
    "01000111", -- 1132 - 0x46c  :   71 - 0x47
    "00100000", -- 1133 - 0x46d  :   32 - 0x20
    "00011001", -- 1134 - 0x46e  :   25 - 0x19
    "00000111", -- 1135 - 0x46f  :    7 - 0x7
    "11100000", -- 1136 - 0x470  :  224 - 0xe0 -- Sprite 0x8e
    "00011000", -- 1137 - 0x471  :   24 - 0x18
    "00000100", -- 1138 - 0x472  :    4 - 0x4
    "11000010", -- 1139 - 0x473  :  194 - 0xc2
    "00110010", -- 1140 - 0x474  :   50 - 0x32
    "00001001", -- 1141 - 0x475  :    9 - 0x9
    "11000101", -- 1142 - 0x476  :  197 - 0xc5
    "00100101", -- 1143 - 0x477  :   37 - 0x25
    "10100101", -- 1144 - 0x478  :  165 - 0xa5 -- Sprite 0x8f
    "01100101", -- 1145 - 0x479  :  101 - 0x65
    "01000101", -- 1146 - 0x47a  :   69 - 0x45
    "10001010", -- 1147 - 0x47b  :  138 - 0x8a
    "10010010", -- 1148 - 0x47c  :  146 - 0x92
    "00100100", -- 1149 - 0x47d  :   36 - 0x24
    "11011000", -- 1150 - 0x47e  :  216 - 0xd8
    "11100000", -- 1151 - 0x47f  :  224 - 0xe0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x90
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00100000", -- 1154 - 0x482  :   32 - 0x20
    "00110000", -- 1155 - 0x483  :   48 - 0x30
    "00101100", -- 1156 - 0x484  :   44 - 0x2c
    "00100010", -- 1157 - 0x485  :   34 - 0x22
    "00010001", -- 1158 - 0x486  :   17 - 0x11
    "00001000", -- 1159 - 0x487  :    8 - 0x8
    "00000100", -- 1160 - 0x488  :    4 - 0x4 -- Sprite 0x91
    "11110010", -- 1161 - 0x489  :  242 - 0xf2
    "11001111", -- 1162 - 0x48a  :  207 - 0xcf
    "00110000", -- 1163 - 0x48b  :   48 - 0x30
    "00001100", -- 1164 - 0x48c  :   12 - 0xc
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "10000000", -- 1166 - 0x48e  :  128 - 0x80
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "01000010", -- 1168 - 0x490  :   66 - 0x42 -- Sprite 0x92
    "10100101", -- 1169 - 0x491  :  165 - 0xa5
    "10100101", -- 1170 - 0x492  :  165 - 0xa5
    "10011001", -- 1171 - 0x493  :  153 - 0x99
    "10011001", -- 1172 - 0x494  :  153 - 0x99
    "10011001", -- 1173 - 0x495  :  153 - 0x99
    "00000001", -- 1174 - 0x496  :    1 - 0x1
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "11111111", -- 1176 - 0x498  :  255 - 0xff -- Sprite 0x93
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "10000001", -- 1179 - 0x49b  :  129 - 0x81
    "11111111", -- 1180 - 0x49c  :  255 - 0xff
    "11111111", -- 1181 - 0x49d  :  255 - 0xff
    "11111111", -- 1182 - 0x49e  :  255 - 0xff
    "10000001", -- 1183 - 0x49f  :  129 - 0x81
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- Sprite 0x94
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000100", -- 1186 - 0x4a2  :    4 - 0x4
    "00001100", -- 1187 - 0x4a3  :   12 - 0xc
    "00110100", -- 1188 - 0x4a4  :   52 - 0x34
    "01000100", -- 1189 - 0x4a5  :   68 - 0x44
    "10001000", -- 1190 - 0x4a6  :  136 - 0x88
    "00010000", -- 1191 - 0x4a7  :   16 - 0x10
    "00100000", -- 1192 - 0x4a8  :   32 - 0x20 -- Sprite 0x95
    "01001111", -- 1193 - 0x4a9  :   79 - 0x4f
    "11110011", -- 1194 - 0x4aa  :  243 - 0xf3
    "00001100", -- 1195 - 0x4ab  :   12 - 0xc
    "00110000", -- 1196 - 0x4ac  :   48 - 0x30
    "11111111", -- 1197 - 0x4ad  :  255 - 0xff
    "00000001", -- 1198 - 0x4ae  :    1 - 0x1
    "11111111", -- 1199 - 0x4af  :  255 - 0xff
    "01111111", -- 1200 - 0x4b0  :  127 - 0x7f -- Sprite 0x96
    "11111111", -- 1201 - 0x4b1  :  255 - 0xff
    "11111111", -- 1202 - 0x4b2  :  255 - 0xff
    "11111111", -- 1203 - 0x4b3  :  255 - 0xff
    "11111011", -- 1204 - 0x4b4  :  251 - 0xfb
    "11111111", -- 1205 - 0x4b5  :  255 - 0xff
    "11111111", -- 1206 - 0x4b6  :  255 - 0xff
    "11111111", -- 1207 - 0x4b7  :  255 - 0xff
    "11111111", -- 1208 - 0x4b8  :  255 - 0xff -- Sprite 0x97
    "11111111", -- 1209 - 0x4b9  :  255 - 0xff
    "11111111", -- 1210 - 0x4ba  :  255 - 0xff
    "11111111", -- 1211 - 0x4bb  :  255 - 0xff
    "11111111", -- 1212 - 0x4bc  :  255 - 0xff
    "11111111", -- 1213 - 0x4bd  :  255 - 0xff
    "11111110", -- 1214 - 0x4be  :  254 - 0xfe
    "11111111", -- 1215 - 0x4bf  :  255 - 0xff
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Sprite 0x98
    "10111111", -- 1217 - 0x4c1  :  191 - 0xbf
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111111", -- 1219 - 0x4c3  :  255 - 0xff
    "11111011", -- 1220 - 0x4c4  :  251 - 0xfb
    "11111111", -- 1221 - 0x4c5  :  255 - 0xff
    "11111111", -- 1222 - 0x4c6  :  255 - 0xff
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "11111111", -- 1224 - 0x4c8  :  255 - 0xff -- Sprite 0x99
    "11111111", -- 1225 - 0x4c9  :  255 - 0xff
    "11111111", -- 1226 - 0x4ca  :  255 - 0xff
    "11111111", -- 1227 - 0x4cb  :  255 - 0xff
    "11111111", -- 1228 - 0x4cc  :  255 - 0xff
    "11111111", -- 1229 - 0x4cd  :  255 - 0xff
    "11111110", -- 1230 - 0x4ce  :  254 - 0xfe
    "11111111", -- 1231 - 0x4cf  :  255 - 0xff
    "11111110", -- 1232 - 0x4d0  :  254 - 0xfe -- Sprite 0x9a
    "11111111", -- 1233 - 0x4d1  :  255 - 0xff
    "11111111", -- 1234 - 0x4d2  :  255 - 0xff
    "11111111", -- 1235 - 0x4d3  :  255 - 0xff
    "11111011", -- 1236 - 0x4d4  :  251 - 0xfb
    "11111111", -- 1237 - 0x4d5  :  255 - 0xff
    "11111111", -- 1238 - 0x4d6  :  255 - 0xff
    "11111111", -- 1239 - 0x4d7  :  255 - 0xff
    "11111111", -- 1240 - 0x4d8  :  255 - 0xff -- Sprite 0x9b
    "11111111", -- 1241 - 0x4d9  :  255 - 0xff
    "11111111", -- 1242 - 0x4da  :  255 - 0xff
    "11111111", -- 1243 - 0x4db  :  255 - 0xff
    "11111111", -- 1244 - 0x4dc  :  255 - 0xff
    "11111111", -- 1245 - 0x4dd  :  255 - 0xff
    "11111111", -- 1246 - 0x4de  :  255 - 0xff
    "11111111", -- 1247 - 0x4df  :  255 - 0xff
    "11111111", -- 1248 - 0x4e0  :  255 - 0xff -- Sprite 0x9c
    "11111111", -- 1249 - 0x4e1  :  255 - 0xff
    "10100000", -- 1250 - 0x4e2  :  160 - 0xa0
    "10010000", -- 1251 - 0x4e3  :  144 - 0x90
    "10001000", -- 1252 - 0x4e4  :  136 - 0x88
    "10000100", -- 1253 - 0x4e5  :  132 - 0x84
    "01101010", -- 1254 - 0x4e6  :  106 - 0x6a
    "00111111", -- 1255 - 0x4e7  :   63 - 0x3f
    "11111111", -- 1256 - 0x4e8  :  255 - 0xff -- Sprite 0x9d
    "11111111", -- 1257 - 0x4e9  :  255 - 0xff
    "00100001", -- 1258 - 0x4ea  :   33 - 0x21
    "00010001", -- 1259 - 0x4eb  :   17 - 0x11
    "00001001", -- 1260 - 0x4ec  :    9 - 0x9
    "00000101", -- 1261 - 0x4ed  :    5 - 0x5
    "10101010", -- 1262 - 0x4ee  :  170 - 0xaa
    "11111100", -- 1263 - 0x4ef  :  252 - 0xfc
    "11111111", -- 1264 - 0x4f0  :  255 - 0xff -- Sprite 0x9e
    "11111111", -- 1265 - 0x4f1  :  255 - 0xff
    "00100000", -- 1266 - 0x4f2  :   32 - 0x20
    "00010000", -- 1267 - 0x4f3  :   16 - 0x10
    "00001000", -- 1268 - 0x4f4  :    8 - 0x8
    "00000100", -- 1269 - 0x4f5  :    4 - 0x4
    "10101010", -- 1270 - 0x4f6  :  170 - 0xaa
    "11111111", -- 1271 - 0x4f7  :  255 - 0xff
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- Sprite 0x9f
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "11111111", -- 1280 - 0x500  :  255 - 0xff -- Sprite 0xa0
    "11010101", -- 1281 - 0x501  :  213 - 0xd5
    "11111111", -- 1282 - 0x502  :  255 - 0xff
    "00000010", -- 1283 - 0x503  :    2 - 0x2
    "00000010", -- 1284 - 0x504  :    2 - 0x2
    "00000010", -- 1285 - 0x505  :    2 - 0x2
    "00000010", -- 1286 - 0x506  :    2 - 0x2
    "00000010", -- 1287 - 0x507  :    2 - 0x2
    "00000010", -- 1288 - 0x508  :    2 - 0x2 -- Sprite 0xa1
    "00000010", -- 1289 - 0x509  :    2 - 0x2
    "00000010", -- 1290 - 0x50a  :    2 - 0x2
    "00000010", -- 1291 - 0x50b  :    2 - 0x2
    "00000010", -- 1292 - 0x50c  :    2 - 0x2
    "00000010", -- 1293 - 0x50d  :    2 - 0x2
    "00000010", -- 1294 - 0x50e  :    2 - 0x2
    "00000010", -- 1295 - 0x50f  :    2 - 0x2
    "11111111", -- 1296 - 0x510  :  255 - 0xff -- Sprite 0xa2
    "01010101", -- 1297 - 0x511  :   85 - 0x55
    "11111111", -- 1298 - 0x512  :  255 - 0xff
    "01000000", -- 1299 - 0x513  :   64 - 0x40
    "01000000", -- 1300 - 0x514  :   64 - 0x40
    "01000000", -- 1301 - 0x515  :   64 - 0x40
    "01000000", -- 1302 - 0x516  :   64 - 0x40
    "01000000", -- 1303 - 0x517  :   64 - 0x40
    "01000000", -- 1304 - 0x518  :   64 - 0x40 -- Sprite 0xa3
    "01000000", -- 1305 - 0x519  :   64 - 0x40
    "01000000", -- 1306 - 0x51a  :   64 - 0x40
    "01000000", -- 1307 - 0x51b  :   64 - 0x40
    "01000000", -- 1308 - 0x51c  :   64 - 0x40
    "01000000", -- 1309 - 0x51d  :   64 - 0x40
    "01000000", -- 1310 - 0x51e  :   64 - 0x40
    "01000000", -- 1311 - 0x51f  :   64 - 0x40
    "00110001", -- 1312 - 0x520  :   49 - 0x31 -- Sprite 0xa4
    "01001000", -- 1313 - 0x521  :   72 - 0x48
    "01000101", -- 1314 - 0x522  :   69 - 0x45
    "10000101", -- 1315 - 0x523  :  133 - 0x85
    "10000011", -- 1316 - 0x524  :  131 - 0x83
    "10000010", -- 1317 - 0x525  :  130 - 0x82
    "01100010", -- 1318 - 0x526  :   98 - 0x62
    "00010010", -- 1319 - 0x527  :   18 - 0x12
    "00110010", -- 1320 - 0x528  :   50 - 0x32 -- Sprite 0xa5
    "00100010", -- 1321 - 0x529  :   34 - 0x22
    "01000010", -- 1322 - 0x52a  :   66 - 0x42
    "01000000", -- 1323 - 0x52b  :   64 - 0x40
    "01000000", -- 1324 - 0x52c  :   64 - 0x40
    "00100000", -- 1325 - 0x52d  :   32 - 0x20
    "00011110", -- 1326 - 0x52e  :   30 - 0x1e
    "00000111", -- 1327 - 0x52f  :    7 - 0x7
    "10000000", -- 1328 - 0x530  :  128 - 0x80 -- Sprite 0xa6
    "11100000", -- 1329 - 0x531  :  224 - 0xe0
    "00111000", -- 1330 - 0x532  :   56 - 0x38
    "00100100", -- 1331 - 0x533  :   36 - 0x24
    "00000100", -- 1332 - 0x534  :    4 - 0x4
    "00001000", -- 1333 - 0x535  :    8 - 0x8
    "00110000", -- 1334 - 0x536  :   48 - 0x30
    "00100000", -- 1335 - 0x537  :   32 - 0x20
    "00110000", -- 1336 - 0x538  :   48 - 0x30 -- Sprite 0xa7
    "00001000", -- 1337 - 0x539  :    8 - 0x8
    "00001000", -- 1338 - 0x53a  :    8 - 0x8
    "00110000", -- 1339 - 0x53b  :   48 - 0x30
    "00100000", -- 1340 - 0x53c  :   32 - 0x20
    "00100000", -- 1341 - 0x53d  :   32 - 0x20
    "00110000", -- 1342 - 0x53e  :   48 - 0x30
    "11110000", -- 1343 - 0x53f  :  240 - 0xf0
    "11111111", -- 1344 - 0x540  :  255 - 0xff -- Sprite 0xa8
    "11010010", -- 1345 - 0x541  :  210 - 0xd2
    "11110100", -- 1346 - 0x542  :  244 - 0xf4
    "11011000", -- 1347 - 0x543  :  216 - 0xd8
    "11111000", -- 1348 - 0x544  :  248 - 0xf8
    "11010100", -- 1349 - 0x545  :  212 - 0xd4
    "11110010", -- 1350 - 0x546  :  242 - 0xf2
    "11010001", -- 1351 - 0x547  :  209 - 0xd1
    "11110001", -- 1352 - 0x548  :  241 - 0xf1 -- Sprite 0xa9
    "11010010", -- 1353 - 0x549  :  210 - 0xd2
    "11110100", -- 1354 - 0x54a  :  244 - 0xf4
    "11011000", -- 1355 - 0x54b  :  216 - 0xd8
    "11111000", -- 1356 - 0x54c  :  248 - 0xf8
    "11010100", -- 1357 - 0x54d  :  212 - 0xd4
    "11110010", -- 1358 - 0x54e  :  242 - 0xf2
    "11111111", -- 1359 - 0x54f  :  255 - 0xff
    "11111111", -- 1360 - 0x550  :  255 - 0xff -- Sprite 0xaa
    "01000010", -- 1361 - 0x551  :   66 - 0x42
    "00100100", -- 1362 - 0x552  :   36 - 0x24
    "00011000", -- 1363 - 0x553  :   24 - 0x18
    "00011000", -- 1364 - 0x554  :   24 - 0x18
    "00100100", -- 1365 - 0x555  :   36 - 0x24
    "01000010", -- 1366 - 0x556  :   66 - 0x42
    "10000001", -- 1367 - 0x557  :  129 - 0x81
    "10000001", -- 1368 - 0x558  :  129 - 0x81 -- Sprite 0xab
    "01000010", -- 1369 - 0x559  :   66 - 0x42
    "00100100", -- 1370 - 0x55a  :   36 - 0x24
    "00011000", -- 1371 - 0x55b  :   24 - 0x18
    "00011000", -- 1372 - 0x55c  :   24 - 0x18
    "00100100", -- 1373 - 0x55d  :   36 - 0x24
    "01000010", -- 1374 - 0x55e  :   66 - 0x42
    "11111111", -- 1375 - 0x55f  :  255 - 0xff
    "11111111", -- 1376 - 0x560  :  255 - 0xff -- Sprite 0xac
    "01001101", -- 1377 - 0x561  :   77 - 0x4d
    "00101111", -- 1378 - 0x562  :   47 - 0x2f
    "00011101", -- 1379 - 0x563  :   29 - 0x1d
    "00011111", -- 1380 - 0x564  :   31 - 0x1f
    "00101101", -- 1381 - 0x565  :   45 - 0x2d
    "01001111", -- 1382 - 0x566  :   79 - 0x4f
    "10001101", -- 1383 - 0x567  :  141 - 0x8d
    "10001111", -- 1384 - 0x568  :  143 - 0x8f -- Sprite 0xad
    "01001101", -- 1385 - 0x569  :   77 - 0x4d
    "00101111", -- 1386 - 0x56a  :   47 - 0x2f
    "00011101", -- 1387 - 0x56b  :   29 - 0x1d
    "00011111", -- 1388 - 0x56c  :   31 - 0x1f
    "00101101", -- 1389 - 0x56d  :   45 - 0x2d
    "01001111", -- 1390 - 0x56e  :   79 - 0x4f
    "11111111", -- 1391 - 0x56f  :  255 - 0xff
    "00000001", -- 1392 - 0x570  :    1 - 0x1 -- Sprite 0xae
    "00000011", -- 1393 - 0x571  :    3 - 0x3
    "00000110", -- 1394 - 0x572  :    6 - 0x6
    "00000111", -- 1395 - 0x573  :    7 - 0x7
    "00000111", -- 1396 - 0x574  :    7 - 0x7
    "00000111", -- 1397 - 0x575  :    7 - 0x7
    "00000110", -- 1398 - 0x576  :    6 - 0x6
    "00000111", -- 1399 - 0x577  :    7 - 0x7
    "00000110", -- 1400 - 0x578  :    6 - 0x6 -- Sprite 0xaf
    "00000110", -- 1401 - 0x579  :    6 - 0x6
    "00001110", -- 1402 - 0x57a  :   14 - 0xe
    "00001111", -- 1403 - 0x57b  :   15 - 0xf
    "00001110", -- 1404 - 0x57c  :   14 - 0xe
    "00011010", -- 1405 - 0x57d  :   26 - 0x1a
    "00011011", -- 1406 - 0x57e  :   27 - 0x1b
    "00001111", -- 1407 - 0x57f  :   15 - 0xf
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Sprite 0xb0
    "11000000", -- 1409 - 0x581  :  192 - 0xc0
    "11110000", -- 1410 - 0x582  :  240 - 0xf0
    "10001000", -- 1411 - 0x583  :  136 - 0x88
    "00010100", -- 1412 - 0x584  :   20 - 0x14
    "01101000", -- 1413 - 0x585  :  104 - 0x68
    "10101000", -- 1414 - 0x586  :  168 - 0xa8
    "00101100", -- 1415 - 0x587  :   44 - 0x2c
    "00000100", -- 1416 - 0x588  :    4 - 0x4 -- Sprite 0xb1
    "00111000", -- 1417 - 0x589  :   56 - 0x38
    "00010000", -- 1418 - 0x58a  :   16 - 0x10
    "10100000", -- 1419 - 0x58b  :  160 - 0xa0
    "01100000", -- 1420 - 0x58c  :   96 - 0x60
    "00100000", -- 1421 - 0x58d  :   32 - 0x20
    "00010000", -- 1422 - 0x58e  :   16 - 0x10
    "10001000", -- 1423 - 0x58f  :  136 - 0x88
    "00001111", -- 1424 - 0x590  :   15 - 0xf -- Sprite 0xb2
    "00011011", -- 1425 - 0x591  :   27 - 0x1b
    "00011011", -- 1426 - 0x592  :   27 - 0x1b
    "00001110", -- 1427 - 0x593  :   14 - 0xe
    "00000110", -- 1428 - 0x594  :    6 - 0x6
    "00001100", -- 1429 - 0x595  :   12 - 0xc
    "00001100", -- 1430 - 0x596  :   12 - 0xc
    "00111111", -- 1431 - 0x597  :   63 - 0x3f
    "01111111", -- 1432 - 0x598  :  127 - 0x7f -- Sprite 0xb3
    "01100000", -- 1433 - 0x599  :   96 - 0x60
    "01100000", -- 1434 - 0x59a  :   96 - 0x60
    "01100000", -- 1435 - 0x59b  :   96 - 0x60
    "01100000", -- 1436 - 0x59c  :   96 - 0x60
    "01100000", -- 1437 - 0x59d  :   96 - 0x60
    "01101010", -- 1438 - 0x59e  :  106 - 0x6a
    "01111111", -- 1439 - 0x59f  :  127 - 0x7f
    "01001000", -- 1440 - 0x5a0  :   72 - 0x48 -- Sprite 0xb4
    "00110000", -- 1441 - 0x5a1  :   48 - 0x30
    "00010000", -- 1442 - 0x5a2  :   16 - 0x10
    "00010000", -- 1443 - 0x5a3  :   16 - 0x10
    "00001000", -- 1444 - 0x5a4  :    8 - 0x8
    "00001000", -- 1445 - 0x5a5  :    8 - 0x8
    "00001000", -- 1446 - 0x5a6  :    8 - 0x8
    "11111100", -- 1447 - 0x5a7  :  252 - 0xfc
    "11111110", -- 1448 - 0x5a8  :  254 - 0xfe -- Sprite 0xb5
    "00000110", -- 1449 - 0x5a9  :    6 - 0x6
    "00000010", -- 1450 - 0x5aa  :    2 - 0x2
    "00000110", -- 1451 - 0x5ab  :    6 - 0x6
    "00000010", -- 1452 - 0x5ac  :    2 - 0x2
    "00000110", -- 1453 - 0x5ad  :    6 - 0x6
    "10101010", -- 1454 - 0x5ae  :  170 - 0xaa
    "11111110", -- 1455 - 0x5af  :  254 - 0xfe
    "11111111", -- 1456 - 0x5b0  :  255 - 0xff -- Sprite 0xb6
    "10000000", -- 1457 - 0x5b1  :  128 - 0x80
    "10000000", -- 1458 - 0x5b2  :  128 - 0x80
    "10000000", -- 1459 - 0x5b3  :  128 - 0x80
    "10000000", -- 1460 - 0x5b4  :  128 - 0x80
    "10000000", -- 1461 - 0x5b5  :  128 - 0x80
    "10010101", -- 1462 - 0x5b6  :  149 - 0x95
    "11111111", -- 1463 - 0x5b7  :  255 - 0xff
    "11111111", -- 1464 - 0x5b8  :  255 - 0xff -- Sprite 0xb7
    "10000100", -- 1465 - 0x5b9  :  132 - 0x84
    "10001100", -- 1466 - 0x5ba  :  140 - 0x8c
    "10000100", -- 1467 - 0x5bb  :  132 - 0x84
    "10001100", -- 1468 - 0x5bc  :  140 - 0x8c
    "10000100", -- 1469 - 0x5bd  :  132 - 0x84
    "10101100", -- 1470 - 0x5be  :  172 - 0xac
    "11111111", -- 1471 - 0x5bf  :  255 - 0xff
    "11111111", -- 1472 - 0x5c0  :  255 - 0xff -- Sprite 0xb8
    "00100001", -- 1473 - 0x5c1  :   33 - 0x21
    "01100001", -- 1474 - 0x5c2  :   97 - 0x61
    "00100011", -- 1475 - 0x5c3  :   35 - 0x23
    "01100001", -- 1476 - 0x5c4  :   97 - 0x61
    "00100011", -- 1477 - 0x5c5  :   35 - 0x23
    "01100101", -- 1478 - 0x5c6  :  101 - 0x65
    "11111111", -- 1479 - 0x5c7  :  255 - 0xff
    "11111111", -- 1480 - 0x5c8  :  255 - 0xff -- Sprite 0xb9
    "00000001", -- 1481 - 0x5c9  :    1 - 0x1
    "00000011", -- 1482 - 0x5ca  :    3 - 0x3
    "00000001", -- 1483 - 0x5cb  :    1 - 0x1
    "00000011", -- 1484 - 0x5cc  :    3 - 0x3
    "00000001", -- 1485 - 0x5cd  :    1 - 0x1
    "10101011", -- 1486 - 0x5ce  :  171 - 0xab
    "11111111", -- 1487 - 0x5cf  :  255 - 0xff
    "11111111", -- 1488 - 0x5d0  :  255 - 0xff -- Sprite 0xba
    "11010101", -- 1489 - 0x5d1  :  213 - 0xd5
    "10101010", -- 1490 - 0x5d2  :  170 - 0xaa
    "11111111", -- 1491 - 0x5d3  :  255 - 0xff
    "10000000", -- 1492 - 0x5d4  :  128 - 0x80
    "10000000", -- 1493 - 0x5d5  :  128 - 0x80
    "10010101", -- 1494 - 0x5d6  :  149 - 0x95
    "11111111", -- 1495 - 0x5d7  :  255 - 0xff
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0 -- Sprite 0xbb
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "11111111", -- 1504 - 0x5e0  :  255 - 0xff -- Sprite 0xbc
    "01010101", -- 1505 - 0x5e1  :   85 - 0x55
    "10101011", -- 1506 - 0x5e2  :  171 - 0xab
    "11111111", -- 1507 - 0x5e3  :  255 - 0xff
    "01100001", -- 1508 - 0x5e4  :   97 - 0x61
    "00100011", -- 1509 - 0x5e5  :   35 - 0x23
    "01100101", -- 1510 - 0x5e6  :  101 - 0x65
    "11111111", -- 1511 - 0x5e7  :  255 - 0xff
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- Sprite 0xbd
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00000000", -- 1514 - 0x5ea  :    0 - 0x0
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "00000000", -- 1516 - 0x5ec  :    0 - 0x0
    "00000000", -- 1517 - 0x5ed  :    0 - 0x0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Sprite 0xbe
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Sprite 0xbf
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0xc0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000000", -- 1542 - 0x606  :    0 - 0x0
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00000000", -- 1544 - 0x608  :    0 - 0x0 -- Sprite 0xc1
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- Sprite 0xc3
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0 -- Sprite 0xc5
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000001", -- 1578 - 0x62a  :    1 - 0x1
    "00000110", -- 1579 - 0x62b  :    6 - 0x6
    "00001010", -- 1580 - 0x62c  :   10 - 0xa
    "00010100", -- 1581 - 0x62d  :   20 - 0x14
    "00010000", -- 1582 - 0x62e  :   16 - 0x10
    "00101000", -- 1583 - 0x62f  :   40 - 0x28
    "00011111", -- 1584 - 0x630  :   31 - 0x1f -- Sprite 0xc6
    "01100000", -- 1585 - 0x631  :   96 - 0x60
    "10100000", -- 1586 - 0x632  :  160 - 0xa0
    "01000000", -- 1587 - 0x633  :   64 - 0x40
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "00000000", -- 1589 - 0x635  :    0 - 0x0
    "00000000", -- 1590 - 0x636  :    0 - 0x0
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00110000", -- 1592 - 0x638  :   48 - 0x30 -- Sprite 0xc7
    "01000000", -- 1593 - 0x639  :   64 - 0x40
    "01100000", -- 1594 - 0x63a  :   96 - 0x60
    "11000000", -- 1595 - 0x63b  :  192 - 0xc0
    "10000000", -- 1596 - 0x63c  :  128 - 0x80
    "10100000", -- 1597 - 0x63d  :  160 - 0xa0
    "11000000", -- 1598 - 0x63e  :  192 - 0xc0
    "10000000", -- 1599 - 0x63f  :  128 - 0x80
    "11111111", -- 1600 - 0x640  :  255 - 0xff -- Sprite 0xc8
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00010100", -- 1608 - 0x648  :   20 - 0x14 -- Sprite 0xc9
    "00101010", -- 1609 - 0x649  :   42 - 0x2a
    "00010110", -- 1610 - 0x64a  :   22 - 0x16
    "00101011", -- 1611 - 0x64b  :   43 - 0x2b
    "00010101", -- 1612 - 0x64c  :   21 - 0x15
    "00101011", -- 1613 - 0x64d  :   43 - 0x2b
    "00010101", -- 1614 - 0x64e  :   21 - 0x15
    "00101011", -- 1615 - 0x64f  :   43 - 0x2b
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0xca
    "00000100", -- 1617 - 0x651  :    4 - 0x4
    "00000100", -- 1618 - 0x652  :    4 - 0x4
    "00000101", -- 1619 - 0x653  :    5 - 0x5
    "00010101", -- 1620 - 0x654  :   21 - 0x15
    "00010101", -- 1621 - 0x655  :   21 - 0x15
    "01010101", -- 1622 - 0x656  :   85 - 0x55
    "01010101", -- 1623 - 0x657  :   85 - 0x55
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- Sprite 0xcb
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00010000", -- 1626 - 0x65a  :   16 - 0x10
    "00010000", -- 1627 - 0x65b  :   16 - 0x10
    "01010001", -- 1628 - 0x65c  :   81 - 0x51
    "01010101", -- 1629 - 0x65d  :   85 - 0x55
    "01010101", -- 1630 - 0x65e  :   85 - 0x55
    "01010101", -- 1631 - 0x65f  :   85 - 0x55
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Sprite 0xcc
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000101", -- 1635 - 0x663  :    5 - 0x5
    "00001111", -- 1636 - 0x664  :   15 - 0xf
    "00000111", -- 1637 - 0x665  :    7 - 0x7
    "00000011", -- 1638 - 0x666  :    3 - 0x3
    "00000001", -- 1639 - 0x667  :    1 - 0x1
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "10000000", -- 1642 - 0x66a  :  128 - 0x80
    "11010000", -- 1643 - 0x66b  :  208 - 0xd0
    "11111000", -- 1644 - 0x66c  :  248 - 0xf8
    "11110000", -- 1645 - 0x66d  :  240 - 0xf0
    "11100000", -- 1646 - 0x66e  :  224 - 0xe0
    "11000000", -- 1647 - 0x66f  :  192 - 0xc0
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "01111000", -- 1651 - 0x673  :  120 - 0x78
    "11001111", -- 1652 - 0x674  :  207 - 0xcf
    "10000000", -- 1653 - 0x675  :  128 - 0x80
    "11001111", -- 1654 - 0x676  :  207 - 0xcf
    "01001000", -- 1655 - 0x677  :   72 - 0x48
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- Sprite 0xcf
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00011110", -- 1659 - 0x67b  :   30 - 0x1e
    "11110011", -- 1660 - 0x67c  :  243 - 0xf3
    "00000001", -- 1661 - 0x67d  :    1 - 0x1
    "11110011", -- 1662 - 0x67e  :  243 - 0xf3
    "00010010", -- 1663 - 0x67f  :   18 - 0x12
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0xd0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- Sprite 0xd1
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00001000", -- 1680 - 0x690  :    8 - 0x8 -- Sprite 0xd2
    "00001100", -- 1681 - 0x691  :   12 - 0xc
    "00001000", -- 1682 - 0x692  :    8 - 0x8
    "00001000", -- 1683 - 0x693  :    8 - 0x8
    "00001010", -- 1684 - 0x694  :   10 - 0xa
    "00001000", -- 1685 - 0x695  :    8 - 0x8
    "00001000", -- 1686 - 0x696  :    8 - 0x8
    "00001100", -- 1687 - 0x697  :   12 - 0xc
    "00010000", -- 1688 - 0x698  :   16 - 0x10 -- Sprite 0xd3
    "00010000", -- 1689 - 0x699  :   16 - 0x10
    "00110000", -- 1690 - 0x69a  :   48 - 0x30
    "00010000", -- 1691 - 0x69b  :   16 - 0x10
    "01010000", -- 1692 - 0x69c  :   80 - 0x50
    "00010000", -- 1693 - 0x69d  :   16 - 0x10
    "00110000", -- 1694 - 0x69e  :   48 - 0x30
    "00010000", -- 1695 - 0x69f  :   16 - 0x10
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0xd4
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "11111000", -- 1704 - 0x6a8  :  248 - 0xf8 -- Sprite 0xd5
    "00000110", -- 1705 - 0x6a9  :    6 - 0x6
    "00000001", -- 1706 - 0x6aa  :    1 - 0x1
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "10000000", -- 1714 - 0x6b2  :  128 - 0x80
    "01100000", -- 1715 - 0x6b3  :   96 - 0x60
    "01010000", -- 1716 - 0x6b4  :   80 - 0x50
    "10101000", -- 1717 - 0x6b5  :  168 - 0xa8
    "01011000", -- 1718 - 0x6b6  :   88 - 0x58
    "00101100", -- 1719 - 0x6b7  :   44 - 0x2c
    "10100000", -- 1720 - 0x6b8  :  160 - 0xa0 -- Sprite 0xd7
    "11000000", -- 1721 - 0x6b9  :  192 - 0xc0
    "10000000", -- 1722 - 0x6ba  :  128 - 0x80
    "01010000", -- 1723 - 0x6bb  :   80 - 0x50
    "01100000", -- 1724 - 0x6bc  :   96 - 0x60
    "00111000", -- 1725 - 0x6bd  :   56 - 0x38
    "00001000", -- 1726 - 0x6be  :    8 - 0x8
    "00000111", -- 1727 - 0x6bf  :    7 - 0x7
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Sprite 0xd8
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000000", -- 1734 - 0x6c6  :    0 - 0x0
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "00010101", -- 1736 - 0x6c8  :   21 - 0x15 -- Sprite 0xd9
    "00101011", -- 1737 - 0x6c9  :   43 - 0x2b
    "00010101", -- 1738 - 0x6ca  :   21 - 0x15
    "00101010", -- 1739 - 0x6cb  :   42 - 0x2a
    "01010110", -- 1740 - 0x6cc  :   86 - 0x56
    "10101100", -- 1741 - 0x6cd  :  172 - 0xac
    "01010000", -- 1742 - 0x6ce  :   80 - 0x50
    "11100000", -- 1743 - 0x6cf  :  224 - 0xe0
    "00000001", -- 1744 - 0x6d0  :    1 - 0x1 -- Sprite 0xda
    "00001101", -- 1745 - 0x6d1  :   13 - 0xd
    "00010011", -- 1746 - 0x6d2  :   19 - 0x13
    "00001101", -- 1747 - 0x6d3  :   13 - 0xd
    "00000001", -- 1748 - 0x6d4  :    1 - 0x1
    "00000001", -- 1749 - 0x6d5  :    1 - 0x1
    "00000001", -- 1750 - 0x6d6  :    1 - 0x1
    "00000001", -- 1751 - 0x6d7  :    1 - 0x1
    "11000000", -- 1752 - 0x6d8  :  192 - 0xc0 -- Sprite 0xdb
    "01000000", -- 1753 - 0x6d9  :   64 - 0x40
    "01000000", -- 1754 - 0x6da  :   64 - 0x40
    "01011000", -- 1755 - 0x6db  :   88 - 0x58
    "01100100", -- 1756 - 0x6dc  :  100 - 0x64
    "01011000", -- 1757 - 0x6dd  :   88 - 0x58
    "01000000", -- 1758 - 0x6de  :   64 - 0x40
    "01000000", -- 1759 - 0x6df  :   64 - 0x40
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Sprite 0xdc
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000110", -- 1763 - 0x6e3  :    6 - 0x6
    "00000111", -- 1764 - 0x6e4  :    7 - 0x7
    "00000111", -- 1765 - 0x6e5  :    7 - 0x7
    "00000111", -- 1766 - 0x6e6  :    7 - 0x7
    "00000011", -- 1767 - 0x6e7  :    3 - 0x3
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- Sprite 0xdd
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "10110000", -- 1771 - 0x6eb  :  176 - 0xb0
    "11110000", -- 1772 - 0x6ec  :  240 - 0xf0
    "11110000", -- 1773 - 0x6ed  :  240 - 0xf0
    "11110000", -- 1774 - 0x6ee  :  240 - 0xf0
    "11100000", -- 1775 - 0x6ef  :  224 - 0xe0
    "11001111", -- 1776 - 0x6f0  :  207 - 0xcf -- Sprite 0xde
    "10000000", -- 1777 - 0x6f1  :  128 - 0x80
    "11001111", -- 1778 - 0x6f2  :  207 - 0xcf
    "01001000", -- 1779 - 0x6f3  :   72 - 0x48
    "01001000", -- 1780 - 0x6f4  :   72 - 0x48
    "01001000", -- 1781 - 0x6f5  :   72 - 0x48
    "01001000", -- 1782 - 0x6f6  :   72 - 0x48
    "01001000", -- 1783 - 0x6f7  :   72 - 0x48
    "11110011", -- 1784 - 0x6f8  :  243 - 0xf3 -- Sprite 0xdf
    "00000001", -- 1785 - 0x6f9  :    1 - 0x1
    "11110011", -- 1786 - 0x6fa  :  243 - 0xf3
    "00010010", -- 1787 - 0x6fb  :   18 - 0x12
    "00010010", -- 1788 - 0x6fc  :   18 - 0x12
    "00010010", -- 1789 - 0x6fd  :   18 - 0x12
    "00010010", -- 1790 - 0x6fe  :   18 - 0x12
    "00010010", -- 1791 - 0x6ff  :   18 - 0x12
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Sprite 0xe0
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0 -- Sprite 0xe1
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0 -- Sprite 0xe2
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000000", -- 1816 - 0x718  :    0 - 0x0 -- Sprite 0xe3
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Sprite 0xe4
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000000", -- 1828 - 0x724  :    0 - 0x0
    "00000000", -- 1829 - 0x725  :    0 - 0x0
    "00000000", -- 1830 - 0x726  :    0 - 0x0
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- Sprite 0xe5
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "00000000", -- 1840 - 0x730  :    0 - 0x0 -- Sprite 0xe6
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "00000000", -- 1845 - 0x735  :    0 - 0x0
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0 -- Sprite 0xe7
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0xe8
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0 -- Sprite 0xe9
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Sprite 0xea
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- Sprite 0xeb
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0 -- Sprite 0xed
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Sprite 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- Sprite 0xef
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- Sprite 0xf1
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Sprite 0xf2
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- Sprite 0xf3
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Sprite 0xf4
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0 -- Sprite 0xf5
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0xf6
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- Sprite 0xf7
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0xf8
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- Sprite 0xf9
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Sprite 0xfa
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- Sprite 0xfb
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0xfc
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "10001110", -- 2018 - 0x7e2  :  142 - 0x8e
    "10001010", -- 2019 - 0x7e3  :  138 - 0x8a
    "10001010", -- 2020 - 0x7e4  :  138 - 0x8a
    "10001010", -- 2021 - 0x7e5  :  138 - 0x8a
    "10001010", -- 2022 - 0x7e6  :  138 - 0x8a
    "11101110", -- 2023 - 0x7e7  :  238 - 0xee
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- Sprite 0xfd
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "01001100", -- 2026 - 0x7ea  :   76 - 0x4c
    "10101010", -- 2027 - 0x7eb  :  170 - 0xaa
    "10101010", -- 2028 - 0x7ec  :  170 - 0xaa
    "11101010", -- 2029 - 0x7ed  :  234 - 0xea
    "10101010", -- 2030 - 0x7ee  :  170 - 0xaa
    "10101100", -- 2031 - 0x7ef  :  172 - 0xac
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Sprite 0xfe
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "11101100", -- 2034 - 0x7f2  :  236 - 0xec
    "01001010", -- 2035 - 0x7f3  :   74 - 0x4a
    "01001010", -- 2036 - 0x7f4  :   74 - 0x4a
    "01001010", -- 2037 - 0x7f5  :   74 - 0x4a
    "01001010", -- 2038 - 0x7f6  :   74 - 0x4a
    "11101010", -- 2039 - 0x7f7  :  234 - 0xea
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Sprite 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "01100000", -- 2042 - 0x7fa  :   96 - 0x60
    "10001000", -- 2043 - 0x7fb  :  136 - 0x88
    "10100000", -- 2044 - 0x7fc  :  160 - 0xa0
    "10100000", -- 2045 - 0x7fd  :  160 - 0xa0
    "10101000", -- 2046 - 0x7fe  :  168 - 0xa8
    "01000000"  -- 2047 - 0x7ff  :   64 - 0x40
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
