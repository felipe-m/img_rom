---   Background Pattern table COLOR PLANE 0
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: lawnmower_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_LAWN_BG_PLN0 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_LAWN_BG_PLN0;

architecture BEHAVIORAL of ROM_PTABLE_LAWN_BG_PLN0 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table COLOR PLANE 0
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Background 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000101", --    8 -  0x8  :    5 - 0x5 -- Background 0x1
    "01010101", --    9 -  0x9  :   85 - 0x55
    "01010101", --   10 -  0xa  :   85 - 0x55
    "01010000", --   11 -  0xb  :   80 - 0x50
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000101", --   16 - 0x10  :    5 - 0x5 -- Background 0x2
    "01010000", --   17 - 0x11  :   80 - 0x50
    "00000101", --   18 - 0x12  :    5 - 0x5
    "01010000", --   19 - 0x13  :   80 - 0x50
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00000000", --   21 - 0x15  :    0 - 0x0
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000101", --   24 - 0x18  :    5 - 0x5 -- Background 0x3
    "01010000", --   25 - 0x19  :   80 - 0x50
    "00000101", --   26 - 0x1a  :    5 - 0x5
    "01010000", --   27 - 0x1b  :   80 - 0x50
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000101", --   32 - 0x20  :    5 - 0x5 -- Background 0x4
    "01010101", --   33 - 0x21  :   85 - 0x55
    "01010101", --   34 - 0x22  :   85 - 0x55
    "01010000", --   35 - 0x23  :   80 - 0x50
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- Background 0x5
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "01010101", --   48 - 0x30  :   85 - 0x55 -- Background 0x6
    "01010101", --   49 - 0x31  :   85 - 0x55
    "01010100", --   50 - 0x32  :   84 - 0x54
    "00000000", --   51 - 0x33  :    0 - 0x0
    "00000000", --   52 - 0x34  :    0 - 0x0
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000000", --   54 - 0x36  :    0 - 0x0
    "00010101", --   55 - 0x37  :   21 - 0x15
    "10101010", --   56 - 0x38  :  170 - 0xaa -- Background 0x7
    "10011010", --   57 - 0x39  :  154 - 0x9a
    "10010100", --   58 - 0x3a  :  148 - 0x94
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00010110", --   63 - 0x3f  :   22 - 0x16
    "01010000", --   64 - 0x40  :   80 - 0x50 -- Background 0x8
    "00000101", --   65 - 0x41  :    5 - 0x5
    "10010100", --   66 - 0x42  :  148 - 0x94
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00010101", --   71 - 0x47  :   21 - 0x15
    "01010000", --   72 - 0x48  :   80 - 0x50 -- Background 0x9
    "00000101", --   73 - 0x49  :    5 - 0x5
    "10010100", --   74 - 0x4a  :  148 - 0x94
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00010110", --   79 - 0x4f  :   22 - 0x16
    "10100110", --   80 - 0x50  :  166 - 0xa6 -- Background 0xa
    "10101010", --   81 - 0x51  :  170 - 0xaa
    "10010100", --   82 - 0x52  :  148 - 0x94
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00010101", --   87 - 0x57  :   21 - 0x15
    "01010101", --   88 - 0x58  :   85 - 0x55 -- Background 0xb
    "01010101", --   89 - 0x59  :   85 - 0x55
    "01010100", --   90 - 0x5a  :   84 - 0x54
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00001110", --   95 - 0x5f  :   14 - 0xe
    "01010101", --   96 - 0x60  :   85 - 0x55 -- Background 0xc
    "01010100", --   97 - 0x61  :   84 - 0x54
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00011010", --  102 - 0x66  :   26 - 0x1a
    "10011101", --  103 - 0x67  :  157 - 0x9d
    "01010101", --  104 - 0x68  :   85 - 0x55 -- Background 0xd
    "01010100", --  105 - 0x69  :   84 - 0x54
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00010111", --  110 - 0x6e  :   23 - 0x17
    "01010101", --  111 - 0x6f  :   85 - 0x55
    "00000101", --  112 - 0x70  :    5 - 0x5 -- Background 0xe
    "01010100", --  113 - 0x71  :   84 - 0x54
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00010101", --  118 - 0x76  :   21 - 0x15
    "01010000", --  119 - 0x77  :   80 - 0x50
    "00000101", --  120 - 0x78  :    5 - 0x5 -- Background 0xf
    "01010100", --  121 - 0x79  :   84 - 0x54
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00010111", --  126 - 0x7e  :   23 - 0x17
    "01010101", --  127 - 0x7f  :   85 - 0x55
    "01010101", --  128 - 0x80  :   85 - 0x55 -- Background 0x10
    "01010100", --  129 - 0x81  :   84 - 0x54
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00011010", --  134 - 0x86  :   26 - 0x1a
    "10011101", --  135 - 0x87  :  157 - 0x9d
    "01010101", --  136 - 0x88  :   85 - 0x55 -- Background 0x11
    "01010100", --  137 - 0x89  :   84 - 0x54
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00001110", --  142 - 0x8e  :   14 - 0xe
    "00000111", --  143 - 0x8f  :    7 - 0x7
    "01010101", --  144 - 0x90  :   85 - 0x55 -- Background 0x12
    "01010101", --  145 - 0x91  :   85 - 0x55
    "01000000", --  146 - 0x92  :   64 - 0x40
    "00000000", --  147 - 0x93  :    0 - 0x0
    "00000000", --  148 - 0x94  :    0 - 0x0
    "00010101", --  149 - 0x95  :   21 - 0x15
    "01010101", --  150 - 0x96  :   85 - 0x55
    "01010101", --  151 - 0x97  :   85 - 0x55
    "01010101", --  152 - 0x98  :   85 - 0x55 -- Background 0x13
    "10101001", --  153 - 0x99  :  169 - 0xa9
    "01000000", --  154 - 0x9a  :   64 - 0x40
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "00010110", --  157 - 0x9d  :   22 - 0x16
    "01010101", --  158 - 0x9e  :   85 - 0x55
    "01101010", --  159 - 0x9f  :  106 - 0x6a
    "01010101", --  160 - 0xa0  :   85 - 0x55 -- Background 0x14
    "01011001", --  161 - 0xa1  :   89 - 0x59
    "01000000", --  162 - 0xa2  :   64 - 0x40
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "00000000", --  164 - 0xa4  :    0 - 0x0
    "00010101", --  165 - 0xa5  :   21 - 0x15
    "01000000", --  166 - 0xa6  :   64 - 0x40
    "01010101", --  167 - 0xa7  :   85 - 0x55
    "01010101", --  168 - 0xa8  :   85 - 0x55 -- Background 0x15
    "01011001", --  169 - 0xa9  :   89 - 0x59
    "01000000", --  170 - 0xaa  :   64 - 0x40
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00010110", --  173 - 0xad  :   22 - 0x16
    "01010101", --  174 - 0xae  :   85 - 0x55
    "01101010", --  175 - 0xaf  :  106 - 0x6a
    "01010101", --  176 - 0xb0  :   85 - 0x55 -- Background 0x16
    "10101001", --  177 - 0xb1  :  169 - 0xa9
    "01000000", --  178 - 0xb2  :   64 - 0x40
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00010101", --  181 - 0xb5  :   21 - 0x15
    "01010101", --  182 - 0xb6  :   85 - 0x55
    "01010101", --  183 - 0xb7  :   85 - 0x55
    "01010101", --  184 - 0xb8  :   85 - 0x55 -- Background 0x17
    "01010101", --  185 - 0xb9  :   85 - 0x55
    "01000000", --  186 - 0xba  :   64 - 0x40
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00010100", --  189 - 0xbd  :   20 - 0x14
    "00000110", --  190 - 0xbe  :    6 - 0x6
    "00001000", --  191 - 0xbf  :    8 - 0x8
    "01010101", --  192 - 0xc0  :   85 - 0x55 -- Background 0x18
    "01000000", --  193 - 0xc1  :   64 - 0x40
    "00000000", --  194 - 0xc2  :    0 - 0x0
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00011010", --  196 - 0xc4  :   26 - 0x1a
    "01010111", --  197 - 0xc5  :   87 - 0x57
    "01010101", --  198 - 0xc6  :   85 - 0x55
    "01011101", --  199 - 0xc7  :   93 - 0x5d
    "01011010", --  200 - 0xc8  :   90 - 0x5a -- Background 0x19
    "01000000", --  201 - 0xc9  :   64 - 0x40
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00010101", --  204 - 0xcc  :   21 - 0x15
    "01010111", --  205 - 0xcd  :   87 - 0x57
    "01011010", --  206 - 0xce  :   90 - 0x5a
    "01011101", --  207 - 0xcf  :   93 - 0x5d
    "01010101", --  208 - 0xd0  :   85 - 0x55 -- Background 0x1a
    "01000000", --  209 - 0xd1  :   64 - 0x40
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00000000", --  211 - 0xd3  :    0 - 0x0
    "00010000", --  212 - 0xd4  :   16 - 0x10
    "00010101", --  213 - 0xd5  :   21 - 0x15
    "01011010", --  214 - 0xd6  :   90 - 0x5a
    "01010101", --  215 - 0xd7  :   85 - 0x55
    "01010101", --  216 - 0xd8  :   85 - 0x55 -- Background 0x1b
    "01000000", --  217 - 0xd9  :   64 - 0x40
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00010101", --  220 - 0xdc  :   21 - 0x15
    "01010111", --  221 - 0xdd  :   87 - 0x57
    "01011010", --  222 - 0xde  :   90 - 0x5a
    "01011101", --  223 - 0xdf  :   93 - 0x5d
    "01011010", --  224 - 0xe0  :   90 - 0x5a -- Background 0x1c
    "01000000", --  225 - 0xe1  :   64 - 0x40
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00011010", --  228 - 0xe4  :   26 - 0x1a
    "01010111", --  229 - 0xe5  :   87 - 0x57
    "01010101", --  230 - 0xe6  :   85 - 0x55
    "01011101", --  231 - 0xe7  :   93 - 0x5d
    "01010101", --  232 - 0xe8  :   85 - 0x55 -- Background 0x1d
    "01000000", --  233 - 0xe9  :   64 - 0x40
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00010100", --  236 - 0xec  :   20 - 0x14
    "00000011", --  237 - 0xed  :    3 - 0x3
    "00001000", --  238 - 0xee  :    8 - 0x8
    "10101101", --  239 - 0xef  :  173 - 0xad
    "01010101", --  240 - 0xf0  :   85 - 0x55 -- Background 0x1e
    "01010000", --  241 - 0xf1  :   80 - 0x50
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "00010101", --  243 - 0xf3  :   21 - 0x15
    "01110101", --  244 - 0xf4  :  117 - 0x75
    "01010101", --  245 - 0xf5  :   85 - 0x55
    "01010111", --  246 - 0xf6  :   87 - 0x57
    "01010101", --  247 - 0xf7  :   85 - 0x55
    "01010101", --  248 - 0xf8  :   85 - 0x55 -- Background 0x1f
    "01010000", --  249 - 0xf9  :   80 - 0x50
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00010101", --  251 - 0xfb  :   21 - 0x15
    "01010111", --  252 - 0xfc  :   87 - 0x57
    "01010101", --  253 - 0xfd  :   85 - 0x55
    "01010101", --  254 - 0xfe  :   85 - 0x55
    "01010101", --  255 - 0xff  :   85 - 0x55
    "01010101", --  256 - 0x100  :   85 - 0x55 -- Background 0x20
    "11010000", --  257 - 0x101  :  208 - 0xd0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00010111", --  259 - 0x103  :   23 - 0x17
    "01010101", --  260 - 0x104  :   85 - 0x55
    "01010101", --  261 - 0x105  :   85 - 0x55
    "00000001", --  262 - 0x106  :    1 - 0x1
    "01010111", --  263 - 0x107  :   87 - 0x57
    "01010101", --  264 - 0x108  :   85 - 0x55 -- Background 0x21
    "01010000", --  265 - 0x109  :   80 - 0x50
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00010101", --  267 - 0x10b  :   21 - 0x15
    "01010101", --  268 - 0x10c  :   85 - 0x55
    "01110101", --  269 - 0x10d  :  117 - 0x75
    "01010101", --  270 - 0x10e  :   85 - 0x55
    "01010101", --  271 - 0x10f  :   85 - 0x55
    "01010101", --  272 - 0x110  :   85 - 0x55 -- Background 0x22
    "01010000", --  273 - 0x111  :   80 - 0x50
    "00000000", --  274 - 0x112  :    0 - 0x0
    "00010101", --  275 - 0x113  :   21 - 0x15
    "01110101", --  276 - 0x114  :  117 - 0x75
    "01010101", --  277 - 0x115  :   85 - 0x55
    "11010101", --  278 - 0x116  :  213 - 0xd5
    "01010101", --  279 - 0x117  :   85 - 0x55
    "01010101", --  280 - 0x118  :   85 - 0x55 -- Background 0x23
    "01010000", --  281 - 0x119  :   80 - 0x50
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00011001", --  283 - 0x11b  :   25 - 0x19
    "00001101", --  284 - 0x11c  :   13 - 0xd
    "00001000", --  285 - 0x11d  :    8 - 0x8
    "11110111", --  286 - 0x11e  :  247 - 0xf7
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "01010000", --  288 - 0x120  :   80 - 0x50 -- Background 0x24
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00011010", --  290 - 0x122  :   26 - 0x1a
    "10101001", --  291 - 0x123  :  169 - 0xa9
    "10101010", --  292 - 0x124  :  170 - 0xaa
    "10011001", --  293 - 0x125  :  153 - 0x99
    "01011001", --  294 - 0x126  :   89 - 0x59
    "10101010", --  295 - 0x127  :  170 - 0xaa
    "10010000", --  296 - 0x128  :  144 - 0x90 -- Background 0x25
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00010101", --  298 - 0x12a  :   21 - 0x15
    "01011001", --  299 - 0x12b  :   89 - 0x59
    "10010101", --  300 - 0x12c  :  149 - 0x95
    "10011001", --  301 - 0x12d  :  153 - 0x99
    "01011001", --  302 - 0x12e  :   89 - 0x59
    "10010101", --  303 - 0x12f  :  149 - 0x95
    "01010000", --  304 - 0x130  :   80 - 0x50 -- Background 0x26
    "00000000", --  305 - 0x131  :    0 - 0x0
    "00010000", --  306 - 0x132  :   16 - 0x10
    "00010101", --  307 - 0x133  :   21 - 0x15
    "01010101", --  308 - 0x134  :   85 - 0x55
    "01010101", --  309 - 0x135  :   85 - 0x55
    "01010101", --  310 - 0x136  :   85 - 0x55
    "01010101", --  311 - 0x137  :   85 - 0x55
    "01010000", --  312 - 0x138  :   80 - 0x50 -- Background 0x27
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00010101", --  314 - 0x13a  :   21 - 0x15
    "01011001", --  315 - 0x13b  :   89 - 0x59
    "10010101", --  316 - 0x13c  :  149 - 0x95
    "10011001", --  317 - 0x13d  :  153 - 0x99
    "01011001", --  318 - 0x13e  :   89 - 0x59
    "10010101", --  319 - 0x13f  :  149 - 0x95
    "10010000", --  320 - 0x140  :  144 - 0x90 -- Background 0x28
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00011010", --  322 - 0x142  :   26 - 0x1a
    "10101001", --  323 - 0x143  :  169 - 0xa9
    "10010101", --  324 - 0x144  :  149 - 0x95
    "10011010", --  325 - 0x145  :  154 - 0x9a
    "10101001", --  326 - 0x146  :  169 - 0xa9
    "10101010", --  327 - 0x147  :  170 - 0xaa
    "01010000", --  328 - 0x148  :   80 - 0x50 -- Background 0x29
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00011001", --  330 - 0x14a  :   25 - 0x19
    "00000011", --  331 - 0x14b  :    3 - 0x3
    "00001000", --  332 - 0x14c  :    8 - 0x8
    "10111110", --  333 - 0x14d  :  190 - 0xbe
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "10000110", --  335 - 0x14f  :  134 - 0x86
    "00000000", --  336 - 0x150  :    0 - 0x0 -- Background 0x2a
    "00010101", --  337 - 0x151  :   21 - 0x15
    "01010111", --  338 - 0x152  :   87 - 0x57
    "01101010", --  339 - 0x153  :  106 - 0x6a
    "01010110", --  340 - 0x154  :   86 - 0x56
    "10100111", --  341 - 0x155  :  167 - 0xa7
    "01010101", --  342 - 0x156  :   85 - 0x55
    "01010000", --  343 - 0x157  :   80 - 0x50
    "00000000", --  344 - 0x158  :    0 - 0x0 -- Background 0x2b
    "00010101", --  345 - 0x159  :   21 - 0x15
    "01010111", --  346 - 0x15a  :   87 - 0x57
    "01010101", --  347 - 0x15b  :   85 - 0x55
    "01110101", --  348 - 0x15c  :  117 - 0x75
    "01010111", --  349 - 0x15d  :   87 - 0x57
    "01010101", --  350 - 0x15e  :   85 - 0x55
    "01010000", --  351 - 0x15f  :   80 - 0x50
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Background 0x2c
    "00010000", --  353 - 0x161  :   16 - 0x10
    "00010101", --  354 - 0x162  :   21 - 0x15
    "01010101", --  355 - 0x163  :   85 - 0x55
    "01110101", --  356 - 0x164  :  117 - 0x75
    "01010101", --  357 - 0x165  :   85 - 0x55
    "01010101", --  358 - 0x166  :   85 - 0x55
    "01010000", --  359 - 0x167  :   80 - 0x50
    "00000000", --  360 - 0x168  :    0 - 0x0 -- Background 0x2d
    "00010101", --  361 - 0x169  :   21 - 0x15
    "01010111", --  362 - 0x16a  :   87 - 0x57
    "01010101", --  363 - 0x16b  :   85 - 0x55
    "01110101", --  364 - 0x16c  :  117 - 0x75
    "01010111", --  365 - 0x16d  :   87 - 0x57
    "01010101", --  366 - 0x16e  :   85 - 0x55
    "01010000", --  367 - 0x16f  :   80 - 0x50
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Background 0x2e
    "00010101", --  369 - 0x171  :   21 - 0x15
    "01010111", --  370 - 0x172  :   87 - 0x57
    "01101010", --  371 - 0x173  :  106 - 0x6a
    "01010110", --  372 - 0x174  :   86 - 0x56
    "10100111", --  373 - 0x175  :  167 - 0xa7
    "01010101", --  374 - 0x176  :   85 - 0x55
    "01010000", --  375 - 0x177  :   80 - 0x50
    "00000000", --  376 - 0x178  :    0 - 0x0 -- Background 0x2f
    "00011001", --  377 - 0x179  :   25 - 0x19
    "00000011", --  378 - 0x17a  :    3 - 0x3
    "00001000", --  379 - 0x17b  :    8 - 0x8
    "11011101", --  380 - 0x17c  :  221 - 0xdd
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "01110011", --  382 - 0x17e  :  115 - 0x73
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00011001", --  384 - 0x180  :   25 - 0x19 -- Background 0x30
    "01100101", --  385 - 0x181  :  101 - 0x65
    "10010110", --  386 - 0x182  :  150 - 0x96
    "10100101", --  387 - 0x183  :  165 - 0xa5
    "01011010", --  388 - 0x184  :   90 - 0x5a
    "10010110", --  389 - 0x185  :  150 - 0x96
    "01011001", --  390 - 0x186  :   89 - 0x59
    "01100100", --  391 - 0x187  :  100 - 0x64
    "00011001", --  392 - 0x188  :   25 - 0x19 -- Background 0x31
    "01100101", --  393 - 0x189  :  101 - 0x65
    "10010110", --  394 - 0x18a  :  150 - 0x96
    "10100101", --  395 - 0x18b  :  165 - 0xa5
    "01011010", --  396 - 0x18c  :   90 - 0x5a
    "10010110", --  397 - 0x18d  :  150 - 0x96
    "01011001", --  398 - 0x18e  :   89 - 0x59
    "01100100", --  399 - 0x18f  :  100 - 0x64
    "00011111", --  400 - 0x190  :   31 - 0x1f -- Background 0x32
    "01111101", --  401 - 0x191  :  125 - 0x7d
    "11010101", --  402 - 0x192  :  213 - 0xd5
    "01010000", --  403 - 0x193  :   80 - 0x50
    "00000101", --  404 - 0x194  :    5 - 0x5
    "01010111", --  405 - 0x195  :   87 - 0x57
    "11111111", --  406 - 0x196  :  255 - 0xff
    "01110100", --  407 - 0x197  :  116 - 0x74
    "00011001", --  408 - 0x198  :   25 - 0x19 -- Background 0x33
    "01100101", --  409 - 0x199  :  101 - 0x65
    "10010110", --  410 - 0x19a  :  150 - 0x96
    "10100101", --  411 - 0x19b  :  165 - 0xa5
    "01011010", --  412 - 0x19c  :   90 - 0x5a
    "10010110", --  413 - 0x19d  :  150 - 0x96
    "01011001", --  414 - 0x19e  :   89 - 0x59
    "01100100", --  415 - 0x19f  :  100 - 0x64
    "00011001", --  416 - 0x1a0  :   25 - 0x19 -- Background 0x34
    "01100101", --  417 - 0x1a1  :  101 - 0x65
    "10010110", --  418 - 0x1a2  :  150 - 0x96
    "10100101", --  419 - 0x1a3  :  165 - 0xa5
    "01011010", --  420 - 0x1a4  :   90 - 0x5a
    "10010110", --  421 - 0x1a5  :  150 - 0x96
    "01011001", --  422 - 0x1a6  :   89 - 0x59
    "01100100", --  423 - 0x1a7  :  100 - 0x64
    "00011110", --  424 - 0x1a8  :   30 - 0x1e -- Background 0x35
    "00001111", --  425 - 0x1a9  :   15 - 0xf
    "00001000", --  426 - 0x1aa  :    8 - 0x8
    "11110111", --  427 - 0x1ab  :  247 - 0xf7
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "01100111", --  429 - 0x1ad  :  103 - 0x67
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00010101", --  431 - 0x1af  :   21 - 0x15
    "01110101", --  432 - 0x1b0  :  117 - 0x75 -- Background 0x36
    "01010110", --  433 - 0x1b1  :   86 - 0x56
    "10100101", --  434 - 0x1b2  :  165 - 0xa5
    "01011010", --  435 - 0x1b3  :   90 - 0x5a
    "10010101", --  436 - 0x1b4  :  149 - 0x95
    "01011101", --  437 - 0x1b5  :   93 - 0x5d
    "11010100", --  438 - 0x1b6  :  212 - 0xd4
    "00010101", --  439 - 0x1b7  :   21 - 0x15
    "01010101", --  440 - 0x1b8  :   85 - 0x55 -- Background 0x37
    "01110101", --  441 - 0x1b9  :  117 - 0x75
    "01010101", --  442 - 0x1ba  :   85 - 0x55
    "01010101", --  443 - 0x1bb  :   85 - 0x55
    "01011101", --  444 - 0x1bc  :   93 - 0x5d
    "01010101", --  445 - 0x1bd  :   85 - 0x55
    "11010100", --  446 - 0x1be  :  212 - 0xd4
    "00010101", --  447 - 0x1bf  :   21 - 0x15
    "01101110", --  448 - 0x1c0  :  110 - 0x6e -- Background 0x38
    "01110101", --  449 - 0x1c1  :  117 - 0x75
    "01010000", --  450 - 0x1c2  :   80 - 0x50
    "00000101", --  451 - 0x1c3  :    5 - 0x5
    "01011101", --  452 - 0x1c4  :   93 - 0x5d
    "10111001", --  453 - 0x1c5  :  185 - 0xb9
    "01010100", --  454 - 0x1c6  :   84 - 0x54
    "00010101", --  455 - 0x1c7  :   21 - 0x15
    "01010101", --  456 - 0x1c8  :   85 - 0x55 -- Background 0x39
    "01110101", --  457 - 0x1c9  :  117 - 0x75
    "01010101", --  458 - 0x1ca  :   85 - 0x55
    "01010101", --  459 - 0x1cb  :   85 - 0x55
    "01011101", --  460 - 0x1cc  :   93 - 0x5d
    "01010101", --  461 - 0x1cd  :   85 - 0x55
    "11010100", --  462 - 0x1ce  :  212 - 0xd4
    "00010101", --  463 - 0x1cf  :   21 - 0x15
    "01110101", --  464 - 0x1d0  :  117 - 0x75 -- Background 0x3a
    "01010101", --  465 - 0x1d1  :   85 - 0x55
    "01101010", --  466 - 0x1d2  :  106 - 0x6a
    "10101001", --  467 - 0x1d3  :  169 - 0xa9
    "01010101", --  468 - 0x1d4  :   85 - 0x55
    "01011101", --  469 - 0x1d5  :   93 - 0x5d
    "11010100", --  470 - 0x1d6  :  212 - 0xd4
    "00010101", --  471 - 0x1d7  :   21 - 0x15
    "00001111", --  472 - 0x1d8  :   15 - 0xf -- Background 0x3b
    "00001000", --  473 - 0x1d9  :    8 - 0x8
    "11111000", --  474 - 0x1da  :  248 - 0xf8
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "01100111", --  476 - 0x1dc  :  103 - 0x67
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Background 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "00000000", --  485 - 0x1e5  :    0 - 0x0
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Background 0x3d
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Background 0x3e
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00000000", --  500 - 0x1f4  :    0 - 0x0
    "00000000", --  501 - 0x1f5  :    0 - 0x0
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- Background 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Background 0x40
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0 -- Background 0x41
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Background 0x42
    "00000000", --  529 - 0x211  :    0 - 0x0
    "00000000", --  530 - 0x212  :    0 - 0x0
    "00000000", --  531 - 0x213  :    0 - 0x0
    "00000000", --  532 - 0x214  :    0 - 0x0
    "00000000", --  533 - 0x215  :    0 - 0x0
    "00000000", --  534 - 0x216  :    0 - 0x0
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00000000", --  536 - 0x218  :    0 - 0x0 -- Background 0x43
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Background 0x44
    "00000000", --  545 - 0x221  :    0 - 0x0
    "00000000", --  546 - 0x222  :    0 - 0x0
    "00000000", --  547 - 0x223  :    0 - 0x0
    "00000000", --  548 - 0x224  :    0 - 0x0
    "00000000", --  549 - 0x225  :    0 - 0x0
    "00000000", --  550 - 0x226  :    0 - 0x0
    "00000000", --  551 - 0x227  :    0 - 0x0
    "00000000", --  552 - 0x228  :    0 - 0x0 -- Background 0x45
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000000", --  560 - 0x230  :    0 - 0x0 -- Background 0x46
    "00000000", --  561 - 0x231  :    0 - 0x0
    "00000000", --  562 - 0x232  :    0 - 0x0
    "00000000", --  563 - 0x233  :    0 - 0x0
    "00000000", --  564 - 0x234  :    0 - 0x0
    "00000000", --  565 - 0x235  :    0 - 0x0
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00000000", --  568 - 0x238  :    0 - 0x0 -- Background 0x47
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Background 0x48
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00000000", --  584 - 0x248  :    0 - 0x0 -- Background 0x49
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000000", --  592 - 0x250  :    0 - 0x0 -- Background 0x4a
    "00000000", --  593 - 0x251  :    0 - 0x0
    "00000000", --  594 - 0x252  :    0 - 0x0
    "00000000", --  595 - 0x253  :    0 - 0x0
    "00000000", --  596 - 0x254  :    0 - 0x0
    "00000000", --  597 - 0x255  :    0 - 0x0
    "00000000", --  598 - 0x256  :    0 - 0x0
    "00000000", --  599 - 0x257  :    0 - 0x0
    "00000000", --  600 - 0x258  :    0 - 0x0 -- Background 0x4b
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Background 0x4c
    "00000000", --  609 - 0x261  :    0 - 0x0
    "00000000", --  610 - 0x262  :    0 - 0x0
    "00000000", --  611 - 0x263  :    0 - 0x0
    "00000000", --  612 - 0x264  :    0 - 0x0
    "00000000", --  613 - 0x265  :    0 - 0x0
    "00000000", --  614 - 0x266  :    0 - 0x0
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0 -- Background 0x4d
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Background 0x4e
    "00000000", --  625 - 0x271  :    0 - 0x0
    "00000000", --  626 - 0x272  :    0 - 0x0
    "00000000", --  627 - 0x273  :    0 - 0x0
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000000", --  629 - 0x275  :    0 - 0x0
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0 -- Background 0x4f
    "00000000", --  633 - 0x279  :    0 - 0x0
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "00000000", --  635 - 0x27b  :    0 - 0x0
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Background 0x50
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Background 0x51
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Background 0x52
    "00000000", --  657 - 0x291  :    0 - 0x0
    "00000000", --  658 - 0x292  :    0 - 0x0
    "00000000", --  659 - 0x293  :    0 - 0x0
    "00000000", --  660 - 0x294  :    0 - 0x0
    "00000000", --  661 - 0x295  :    0 - 0x0
    "00000000", --  662 - 0x296  :    0 - 0x0
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Background 0x53
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Background 0x54
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "00000000", --  674 - 0x2a2  :    0 - 0x0
    "00000000", --  675 - 0x2a3  :    0 - 0x0
    "00000000", --  676 - 0x2a4  :    0 - 0x0
    "00000000", --  677 - 0x2a5  :    0 - 0x0
    "00000000", --  678 - 0x2a6  :    0 - 0x0
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- Background 0x55
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "00000000", --  686 - 0x2ae  :    0 - 0x0
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "00000000", --  688 - 0x2b0  :    0 - 0x0 -- Background 0x56
    "00000000", --  689 - 0x2b1  :    0 - 0x0
    "00000000", --  690 - 0x2b2  :    0 - 0x0
    "00000000", --  691 - 0x2b3  :    0 - 0x0
    "00000000", --  692 - 0x2b4  :    0 - 0x0
    "00000000", --  693 - 0x2b5  :    0 - 0x0
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "00000000", --  696 - 0x2b8  :    0 - 0x0 -- Background 0x57
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Background 0x58
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "00000000", --  707 - 0x2c3  :    0 - 0x0
    "00000000", --  708 - 0x2c4  :    0 - 0x0
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0 -- Background 0x59
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Background 0x5a
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Background 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Background 0x5c
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- Background 0x5d
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Background 0x5e
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00000000", --  754 - 0x2f2  :    0 - 0x0
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "00000000", --  756 - 0x2f4  :    0 - 0x0
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- Background 0x5f
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "00000000", --  764 - 0x2fc  :    0 - 0x0
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Background 0x60
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00000000", --  770 - 0x302  :    0 - 0x0
    "00000000", --  771 - 0x303  :    0 - 0x0
    "00000000", --  772 - 0x304  :    0 - 0x0
    "00000000", --  773 - 0x305  :    0 - 0x0
    "00000000", --  774 - 0x306  :    0 - 0x0
    "00000000", --  775 - 0x307  :    0 - 0x0
    "00000000", --  776 - 0x308  :    0 - 0x0 -- Background 0x61
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000000", --  779 - 0x30b  :    0 - 0x0
    "00000000", --  780 - 0x30c  :    0 - 0x0
    "00000000", --  781 - 0x30d  :    0 - 0x0
    "00000000", --  782 - 0x30e  :    0 - 0x0
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Background 0x62
    "00000000", --  785 - 0x311  :    0 - 0x0
    "00000000", --  786 - 0x312  :    0 - 0x0
    "00000000", --  787 - 0x313  :    0 - 0x0
    "00000000", --  788 - 0x314  :    0 - 0x0
    "00000000", --  789 - 0x315  :    0 - 0x0
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0 -- Background 0x63
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Background 0x64
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "00000000", --  804 - 0x324  :    0 - 0x0
    "00000000", --  805 - 0x325  :    0 - 0x0
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0 -- Background 0x65
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "00000000", --  813 - 0x32d  :    0 - 0x0
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Background 0x66
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000000", --  818 - 0x332  :    0 - 0x0
    "00000000", --  819 - 0x333  :    0 - 0x0
    "00000000", --  820 - 0x334  :    0 - 0x0
    "00000000", --  821 - 0x335  :    0 - 0x0
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000000", --  824 - 0x338  :    0 - 0x0 -- Background 0x67
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Background 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Background 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Background 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0 -- Background 0x6b
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Background 0x6c
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "00000000", --  868 - 0x364  :    0 - 0x0
    "00000000", --  869 - 0x365  :    0 - 0x0
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Background 0x6d
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Background 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00000000", --  888 - 0x378  :    0 - 0x0 -- Background 0x6f
    "00000000", --  889 - 0x379  :    0 - 0x0
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Background 0x70
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0 -- Background 0x71
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Background 0x72
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0 -- Background 0x73
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Background 0x74
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- Background 0x75
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Background 0x76
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- Background 0x77
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Background 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Background 0x79
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Background 0x7a
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Background 0x7b
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Background 0x7c
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Background 0x7d
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- Background 0x7f
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "10111111", -- 1024 - 0x400  :  191 - 0xbf -- Background 0x80
    "11110111", -- 1025 - 0x401  :  247 - 0xf7
    "11111101", -- 1026 - 0x402  :  253 - 0xfd
    "11011111", -- 1027 - 0x403  :  223 - 0xdf
    "11111011", -- 1028 - 0x404  :  251 - 0xfb
    "10111111", -- 1029 - 0x405  :  191 - 0xbf
    "11111110", -- 1030 - 0x406  :  254 - 0xfe
    "11101111", -- 1031 - 0x407  :  239 - 0xef
    "11111111", -- 1032 - 0x408  :  255 - 0xff -- Background 0x81
    "11101110", -- 1033 - 0x409  :  238 - 0xee
    "11111111", -- 1034 - 0x40a  :  255 - 0xff
    "11011111", -- 1035 - 0x40b  :  223 - 0xdf
    "01110111", -- 1036 - 0x40c  :  119 - 0x77
    "11111101", -- 1037 - 0x40d  :  253 - 0xfd
    "11011111", -- 1038 - 0x40e  :  223 - 0xdf
    "10111111", -- 1039 - 0x40f  :  191 - 0xbf
    "11111110", -- 1040 - 0x410  :  254 - 0xfe -- Background 0x82
    "11101111", -- 1041 - 0x411  :  239 - 0xef
    "10111111", -- 1042 - 0x412  :  191 - 0xbf
    "11110111", -- 1043 - 0x413  :  247 - 0xf7
    "11111101", -- 1044 - 0x414  :  253 - 0xfd
    "11011111", -- 1045 - 0x415  :  223 - 0xdf
    "11111011", -- 1046 - 0x416  :  251 - 0xfb
    "10111111", -- 1047 - 0x417  :  191 - 0xbf
    "11101111", -- 1048 - 0x418  :  239 - 0xef -- Background 0x83
    "11111111", -- 1049 - 0x419  :  255 - 0xff
    "10111011", -- 1050 - 0x41a  :  187 - 0xbb
    "11111111", -- 1051 - 0x41b  :  255 - 0xff
    "11110111", -- 1052 - 0x41c  :  247 - 0xf7
    "11011101", -- 1053 - 0x41d  :  221 - 0xdd
    "01111111", -- 1054 - 0x41e  :  127 - 0x7f
    "11110111", -- 1055 - 0x41f  :  247 - 0xf7
    "11111111", -- 1056 - 0x420  :  255 - 0xff -- Background 0x84
    "11101110", -- 1057 - 0x421  :  238 - 0xee
    "11111011", -- 1058 - 0x422  :  251 - 0xfb
    "10111111", -- 1059 - 0x423  :  191 - 0xbf
    "01111111", -- 1060 - 0x424  :  127 - 0x7f
    "11101101", -- 1061 - 0x425  :  237 - 0xed
    "11111111", -- 1062 - 0x426  :  255 - 0xff
    "10111111", -- 1063 - 0x427  :  191 - 0xbf
    "11111111", -- 1064 - 0x428  :  255 - 0xff -- Background 0x85
    "10111111", -- 1065 - 0x429  :  191 - 0xbf
    "01111101", -- 1066 - 0x42a  :  125 - 0x7d
    "11110111", -- 1067 - 0x42b  :  247 - 0xf7
    "11011011", -- 1068 - 0x42c  :  219 - 0xdb
    "11111101", -- 1069 - 0x42d  :  253 - 0xfd
    "01111110", -- 1070 - 0x42e  :  126 - 0x7e
    "11111011", -- 1071 - 0x42f  :  251 - 0xfb
    "11111111", -- 1072 - 0x430  :  255 - 0xff -- Background 0x86
    "11110111", -- 1073 - 0x431  :  247 - 0xf7
    "11111111", -- 1074 - 0x432  :  255 - 0xff
    "11011101", -- 1075 - 0x433  :  221 - 0xdd
    "01111111", -- 1076 - 0x434  :  127 - 0x7f
    "11110111", -- 1077 - 0x435  :  247 - 0xf7
    "11101111", -- 1078 - 0x436  :  239 - 0xef
    "10111101", -- 1079 - 0x437  :  189 - 0xbd
    "01011111", -- 1080 - 0x438  :   95 - 0x5f -- Background 0x87
    "11111101", -- 1081 - 0x439  :  253 - 0xfd
    "11110110", -- 1082 - 0x43a  :  246 - 0xf6
    "01111111", -- 1083 - 0x43b  :  127 - 0x7f
    "10011111", -- 1084 - 0x43c  :  159 - 0x9f
    "11111110", -- 1085 - 0x43d  :  254 - 0xfe
    "11111111", -- 1086 - 0x43e  :  255 - 0xff
    "11101111", -- 1087 - 0x43f  :  239 - 0xef
    "11111111", -- 1088 - 0x440  :  255 - 0xff -- Background 0x88
    "10011111", -- 1089 - 0x441  :  159 - 0x9f
    "10111111", -- 1090 - 0x442  :  191 - 0xbf
    "11111111", -- 1091 - 0x443  :  255 - 0xff
    "11110011", -- 1092 - 0x444  :  243 - 0xf3
    "11110011", -- 1093 - 0x445  :  243 - 0xf3
    "11111111", -- 1094 - 0x446  :  255 - 0xff
    "11111111", -- 1095 - 0x447  :  255 - 0xff
    "11111111", -- 1096 - 0x448  :  255 - 0xff -- Background 0x89
    "10011111", -- 1097 - 0x449  :  159 - 0x9f
    "10111111", -- 1098 - 0x44a  :  191 - 0xbf
    "11110011", -- 1099 - 0x44b  :  243 - 0xf3
    "11110011", -- 1100 - 0x44c  :  243 - 0xf3
    "11111111", -- 1101 - 0x44d  :  255 - 0xff
    "11111111", -- 1102 - 0x44e  :  255 - 0xff
    "11111111", -- 1103 - 0x44f  :  255 - 0xff
    "10111111", -- 1104 - 0x450  :  191 - 0xbf -- Background 0x8a
    "11110111", -- 1105 - 0x451  :  247 - 0xf7
    "11111101", -- 1106 - 0x452  :  253 - 0xfd
    "11111111", -- 1107 - 0x453  :  255 - 0xff
    "11111011", -- 1108 - 0x454  :  251 - 0xfb
    "10111111", -- 1109 - 0x455  :  191 - 0xbf
    "11111110", -- 1110 - 0x456  :  254 - 0xfe
    "11101111", -- 1111 - 0x457  :  239 - 0xef
    "10111111", -- 1112 - 0x458  :  191 - 0xbf -- Background 0x8b
    "11111111", -- 1113 - 0x459  :  255 - 0xff
    "11101110", -- 1114 - 0x45a  :  238 - 0xee
    "11111111", -- 1115 - 0x45b  :  255 - 0xff
    "11011111", -- 1116 - 0x45c  :  223 - 0xdf
    "01111101", -- 1117 - 0x45d  :  125 - 0x7d
    "11111111", -- 1118 - 0x45e  :  255 - 0xff
    "11011111", -- 1119 - 0x45f  :  223 - 0xdf
    "11111111", -- 1120 - 0x460  :  255 - 0xff -- Background 0x8c
    "11111000", -- 1121 - 0x461  :  248 - 0xf8
    "11100010", -- 1122 - 0x462  :  226 - 0xe2
    "11010111", -- 1123 - 0x463  :  215 - 0xd7
    "11001111", -- 1124 - 0x464  :  207 - 0xcf
    "10011111", -- 1125 - 0x465  :  159 - 0x9f
    "10111110", -- 1126 - 0x466  :  190 - 0xbe
    "10011101", -- 1127 - 0x467  :  157 - 0x9d
    "11111111", -- 1128 - 0x468  :  255 - 0xff -- Background 0x8d
    "00011111", -- 1129 - 0x469  :   31 - 0x1f
    "10100111", -- 1130 - 0x46a  :  167 - 0xa7
    "11000011", -- 1131 - 0x46b  :  195 - 0xc3
    "11100011", -- 1132 - 0x46c  :  227 - 0xe3
    "01000001", -- 1133 - 0x46d  :   65 - 0x41
    "10100001", -- 1134 - 0x46e  :  161 - 0xa1
    "00000001", -- 1135 - 0x46f  :    1 - 0x1
    "10111110", -- 1136 - 0x470  :  190 - 0xbe -- Background 0x8e
    "11111111", -- 1137 - 0x471  :  255 - 0xff
    "11011111", -- 1138 - 0x472  :  223 - 0xdf
    "11111111", -- 1139 - 0x473  :  255 - 0xff
    "11101111", -- 1140 - 0x474  :  239 - 0xef
    "11111111", -- 1141 - 0x475  :  255 - 0xff
    "11110111", -- 1142 - 0x476  :  247 - 0xf7
    "11111111", -- 1143 - 0x477  :  255 - 0xff
    "01111101", -- 1144 - 0x478  :  125 - 0x7d -- Background 0x8f
    "11111111", -- 1145 - 0x479  :  255 - 0xff
    "11111011", -- 1146 - 0x47a  :  251 - 0xfb
    "11111111", -- 1147 - 0x47b  :  255 - 0xff
    "11110111", -- 1148 - 0x47c  :  247 - 0xf7
    "11111111", -- 1149 - 0x47d  :  255 - 0xff
    "11101111", -- 1150 - 0x47e  :  239 - 0xef
    "11111111", -- 1151 - 0x47f  :  255 - 0xff
    "10111110", -- 1152 - 0x480  :  190 - 0xbe -- Background 0x90
    "11110111", -- 1153 - 0x481  :  247 - 0xf7
    "11111111", -- 1154 - 0x482  :  255 - 0xff
    "11011111", -- 1155 - 0x483  :  223 - 0xdf
    "11111011", -- 1156 - 0x484  :  251 - 0xfb
    "11111110", -- 1157 - 0x485  :  254 - 0xfe
    "10111111", -- 1158 - 0x486  :  191 - 0xbf
    "11110111", -- 1159 - 0x487  :  247 - 0xf7
    "11101110", -- 1160 - 0x488  :  238 - 0xee -- Background 0x91
    "11111111", -- 1161 - 0x489  :  255 - 0xff
    "01111011", -- 1162 - 0x48a  :  123 - 0x7b
    "11111101", -- 1163 - 0x48b  :  253 - 0xfd
    "11101111", -- 1164 - 0x48c  :  239 - 0xef
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "10111101", -- 1166 - 0x48e  :  189 - 0xbd
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "11111011", -- 1168 - 0x490  :  251 - 0xfb -- Background 0x92
    "10111111", -- 1169 - 0x491  :  191 - 0xbf
    "11101111", -- 1170 - 0x492  :  239 - 0xef
    "11111101", -- 1171 - 0x493  :  253 - 0xfd
    "11111111", -- 1172 - 0x494  :  255 - 0xff
    "10111111", -- 1173 - 0x495  :  191 - 0xbf
    "11111011", -- 1174 - 0x496  :  251 - 0xfb
    "11011111", -- 1175 - 0x497  :  223 - 0xdf
    "10111101", -- 1176 - 0x498  :  189 - 0xbd -- Background 0x93
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "01110111", -- 1178 - 0x49a  :  119 - 0x77
    "11111110", -- 1179 - 0x49b  :  254 - 0xfe
    "11011111", -- 1180 - 0x49c  :  223 - 0xdf
    "11111011", -- 1181 - 0x49d  :  251 - 0xfb
    "11101111", -- 1182 - 0x49e  :  239 - 0xef
    "01111111", -- 1183 - 0x49f  :  127 - 0x7f
    "01111111", -- 1184 - 0x4a0  :  127 - 0x7f -- Background 0x94
    "11110111", -- 1185 - 0x4a1  :  247 - 0xf7
    "11011101", -- 1186 - 0x4a2  :  221 - 0xdd
    "01111011", -- 1187 - 0x4a3  :  123 - 0x7b
    "11111111", -- 1188 - 0x4a4  :  255 - 0xff
    "11101110", -- 1189 - 0x4a5  :  238 - 0xee
    "10111011", -- 1190 - 0x4a6  :  187 - 0xbb
    "11111101", -- 1191 - 0x4a7  :  253 - 0xfd
    "11010111", -- 1192 - 0x4a8  :  215 - 0xd7 -- Background 0x95
    "01111111", -- 1193 - 0x4a9  :  127 - 0x7f
    "11111101", -- 1194 - 0x4aa  :  253 - 0xfd
    "11101110", -- 1195 - 0x4ab  :  238 - 0xee
    "11110111", -- 1196 - 0x4ac  :  247 - 0xf7
    "10111011", -- 1197 - 0x4ad  :  187 - 0xbb
    "11101111", -- 1198 - 0x4ae  :  239 - 0xef
    "11110111", -- 1199 - 0x4af  :  247 - 0xf7
    "10111111", -- 1200 - 0x4b0  :  191 - 0xbf -- Background 0x96
    "11101110", -- 1201 - 0x4b1  :  238 - 0xee
    "11011011", -- 1202 - 0x4b2  :  219 - 0xdb
    "11111111", -- 1203 - 0x4b3  :  255 - 0xff
    "01110111", -- 1204 - 0x4b4  :  119 - 0x77
    "11011101", -- 1205 - 0x4b5  :  221 - 0xdd
    "11101111", -- 1206 - 0x4b6  :  239 - 0xef
    "11111011", -- 1207 - 0x4b7  :  251 - 0xfb
    "11111101", -- 1208 - 0x4b8  :  253 - 0xfd -- Background 0x97
    "11101110", -- 1209 - 0x4b9  :  238 - 0xee
    "11111011", -- 1210 - 0x4ba  :  251 - 0xfb
    "11111101", -- 1211 - 0x4bb  :  253 - 0xfd
    "11110101", -- 1212 - 0x4bc  :  245 - 0xf5
    "11011111", -- 1213 - 0x4bd  :  223 - 0xdf
    "01111111", -- 1214 - 0x4be  :  127 - 0x7f
    "10111011", -- 1215 - 0x4bf  :  187 - 0xbb
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Background 0x98
    "10011111", -- 1217 - 0x4c1  :  159 - 0x9f
    "10111111", -- 1218 - 0x4c2  :  191 - 0xbf
    "11110011", -- 1219 - 0x4c3  :  243 - 0xf3
    "11110011", -- 1220 - 0x4c4  :  243 - 0xf3
    "11111111", -- 1221 - 0x4c5  :  255 - 0xff
    "11111111", -- 1222 - 0x4c6  :  255 - 0xff
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "11111111", -- 1224 - 0x4c8  :  255 - 0xff -- Background 0x99
    "10011111", -- 1225 - 0x4c9  :  159 - 0x9f
    "10111111", -- 1226 - 0x4ca  :  191 - 0xbf
    "11111111", -- 1227 - 0x4cb  :  255 - 0xff
    "11110011", -- 1228 - 0x4cc  :  243 - 0xf3
    "11110011", -- 1229 - 0x4cd  :  243 - 0xf3
    "11111111", -- 1230 - 0x4ce  :  255 - 0xff
    "11111111", -- 1231 - 0x4cf  :  255 - 0xff
    "10111111", -- 1232 - 0x4d0  :  191 - 0xbf -- Background 0x9a
    "11110111", -- 1233 - 0x4d1  :  247 - 0xf7
    "11111111", -- 1234 - 0x4d2  :  255 - 0xff
    "11011111", -- 1235 - 0x4d3  :  223 - 0xdf
    "11111011", -- 1236 - 0x4d4  :  251 - 0xfb
    "11111111", -- 1237 - 0x4d5  :  255 - 0xff
    "10111111", -- 1238 - 0x4d6  :  191 - 0xbf
    "11110111", -- 1239 - 0x4d7  :  247 - 0xf7
    "11011111", -- 1240 - 0x4d8  :  223 - 0xdf -- Background 0x9b
    "11111111", -- 1241 - 0x4d9  :  255 - 0xff
    "01111011", -- 1242 - 0x4da  :  123 - 0x7b
    "11111111", -- 1243 - 0x4db  :  255 - 0xff
    "11101111", -- 1244 - 0x4dc  :  239 - 0xef
    "11111101", -- 1245 - 0x4dd  :  253 - 0xfd
    "10111111", -- 1246 - 0x4de  :  191 - 0xbf
    "11111111", -- 1247 - 0x4df  :  255 - 0xff
    "10111010", -- 1248 - 0x4e0  :  186 - 0xba -- Background 0x9c
    "10011100", -- 1249 - 0x4e1  :  156 - 0x9c
    "10101010", -- 1250 - 0x4e2  :  170 - 0xaa
    "11000000", -- 1251 - 0x4e3  :  192 - 0xc0
    "11000000", -- 1252 - 0x4e4  :  192 - 0xc0
    "11100000", -- 1253 - 0x4e5  :  224 - 0xe0
    "11111000", -- 1254 - 0x4e6  :  248 - 0xf8
    "11111111", -- 1255 - 0x4e7  :  255 - 0xff
    "00000001", -- 1256 - 0x4e8  :    1 - 0x1 -- Background 0x9d
    "00000001", -- 1257 - 0x4e9  :    1 - 0x1
    "00000001", -- 1258 - 0x4ea  :    1 - 0x1
    "00000011", -- 1259 - 0x4eb  :    3 - 0x3
    "00000011", -- 1260 - 0x4ec  :    3 - 0x3
    "00000111", -- 1261 - 0x4ed  :    7 - 0x7
    "00011111", -- 1262 - 0x4ee  :   31 - 0x1f
    "11111111", -- 1263 - 0x4ef  :  255 - 0xff
    "01111101", -- 1264 - 0x4f0  :  125 - 0x7d -- Background 0x9e
    "11111111", -- 1265 - 0x4f1  :  255 - 0xff
    "11111011", -- 1266 - 0x4f2  :  251 - 0xfb
    "11111111", -- 1267 - 0x4f3  :  255 - 0xff
    "11111111", -- 1268 - 0x4f4  :  255 - 0xff
    "11111011", -- 1269 - 0x4f5  :  251 - 0xfb
    "11111111", -- 1270 - 0x4f6  :  255 - 0xff
    "01111101", -- 1271 - 0x4f7  :  125 - 0x7d
    "11111111", -- 1272 - 0x4f8  :  255 - 0xff -- Background 0x9f
    "11111111", -- 1273 - 0x4f9  :  255 - 0xff
    "10111101", -- 1274 - 0x4fa  :  189 - 0xbd
    "11111111", -- 1275 - 0x4fb  :  255 - 0xff
    "11111111", -- 1276 - 0x4fc  :  255 - 0xff
    "11111111", -- 1277 - 0x4fd  :  255 - 0xff
    "11111111", -- 1278 - 0x4fe  :  255 - 0xff
    "10111101", -- 1279 - 0x4ff  :  189 - 0xbd
    "11101111", -- 1280 - 0x500  :  239 - 0xef -- Background 0xa0
    "11000111", -- 1281 - 0x501  :  199 - 0xc7
    "10000011", -- 1282 - 0x502  :  131 - 0x83
    "00000111", -- 1283 - 0x503  :    7 - 0x7
    "10001111", -- 1284 - 0x504  :  143 - 0x8f
    "11011101", -- 1285 - 0x505  :  221 - 0xdd
    "11111010", -- 1286 - 0x506  :  250 - 0xfa
    "11111101", -- 1287 - 0x507  :  253 - 0xfd
    "11101111", -- 1288 - 0x508  :  239 - 0xef -- Background 0xa1
    "11000111", -- 1289 - 0x509  :  199 - 0xc7
    "10000011", -- 1290 - 0x50a  :  131 - 0x83
    "00011111", -- 1291 - 0x50b  :   31 - 0x1f
    "10010000", -- 1292 - 0x50c  :  144 - 0x90
    "11010100", -- 1293 - 0x50d  :  212 - 0xd4
    "11110011", -- 1294 - 0x50e  :  243 - 0xf3
    "11110010", -- 1295 - 0x50f  :  242 - 0xf2
    "11101111", -- 1296 - 0x510  :  239 - 0xef -- Background 0xa2
    "11000111", -- 1297 - 0x511  :  199 - 0xc7
    "10000011", -- 1298 - 0x512  :  131 - 0x83
    "11111111", -- 1299 - 0x513  :  255 - 0xff
    "00000000", -- 1300 - 0x514  :    0 - 0x0
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "01010101", -- 1302 - 0x516  :   85 - 0x55
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "11110000", -- 1304 - 0x518  :  240 - 0xf0 -- Background 0xa3
    "11010010", -- 1305 - 0x519  :  210 - 0xd2
    "10010000", -- 1306 - 0x51a  :  144 - 0x90
    "00010010", -- 1307 - 0x51b  :   18 - 0x12
    "10010000", -- 1308 - 0x51c  :  144 - 0x90
    "11010010", -- 1309 - 0x51d  :  210 - 0xd2
    "11110000", -- 1310 - 0x51e  :  240 - 0xf0
    "11110010", -- 1311 - 0x51f  :  242 - 0xf2
    "11110000", -- 1312 - 0x520  :  240 - 0xf0 -- Background 0xa4
    "11010011", -- 1313 - 0x521  :  211 - 0xd3
    "10010100", -- 1314 - 0x522  :  148 - 0x94
    "00011000", -- 1315 - 0x523  :   24 - 0x18
    "10011111", -- 1316 - 0x524  :  159 - 0x9f
    "11011101", -- 1317 - 0x525  :  221 - 0xdd
    "11111010", -- 1318 - 0x526  :  250 - 0xfa
    "11111101", -- 1319 - 0x527  :  253 - 0xfd
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- Background 0xa5
    "11111111", -- 1321 - 0x529  :  255 - 0xff
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "11111111", -- 1324 - 0x52c  :  255 - 0xff
    "11011101", -- 1325 - 0x52d  :  221 - 0xdd
    "11111010", -- 1326 - 0x52e  :  250 - 0xfa
    "11111101", -- 1327 - 0x52f  :  253 - 0xfd
    "11101111", -- 1328 - 0x530  :  239 - 0xef -- Background 0xa6
    "11000111", -- 1329 - 0x531  :  199 - 0xc7
    "10000011", -- 1330 - 0x532  :  131 - 0x83
    "11111111", -- 1331 - 0x533  :  255 - 0xff
    "00011111", -- 1332 - 0x534  :   31 - 0x1f
    "00101101", -- 1333 - 0x535  :   45 - 0x2d
    "01001010", -- 1334 - 0x536  :   74 - 0x4a
    "01001101", -- 1335 - 0x537  :   77 - 0x4d
    "01001111", -- 1336 - 0x538  :   79 - 0x4f -- Background 0xa7
    "01001111", -- 1337 - 0x539  :   79 - 0x4f
    "01001011", -- 1338 - 0x53a  :   75 - 0x4b
    "01001111", -- 1339 - 0x53b  :   79 - 0x4f
    "01001111", -- 1340 - 0x53c  :   79 - 0x4f
    "01001101", -- 1341 - 0x53d  :   77 - 0x4d
    "01001010", -- 1342 - 0x53e  :   74 - 0x4a
    "01001101", -- 1343 - 0x53f  :   77 - 0x4d
    "01001111", -- 1344 - 0x540  :   79 - 0x4f -- Background 0xa8
    "11001111", -- 1345 - 0x541  :  207 - 0xcf
    "00001011", -- 1346 - 0x542  :   11 - 0xb
    "00001111", -- 1347 - 0x543  :   15 - 0xf
    "11111111", -- 1348 - 0x544  :  255 - 0xff
    "11011101", -- 1349 - 0x545  :  221 - 0xdd
    "11111010", -- 1350 - 0x546  :  250 - 0xfa
    "11111101", -- 1351 - 0x547  :  253 - 0xfd
    "11111111", -- 1352 - 0x548  :  255 - 0xff -- Background 0xa9
    "11111111", -- 1353 - 0x549  :  255 - 0xff
    "11111111", -- 1354 - 0x54a  :  255 - 0xff
    "11111111", -- 1355 - 0x54b  :  255 - 0xff
    "11111111", -- 1356 - 0x54c  :  255 - 0xff
    "11111111", -- 1357 - 0x54d  :  255 - 0xff
    "11111111", -- 1358 - 0x54e  :  255 - 0xff
    "11111111", -- 1359 - 0x54f  :  255 - 0xff
    "11111111", -- 1360 - 0x550  :  255 - 0xff -- Background 0xaa
    "11111111", -- 1361 - 0x551  :  255 - 0xff
    "10101111", -- 1362 - 0x552  :  175 - 0xaf
    "01010111", -- 1363 - 0x553  :   87 - 0x57
    "10001111", -- 1364 - 0x554  :  143 - 0x8f
    "11011101", -- 1365 - 0x555  :  221 - 0xdd
    "11111010", -- 1366 - 0x556  :  250 - 0xfa
    "11111101", -- 1367 - 0x557  :  253 - 0xfd
    "11111111", -- 1368 - 0x558  :  255 - 0xff -- Background 0xab
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Background 0xac
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "00000000", -- 1380 - 0x564  :    0 - 0x0
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0 -- Background 0xad
    "11111111", -- 1385 - 0x569  :  255 - 0xff
    "00000000", -- 1386 - 0x56a  :    0 - 0x0
    "11111111", -- 1387 - 0x56b  :  255 - 0xff
    "11111111", -- 1388 - 0x56c  :  255 - 0xff
    "11111111", -- 1389 - 0x56d  :  255 - 0xff
    "11111111", -- 1390 - 0x56e  :  255 - 0xff
    "11111111", -- 1391 - 0x56f  :  255 - 0xff
    "11111111", -- 1392 - 0x570  :  255 - 0xff -- Background 0xae
    "11111111", -- 1393 - 0x571  :  255 - 0xff
    "11111111", -- 1394 - 0x572  :  255 - 0xff
    "11111111", -- 1395 - 0x573  :  255 - 0xff
    "11111111", -- 1396 - 0x574  :  255 - 0xff
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "11111111", -- 1398 - 0x576  :  255 - 0xff
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "11111111", -- 1400 - 0x578  :  255 - 0xff -- Background 0xaf
    "11111111", -- 1401 - 0x579  :  255 - 0xff
    "11111111", -- 1402 - 0x57a  :  255 - 0xff
    "11111111", -- 1403 - 0x57b  :  255 - 0xff
    "11111111", -- 1404 - 0x57c  :  255 - 0xff
    "11111111", -- 1405 - 0x57d  :  255 - 0xff
    "11111111", -- 1406 - 0x57e  :  255 - 0xff
    "11111111", -- 1407 - 0x57f  :  255 - 0xff
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Background 0xb0
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "00011111", -- 1410 - 0x582  :   31 - 0x1f
    "00010000", -- 1411 - 0x583  :   16 - 0x10
    "00010000", -- 1412 - 0x584  :   16 - 0x10
    "00010000", -- 1413 - 0x585  :   16 - 0x10
    "00010000", -- 1414 - 0x586  :   16 - 0x10
    "00010000", -- 1415 - 0x587  :   16 - 0x10
    "00000000", -- 1416 - 0x588  :    0 - 0x0 -- Background 0xb1
    "00000000", -- 1417 - 0x589  :    0 - 0x0
    "11111000", -- 1418 - 0x58a  :  248 - 0xf8
    "00001000", -- 1419 - 0x58b  :    8 - 0x8
    "00001000", -- 1420 - 0x58c  :    8 - 0x8
    "00001000", -- 1421 - 0x58d  :    8 - 0x8
    "00001000", -- 1422 - 0x58e  :    8 - 0x8
    "00001000", -- 1423 - 0x58f  :    8 - 0x8
    "00010000", -- 1424 - 0x590  :   16 - 0x10 -- Background 0xb2
    "00010000", -- 1425 - 0x591  :   16 - 0x10
    "00010000", -- 1426 - 0x592  :   16 - 0x10
    "00010000", -- 1427 - 0x593  :   16 - 0x10
    "00010000", -- 1428 - 0x594  :   16 - 0x10
    "00011111", -- 1429 - 0x595  :   31 - 0x1f
    "00011111", -- 1430 - 0x596  :   31 - 0x1f
    "00001111", -- 1431 - 0x597  :   15 - 0xf
    "00001000", -- 1432 - 0x598  :    8 - 0x8 -- Background 0xb3
    "00001000", -- 1433 - 0x599  :    8 - 0x8
    "00001000", -- 1434 - 0x59a  :    8 - 0x8
    "00001000", -- 1435 - 0x59b  :    8 - 0x8
    "00001000", -- 1436 - 0x59c  :    8 - 0x8
    "11111000", -- 1437 - 0x59d  :  248 - 0xf8
    "11111000", -- 1438 - 0x59e  :  248 - 0xf8
    "11110000", -- 1439 - 0x59f  :  240 - 0xf0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0 -- Background 0xb4
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "00000000", -- 1442 - 0x5a2  :    0 - 0x0
    "00111111", -- 1443 - 0x5a3  :   63 - 0x3f
    "01100000", -- 1444 - 0x5a4  :   96 - 0x60
    "01100000", -- 1445 - 0x5a5  :   96 - 0x60
    "01100000", -- 1446 - 0x5a6  :   96 - 0x60
    "01100000", -- 1447 - 0x5a7  :   96 - 0x60
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0 -- Background 0xb5
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "00000000", -- 1450 - 0x5aa  :    0 - 0x0
    "11111100", -- 1451 - 0x5ab  :  252 - 0xfc
    "00000110", -- 1452 - 0x5ac  :    6 - 0x6
    "00000110", -- 1453 - 0x5ad  :    6 - 0x6
    "00000110", -- 1454 - 0x5ae  :    6 - 0x6
    "00000110", -- 1455 - 0x5af  :    6 - 0x6
    "01100000", -- 1456 - 0x5b0  :   96 - 0x60 -- Background 0xb6
    "01100000", -- 1457 - 0x5b1  :   96 - 0x60
    "01100000", -- 1458 - 0x5b2  :   96 - 0x60
    "01100000", -- 1459 - 0x5b3  :   96 - 0x60
    "01111111", -- 1460 - 0x5b4  :  127 - 0x7f
    "01111111", -- 1461 - 0x5b5  :  127 - 0x7f
    "00111111", -- 1462 - 0x5b6  :   63 - 0x3f
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000110", -- 1464 - 0x5b8  :    6 - 0x6 -- Background 0xb7
    "00000110", -- 1465 - 0x5b9  :    6 - 0x6
    "00000110", -- 1466 - 0x5ba  :    6 - 0x6
    "00000110", -- 1467 - 0x5bb  :    6 - 0x6
    "11111110", -- 1468 - 0x5bc  :  254 - 0xfe
    "11111110", -- 1469 - 0x5bd  :  254 - 0xfe
    "11111100", -- 1470 - 0x5be  :  252 - 0xfc
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "01100000", -- 1472 - 0x5c0  :   96 - 0x60 -- Background 0xb8
    "11110000", -- 1473 - 0x5c1  :  240 - 0xf0
    "11000011", -- 1474 - 0x5c2  :  195 - 0xc3
    "10000111", -- 1475 - 0x5c3  :  135 - 0x87
    "00000110", -- 1476 - 0x5c4  :    6 - 0x6
    "00000100", -- 1477 - 0x5c5  :    4 - 0x4
    "00000100", -- 1478 - 0x5c6  :    4 - 0x4
    "00000111", -- 1479 - 0x5c7  :    7 - 0x7
    "00000110", -- 1480 - 0x5c8  :    6 - 0x6 -- Background 0xb9
    "00001111", -- 1481 - 0x5c9  :   15 - 0xf
    "10000111", -- 1482 - 0x5ca  :  135 - 0x87
    "11000001", -- 1483 - 0x5cb  :  193 - 0xc1
    "00100011", -- 1484 - 0x5cc  :   35 - 0x23
    "00101110", -- 1485 - 0x5cd  :   46 - 0x2e
    "01100000", -- 1486 - 0x5ce  :   96 - 0x60
    "11100001", -- 1487 - 0x5cf  :  225 - 0xe1
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Background 0xba
    "11001000", -- 1489 - 0x5d1  :  200 - 0xc8
    "11111000", -- 1490 - 0x5d2  :  248 - 0xf8
    "10110000", -- 1491 - 0x5d3  :  176 - 0xb0
    "00010000", -- 1492 - 0x5d4  :   16 - 0x10
    "00110000", -- 1493 - 0x5d5  :   48 - 0x30
    "11001000", -- 1494 - 0x5d6  :  200 - 0xc8
    "11111000", -- 1495 - 0x5d7  :  248 - 0xf8
    "00000111", -- 1496 - 0x5d8  :    7 - 0x7 -- Background 0xbb
    "00000011", -- 1497 - 0x5d9  :    3 - 0x3
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "01100000", -- 1499 - 0x5db  :   96 - 0x60
    "11110000", -- 1500 - 0x5dc  :  240 - 0xf0
    "11010000", -- 1501 - 0x5dd  :  208 - 0xd0
    "10010000", -- 1502 - 0x5de  :  144 - 0x90
    "01100000", -- 1503 - 0x5df  :   96 - 0x60
    "11100001", -- 1504 - 0x5e0  :  225 - 0xe1 -- Background 0xbc
    "11000011", -- 1505 - 0x5e1  :  195 - 0xc3
    "00001110", -- 1506 - 0x5e2  :   14 - 0xe
    "00000110", -- 1507 - 0x5e3  :    6 - 0x6
    "00001111", -- 1508 - 0x5e4  :   15 - 0xf
    "00001101", -- 1509 - 0x5e5  :   13 - 0xd
    "00001001", -- 1510 - 0x5e6  :    9 - 0x9
    "00000110", -- 1511 - 0x5e7  :    6 - 0x6
    "11100000", -- 1512 - 0x5e8  :  224 - 0xe0 -- Background 0xbd
    "01100000", -- 1513 - 0x5e9  :   96 - 0x60
    "11100011", -- 1514 - 0x5ea  :  227 - 0xe3
    "11100111", -- 1515 - 0x5eb  :  231 - 0xe7
    "00000110", -- 1516 - 0x5ec  :    6 - 0x6
    "00000100", -- 1517 - 0x5ed  :    4 - 0x4
    "00000100", -- 1518 - 0x5ee  :    4 - 0x4
    "00000111", -- 1519 - 0x5ef  :    7 - 0x7
    "00000111", -- 1520 - 0x5f0  :    7 - 0x7 -- Background 0xbe
    "00000011", -- 1521 - 0x5f1  :    3 - 0x3
    "10000111", -- 1522 - 0x5f2  :  135 - 0x87
    "11000111", -- 1523 - 0x5f3  :  199 - 0xc7
    "00100000", -- 1524 - 0x5f4  :   32 - 0x20
    "00100000", -- 1525 - 0x5f5  :   32 - 0x20
    "01100000", -- 1526 - 0x5f6  :   96 - 0x60
    "11100000", -- 1527 - 0x5f7  :  224 - 0xe0
    "00000111", -- 1528 - 0x5f8  :    7 - 0x7 -- Background 0xbf
    "00000011", -- 1529 - 0x5f9  :    3 - 0x3
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00001100", -- 1531 - 0x5fb  :   12 - 0xc
    "11101100", -- 1532 - 0x5fc  :  236 - 0xec
    "01100100", -- 1533 - 0x5fd  :  100 - 0x64
    "11101100", -- 1534 - 0x5fe  :  236 - 0xec
    "11101101", -- 1535 - 0x5ff  :  237 - 0xed
    "11100000", -- 1536 - 0x600  :  224 - 0xe0 -- Background 0xc0
    "11000000", -- 1537 - 0x601  :  192 - 0xc0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00110000", -- 1539 - 0x603  :   48 - 0x30
    "00110111", -- 1540 - 0x604  :   55 - 0x37
    "00010011", -- 1541 - 0x605  :   19 - 0x13
    "00110111", -- 1542 - 0x606  :   55 - 0x37
    "01110111", -- 1543 - 0x607  :  119 - 0x77
    "00001111", -- 1544 - 0x608  :   15 - 0xf -- Background 0xc1
    "00001100", -- 1545 - 0x609  :   12 - 0xc
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "11110000", -- 1552 - 0x610  :  240 - 0xf0 -- Background 0xc2
    "00110000", -- 1553 - 0x611  :   48 - 0x30
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- Background 0xc3
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000100", -- 1563 - 0x61b  :    4 - 0x4
    "00001101", -- 1564 - 0x61c  :   13 - 0xd
    "00001111", -- 1565 - 0x61d  :   15 - 0xf
    "00001100", -- 1566 - 0x61e  :   12 - 0xc
    "00001100", -- 1567 - 0x61f  :   12 - 0xc
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Background 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00010000", -- 1571 - 0x623  :   16 - 0x10
    "01110000", -- 1572 - 0x624  :  112 - 0x70
    "11110000", -- 1573 - 0x625  :  240 - 0xf0
    "00110000", -- 1574 - 0x626  :   48 - 0x30
    "00110000", -- 1575 - 0x627  :   48 - 0x30
    "11100100", -- 1576 - 0x628  :  228 - 0xe4 -- Background 0xc5
    "00100100", -- 1577 - 0x629  :   36 - 0x24
    "11100100", -- 1578 - 0x62a  :  228 - 0xe4
    "11101111", -- 1579 - 0x62b  :  239 - 0xef
    "00000111", -- 1580 - 0x62c  :    7 - 0x7
    "00000110", -- 1581 - 0x62d  :    6 - 0x6
    "00000100", -- 1582 - 0x62e  :    4 - 0x4
    "00000100", -- 1583 - 0x62f  :    4 - 0x4
    "00010111", -- 1584 - 0x630  :   23 - 0x17 -- Background 0xc6
    "00010001", -- 1585 - 0x631  :   17 - 0x11
    "00010111", -- 1586 - 0x632  :   23 - 0x17
    "10110111", -- 1587 - 0x633  :  183 - 0xb7
    "11000000", -- 1588 - 0x634  :  192 - 0xc0
    "00100000", -- 1589 - 0x635  :   32 - 0x20
    "00100000", -- 1590 - 0x636  :   32 - 0x20
    "01100000", -- 1591 - 0x637  :   96 - 0x60
    "00000111", -- 1592 - 0x638  :    7 - 0x7 -- Background 0xc7
    "00000111", -- 1593 - 0x639  :    7 - 0x7
    "00000011", -- 1594 - 0x63a  :    3 - 0x3
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "11100000", -- 1596 - 0x63c  :  224 - 0xe0
    "00100000", -- 1597 - 0x63d  :   32 - 0x20
    "11100000", -- 1598 - 0x63e  :  224 - 0xe0
    "11100000", -- 1599 - 0x63f  :  224 - 0xe0
    "11100000", -- 1600 - 0x640  :  224 - 0xe0 -- Background 0xc8
    "11100000", -- 1601 - 0x641  :  224 - 0xe0
    "11000000", -- 1602 - 0x642  :  192 - 0xc0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000111", -- 1604 - 0x644  :    7 - 0x7
    "00000001", -- 1605 - 0x645  :    1 - 0x1
    "00000111", -- 1606 - 0x646  :    7 - 0x7
    "00000111", -- 1607 - 0x647  :    7 - 0x7
    "00000001", -- 1608 - 0x648  :    1 - 0x1 -- Background 0xc9
    "00010011", -- 1609 - 0x649  :   19 - 0x13
    "00011111", -- 1610 - 0x64a  :   31 - 0x1f
    "00001101", -- 1611 - 0x64b  :   13 - 0xd
    "00000100", -- 1612 - 0x64c  :    4 - 0x4
    "00001100", -- 1613 - 0x64d  :   12 - 0xc
    "00010011", -- 1614 - 0x64e  :   19 - 0x13
    "00011111", -- 1615 - 0x64f  :   31 - 0x1f
    "01100000", -- 1616 - 0x650  :   96 - 0x60 -- Background 0xca
    "01110000", -- 1617 - 0x651  :  112 - 0x70
    "10100011", -- 1618 - 0x652  :  163 - 0xa3
    "10000111", -- 1619 - 0x653  :  135 - 0x87
    "11000110", -- 1620 - 0x654  :  198 - 0xc6
    "01110100", -- 1621 - 0x655  :  116 - 0x74
    "00000100", -- 1622 - 0x656  :    4 - 0x4
    "10000111", -- 1623 - 0x657  :  135 - 0x87
    "00000110", -- 1624 - 0x658  :    6 - 0x6 -- Background 0xcb
    "00001111", -- 1625 - 0x659  :   15 - 0xf
    "10000011", -- 1626 - 0x65a  :  131 - 0x83
    "11000001", -- 1627 - 0x65b  :  193 - 0xc1
    "00100000", -- 1628 - 0x65c  :   32 - 0x20
    "00100000", -- 1629 - 0x65d  :   32 - 0x20
    "01100000", -- 1630 - 0x65e  :   96 - 0x60
    "11100000", -- 1631 - 0x65f  :  224 - 0xe0
    "10000111", -- 1632 - 0x660  :  135 - 0x87 -- Background 0xcc
    "01000011", -- 1633 - 0x661  :   67 - 0x43
    "00110000", -- 1634 - 0x662  :   48 - 0x30
    "01100000", -- 1635 - 0x663  :   96 - 0x60
    "11110000", -- 1636 - 0x664  :  240 - 0xf0
    "11010000", -- 1637 - 0x665  :  208 - 0xd0
    "10010000", -- 1638 - 0x666  :  144 - 0x90
    "01100000", -- 1639 - 0x667  :   96 - 0x60
    "11100000", -- 1640 - 0x668  :  224 - 0xe0 -- Background 0xcd
    "11000000", -- 1641 - 0x669  :  192 - 0xc0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000110", -- 1643 - 0x66b  :    6 - 0x6
    "00001111", -- 1644 - 0x66c  :   15 - 0xf
    "00001101", -- 1645 - 0x66d  :   13 - 0xd
    "00001001", -- 1646 - 0x66e  :    9 - 0x9
    "00000110", -- 1647 - 0x66f  :    6 - 0x6
    "11111100", -- 1648 - 0x670  :  252 - 0xfc -- Background 0xce
    "11000000", -- 1649 - 0x671  :  192 - 0xc0
    "11010001", -- 1650 - 0x672  :  209 - 0xd1
    "11000010", -- 1651 - 0x673  :  194 - 0xc2
    "10011110", -- 1652 - 0x674  :  158 - 0x9e
    "10111111", -- 1653 - 0x675  :  191 - 0xbf
    "10110000", -- 1654 - 0x676  :  176 - 0xb0
    "10110011", -- 1655 - 0x677  :  179 - 0xb3
    "00000111", -- 1656 - 0x678  :    7 - 0x7 -- Background 0xcf
    "11110011", -- 1657 - 0x679  :  243 - 0xf3
    "00001011", -- 1658 - 0x67a  :   11 - 0xb
    "01111011", -- 1659 - 0x67b  :  123 - 0x7b
    "01111011", -- 1660 - 0x67c  :  123 - 0x7b
    "11111001", -- 1661 - 0x67d  :  249 - 0xf9
    "00001101", -- 1662 - 0x67e  :   13 - 0xd
    "11101101", -- 1663 - 0x67f  :  237 - 0xed
    "11111111", -- 1664 - 0x680  :  255 - 0xff -- Background 0xd0
    "11111111", -- 1665 - 0x681  :  255 - 0xff
    "11111111", -- 1666 - 0x682  :  255 - 0xff
    "11111111", -- 1667 - 0x683  :  255 - 0xff
    "11101110", -- 1668 - 0x684  :  238 - 0xee
    "11101110", -- 1669 - 0x685  :  238 - 0xee
    "11101110", -- 1670 - 0x686  :  238 - 0xee
    "11101110", -- 1671 - 0x687  :  238 - 0xee
    "11111111", -- 1672 - 0x688  :  255 - 0xff -- Background 0xd1
    "11111111", -- 1673 - 0x689  :  255 - 0xff
    "11111111", -- 1674 - 0x68a  :  255 - 0xff
    "11111011", -- 1675 - 0x68b  :  251 - 0xfb
    "11111011", -- 1676 - 0x68c  :  251 - 0xfb
    "11111011", -- 1677 - 0x68d  :  251 - 0xfb
    "11111011", -- 1678 - 0x68e  :  251 - 0xfb
    "11111011", -- 1679 - 0x68f  :  251 - 0xfb
    "11111111", -- 1680 - 0x690  :  255 - 0xff -- Background 0xd2
    "11111111", -- 1681 - 0x691  :  255 - 0xff
    "11111111", -- 1682 - 0x692  :  255 - 0xff
    "11111111", -- 1683 - 0x693  :  255 - 0xff
    "11101110", -- 1684 - 0x694  :  238 - 0xee
    "10001110", -- 1685 - 0x695  :  142 - 0x8e
    "11111110", -- 1686 - 0x696  :  254 - 0xfe
    "11111110", -- 1687 - 0x697  :  254 - 0xfe
    "11111111", -- 1688 - 0x698  :  255 - 0xff -- Background 0xd3
    "11111111", -- 1689 - 0x699  :  255 - 0xff
    "11111111", -- 1690 - 0x69a  :  255 - 0xff
    "11111111", -- 1691 - 0x69b  :  255 - 0xff
    "11101110", -- 1692 - 0x69c  :  238 - 0xee
    "10001110", -- 1693 - 0x69d  :  142 - 0x8e
    "11111100", -- 1694 - 0x69e  :  252 - 0xfc
    "11111101", -- 1695 - 0x69f  :  253 - 0xfd
    "11111111", -- 1696 - 0x6a0  :  255 - 0xff -- Background 0xd4
    "11111111", -- 1697 - 0x6a1  :  255 - 0xff
    "11111111", -- 1698 - 0x6a2  :  255 - 0xff
    "11111110", -- 1699 - 0x6a3  :  254 - 0xfe
    "11101110", -- 1700 - 0x6a4  :  238 - 0xee
    "11101110", -- 1701 - 0x6a5  :  238 - 0xee
    "11101110", -- 1702 - 0x6a6  :  238 - 0xee
    "11101110", -- 1703 - 0x6a7  :  238 - 0xee
    "11111111", -- 1704 - 0x6a8  :  255 - 0xff -- Background 0xd5
    "11111111", -- 1705 - 0x6a9  :  255 - 0xff
    "11111111", -- 1706 - 0x6aa  :  255 - 0xff
    "11111101", -- 1707 - 0x6ab  :  253 - 0xfd
    "11100001", -- 1708 - 0x6ac  :  225 - 0xe1
    "11101111", -- 1709 - 0x6ad  :  239 - 0xef
    "11111111", -- 1710 - 0x6ae  :  255 - 0xff
    "11111111", -- 1711 - 0x6af  :  255 - 0xff
    "11111111", -- 1712 - 0x6b0  :  255 - 0xff -- Background 0xd6
    "11111111", -- 1713 - 0x6b1  :  255 - 0xff
    "11111111", -- 1714 - 0x6b2  :  255 - 0xff
    "11111101", -- 1715 - 0x6b3  :  253 - 0xfd
    "11100001", -- 1716 - 0x6b4  :  225 - 0xe1
    "11101111", -- 1717 - 0x6b5  :  239 - 0xef
    "11111111", -- 1718 - 0x6b6  :  255 - 0xff
    "11111111", -- 1719 - 0x6b7  :  255 - 0xff
    "11111111", -- 1720 - 0x6b8  :  255 - 0xff -- Background 0xd7
    "11111111", -- 1721 - 0x6b9  :  255 - 0xff
    "11111111", -- 1722 - 0x6ba  :  255 - 0xff
    "11111110", -- 1723 - 0x6bb  :  254 - 0xfe
    "11101110", -- 1724 - 0x6bc  :  238 - 0xee
    "10001110", -- 1725 - 0x6bd  :  142 - 0x8e
    "11111110", -- 1726 - 0x6be  :  254 - 0xfe
    "11111100", -- 1727 - 0x6bf  :  252 - 0xfc
    "11111111", -- 1728 - 0x6c0  :  255 - 0xff -- Background 0xd8
    "11111111", -- 1729 - 0x6c1  :  255 - 0xff
    "11111111", -- 1730 - 0x6c2  :  255 - 0xff
    "11111111", -- 1731 - 0x6c3  :  255 - 0xff
    "11101110", -- 1732 - 0x6c4  :  238 - 0xee
    "11101110", -- 1733 - 0x6c5  :  238 - 0xee
    "11111100", -- 1734 - 0x6c6  :  252 - 0xfc
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "11111111", -- 1736 - 0x6c8  :  255 - 0xff -- Background 0xd9
    "11111111", -- 1737 - 0x6c9  :  255 - 0xff
    "11111111", -- 1738 - 0x6ca  :  255 - 0xff
    "11111111", -- 1739 - 0x6cb  :  255 - 0xff
    "11101110", -- 1740 - 0x6cc  :  238 - 0xee
    "11101110", -- 1741 - 0x6cd  :  238 - 0xee
    "11101110", -- 1742 - 0x6ce  :  238 - 0xee
    "11101110", -- 1743 - 0x6cf  :  238 - 0xee
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Background 0xda
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "10000000", -- 1747 - 0x6d3  :  128 - 0x80
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000100", -- 1750 - 0x6d6  :    4 - 0x4
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0 -- Background 0xdb
    "00000100", -- 1753 - 0x6d9  :    4 - 0x4
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "00010001", -- 1755 - 0x6db  :   17 - 0x11
    "00000000", -- 1756 - 0x6dc  :    0 - 0x0
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00100000", -- 1759 - 0x6df  :   32 - 0x20
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00100000", -- 1763 - 0x6e3  :   32 - 0x20
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000100", -- 1767 - 0x6e7  :    4 - 0x4
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- Background 0xdd
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00010001", -- 1770 - 0x6ea  :   17 - 0x11
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "10000000", -- 1773 - 0x6ed  :  128 - 0x80
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "10110011", -- 1776 - 0x6f0  :  179 - 0xb3 -- Background 0xde
    "10110011", -- 1777 - 0x6f1  :  179 - 0xb3
    "10110011", -- 1778 - 0x6f2  :  179 - 0xb3
    "10110011", -- 1779 - 0x6f3  :  179 - 0xb3
    "10110000", -- 1780 - 0x6f4  :  176 - 0xb0
    "10101111", -- 1781 - 0x6f5  :  175 - 0xaf
    "10011111", -- 1782 - 0x6f6  :  159 - 0x9f
    "11000000", -- 1783 - 0x6f7  :  192 - 0xc0
    "11101101", -- 1784 - 0x6f8  :  237 - 0xed -- Background 0xdf
    "11001101", -- 1785 - 0x6f9  :  205 - 0xcd
    "11001101", -- 1786 - 0x6fa  :  205 - 0xcd
    "00001101", -- 1787 - 0x6fb  :   13 - 0xd
    "00001101", -- 1788 - 0x6fc  :   13 - 0xd
    "11111101", -- 1789 - 0x6fd  :  253 - 0xfd
    "11111101", -- 1790 - 0x6fe  :  253 - 0xfd
    "00000011", -- 1791 - 0x6ff  :    3 - 0x3
    "11101110", -- 1792 - 0x700  :  238 - 0xee -- Background 0xe0
    "11101110", -- 1793 - 0x701  :  238 - 0xee
    "11101110", -- 1794 - 0x702  :  238 - 0xee
    "11101110", -- 1795 - 0x703  :  238 - 0xee
    "11111110", -- 1796 - 0x704  :  254 - 0xfe
    "11111100", -- 1797 - 0x705  :  252 - 0xfc
    "11000001", -- 1798 - 0x706  :  193 - 0xc1
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "11111011", -- 1800 - 0x708  :  251 - 0xfb -- Background 0xe1
    "11111011", -- 1801 - 0x709  :  251 - 0xfb
    "11111011", -- 1802 - 0x70a  :  251 - 0xfb
    "11111011", -- 1803 - 0x70b  :  251 - 0xfb
    "11111111", -- 1804 - 0x70c  :  255 - 0xff
    "11111101", -- 1805 - 0x70d  :  253 - 0xfd
    "11000001", -- 1806 - 0x70e  :  193 - 0xc1
    "11111111", -- 1807 - 0x70f  :  255 - 0xff
    "11111100", -- 1808 - 0x710  :  252 - 0xfc -- Background 0xe2
    "11100001", -- 1809 - 0x711  :  225 - 0xe1
    "11101111", -- 1810 - 0x712  :  239 - 0xef
    "11101111", -- 1811 - 0x713  :  239 - 0xef
    "11111111", -- 1812 - 0x714  :  255 - 0xff
    "11111110", -- 1813 - 0x715  :  254 - 0xfe
    "10000000", -- 1814 - 0x716  :  128 - 0x80
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "11101110", -- 1816 - 0x718  :  238 - 0xee -- Background 0xe3
    "11111110", -- 1817 - 0x719  :  254 - 0xfe
    "11111110", -- 1818 - 0x71a  :  254 - 0xfe
    "11111110", -- 1819 - 0x71b  :  254 - 0xfe
    "11111110", -- 1820 - 0x71c  :  254 - 0xfe
    "11111100", -- 1821 - 0x71d  :  252 - 0xfc
    "11000001", -- 1822 - 0x71e  :  193 - 0xc1
    "11111111", -- 1823 - 0x71f  :  255 - 0xff
    "11101110", -- 1824 - 0x720  :  238 - 0xee -- Background 0xe4
    "11101110", -- 1825 - 0x721  :  238 - 0xee
    "11111110", -- 1826 - 0x722  :  254 - 0xfe
    "11111110", -- 1827 - 0x723  :  254 - 0xfe
    "10001110", -- 1828 - 0x724  :  142 - 0x8e
    "11111110", -- 1829 - 0x725  :  254 - 0xfe
    "11111000", -- 1830 - 0x726  :  248 - 0xf8
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "10001110", -- 1832 - 0x728  :  142 - 0x8e -- Background 0xe5
    "11111110", -- 1833 - 0x729  :  254 - 0xfe
    "11111110", -- 1834 - 0x72a  :  254 - 0xfe
    "11111110", -- 1835 - 0x72b  :  254 - 0xfe
    "11111110", -- 1836 - 0x72c  :  254 - 0xfe
    "11111100", -- 1837 - 0x72d  :  252 - 0xfc
    "11000001", -- 1838 - 0x72e  :  193 - 0xc1
    "11111111", -- 1839 - 0x72f  :  255 - 0xff
    "11101110", -- 1840 - 0x730  :  238 - 0xee -- Background 0xe6
    "11101110", -- 1841 - 0x731  :  238 - 0xee
    "11101110", -- 1842 - 0x732  :  238 - 0xee
    "11101110", -- 1843 - 0x733  :  238 - 0xee
    "11111110", -- 1844 - 0x734  :  254 - 0xfe
    "11111100", -- 1845 - 0x735  :  252 - 0xfc
    "11000001", -- 1846 - 0x736  :  193 - 0xc1
    "11111111", -- 1847 - 0x737  :  255 - 0xff
    "11111101", -- 1848 - 0x738  :  253 - 0xfd -- Background 0xe7
    "11111101", -- 1849 - 0x739  :  253 - 0xfd
    "11111001", -- 1850 - 0x73a  :  249 - 0xf9
    "11111011", -- 1851 - 0x73b  :  251 - 0xfb
    "11111011", -- 1852 - 0x73c  :  251 - 0xfb
    "11111011", -- 1853 - 0x73d  :  251 - 0xfb
    "11100011", -- 1854 - 0x73e  :  227 - 0xe3
    "11111111", -- 1855 - 0x73f  :  255 - 0xff
    "11101110", -- 1856 - 0x740  :  238 - 0xee -- Background 0xe8
    "11101110", -- 1857 - 0x741  :  238 - 0xee
    "11101110", -- 1858 - 0x742  :  238 - 0xee
    "11101110", -- 1859 - 0x743  :  238 - 0xee
    "11111110", -- 1860 - 0x744  :  254 - 0xfe
    "11111100", -- 1861 - 0x745  :  252 - 0xfc
    "11000001", -- 1862 - 0x746  :  193 - 0xc1
    "11111111", -- 1863 - 0x747  :  255 - 0xff
    "11111110", -- 1864 - 0x748  :  254 - 0xfe -- Background 0xe9
    "11111110", -- 1865 - 0x749  :  254 - 0xfe
    "11001110", -- 1866 - 0x74a  :  206 - 0xce
    "11111110", -- 1867 - 0x74b  :  254 - 0xfe
    "11111110", -- 1868 - 0x74c  :  254 - 0xfe
    "11111100", -- 1869 - 0x74d  :  252 - 0xfc
    "11000001", -- 1870 - 0x74e  :  193 - 0xc1
    "11111111", -- 1871 - 0x74f  :  255 - 0xff
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Background 0xea
    "01110000", -- 1873 - 0x751  :  112 - 0x70
    "00111000", -- 1874 - 0x752  :   56 - 0x38
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000010", -- 1876 - 0x754  :    2 - 0x2
    "00000111", -- 1877 - 0x755  :    7 - 0x7
    "00000011", -- 1878 - 0x756  :    3 - 0x3
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- Background 0xeb
    "00001100", -- 1881 - 0x759  :   12 - 0xc
    "00000110", -- 1882 - 0x75a  :    6 - 0x6
    "00000110", -- 1883 - 0x75b  :    6 - 0x6
    "01100000", -- 1884 - 0x75c  :   96 - 0x60
    "01110000", -- 1885 - 0x75d  :  112 - 0x70
    "00110000", -- 1886 - 0x75e  :   48 - 0x30
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Background 0xec
    "11000000", -- 1889 - 0x761  :  192 - 0xc0
    "11100000", -- 1890 - 0x762  :  224 - 0xe0
    "01100000", -- 1891 - 0x763  :   96 - 0x60
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00001100", -- 1893 - 0x765  :   12 - 0xc
    "00001110", -- 1894 - 0x766  :   14 - 0xe
    "00000110", -- 1895 - 0x767  :    6 - 0x6
    "01100000", -- 1896 - 0x768  :   96 - 0x60 -- Background 0xed
    "01110000", -- 1897 - 0x769  :  112 - 0x70
    "00110000", -- 1898 - 0x76a  :   48 - 0x30
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00001100", -- 1901 - 0x76d  :   12 - 0xc
    "00001110", -- 1902 - 0x76e  :   14 - 0xe
    "00000110", -- 1903 - 0x76f  :    6 - 0x6
    "11111111", -- 1904 - 0x770  :  255 - 0xff -- Background 0xee
    "11111111", -- 1905 - 0x771  :  255 - 0xff
    "10111101", -- 1906 - 0x772  :  189 - 0xbd
    "11111111", -- 1907 - 0x773  :  255 - 0xff
    "11111111", -- 1908 - 0x774  :  255 - 0xff
    "11111011", -- 1909 - 0x775  :  251 - 0xfb
    "11111111", -- 1910 - 0x776  :  255 - 0xff
    "11111111", -- 1911 - 0x777  :  255 - 0xff
    "11111111", -- 1912 - 0x778  :  255 - 0xff -- Background 0xef
    "11111111", -- 1913 - 0x779  :  255 - 0xff
    "11111011", -- 1914 - 0x77a  :  251 - 0xfb
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "11011111", -- 1916 - 0x77c  :  223 - 0xdf
    "11111111", -- 1917 - 0x77d  :  255 - 0xff
    "11111111", -- 1918 - 0x77e  :  255 - 0xff
    "11111111", -- 1919 - 0x77f  :  255 - 0xff
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- Background 0xf1
    "10000000", -- 1929 - 0x789  :  128 - 0x80
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Background 0xf2
    "11000000", -- 1937 - 0x791  :  192 - 0xc0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- Background 0xf3
    "11100000", -- 1945 - 0x799  :  224 - 0xe0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Background 0xf4
    "11110000", -- 1953 - 0x7a1  :  240 - 0xf0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0 -- Background 0xf5
    "11111000", -- 1961 - 0x7a9  :  248 - 0xf8
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Background 0xf6
    "11111100", -- 1969 - 0x7b1  :  252 - 0xfc
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- Background 0xf7
    "11111110", -- 1977 - 0x7b9  :  254 - 0xfe
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Background 0xf8
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "11111111", -- 1992 - 0x7c8  :  255 - 0xff -- Background 0xf9
    "11111111", -- 1993 - 0x7c9  :  255 - 0xff
    "11111111", -- 1994 - 0x7ca  :  255 - 0xff
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "10000000", -- 1996 - 0x7cc  :  128 - 0x80
    "10000000", -- 1997 - 0x7cd  :  128 - 0x80
    "11000000", -- 1998 - 0x7ce  :  192 - 0xc0
    "11000000", -- 1999 - 0x7cf  :  192 - 0xc0
    "11111111", -- 2000 - 0x7d0  :  255 - 0xff -- Background 0xfa
    "11111111", -- 2001 - 0x7d1  :  255 - 0xff
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "11111111", -- 2008 - 0x7d8  :  255 - 0xff -- Background 0xfb
    "11111111", -- 2009 - 0x7d9  :  255 - 0xff
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111111", -- 2011 - 0x7db  :  255 - 0xff
    "00000001", -- 2012 - 0x7dc  :    1 - 0x1
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000010", -- 2014 - 0x7de  :    2 - 0x2
    "00000010", -- 2015 - 0x7df  :    2 - 0x2
    "11000000", -- 2016 - 0x7e0  :  192 - 0xc0 -- Background 0xfc
    "11000000", -- 2017 - 0x7e1  :  192 - 0xc0
    "10000000", -- 2018 - 0x7e2  :  128 - 0x80
    "10000000", -- 2019 - 0x7e3  :  128 - 0x80
    "11000000", -- 2020 - 0x7e4  :  192 - 0xc0
    "11111111", -- 2021 - 0x7e5  :  255 - 0xff
    "11111111", -- 2022 - 0x7e6  :  255 - 0xff
    "11111111", -- 2023 - 0x7e7  :  255 - 0xff
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- Background 0xfd
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "11111111", -- 2029 - 0x7ed  :  255 - 0xff
    "11111111", -- 2030 - 0x7ee  :  255 - 0xff
    "11111111", -- 2031 - 0x7ef  :  255 - 0xff
    "00000010", -- 2032 - 0x7f0  :    2 - 0x2 -- Background 0xfe
    "00000010", -- 2033 - 0x7f1  :    2 - 0x2
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "11111111", -- 2037 - 0x7f5  :  255 - 0xff
    "11111111", -- 2038 - 0x7f6  :  255 - 0xff
    "11111111", -- 2039 - 0x7f7  :  255 - 0xff
    "11111111", -- 2040 - 0x7f8  :  255 - 0xff -- Background 0xff
    "11111111", -- 2041 - 0x7f9  :  255 - 0xff
    "11111111", -- 2042 - 0x7fa  :  255 - 0xff
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111111", -- 2044 - 0x7fc  :  255 - 0xff
    "11111111", -- 2045 - 0x7fd  :  255 - 0xff
    "11111111", -- 2046 - 0x7fe  :  255 - 0xff
    "11111111"  -- 2047 - 0x7ff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
