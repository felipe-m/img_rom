//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables
//- Only the first Name Table: 1KiB


//-  Original memory dump file name: lawnmower_ntable_start.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_NTABLE0_LAWN_START
  (
     input     clk,   // clock
     input      [10-1:0] addr,  //1024 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      10'h0: dout <= 8'b10000100; //    0 : 132 - 0x84 -- line 0x0
      10'h1: dout <= 8'b10000101; //    1 : 133 - 0x85
      10'h2: dout <= 8'b10000100; //    2 : 132 - 0x84
      10'h3: dout <= 8'b10000101; //    3 : 133 - 0x85
      10'h4: dout <= 8'b10000111; //    4 : 135 - 0x87
      10'h5: dout <= 8'b10000101; //    5 : 133 - 0x85
      10'h6: dout <= 8'b10000100; //    6 : 132 - 0x84
      10'h7: dout <= 8'b10000111; //    7 : 135 - 0x87
      10'h8: dout <= 8'b10000100; //    8 : 132 - 0x84
      10'h9: dout <= 8'b10000101; //    9 : 133 - 0x85
      10'hA: dout <= 8'b10000100; //   10 : 132 - 0x84
      10'hB: dout <= 8'b10000101; //   11 : 133 - 0x85
      10'hC: dout <= 8'b10000100; //   12 : 132 - 0x84
      10'hD: dout <= 8'b10000110; //   13 : 134 - 0x86
      10'hE: dout <= 8'b10000100; //   14 : 132 - 0x84
      10'hF: dout <= 8'b10010110; //   15 : 150 - 0x96
      10'h10: dout <= 8'b10000111; //   16 : 135 - 0x87
      10'h11: dout <= 8'b10000101; //   17 : 133 - 0x85
      10'h12: dout <= 8'b10000100; //   18 : 132 - 0x84
      10'h13: dout <= 8'b10010111; //   19 : 151 - 0x97
      10'h14: dout <= 8'b10000100; //   20 : 132 - 0x84
      10'h15: dout <= 8'b10000101; //   21 : 133 - 0x85
      10'h16: dout <= 8'b10000100; //   22 : 132 - 0x84
      10'h17: dout <= 8'b10000101; //   23 : 133 - 0x85
      10'h18: dout <= 8'b10000100; //   24 : 132 - 0x84
      10'h19: dout <= 8'b10000111; //   25 : 135 - 0x87
      10'h1A: dout <= 8'b10000100; //   26 : 132 - 0x84
      10'h1B: dout <= 8'b10000101; //   27 : 133 - 0x85
      10'h1C: dout <= 8'b10000110; //   28 : 134 - 0x86
      10'h1D: dout <= 8'b10000101; //   29 : 133 - 0x85
      10'h1E: dout <= 8'b10000100; //   30 : 132 - 0x84
      10'h1F: dout <= 8'b10000101; //   31 : 133 - 0x85
      10'h20: dout <= 8'b10010100; //   32 : 148 - 0x94 -- line 0x1
      10'h21: dout <= 8'b10000111; //   33 : 135 - 0x87
      10'h22: dout <= 8'b10010100; //   34 : 148 - 0x94
      10'h23: dout <= 8'b10000110; //   35 : 134 - 0x86
      10'h24: dout <= 8'b10010100; //   36 : 148 - 0x94
      10'h25: dout <= 8'b10010101; //   37 : 149 - 0x95
      10'h26: dout <= 8'b10010110; //   38 : 150 - 0x96
      10'h27: dout <= 8'b10010101; //   39 : 149 - 0x95
      10'h28: dout <= 8'b10010100; //   40 : 148 - 0x94
      10'h29: dout <= 8'b10010101; //   41 : 149 - 0x95
      10'h2A: dout <= 8'b10010100; //   42 : 148 - 0x94
      10'h2B: dout <= 8'b10010111; //   43 : 151 - 0x97
      10'h2C: dout <= 8'b10010100; //   44 : 148 - 0x94
      10'h2D: dout <= 8'b10010101; //   45 : 149 - 0x95
      10'h2E: dout <= 8'b10010100; //   46 : 148 - 0x94
      10'h2F: dout <= 8'b10010101; //   47 : 149 - 0x95
      10'h30: dout <= 8'b10010100; //   48 : 148 - 0x94
      10'h31: dout <= 8'b10000110; //   49 : 134 - 0x86
      10'h32: dout <= 8'b10010100; //   50 : 148 - 0x94
      10'h33: dout <= 8'b10010101; //   51 : 149 - 0x95
      10'h34: dout <= 8'b10010100; //   52 : 148 - 0x94
      10'h35: dout <= 8'b10010101; //   53 : 149 - 0x95
      10'h36: dout <= 8'b10010110; //   54 : 150 - 0x96
      10'h37: dout <= 8'b10010101; //   55 : 149 - 0x95
      10'h38: dout <= 8'b10000110; //   56 : 134 - 0x86
      10'h39: dout <= 8'b10010101; //   57 : 149 - 0x95
      10'h3A: dout <= 8'b10010100; //   58 : 148 - 0x94
      10'h3B: dout <= 8'b10010111; //   59 : 151 - 0x97
      10'h3C: dout <= 8'b10010100; //   60 : 148 - 0x94
      10'h3D: dout <= 8'b10000111; //   61 : 135 - 0x87
      10'h3E: dout <= 8'b10010100; //   62 : 148 - 0x94
      10'h3F: dout <= 8'b10010101; //   63 : 149 - 0x95
      10'h40: dout <= 8'b10000010; //   64 : 130 - 0x82 -- line 0x2
      10'h41: dout <= 8'b10000011; //   65 : 131 - 0x83
      10'h42: dout <= 8'b10000010; //   66 : 130 - 0x82
      10'h43: dout <= 8'b10000011; //   67 : 131 - 0x83
      10'h44: dout <= 8'b10000010; //   68 : 130 - 0x82
      10'h45: dout <= 8'b10010001; //   69 : 145 - 0x91
      10'h46: dout <= 8'b10010000; //   70 : 144 - 0x90
      10'h47: dout <= 8'b10000011; //   71 : 131 - 0x83
      10'h48: dout <= 8'b10000010; //   72 : 130 - 0x82
      10'h49: dout <= 8'b10010001; //   73 : 145 - 0x91
      10'h4A: dout <= 8'b10010010; //   74 : 146 - 0x92
      10'h4B: dout <= 8'b10000011; //   75 : 131 - 0x83
      10'h4C: dout <= 8'b10000010; //   76 : 130 - 0x82
      10'h4D: dout <= 8'b10000011; //   77 : 131 - 0x83
      10'h4E: dout <= 8'b10000010; //   78 : 130 - 0x82
      10'h4F: dout <= 8'b10000001; //   79 : 129 - 0x81
      10'h50: dout <= 8'b10000010; //   80 : 130 - 0x82
      10'h51: dout <= 8'b10000011; //   81 : 131 - 0x83
      10'h52: dout <= 8'b10000010; //   82 : 130 - 0x82
      10'h53: dout <= 8'b10000011; //   83 : 131 - 0x83
      10'h54: dout <= 8'b10000010; //   84 : 130 - 0x82
      10'h55: dout <= 8'b10000011; //   85 : 131 - 0x83
      10'h56: dout <= 8'b10000010; //   86 : 130 - 0x82
      10'h57: dout <= 8'b10000011; //   87 : 131 - 0x83
      10'h58: dout <= 8'b10000001; //   88 : 129 - 0x81
      10'h59: dout <= 8'b10000011; //   89 : 131 - 0x83
      10'h5A: dout <= 8'b10010000; //   90 : 144 - 0x90
      10'h5B: dout <= 8'b10010011; //   91 : 147 - 0x93
      10'h5C: dout <= 8'b10000010; //   92 : 130 - 0x82
      10'h5D: dout <= 8'b10010000; //   93 : 144 - 0x90
      10'h5E: dout <= 8'b10010010; //   94 : 146 - 0x92
      10'h5F: dout <= 8'b10000011; //   95 : 131 - 0x83
      10'h60: dout <= 8'b01001001; //   96 :  73 - 0x49 -- line 0x3
      10'h61: dout <= 8'b01001001; //   97 :  73 - 0x49
      10'h62: dout <= 8'b01001001; //   98 :  73 - 0x49
      10'h63: dout <= 8'b01001001; //   99 :  73 - 0x49
      10'h64: dout <= 8'b01001001; //  100 :  73 - 0x49
      10'h65: dout <= 8'b01001001; //  101 :  73 - 0x49
      10'h66: dout <= 8'b01001001; //  102 :  73 - 0x49
      10'h67: dout <= 8'b01001001; //  103 :  73 - 0x49
      10'h68: dout <= 8'b01001001; //  104 :  73 - 0x49
      10'h69: dout <= 8'b01001001; //  105 :  73 - 0x49
      10'h6A: dout <= 8'b01001001; //  106 :  73 - 0x49
      10'h6B: dout <= 8'b01001001; //  107 :  73 - 0x49
      10'h6C: dout <= 8'b01001001; //  108 :  73 - 0x49
      10'h6D: dout <= 8'b01001001; //  109 :  73 - 0x49
      10'h6E: dout <= 8'b01001001; //  110 :  73 - 0x49
      10'h6F: dout <= 8'b01001001; //  111 :  73 - 0x49
      10'h70: dout <= 8'b01001001; //  112 :  73 - 0x49
      10'h71: dout <= 8'b01001001; //  113 :  73 - 0x49
      10'h72: dout <= 8'b01001001; //  114 :  73 - 0x49
      10'h73: dout <= 8'b01001001; //  115 :  73 - 0x49
      10'h74: dout <= 8'b01001001; //  116 :  73 - 0x49
      10'h75: dout <= 8'b01001001; //  117 :  73 - 0x49
      10'h76: dout <= 8'b01001001; //  118 :  73 - 0x49
      10'h77: dout <= 8'b01001001; //  119 :  73 - 0x49
      10'h78: dout <= 8'b01001001; //  120 :  73 - 0x49
      10'h79: dout <= 8'b01001001; //  121 :  73 - 0x49
      10'h7A: dout <= 8'b01001001; //  122 :  73 - 0x49
      10'h7B: dout <= 8'b01001001; //  123 :  73 - 0x49
      10'h7C: dout <= 8'b01001001; //  124 :  73 - 0x49
      10'h7D: dout <= 8'b01001001; //  125 :  73 - 0x49
      10'h7E: dout <= 8'b01001001; //  126 :  73 - 0x49
      10'h7F: dout <= 8'b01001001; //  127 :  73 - 0x49
      10'h80: dout <= 8'b00000000; //  128 :   0 - 0x0 -- line 0x4
      10'h81: dout <= 8'b00000000; //  129 :   0 - 0x0
      10'h82: dout <= 8'b00000000; //  130 :   0 - 0x0
      10'h83: dout <= 8'b00000000; //  131 :   0 - 0x0
      10'h84: dout <= 8'b00000001; //  132 :   1 - 0x1
      10'h85: dout <= 8'b00000010; //  133 :   2 - 0x2
      10'h86: dout <= 8'b00000010; //  134 :   2 - 0x2
      10'h87: dout <= 8'b00000011; //  135 :   3 - 0x3
      10'h88: dout <= 8'b00000000; //  136 :   0 - 0x0
      10'h89: dout <= 8'b00000000; //  137 :   0 - 0x0
      10'h8A: dout <= 8'b00000000; //  138 :   0 - 0x0
      10'h8B: dout <= 8'b00000100; //  139 :   4 - 0x4
      10'h8C: dout <= 8'b00000010; //  140 :   2 - 0x2
      10'h8D: dout <= 8'b00000010; //  141 :   2 - 0x2
      10'h8E: dout <= 8'b00000010; //  142 :   2 - 0x2
      10'h8F: dout <= 8'b00000101; //  143 :   5 - 0x5
      10'h90: dout <= 8'b00000001; //  144 :   1 - 0x1
      10'h91: dout <= 8'b00000010; //  145 :   2 - 0x2
      10'h92: dout <= 8'b00000010; //  146 :   2 - 0x2
      10'h93: dout <= 8'b00000110; //  147 :   6 - 0x6
      10'h94: dout <= 8'b00000010; //  148 :   2 - 0x2
      10'h95: dout <= 8'b00000010; //  149 :   2 - 0x2
      10'h96: dout <= 8'b00000110; //  150 :   6 - 0x6
      10'h97: dout <= 8'b00000010; //  151 :   2 - 0x2
      10'h98: dout <= 8'b00000010; //  152 :   2 - 0x2
      10'h99: dout <= 8'b00000111; //  153 :   7 - 0x7
      10'h9A: dout <= 8'b00000010; //  154 :   2 - 0x2
      10'h9B: dout <= 8'b00000010; //  155 :   2 - 0x2
      10'h9C: dout <= 8'b00000011; //  156 :   3 - 0x3
      10'h9D: dout <= 8'b00000000; //  157 :   0 - 0x0
      10'h9E: dout <= 8'b00000000; //  158 :   0 - 0x0
      10'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      10'hA0: dout <= 8'b00000000; //  160 :   0 - 0x0 -- line 0x5
      10'hA1: dout <= 8'b00000000; //  161 :   0 - 0x0
      10'hA2: dout <= 8'b00000000; //  162 :   0 - 0x0
      10'hA3: dout <= 8'b00000000; //  163 :   0 - 0x0
      10'hA4: dout <= 8'b00001000; //  164 :   8 - 0x8
      10'hA5: dout <= 8'b00001001; //  165 :   9 - 0x9
      10'hA6: dout <= 8'b00001001; //  166 :   9 - 0x9
      10'hA7: dout <= 8'b00001010; //  167 :  10 - 0xa
      10'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0
      10'hA9: dout <= 8'b00000000; //  169 :   0 - 0x0
      10'hAA: dout <= 8'b00001011; //  170 :  11 - 0xb
      10'hAB: dout <= 8'b00001100; //  171 :  12 - 0xc
      10'hAC: dout <= 8'b00001001; //  172 :   9 - 0x9
      10'hAD: dout <= 8'b00001001; //  173 :   9 - 0x9
      10'hAE: dout <= 8'b00001001; //  174 :   9 - 0x9
      10'hAF: dout <= 8'b00001101; //  175 :  13 - 0xd
      10'hB0: dout <= 8'b00001110; //  176 :  14 - 0xe
      10'hB1: dout <= 8'b00001001; //  177 :   9 - 0x9
      10'hB2: dout <= 8'b00001001; //  178 :   9 - 0x9
      10'hB3: dout <= 8'b00001111; //  179 :  15 - 0xf
      10'hB4: dout <= 8'b00001001; //  180 :   9 - 0x9
      10'hB5: dout <= 8'b00001001; //  181 :   9 - 0x9
      10'hB6: dout <= 8'b00001111; //  182 :  15 - 0xf
      10'hB7: dout <= 8'b00001001; //  183 :   9 - 0x9
      10'hB8: dout <= 8'b00001001; //  184 :   9 - 0x9
      10'hB9: dout <= 8'b00010000; //  185 :  16 - 0x10
      10'hBA: dout <= 8'b00001001; //  186 :   9 - 0x9
      10'hBB: dout <= 8'b00001001; //  187 :   9 - 0x9
      10'hBC: dout <= 8'b00001010; //  188 :  10 - 0xa
      10'hBD: dout <= 8'b00000000; //  189 :   0 - 0x0
      10'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      10'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      10'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- line 0x6
      10'hC1: dout <= 8'b00000000; //  193 :   0 - 0x0
      10'hC2: dout <= 8'b00000000; //  194 :   0 - 0x0
      10'hC3: dout <= 8'b00000000; //  195 :   0 - 0x0
      10'hC4: dout <= 8'b00001000; //  196 :   8 - 0x8
      10'hC5: dout <= 8'b00001001; //  197 :   9 - 0x9
      10'hC6: dout <= 8'b00001001; //  198 :   9 - 0x9
      10'hC7: dout <= 8'b00001010; //  199 :  10 - 0xa
      10'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0
      10'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      10'hCA: dout <= 8'b00001000; //  202 :   8 - 0x8
      10'hCB: dout <= 8'b00001001; //  203 :   9 - 0x9
      10'hCC: dout <= 8'b00001001; //  204 :   9 - 0x9
      10'hCD: dout <= 8'b00010001; //  205 :  17 - 0x11
      10'hCE: dout <= 8'b00001001; //  206 :   9 - 0x9
      10'hCF: dout <= 8'b00001001; //  207 :   9 - 0x9
      10'hD0: dout <= 8'b00001111; //  208 :  15 - 0xf
      10'hD1: dout <= 8'b00001001; //  209 :   9 - 0x9
      10'hD2: dout <= 8'b00001001; //  210 :   9 - 0x9
      10'hD3: dout <= 8'b00001111; //  211 :  15 - 0xf
      10'hD4: dout <= 8'b00001001; //  212 :   9 - 0x9
      10'hD5: dout <= 8'b00001001; //  213 :   9 - 0x9
      10'hD6: dout <= 8'b00001111; //  214 :  15 - 0xf
      10'hD7: dout <= 8'b00001001; //  215 :   9 - 0x9
      10'hD8: dout <= 8'b00001001; //  216 :   9 - 0x9
      10'hD9: dout <= 8'b00010010; //  217 :  18 - 0x12
      10'hDA: dout <= 8'b00001001; //  218 :   9 - 0x9
      10'hDB: dout <= 8'b00001001; //  219 :   9 - 0x9
      10'hDC: dout <= 8'b00001010; //  220 :  10 - 0xa
      10'hDD: dout <= 8'b00000000; //  221 :   0 - 0x0
      10'hDE: dout <= 8'b00000000; //  222 :   0 - 0x0
      10'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      10'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- line 0x7
      10'hE1: dout <= 8'b00000000; //  225 :   0 - 0x0
      10'hE2: dout <= 8'b00000000; //  226 :   0 - 0x0
      10'hE3: dout <= 8'b00000000; //  227 :   0 - 0x0
      10'hE4: dout <= 8'b00001000; //  228 :   8 - 0x8
      10'hE5: dout <= 8'b00001001; //  229 :   9 - 0x9
      10'hE6: dout <= 8'b00001001; //  230 :   9 - 0x9
      10'hE7: dout <= 8'b00001010; //  231 :  10 - 0xa
      10'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0
      10'hE9: dout <= 8'b00000000; //  233 :   0 - 0x0
      10'hEA: dout <= 8'b00001000; //  234 :   8 - 0x8
      10'hEB: dout <= 8'b00001001; //  235 :   9 - 0x9
      10'hEC: dout <= 8'b00001001; //  236 :   9 - 0x9
      10'hED: dout <= 8'b00001111; //  237 :  15 - 0xf
      10'hEE: dout <= 8'b00001001; //  238 :   9 - 0x9
      10'hEF: dout <= 8'b00001001; //  239 :   9 - 0x9
      10'hF0: dout <= 8'b00001111; //  240 :  15 - 0xf
      10'hF1: dout <= 8'b00001001; //  241 :   9 - 0x9
      10'hF2: dout <= 8'b00001001; //  242 :   9 - 0x9
      10'hF3: dout <= 8'b00010011; //  243 :  19 - 0x13
      10'hF4: dout <= 8'b00001001; //  244 :   9 - 0x9
      10'hF5: dout <= 8'b00001001; //  245 :   9 - 0x9
      10'hF6: dout <= 8'b00001111; //  246 :  15 - 0xf
      10'hF7: dout <= 8'b00001001; //  247 :   9 - 0x9
      10'hF8: dout <= 8'b00001001; //  248 :   9 - 0x9
      10'hF9: dout <= 8'b00010100; //  249 :  20 - 0x14
      10'hFA: dout <= 8'b00001001; //  250 :   9 - 0x9
      10'hFB: dout <= 8'b00001001; //  251 :   9 - 0x9
      10'hFC: dout <= 8'b00001010; //  252 :  10 - 0xa
      10'hFD: dout <= 8'b00000000; //  253 :   0 - 0x0
      10'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      10'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      10'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- line 0x8
      10'h101: dout <= 8'b00000000; //  257 :   0 - 0x0
      10'h102: dout <= 8'b00000000; //  258 :   0 - 0x0
      10'h103: dout <= 8'b00000000; //  259 :   0 - 0x0
      10'h104: dout <= 8'b00001000; //  260 :   8 - 0x8
      10'h105: dout <= 8'b00001001; //  261 :   9 - 0x9
      10'h106: dout <= 8'b00001001; //  262 :   9 - 0x9
      10'h107: dout <= 8'b00001010; //  263 :  10 - 0xa
      10'h108: dout <= 8'b00000000; //  264 :   0 - 0x0
      10'h109: dout <= 8'b00000000; //  265 :   0 - 0x0
      10'h10A: dout <= 8'b00001000; //  266 :   8 - 0x8
      10'h10B: dout <= 8'b00001001; //  267 :   9 - 0x9
      10'h10C: dout <= 8'b00001001; //  268 :   9 - 0x9
      10'h10D: dout <= 8'b00010101; //  269 :  21 - 0x15
      10'h10E: dout <= 8'b00001001; //  270 :   9 - 0x9
      10'h10F: dout <= 8'b00001001; //  271 :   9 - 0x9
      10'h110: dout <= 8'b00001111; //  272 :  15 - 0xf
      10'h111: dout <= 8'b00001001; //  273 :   9 - 0x9
      10'h112: dout <= 8'b00001001; //  274 :   9 - 0x9
      10'h113: dout <= 8'b00010110; //  275 :  22 - 0x16
      10'h114: dout <= 8'b00001001; //  276 :   9 - 0x9
      10'h115: dout <= 8'b00001001; //  277 :   9 - 0x9
      10'h116: dout <= 8'b00001111; //  278 :  15 - 0xf
      10'h117: dout <= 8'b00001001; //  279 :   9 - 0x9
      10'h118: dout <= 8'b00001001; //  280 :   9 - 0x9
      10'h119: dout <= 8'b00010111; //  281 :  23 - 0x17
      10'h11A: dout <= 8'b00001001; //  282 :   9 - 0x9
      10'h11B: dout <= 8'b00001001; //  283 :   9 - 0x9
      10'h11C: dout <= 8'b00001010; //  284 :  10 - 0xa
      10'h11D: dout <= 8'b00000000; //  285 :   0 - 0x0
      10'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      10'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      10'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- line 0x9
      10'h121: dout <= 8'b00000000; //  289 :   0 - 0x0
      10'h122: dout <= 8'b00000000; //  290 :   0 - 0x0
      10'h123: dout <= 8'b00000000; //  291 :   0 - 0x0
      10'h124: dout <= 8'b00001000; //  292 :   8 - 0x8
      10'h125: dout <= 8'b00001001; //  293 :   9 - 0x9
      10'h126: dout <= 8'b00001001; //  294 :   9 - 0x9
      10'h127: dout <= 8'b00011000; //  295 :  24 - 0x18
      10'h128: dout <= 8'b00000010; //  296 :   2 - 0x2
      10'h129: dout <= 8'b00000010; //  297 :   2 - 0x2
      10'h12A: dout <= 8'b00011001; //  298 :  25 - 0x19
      10'h12B: dout <= 8'b00001001; //  299 :   9 - 0x9
      10'h12C: dout <= 8'b00001001; //  300 :   9 - 0x9
      10'h12D: dout <= 8'b00001001; //  301 :   9 - 0x9
      10'h12E: dout <= 8'b00001001; //  302 :   9 - 0x9
      10'h12F: dout <= 8'b00001001; //  303 :   9 - 0x9
      10'h130: dout <= 8'b00001111; //  304 :  15 - 0xf
      10'h131: dout <= 8'b00001001; //  305 :   9 - 0x9
      10'h132: dout <= 8'b00001001; //  306 :   9 - 0x9
      10'h133: dout <= 8'b00011010; //  307 :  26 - 0x1a
      10'h134: dout <= 8'b00001001; //  308 :   9 - 0x9
      10'h135: dout <= 8'b00001001; //  309 :   9 - 0x9
      10'h136: dout <= 8'b00001111; //  310 :  15 - 0xf
      10'h137: dout <= 8'b00001001; //  311 :   9 - 0x9
      10'h138: dout <= 8'b00001001; //  312 :   9 - 0x9
      10'h139: dout <= 8'b00001111; //  313 :  15 - 0xf
      10'h13A: dout <= 8'b00001001; //  314 :   9 - 0x9
      10'h13B: dout <= 8'b00001001; //  315 :   9 - 0x9
      10'h13C: dout <= 8'b00001010; //  316 :  10 - 0xa
      10'h13D: dout <= 8'b00000000; //  317 :   0 - 0x0
      10'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      10'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      10'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- line 0xa
      10'h141: dout <= 8'b00000000; //  321 :   0 - 0x0
      10'h142: dout <= 8'b00000000; //  322 :   0 - 0x0
      10'h143: dout <= 8'b00000000; //  323 :   0 - 0x0
      10'h144: dout <= 8'b00001000; //  324 :   8 - 0x8
      10'h145: dout <= 8'b00001001; //  325 :   9 - 0x9
      10'h146: dout <= 8'b00001001; //  326 :   9 - 0x9
      10'h147: dout <= 8'b00001001; //  327 :   9 - 0x9
      10'h148: dout <= 8'b00001001; //  328 :   9 - 0x9
      10'h149: dout <= 8'b00001001; //  329 :   9 - 0x9
      10'h14A: dout <= 8'b00001111; //  330 :  15 - 0xf
      10'h14B: dout <= 8'b00001001; //  331 :   9 - 0x9
      10'h14C: dout <= 8'b00001001; //  332 :   9 - 0x9
      10'h14D: dout <= 8'b00011011; //  333 :  27 - 0x1b
      10'h14E: dout <= 8'b00001001; //  334 :   9 - 0x9
      10'h14F: dout <= 8'b00001001; //  335 :   9 - 0x9
      10'h150: dout <= 8'b00001111; //  336 :  15 - 0xf
      10'h151: dout <= 8'b00001001; //  337 :   9 - 0x9
      10'h152: dout <= 8'b00011100; //  338 :  28 - 0x1c
      10'h153: dout <= 8'b00011101; //  339 :  29 - 0x1d
      10'h154: dout <= 8'b00011110; //  340 :  30 - 0x1e
      10'h155: dout <= 8'b00001001; //  341 :   9 - 0x9
      10'h156: dout <= 8'b00001111; //  342 :  15 - 0xf
      10'h157: dout <= 8'b00001001; //  343 :   9 - 0x9
      10'h158: dout <= 8'b00001001; //  344 :   9 - 0x9
      10'h159: dout <= 8'b00001111; //  345 :  15 - 0xf
      10'h15A: dout <= 8'b00001001; //  346 :   9 - 0x9
      10'h15B: dout <= 8'b00001001; //  347 :   9 - 0x9
      10'h15C: dout <= 8'b00001010; //  348 :  10 - 0xa
      10'h15D: dout <= 8'b00000000; //  349 :   0 - 0x0
      10'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      10'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      10'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- line 0xb
      10'h161: dout <= 8'b00000000; //  353 :   0 - 0x0
      10'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      10'h163: dout <= 8'b00000000; //  355 :   0 - 0x0
      10'h164: dout <= 8'b00011111; //  356 :  31 - 0x1f
      10'h165: dout <= 8'b00100000; //  357 :  32 - 0x20
      10'h166: dout <= 8'b00100000; //  358 :  32 - 0x20
      10'h167: dout <= 8'b00100000; //  359 :  32 - 0x20
      10'h168: dout <= 8'b00100000; //  360 :  32 - 0x20
      10'h169: dout <= 8'b00100000; //  361 :  32 - 0x20
      10'h16A: dout <= 8'b00100001; //  362 :  33 - 0x21
      10'h16B: dout <= 8'b00100000; //  363 :  32 - 0x20
      10'h16C: dout <= 8'b00100000; //  364 :  32 - 0x20
      10'h16D: dout <= 8'b00100001; //  365 :  33 - 0x21
      10'h16E: dout <= 8'b00100000; //  366 :  32 - 0x20
      10'h16F: dout <= 8'b00100000; //  367 :  32 - 0x20
      10'h170: dout <= 8'b00100001; //  368 :  33 - 0x21
      10'h171: dout <= 8'b00100000; //  369 :  32 - 0x20
      10'h172: dout <= 8'b00100010; //  370 :  34 - 0x22
      10'h173: dout <= 8'b00000000; //  371 :   0 - 0x0
      10'h174: dout <= 8'b00100011; //  372 :  35 - 0x23
      10'h175: dout <= 8'b00100000; //  373 :  32 - 0x20
      10'h176: dout <= 8'b00100001; //  374 :  33 - 0x21
      10'h177: dout <= 8'b00100000; //  375 :  32 - 0x20
      10'h178: dout <= 8'b00100000; //  376 :  32 - 0x20
      10'h179: dout <= 8'b00100001; //  377 :  33 - 0x21
      10'h17A: dout <= 8'b00100000; //  378 :  32 - 0x20
      10'h17B: dout <= 8'b00100000; //  379 :  32 - 0x20
      10'h17C: dout <= 8'b00100100; //  380 :  36 - 0x24
      10'h17D: dout <= 8'b00000000; //  381 :   0 - 0x0
      10'h17E: dout <= 8'b00000000; //  382 :   0 - 0x0
      10'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      10'h180: dout <= 8'b00000000; //  384 :   0 - 0x0 -- line 0xc
      10'h181: dout <= 8'b00000001; //  385 :   1 - 0x1
      10'h182: dout <= 8'b00000010; //  386 :   2 - 0x2
      10'h183: dout <= 8'b00100101; //  387 :  37 - 0x25
      10'h184: dout <= 8'b00000000; //  388 :   0 - 0x0
      10'h185: dout <= 8'b00100110; //  389 :  38 - 0x26
      10'h186: dout <= 8'b00000010; //  390 :   2 - 0x2
      10'h187: dout <= 8'b00000011; //  391 :   3 - 0x3
      10'h188: dout <= 8'b00000100; //  392 :   4 - 0x4
      10'h189: dout <= 8'b00000010; //  393 :   2 - 0x2
      10'h18A: dout <= 8'b00000010; //  394 :   2 - 0x2
      10'h18B: dout <= 8'b00000010; //  395 :   2 - 0x2
      10'h18C: dout <= 8'b00000101; //  396 :   5 - 0x5
      10'h18D: dout <= 8'b00000001; //  397 :   1 - 0x1
      10'h18E: dout <= 8'b00000010; //  398 :   2 - 0x2
      10'h18F: dout <= 8'b00000010; //  399 :   2 - 0x2
      10'h190: dout <= 8'b00000110; //  400 :   6 - 0x6
      10'h191: dout <= 8'b00000010; //  401 :   2 - 0x2
      10'h192: dout <= 8'b00000010; //  402 :   2 - 0x2
      10'h193: dout <= 8'b00000110; //  403 :   6 - 0x6
      10'h194: dout <= 8'b00000010; //  404 :   2 - 0x2
      10'h195: dout <= 8'b00000010; //  405 :   2 - 0x2
      10'h196: dout <= 8'b00000010; //  406 :   2 - 0x2
      10'h197: dout <= 8'b00000010; //  407 :   2 - 0x2
      10'h198: dout <= 8'b00000010; //  408 :   2 - 0x2
      10'h199: dout <= 8'b00000110; //  409 :   6 - 0x6
      10'h19A: dout <= 8'b00000010; //  410 :   2 - 0x2
      10'h19B: dout <= 8'b00000010; //  411 :   2 - 0x2
      10'h19C: dout <= 8'b00000010; //  412 :   2 - 0x2
      10'h19D: dout <= 8'b00000010; //  413 :   2 - 0x2
      10'h19E: dout <= 8'b00000101; //  414 :   5 - 0x5
      10'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      10'h1A0: dout <= 8'b00000000; //  416 :   0 - 0x0 -- line 0xd
      10'h1A1: dout <= 8'b00001000; //  417 :   8 - 0x8
      10'h1A2: dout <= 8'b00001001; //  418 :   9 - 0x9
      10'h1A3: dout <= 8'b00100111; //  419 :  39 - 0x27
      10'h1A4: dout <= 8'b00101000; //  420 :  40 - 0x28
      10'h1A5: dout <= 8'b00101001; //  421 :  41 - 0x29
      10'h1A6: dout <= 8'b00001001; //  422 :   9 - 0x9
      10'h1A7: dout <= 8'b00101010; //  423 :  42 - 0x2a
      10'h1A8: dout <= 8'b00001100; //  424 :  12 - 0xc
      10'h1A9: dout <= 8'b00001001; //  425 :   9 - 0x9
      10'h1AA: dout <= 8'b00001001; //  426 :   9 - 0x9
      10'h1AB: dout <= 8'b00001001; //  427 :   9 - 0x9
      10'h1AC: dout <= 8'b00001101; //  428 :  13 - 0xd
      10'h1AD: dout <= 8'b00001110; //  429 :  14 - 0xe
      10'h1AE: dout <= 8'b00001001; //  430 :   9 - 0x9
      10'h1AF: dout <= 8'b00001001; //  431 :   9 - 0x9
      10'h1B0: dout <= 8'b00001111; //  432 :  15 - 0xf
      10'h1B1: dout <= 8'b00001001; //  433 :   9 - 0x9
      10'h1B2: dout <= 8'b00001001; //  434 :   9 - 0x9
      10'h1B3: dout <= 8'b00001111; //  435 :  15 - 0xf
      10'h1B4: dout <= 8'b00001001; //  436 :   9 - 0x9
      10'h1B5: dout <= 8'b00001001; //  437 :   9 - 0x9
      10'h1B6: dout <= 8'b00001001; //  438 :   9 - 0x9
      10'h1B7: dout <= 8'b00001001; //  439 :   9 - 0x9
      10'h1B8: dout <= 8'b00001001; //  440 :   9 - 0x9
      10'h1B9: dout <= 8'b00001111; //  441 :  15 - 0xf
      10'h1BA: dout <= 8'b00001001; //  442 :   9 - 0x9
      10'h1BB: dout <= 8'b00001001; //  443 :   9 - 0x9
      10'h1BC: dout <= 8'b00001001; //  444 :   9 - 0x9
      10'h1BD: dout <= 8'b00001001; //  445 :   9 - 0x9
      10'h1BE: dout <= 8'b00001101; //  446 :  13 - 0xd
      10'h1BF: dout <= 8'b00101011; //  447 :  43 - 0x2b
      10'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- line 0xe
      10'h1C1: dout <= 8'b00001000; //  449 :   8 - 0x8
      10'h1C2: dout <= 8'b00001001; //  450 :   9 - 0x9
      10'h1C3: dout <= 8'b00001001; //  451 :   9 - 0x9
      10'h1C4: dout <= 8'b00101100; //  452 :  44 - 0x2c
      10'h1C5: dout <= 8'b00001001; //  453 :   9 - 0x9
      10'h1C6: dout <= 8'b00001001; //  454 :   9 - 0x9
      10'h1C7: dout <= 8'b00001111; //  455 :  15 - 0xf
      10'h1C8: dout <= 8'b00001001; //  456 :   9 - 0x9
      10'h1C9: dout <= 8'b00001001; //  457 :   9 - 0x9
      10'h1CA: dout <= 8'b00010001; //  458 :  17 - 0x11
      10'h1CB: dout <= 8'b00001001; //  459 :   9 - 0x9
      10'h1CC: dout <= 8'b00001001; //  460 :   9 - 0x9
      10'h1CD: dout <= 8'b00001111; //  461 :  15 - 0xf
      10'h1CE: dout <= 8'b00001001; //  462 :   9 - 0x9
      10'h1CF: dout <= 8'b00001001; //  463 :   9 - 0x9
      10'h1D0: dout <= 8'b00001111; //  464 :  15 - 0xf
      10'h1D1: dout <= 8'b00001001; //  465 :   9 - 0x9
      10'h1D2: dout <= 8'b00001001; //  466 :   9 - 0x9
      10'h1D3: dout <= 8'b00001111; //  467 :  15 - 0xf
      10'h1D4: dout <= 8'b00001001; //  468 :   9 - 0x9
      10'h1D5: dout <= 8'b00001001; //  469 :   9 - 0x9
      10'h1D6: dout <= 8'b00101101; //  470 :  45 - 0x2d
      10'h1D7: dout <= 8'b00100000; //  471 :  32 - 0x20
      10'h1D8: dout <= 8'b00100000; //  472 :  32 - 0x20
      10'h1D9: dout <= 8'b00101110; //  473 :  46 - 0x2e
      10'h1DA: dout <= 8'b00001001; //  474 :   9 - 0x9
      10'h1DB: dout <= 8'b00001001; //  475 :   9 - 0x9
      10'h1DC: dout <= 8'b00101111; //  476 :  47 - 0x2f
      10'h1DD: dout <= 8'b00001001; //  477 :   9 - 0x9
      10'h1DE: dout <= 8'b00001001; //  478 :   9 - 0x9
      10'h1DF: dout <= 8'b00001010; //  479 :  10 - 0xa
      10'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- line 0xf
      10'h1E1: dout <= 8'b00001000; //  481 :   8 - 0x8
      10'h1E2: dout <= 8'b00001001; //  482 :   9 - 0x9
      10'h1E3: dout <= 8'b00001001; //  483 :   9 - 0x9
      10'h1E4: dout <= 8'b00110000; //  484 :  48 - 0x30
      10'h1E5: dout <= 8'b00001001; //  485 :   9 - 0x9
      10'h1E6: dout <= 8'b00001001; //  486 :   9 - 0x9
      10'h1E7: dout <= 8'b00001111; //  487 :  15 - 0xf
      10'h1E8: dout <= 8'b00001001; //  488 :   9 - 0x9
      10'h1E9: dout <= 8'b00001001; //  489 :   9 - 0x9
      10'h1EA: dout <= 8'b00001111; //  490 :  15 - 0xf
      10'h1EB: dout <= 8'b00001001; //  491 :   9 - 0x9
      10'h1EC: dout <= 8'b00001001; //  492 :   9 - 0x9
      10'h1ED: dout <= 8'b00001111; //  493 :  15 - 0xf
      10'h1EE: dout <= 8'b00001001; //  494 :   9 - 0x9
      10'h1EF: dout <= 8'b00001001; //  495 :   9 - 0x9
      10'h1F0: dout <= 8'b00010011; //  496 :  19 - 0x13
      10'h1F1: dout <= 8'b00001001; //  497 :   9 - 0x9
      10'h1F2: dout <= 8'b00001001; //  498 :   9 - 0x9
      10'h1F3: dout <= 8'b00001111; //  499 :  15 - 0xf
      10'h1F4: dout <= 8'b00001001; //  500 :   9 - 0x9
      10'h1F5: dout <= 8'b00001001; //  501 :   9 - 0x9
      10'h1F6: dout <= 8'b00110001; //  502 :  49 - 0x31
      10'h1F7: dout <= 8'b00110010; //  503 :  50 - 0x32
      10'h1F8: dout <= 8'b00110011; //  504 :  51 - 0x33
      10'h1F9: dout <= 8'b00001000; //  505 :   8 - 0x8
      10'h1FA: dout <= 8'b00001001; //  506 :   9 - 0x9
      10'h1FB: dout <= 8'b00001001; //  507 :   9 - 0x9
      10'h1FC: dout <= 8'b00001111; //  508 :  15 - 0xf
      10'h1FD: dout <= 8'b00001001; //  509 :   9 - 0x9
      10'h1FE: dout <= 8'b00001001; //  510 :   9 - 0x9
      10'h1FF: dout <= 8'b00001010; //  511 :  10 - 0xa
      10'h200: dout <= 8'b00000000; //  512 :   0 - 0x0 -- line 0x10
      10'h201: dout <= 8'b00001000; //  513 :   8 - 0x8
      10'h202: dout <= 8'b00001001; //  514 :   9 - 0x9
      10'h203: dout <= 8'b00001001; //  515 :   9 - 0x9
      10'h204: dout <= 8'b00110100; //  516 :  52 - 0x34
      10'h205: dout <= 8'b00001001; //  517 :   9 - 0x9
      10'h206: dout <= 8'b00001001; //  518 :   9 - 0x9
      10'h207: dout <= 8'b00001111; //  519 :  15 - 0xf
      10'h208: dout <= 8'b00001001; //  520 :   9 - 0x9
      10'h209: dout <= 8'b00001001; //  521 :   9 - 0x9
      10'h20A: dout <= 8'b00001111; //  522 :  15 - 0xf
      10'h20B: dout <= 8'b00001001; //  523 :   9 - 0x9
      10'h20C: dout <= 8'b00001001; //  524 :   9 - 0x9
      10'h20D: dout <= 8'b00001111; //  525 :  15 - 0xf
      10'h20E: dout <= 8'b00001001; //  526 :   9 - 0x9
      10'h20F: dout <= 8'b00001001; //  527 :   9 - 0x9
      10'h210: dout <= 8'b00010110; //  528 :  22 - 0x16
      10'h211: dout <= 8'b00001001; //  529 :   9 - 0x9
      10'h212: dout <= 8'b00001001; //  530 :   9 - 0x9
      10'h213: dout <= 8'b00001111; //  531 :  15 - 0xf
      10'h214: dout <= 8'b00001001; //  532 :   9 - 0x9
      10'h215: dout <= 8'b00001001; //  533 :   9 - 0x9
      10'h216: dout <= 8'b00110101; //  534 :  53 - 0x35
      10'h217: dout <= 8'b00110110; //  535 :  54 - 0x36
      10'h218: dout <= 8'b00110111; //  536 :  55 - 0x37
      10'h219: dout <= 8'b00001000; //  537 :   8 - 0x8
      10'h21A: dout <= 8'b00001001; //  538 :   9 - 0x9
      10'h21B: dout <= 8'b00001001; //  539 :   9 - 0x9
      10'h21C: dout <= 8'b00111000; //  540 :  56 - 0x38
      10'h21D: dout <= 8'b00001001; //  541 :   9 - 0x9
      10'h21E: dout <= 8'b00111001; //  542 :  57 - 0x39
      10'h21F: dout <= 8'b00001010; //  543 :  10 - 0xa
      10'h220: dout <= 8'b00000000; //  544 :   0 - 0x0 -- line 0x11
      10'h221: dout <= 8'b00001000; //  545 :   8 - 0x8
      10'h222: dout <= 8'b00001001; //  546 :   9 - 0x9
      10'h223: dout <= 8'b00001001; //  547 :   9 - 0x9
      10'h224: dout <= 8'b00001111; //  548 :  15 - 0xf
      10'h225: dout <= 8'b00001001; //  549 :   9 - 0x9
      10'h226: dout <= 8'b00001001; //  550 :   9 - 0x9
      10'h227: dout <= 8'b00001111; //  551 :  15 - 0xf
      10'h228: dout <= 8'b00001001; //  552 :   9 - 0x9
      10'h229: dout <= 8'b00001001; //  553 :   9 - 0x9
      10'h22A: dout <= 8'b00111010; //  554 :  58 - 0x3a
      10'h22B: dout <= 8'b00001001; //  555 :   9 - 0x9
      10'h22C: dout <= 8'b00001001; //  556 :   9 - 0x9
      10'h22D: dout <= 8'b00001111; //  557 :  15 - 0xf
      10'h22E: dout <= 8'b00001001; //  558 :   9 - 0x9
      10'h22F: dout <= 8'b00001001; //  559 :   9 - 0x9
      10'h230: dout <= 8'b00011010; //  560 :  26 - 0x1a
      10'h231: dout <= 8'b00001001; //  561 :   9 - 0x9
      10'h232: dout <= 8'b00001001; //  562 :   9 - 0x9
      10'h233: dout <= 8'b00001111; //  563 :  15 - 0xf
      10'h234: dout <= 8'b00001001; //  564 :   9 - 0x9
      10'h235: dout <= 8'b00001001; //  565 :   9 - 0x9
      10'h236: dout <= 8'b00111011; //  566 :  59 - 0x3b
      10'h237: dout <= 8'b00111100; //  567 :  60 - 0x3c
      10'h238: dout <= 8'b00111101; //  568 :  61 - 0x3d
      10'h239: dout <= 8'b00011001; //  569 :  25 - 0x19
      10'h23A: dout <= 8'b00001001; //  570 :   9 - 0x9
      10'h23B: dout <= 8'b00001001; //  571 :   9 - 0x9
      10'h23C: dout <= 8'b00001001; //  572 :   9 - 0x9
      10'h23D: dout <= 8'b00001001; //  573 :   9 - 0x9
      10'h23E: dout <= 8'b00111110; //  574 :  62 - 0x3e
      10'h23F: dout <= 8'b00111111; //  575 :  63 - 0x3f
      10'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- line 0x12
      10'h241: dout <= 8'b00001000; //  577 :   8 - 0x8
      10'h242: dout <= 8'b00001001; //  578 :   9 - 0x9
      10'h243: dout <= 8'b00001001; //  579 :   9 - 0x9
      10'h244: dout <= 8'b00001111; //  580 :  15 - 0xf
      10'h245: dout <= 8'b00001001; //  581 :   9 - 0x9
      10'h246: dout <= 8'b00001001; //  582 :   9 - 0x9
      10'h247: dout <= 8'b01000000; //  583 :  64 - 0x40
      10'h248: dout <= 8'b01000001; //  584 :  65 - 0x41
      10'h249: dout <= 8'b00001001; //  585 :   9 - 0x9
      10'h24A: dout <= 8'b00001001; //  586 :   9 - 0x9
      10'h24B: dout <= 8'b00001001; //  587 :   9 - 0x9
      10'h24C: dout <= 8'b01000010; //  588 :  66 - 0x42
      10'h24D: dout <= 8'b01000011; //  589 :  67 - 0x43
      10'h24E: dout <= 8'b00001001; //  590 :   9 - 0x9
      10'h24F: dout <= 8'b00011100; //  591 :  28 - 0x1c
      10'h250: dout <= 8'b00011101; //  592 :  29 - 0x1d
      10'h251: dout <= 8'b00011110; //  593 :  30 - 0x1e
      10'h252: dout <= 8'b00001001; //  594 :   9 - 0x9
      10'h253: dout <= 8'b00001111; //  595 :  15 - 0xf
      10'h254: dout <= 8'b00001001; //  596 :   9 - 0x9
      10'h255: dout <= 8'b00001001; //  597 :   9 - 0x9
      10'h256: dout <= 8'b00001001; //  598 :   9 - 0x9
      10'h257: dout <= 8'b00001001; //  599 :   9 - 0x9
      10'h258: dout <= 8'b00001001; //  600 :   9 - 0x9
      10'h259: dout <= 8'b00001111; //  601 :  15 - 0xf
      10'h25A: dout <= 8'b00001001; //  602 :   9 - 0x9
      10'h25B: dout <= 8'b00001001; //  603 :   9 - 0x9
      10'h25C: dout <= 8'b00101111; //  604 :  47 - 0x2f
      10'h25D: dout <= 8'b00001001; //  605 :   9 - 0x9
      10'h25E: dout <= 8'b01000100; //  606 :  68 - 0x44
      10'h25F: dout <= 8'b01000101; //  607 :  69 - 0x45
      10'h260: dout <= 8'b00000000; //  608 :   0 - 0x0 -- line 0x13
      10'h261: dout <= 8'b00011111; //  609 :  31 - 0x1f
      10'h262: dout <= 8'b00100000; //  610 :  32 - 0x20
      10'h263: dout <= 8'b00100000; //  611 :  32 - 0x20
      10'h264: dout <= 8'b00100001; //  612 :  33 - 0x21
      10'h265: dout <= 8'b00100000; //  613 :  32 - 0x20
      10'h266: dout <= 8'b00100000; //  614 :  32 - 0x20
      10'h267: dout <= 8'b00100100; //  615 :  36 - 0x24
      10'h268: dout <= 8'b01000110; //  616 :  70 - 0x46
      10'h269: dout <= 8'b00100000; //  617 :  32 - 0x20
      10'h26A: dout <= 8'b00100000; //  618 :  32 - 0x20
      10'h26B: dout <= 8'b00100000; //  619 :  32 - 0x20
      10'h26C: dout <= 8'b01000111; //  620 :  71 - 0x47
      10'h26D: dout <= 8'b01001000; //  621 :  72 - 0x48
      10'h26E: dout <= 8'b00100000; //  622 :  32 - 0x20
      10'h26F: dout <= 8'b00100010; //  623 :  34 - 0x22
      10'h270: dout <= 8'b00000000; //  624 :   0 - 0x0
      10'h271: dout <= 8'b00100011; //  625 :  35 - 0x23
      10'h272: dout <= 8'b00100000; //  626 :  32 - 0x20
      10'h273: dout <= 8'b00100001; //  627 :  33 - 0x21
      10'h274: dout <= 8'b00100000; //  628 :  32 - 0x20
      10'h275: dout <= 8'b00100000; //  629 :  32 - 0x20
      10'h276: dout <= 8'b00100000; //  630 :  32 - 0x20
      10'h277: dout <= 8'b00100000; //  631 :  32 - 0x20
      10'h278: dout <= 8'b00100000; //  632 :  32 - 0x20
      10'h279: dout <= 8'b00100001; //  633 :  33 - 0x21
      10'h27A: dout <= 8'b00100000; //  634 :  32 - 0x20
      10'h27B: dout <= 8'b00100000; //  635 :  32 - 0x20
      10'h27C: dout <= 8'b00100001; //  636 :  33 - 0x21
      10'h27D: dout <= 8'b00100000; //  637 :  32 - 0x20
      10'h27E: dout <= 8'b00100000; //  638 :  32 - 0x20
      10'h27F: dout <= 8'b00100100; //  639 :  36 - 0x24
      10'h280: dout <= 8'b00000000; //  640 :   0 - 0x0 -- line 0x14
      10'h281: dout <= 8'b00000000; //  641 :   0 - 0x0
      10'h282: dout <= 8'b00000000; //  642 :   0 - 0x0
      10'h283: dout <= 8'b00000000; //  643 :   0 - 0x0
      10'h284: dout <= 8'b00000000; //  644 :   0 - 0x0
      10'h285: dout <= 8'b00000000; //  645 :   0 - 0x0
      10'h286: dout <= 8'b00000000; //  646 :   0 - 0x0
      10'h287: dout <= 8'b00000000; //  647 :   0 - 0x0
      10'h288: dout <= 8'b00000000; //  648 :   0 - 0x0
      10'h289: dout <= 8'b00000000; //  649 :   0 - 0x0
      10'h28A: dout <= 8'b00000000; //  650 :   0 - 0x0
      10'h28B: dout <= 8'b00000000; //  651 :   0 - 0x0
      10'h28C: dout <= 8'b00000000; //  652 :   0 - 0x0
      10'h28D: dout <= 8'b00000000; //  653 :   0 - 0x0
      10'h28E: dout <= 8'b00000000; //  654 :   0 - 0x0
      10'h28F: dout <= 8'b00000000; //  655 :   0 - 0x0
      10'h290: dout <= 8'b00000000; //  656 :   0 - 0x0
      10'h291: dout <= 8'b00000000; //  657 :   0 - 0x0
      10'h292: dout <= 8'b00000000; //  658 :   0 - 0x0
      10'h293: dout <= 8'b00000000; //  659 :   0 - 0x0
      10'h294: dout <= 8'b00000000; //  660 :   0 - 0x0
      10'h295: dout <= 8'b00000000; //  661 :   0 - 0x0
      10'h296: dout <= 8'b00000000; //  662 :   0 - 0x0
      10'h297: dout <= 8'b00000000; //  663 :   0 - 0x0
      10'h298: dout <= 8'b00000000; //  664 :   0 - 0x0
      10'h299: dout <= 8'b00000000; //  665 :   0 - 0x0
      10'h29A: dout <= 8'b00000000; //  666 :   0 - 0x0
      10'h29B: dout <= 8'b00000000; //  667 :   0 - 0x0
      10'h29C: dout <= 8'b00000000; //  668 :   0 - 0x0
      10'h29D: dout <= 8'b00000000; //  669 :   0 - 0x0
      10'h29E: dout <= 8'b00000000; //  670 :   0 - 0x0
      10'h29F: dout <= 8'b00000000; //  671 :   0 - 0x0
      10'h2A0: dout <= 8'b00000000; //  672 :   0 - 0x0 -- line 0x15
      10'h2A1: dout <= 8'b00000000; //  673 :   0 - 0x0
      10'h2A2: dout <= 8'b00000000; //  674 :   0 - 0x0
      10'h2A3: dout <= 8'b00000000; //  675 :   0 - 0x0
      10'h2A4: dout <= 8'b00000000; //  676 :   0 - 0x0
      10'h2A5: dout <= 8'b00000000; //  677 :   0 - 0x0
      10'h2A6: dout <= 8'b00000000; //  678 :   0 - 0x0
      10'h2A7: dout <= 8'b00000000; //  679 :   0 - 0x0
      10'h2A8: dout <= 8'b00000000; //  680 :   0 - 0x0
      10'h2A9: dout <= 8'b00000000; //  681 :   0 - 0x0
      10'h2AA: dout <= 8'b00000000; //  682 :   0 - 0x0
      10'h2AB: dout <= 8'b01010000; //  683 :  80 - 0x50
      10'h2AC: dout <= 8'b01010001; //  684 :  81 - 0x51
      10'h2AD: dout <= 8'b01010010; //  685 :  82 - 0x52
      10'h2AE: dout <= 8'b01010011; //  686 :  83 - 0x53
      10'h2AF: dout <= 8'b01010011; //  687 :  83 - 0x53
      10'h2B0: dout <= 8'b00000000; //  688 :   0 - 0x0
      10'h2B1: dout <= 8'b01010011; //  689 :  83 - 0x53
      10'h2B2: dout <= 8'b01010100; //  690 :  84 - 0x54
      10'h2B3: dout <= 8'b01010101; //  691 :  85 - 0x55
      10'h2B4: dout <= 8'b01010001; //  692 :  81 - 0x51
      10'h2B5: dout <= 8'b01010100; //  693 :  84 - 0x54
      10'h2B6: dout <= 8'b00000000; //  694 :   0 - 0x0
      10'h2B7: dout <= 8'b00000000; //  695 :   0 - 0x0
      10'h2B8: dout <= 8'b00000000; //  696 :   0 - 0x0
      10'h2B9: dout <= 8'b00000000; //  697 :   0 - 0x0
      10'h2BA: dout <= 8'b00000000; //  698 :   0 - 0x0
      10'h2BB: dout <= 8'b00000000; //  699 :   0 - 0x0
      10'h2BC: dout <= 8'b00000000; //  700 :   0 - 0x0
      10'h2BD: dout <= 8'b00000000; //  701 :   0 - 0x0
      10'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      10'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      10'h2C0: dout <= 8'b00000000; //  704 :   0 - 0x0 -- line 0x16
      10'h2C1: dout <= 8'b00000000; //  705 :   0 - 0x0
      10'h2C2: dout <= 8'b00000000; //  706 :   0 - 0x0
      10'h2C3: dout <= 8'b00000000; //  707 :   0 - 0x0
      10'h2C4: dout <= 8'b00000000; //  708 :   0 - 0x0
      10'h2C5: dout <= 8'b00000000; //  709 :   0 - 0x0
      10'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      10'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      10'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0
      10'h2C9: dout <= 8'b00000000; //  713 :   0 - 0x0
      10'h2CA: dout <= 8'b00000000; //  714 :   0 - 0x0
      10'h2CB: dout <= 8'b01100000; //  715 :  96 - 0x60
      10'h2CC: dout <= 8'b01100001; //  716 :  97 - 0x61
      10'h2CD: dout <= 8'b01100010; //  717 :  98 - 0x62
      10'h2CE: dout <= 8'b01100011; //  718 :  99 - 0x63
      10'h2CF: dout <= 8'b01100011; //  719 :  99 - 0x63
      10'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0
      10'h2D1: dout <= 8'b01100011; //  721 :  99 - 0x63
      10'h2D2: dout <= 8'b01100100; //  722 : 100 - 0x64
      10'h2D3: dout <= 8'b01100101; //  723 : 101 - 0x65
      10'h2D4: dout <= 8'b01100001; //  724 :  97 - 0x61
      10'h2D5: dout <= 8'b01100100; //  725 : 100 - 0x64
      10'h2D6: dout <= 8'b00000000; //  726 :   0 - 0x0
      10'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      10'h2D8: dout <= 8'b00000000; //  728 :   0 - 0x0
      10'h2D9: dout <= 8'b00000000; //  729 :   0 - 0x0
      10'h2DA: dout <= 8'b00000000; //  730 :   0 - 0x0
      10'h2DB: dout <= 8'b00000000; //  731 :   0 - 0x0
      10'h2DC: dout <= 8'b00000000; //  732 :   0 - 0x0
      10'h2DD: dout <= 8'b00000000; //  733 :   0 - 0x0
      10'h2DE: dout <= 8'b00000000; //  734 :   0 - 0x0
      10'h2DF: dout <= 8'b00000000; //  735 :   0 - 0x0
      10'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- line 0x17
      10'h2E1: dout <= 8'b00000000; //  737 :   0 - 0x0
      10'h2E2: dout <= 8'b00000000; //  738 :   0 - 0x0
      10'h2E3: dout <= 8'b00000000; //  739 :   0 - 0x0
      10'h2E4: dout <= 8'b00000000; //  740 :   0 - 0x0
      10'h2E5: dout <= 8'b00000000; //  741 :   0 - 0x0
      10'h2E6: dout <= 8'b00000000; //  742 :   0 - 0x0
      10'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      10'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0
      10'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      10'h2EA: dout <= 8'b00000000; //  746 :   0 - 0x0
      10'h2EB: dout <= 8'b00000000; //  747 :   0 - 0x0
      10'h2EC: dout <= 8'b00000000; //  748 :   0 - 0x0
      10'h2ED: dout <= 8'b00000000; //  749 :   0 - 0x0
      10'h2EE: dout <= 8'b00000000; //  750 :   0 - 0x0
      10'h2EF: dout <= 8'b00000000; //  751 :   0 - 0x0
      10'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0
      10'h2F1: dout <= 8'b00000000; //  753 :   0 - 0x0
      10'h2F2: dout <= 8'b00000000; //  754 :   0 - 0x0
      10'h2F3: dout <= 8'b00000000; //  755 :   0 - 0x0
      10'h2F4: dout <= 8'b00000000; //  756 :   0 - 0x0
      10'h2F5: dout <= 8'b00000000; //  757 :   0 - 0x0
      10'h2F6: dout <= 8'b00000000; //  758 :   0 - 0x0
      10'h2F7: dout <= 8'b00000000; //  759 :   0 - 0x0
      10'h2F8: dout <= 8'b00000000; //  760 :   0 - 0x0
      10'h2F9: dout <= 8'b00000000; //  761 :   0 - 0x0
      10'h2FA: dout <= 8'b00000000; //  762 :   0 - 0x0
      10'h2FB: dout <= 8'b00000000; //  763 :   0 - 0x0
      10'h2FC: dout <= 8'b00000000; //  764 :   0 - 0x0
      10'h2FD: dout <= 8'b00000000; //  765 :   0 - 0x0
      10'h2FE: dout <= 8'b00000000; //  766 :   0 - 0x0
      10'h2FF: dout <= 8'b00000000; //  767 :   0 - 0x0
      10'h300: dout <= 8'b00000000; //  768 :   0 - 0x0 -- line 0x18
      10'h301: dout <= 8'b00000000; //  769 :   0 - 0x0
      10'h302: dout <= 8'b00000000; //  770 :   0 - 0x0
      10'h303: dout <= 8'b00000000; //  771 :   0 - 0x0
      10'h304: dout <= 8'b00000000; //  772 :   0 - 0x0
      10'h305: dout <= 8'b00000000; //  773 :   0 - 0x0
      10'h306: dout <= 8'b00000000; //  774 :   0 - 0x0
      10'h307: dout <= 8'b00000000; //  775 :   0 - 0x0
      10'h308: dout <= 8'b00000000; //  776 :   0 - 0x0
      10'h309: dout <= 8'b00000000; //  777 :   0 - 0x0
      10'h30A: dout <= 8'b00000000; //  778 :   0 - 0x0
      10'h30B: dout <= 8'b00000000; //  779 :   0 - 0x0
      10'h30C: dout <= 8'b00000000; //  780 :   0 - 0x0
      10'h30D: dout <= 8'b00000000; //  781 :   0 - 0x0
      10'h30E: dout <= 8'b00000000; //  782 :   0 - 0x0
      10'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      10'h310: dout <= 8'b00000000; //  784 :   0 - 0x0
      10'h311: dout <= 8'b00000000; //  785 :   0 - 0x0
      10'h312: dout <= 8'b00000000; //  786 :   0 - 0x0
      10'h313: dout <= 8'b00000000; //  787 :   0 - 0x0
      10'h314: dout <= 8'b00000000; //  788 :   0 - 0x0
      10'h315: dout <= 8'b00000000; //  789 :   0 - 0x0
      10'h316: dout <= 8'b00000000; //  790 :   0 - 0x0
      10'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      10'h318: dout <= 8'b00000000; //  792 :   0 - 0x0
      10'h319: dout <= 8'b00000000; //  793 :   0 - 0x0
      10'h31A: dout <= 8'b00000000; //  794 :   0 - 0x0
      10'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      10'h31C: dout <= 8'b00000000; //  796 :   0 - 0x0
      10'h31D: dout <= 8'b00000000; //  797 :   0 - 0x0
      10'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      10'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      10'h320: dout <= 8'b10010010; //  800 : 146 - 0x92 -- line 0x19
      10'h321: dout <= 8'b10010011; //  801 : 147 - 0x93
      10'h322: dout <= 8'b10010010; //  802 : 146 - 0x92
      10'h323: dout <= 8'b10000011; //  803 : 131 - 0x83
      10'h324: dout <= 8'b10010010; //  804 : 146 - 0x92
      10'h325: dout <= 8'b10010011; //  805 : 147 - 0x93
      10'h326: dout <= 8'b10000010; //  806 : 130 - 0x82
      10'h327: dout <= 8'b10010011; //  807 : 147 - 0x93
      10'h328: dout <= 8'b10010010; //  808 : 146 - 0x92
      10'h329: dout <= 8'b10010010; //  809 : 146 - 0x92
      10'h32A: dout <= 8'b10010011; //  810 : 147 - 0x93
      10'h32B: dout <= 8'b10010000; //  811 : 144 - 0x90
      10'h32C: dout <= 8'b10010010; //  812 : 146 - 0x92
      10'h32D: dout <= 8'b10000010; //  813 : 130 - 0x82
      10'h32E: dout <= 8'b10010000; //  814 : 144 - 0x90
      10'h32F: dout <= 8'b10010011; //  815 : 147 - 0x93
      10'h330: dout <= 8'b10010010; //  816 : 146 - 0x92
      10'h331: dout <= 8'b10010011; //  817 : 147 - 0x93
      10'h332: dout <= 8'b10000011; //  818 : 131 - 0x83
      10'h333: dout <= 8'b10010011; //  819 : 147 - 0x93
      10'h334: dout <= 8'b10010011; //  820 : 147 - 0x93
      10'h335: dout <= 8'b10010000; //  821 : 144 - 0x90
      10'h336: dout <= 8'b10010010; //  822 : 146 - 0x92
      10'h337: dout <= 8'b10010011; //  823 : 147 - 0x93
      10'h338: dout <= 8'b10010010; //  824 : 146 - 0x92
      10'h339: dout <= 8'b01001010; //  825 :  74 - 0x4a
      10'h33A: dout <= 8'b01001011; //  826 :  75 - 0x4b
      10'h33B: dout <= 8'b01001100; //  827 :  76 - 0x4c
      10'h33C: dout <= 8'b01001101; //  828 :  77 - 0x4d
      10'h33D: dout <= 8'b01001110; //  829 :  78 - 0x4e
      10'h33E: dout <= 8'b01001111; //  830 :  79 - 0x4f
      10'h33F: dout <= 8'b10010010; //  831 : 146 - 0x92
      10'h340: dout <= 8'b10000100; //  832 : 132 - 0x84 -- line 0x1a
      10'h341: dout <= 8'b10000101; //  833 : 133 - 0x85
      10'h342: dout <= 8'b10000100; //  834 : 132 - 0x84
      10'h343: dout <= 8'b10000101; //  835 : 133 - 0x85
      10'h344: dout <= 8'b10000100; //  836 : 132 - 0x84
      10'h345: dout <= 8'b10000101; //  837 : 133 - 0x85
      10'h346: dout <= 8'b10000100; //  838 : 132 - 0x84
      10'h347: dout <= 8'b10000101; //  839 : 133 - 0x85
      10'h348: dout <= 8'b10000100; //  840 : 132 - 0x84
      10'h349: dout <= 8'b10000101; //  841 : 133 - 0x85
      10'h34A: dout <= 8'b10000100; //  842 : 132 - 0x84
      10'h34B: dout <= 8'b10000101; //  843 : 133 - 0x85
      10'h34C: dout <= 8'b10000100; //  844 : 132 - 0x84
      10'h34D: dout <= 8'b10000101; //  845 : 133 - 0x85
      10'h34E: dout <= 8'b10000100; //  846 : 132 - 0x84
      10'h34F: dout <= 8'b10000101; //  847 : 133 - 0x85
      10'h350: dout <= 8'b10000100; //  848 : 132 - 0x84
      10'h351: dout <= 8'b10000101; //  849 : 133 - 0x85
      10'h352: dout <= 8'b10000100; //  850 : 132 - 0x84
      10'h353: dout <= 8'b10000101; //  851 : 133 - 0x85
      10'h354: dout <= 8'b10000100; //  852 : 132 - 0x84
      10'h355: dout <= 8'b10000101; //  853 : 133 - 0x85
      10'h356: dout <= 8'b10000100; //  854 : 132 - 0x84
      10'h357: dout <= 8'b10000101; //  855 : 133 - 0x85
      10'h358: dout <= 8'b10000100; //  856 : 132 - 0x84
      10'h359: dout <= 8'b10000101; //  857 : 133 - 0x85
      10'h35A: dout <= 8'b10000100; //  858 : 132 - 0x84
      10'h35B: dout <= 8'b10000101; //  859 : 133 - 0x85
      10'h35C: dout <= 8'b10000100; //  860 : 132 - 0x84
      10'h35D: dout <= 8'b10000101; //  861 : 133 - 0x85
      10'h35E: dout <= 8'b10000100; //  862 : 132 - 0x84
      10'h35F: dout <= 8'b10000101; //  863 : 133 - 0x85
      10'h360: dout <= 8'b10010100; //  864 : 148 - 0x94 -- line 0x1b
      10'h361: dout <= 8'b10010111; //  865 : 151 - 0x97
      10'h362: dout <= 8'b10010100; //  866 : 148 - 0x94
      10'h363: dout <= 8'b10010101; //  867 : 149 - 0x95
      10'h364: dout <= 8'b10010100; //  868 : 148 - 0x94
      10'h365: dout <= 8'b10000111; //  869 : 135 - 0x87
      10'h366: dout <= 8'b10010111; //  870 : 151 - 0x97
      10'h367: dout <= 8'b10010111; //  871 : 151 - 0x97
      10'h368: dout <= 8'b10010100; //  872 : 148 - 0x94
      10'h369: dout <= 8'b10000110; //  873 : 134 - 0x86
      10'h36A: dout <= 8'b10010100; //  874 : 148 - 0x94
      10'h36B: dout <= 8'b10010101; //  875 : 149 - 0x95
      10'h36C: dout <= 8'b10010110; //  876 : 150 - 0x96
      10'h36D: dout <= 8'b10010101; //  877 : 149 - 0x95
      10'h36E: dout <= 8'b10010100; //  878 : 148 - 0x94
      10'h36F: dout <= 8'b10010101; //  879 : 149 - 0x95
      10'h370: dout <= 8'b10000111; //  880 : 135 - 0x87
      10'h371: dout <= 8'b10010111; //  881 : 151 - 0x97
      10'h372: dout <= 8'b10010100; //  882 : 148 - 0x94
      10'h373: dout <= 8'b10000111; //  883 : 135 - 0x87
      10'h374: dout <= 8'b10010110; //  884 : 150 - 0x96
      10'h375: dout <= 8'b10000110; //  885 : 134 - 0x86
      10'h376: dout <= 8'b10010100; //  886 : 148 - 0x94
      10'h377: dout <= 8'b10010101; //  887 : 149 - 0x95
      10'h378: dout <= 8'b10000111; //  888 : 135 - 0x87
      10'h379: dout <= 8'b10010101; //  889 : 149 - 0x95
      10'h37A: dout <= 8'b10010100; //  890 : 148 - 0x94
      10'h37B: dout <= 8'b10010111; //  891 : 151 - 0x97
      10'h37C: dout <= 8'b10010100; //  892 : 148 - 0x94
      10'h37D: dout <= 8'b10000110; //  893 : 134 - 0x86
      10'h37E: dout <= 8'b10010100; //  894 : 148 - 0x94
      10'h37F: dout <= 8'b10010101; //  895 : 149 - 0x95
      10'h380: dout <= 8'b10000100; //  896 : 132 - 0x84 -- line 0x1c
      10'h381: dout <= 8'b10000101; //  897 : 133 - 0x85
      10'h382: dout <= 8'b10010110; //  898 : 150 - 0x96
      10'h383: dout <= 8'b10000101; //  899 : 133 - 0x85
      10'h384: dout <= 8'b10000111; //  900 : 135 - 0x87
      10'h385: dout <= 8'b10010111; //  901 : 151 - 0x97
      10'h386: dout <= 8'b10000100; //  902 : 132 - 0x84
      10'h387: dout <= 8'b10000101; //  903 : 133 - 0x85
      10'h388: dout <= 8'b10000100; //  904 : 132 - 0x84
      10'h389: dout <= 8'b10000101; //  905 : 133 - 0x85
      10'h38A: dout <= 8'b10000100; //  906 : 132 - 0x84
      10'h38B: dout <= 8'b10000111; //  907 : 135 - 0x87
      10'h38C: dout <= 8'b10000100; //  908 : 132 - 0x84
      10'h38D: dout <= 8'b10000110; //  909 : 134 - 0x86
      10'h38E: dout <= 8'b10000100; //  910 : 132 - 0x84
      10'h38F: dout <= 8'b10000101; //  911 : 133 - 0x85
      10'h390: dout <= 8'b10000100; //  912 : 132 - 0x84
      10'h391: dout <= 8'b10000101; //  913 : 133 - 0x85
      10'h392: dout <= 8'b10000100; //  914 : 132 - 0x84
      10'h393: dout <= 8'b10000101; //  915 : 133 - 0x85
      10'h394: dout <= 8'b10000100; //  916 : 132 - 0x84
      10'h395: dout <= 8'b10000101; //  917 : 133 - 0x85
      10'h396: dout <= 8'b10010111; //  918 : 151 - 0x97
      10'h397: dout <= 8'b10000101; //  919 : 133 - 0x85
      10'h398: dout <= 8'b10000100; //  920 : 132 - 0x84
      10'h399: dout <= 8'b10010111; //  921 : 151 - 0x97
      10'h39A: dout <= 8'b10000111; //  922 : 135 - 0x87
      10'h39B: dout <= 8'b10000101; //  923 : 133 - 0x85
      10'h39C: dout <= 8'b10000110; //  924 : 134 - 0x86
      10'h39D: dout <= 8'b10000111; //  925 : 135 - 0x87
      10'h39E: dout <= 8'b10000100; //  926 : 132 - 0x84
      10'h39F: dout <= 8'b10000101; //  927 : 133 - 0x85
      10'h3A0: dout <= 8'b10010100; //  928 : 148 - 0x94 -- line 0x1d
      10'h3A1: dout <= 8'b10010101; //  929 : 149 - 0x95
      10'h3A2: dout <= 8'b10010100; //  930 : 148 - 0x94
      10'h3A3: dout <= 8'b10010101; //  931 : 149 - 0x95
      10'h3A4: dout <= 8'b10010100; //  932 : 148 - 0x94
      10'h3A5: dout <= 8'b10000110; //  933 : 134 - 0x86
      10'h3A6: dout <= 8'b10010100; //  934 : 148 - 0x94
      10'h3A7: dout <= 8'b10010101; //  935 : 149 - 0x95
      10'h3A8: dout <= 8'b10010100; //  936 : 148 - 0x94
      10'h3A9: dout <= 8'b10010101; //  937 : 149 - 0x95
      10'h3AA: dout <= 8'b10010100; //  938 : 148 - 0x94
      10'h3AB: dout <= 8'b10010101; //  939 : 149 - 0x95
      10'h3AC: dout <= 8'b10010100; //  940 : 148 - 0x94
      10'h3AD: dout <= 8'b10010111; //  941 : 151 - 0x97
      10'h3AE: dout <= 8'b10010110; //  942 : 150 - 0x96
      10'h3AF: dout <= 8'b10010101; //  943 : 149 - 0x95
      10'h3B0: dout <= 8'b10010100; //  944 : 148 - 0x94
      10'h3B1: dout <= 8'b10010101; //  945 : 149 - 0x95
      10'h3B2: dout <= 8'b10010100; //  946 : 148 - 0x94
      10'h3B3: dout <= 8'b10010101; //  947 : 149 - 0x95
      10'h3B4: dout <= 8'b10010100; //  948 : 148 - 0x94
      10'h3B5: dout <= 8'b10010101; //  949 : 149 - 0x95
      10'h3B6: dout <= 8'b10010100; //  950 : 148 - 0x94
      10'h3B7: dout <= 8'b10010101; //  951 : 149 - 0x95
      10'h3B8: dout <= 8'b10000110; //  952 : 134 - 0x86
      10'h3B9: dout <= 8'b10010101; //  953 : 149 - 0x95
      10'h3BA: dout <= 8'b10010100; //  954 : 148 - 0x94
      10'h3BB: dout <= 8'b10010101; //  955 : 149 - 0x95
      10'h3BC: dout <= 8'b10010100; //  956 : 148 - 0x94
      10'h3BD: dout <= 8'b10010101; //  957 : 149 - 0x95
      10'h3BE: dout <= 8'b10010100; //  958 : 148 - 0x94
      10'h3BF: dout <= 8'b10010101; //  959 : 149 - 0x95
        //-- Attribute Table 0----
      10'h3C0: dout <= 8'b10101010; //  960 : 170 - 0xaa
      10'h3C1: dout <= 8'b10101010; //  961 : 170 - 0xaa
      10'h3C2: dout <= 8'b10101010; //  962 : 170 - 0xaa
      10'h3C3: dout <= 8'b10101010; //  963 : 170 - 0xaa
      10'h3C4: dout <= 8'b10101010; //  964 : 170 - 0xaa
      10'h3C5: dout <= 8'b10101010; //  965 : 170 - 0xaa
      10'h3C6: dout <= 8'b10101010; //  966 : 170 - 0xaa
      10'h3C7: dout <= 8'b10101010; //  967 : 170 - 0xaa
      10'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0
      10'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      10'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      10'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      10'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      10'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      10'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      10'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      10'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0
      10'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      10'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      10'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      10'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      10'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      10'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      10'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      10'h3D8: dout <= 8'b01010101; //  984 :  85 - 0x55
      10'h3D9: dout <= 8'b01010101; //  985 :  85 - 0x55
      10'h3DA: dout <= 8'b01010101; //  986 :  85 - 0x55
      10'h3DB: dout <= 8'b01010101; //  987 :  85 - 0x55
      10'h3DC: dout <= 8'b01010101; //  988 :  85 - 0x55
      10'h3DD: dout <= 8'b01010101; //  989 :  85 - 0x55
      10'h3DE: dout <= 8'b01010101; //  990 :  85 - 0x55
      10'h3DF: dout <= 8'b01010101; //  991 :  85 - 0x55
      10'h3E0: dout <= 8'b01010101; //  992 :  85 - 0x55
      10'h3E1: dout <= 8'b01010101; //  993 :  85 - 0x55
      10'h3E2: dout <= 8'b01010101; //  994 :  85 - 0x55
      10'h3E3: dout <= 8'b01010101; //  995 :  85 - 0x55
      10'h3E4: dout <= 8'b01010101; //  996 :  85 - 0x55
      10'h3E5: dout <= 8'b01010101; //  997 :  85 - 0x55
      10'h3E6: dout <= 8'b01010101; //  998 :  85 - 0x55
      10'h3E7: dout <= 8'b01010101; //  999 :  85 - 0x55
      10'h3E8: dout <= 8'b00000101; // 1000 :   5 - 0x5
      10'h3E9: dout <= 8'b10000101; // 1001 : 133 - 0x85
      10'h3EA: dout <= 8'b11101101; // 1002 : 237 - 0xed
      10'h3EB: dout <= 8'b11111111; // 1003 : 255 - 0xff
      10'h3EC: dout <= 8'b11111111; // 1004 : 255 - 0xff
      10'h3ED: dout <= 8'b00110111; // 1005 :  55 - 0x37
      10'h3EE: dout <= 8'b00000101; // 1006 :   5 - 0x5
      10'h3EF: dout <= 8'b00000101; // 1007 :   5 - 0x5
      10'h3F0: dout <= 8'b10101010; // 1008 : 170 - 0xaa
      10'h3F1: dout <= 8'b10101010; // 1009 : 170 - 0xaa
      10'h3F2: dout <= 8'b10101010; // 1010 : 170 - 0xaa
      10'h3F3: dout <= 8'b10101010; // 1011 : 170 - 0xaa
      10'h3F4: dout <= 8'b10101010; // 1012 : 170 - 0xaa
      10'h3F5: dout <= 8'b10101010; // 1013 : 170 - 0xaa
      10'h3F6: dout <= 8'b10101010; // 1014 : 170 - 0xaa
      10'h3F7: dout <= 8'b10101010; // 1015 : 170 - 0xaa
      10'h3F8: dout <= 8'b00001010; // 1016 :  10 - 0xa
      10'h3F9: dout <= 8'b00001010; // 1017 :  10 - 0xa
      10'h3FA: dout <= 8'b00001010; // 1018 :  10 - 0xa
      10'h3FB: dout <= 8'b00001010; // 1019 :  10 - 0xa
      10'h3FC: dout <= 8'b00001010; // 1020 :  10 - 0xa
      10'h3FD: dout <= 8'b00001010; // 1021 :  10 - 0xa
      10'h3FE: dout <= 8'b00001010; // 1022 :  10 - 0xa
      10'h3FF: dout <= 8'b00001010; // 1023 :  10 - 0xa
    endcase
  end

endmodule
