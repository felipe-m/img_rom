--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables


---  Original memory dump file name: nova_ntable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_NOVA_00 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_NOVA_00;

architecture BEHAVIORAL of ROM_NTABLE_NOVA_00 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "00110000", --    0 -  0x0  :   48 - 0x30 -- line 0x0
    "00111111", --    1 -  0x1  :   63 - 0x3f
    "00110000", --    2 -  0x2  :   48 - 0x30
    "00111111", --    3 -  0x3  :   63 - 0x3f
    "00110000", --    4 -  0x4  :   48 - 0x30
    "00111111", --    5 -  0x5  :   63 - 0x3f
    "00110000", --    6 -  0x6  :   48 - 0x30
    "00111111", --    7 -  0x7  :   63 - 0x3f
    "00110000", --    8 -  0x8  :   48 - 0x30
    "00111111", --    9 -  0x9  :   63 - 0x3f
    "00110000", --   10 -  0xa  :   48 - 0x30
    "00111111", --   11 -  0xb  :   63 - 0x3f
    "00110000", --   12 -  0xc  :   48 - 0x30
    "00111111", --   13 -  0xd  :   63 - 0x3f
    "00110000", --   14 -  0xe  :   48 - 0x30
    "00111111", --   15 -  0xf  :   63 - 0x3f
    "00110000", --   16 - 0x10  :   48 - 0x30
    "00111111", --   17 - 0x11  :   63 - 0x3f
    "00110000", --   18 - 0x12  :   48 - 0x30
    "00111111", --   19 - 0x13  :   63 - 0x3f
    "01110000", --   20 - 0x14  :  112 - 0x70
    "01110001", --   21 - 0x15  :  113 - 0x71
    "01110001", --   22 - 0x16  :  113 - 0x71
    "01110001", --   23 - 0x17  :  113 - 0x71
    "01110001", --   24 - 0x18  :  113 - 0x71
    "01110001", --   25 - 0x19  :  113 - 0x71
    "01110001", --   26 - 0x1a  :  113 - 0x71
    "01110001", --   27 - 0x1b  :  113 - 0x71
    "01110001", --   28 - 0x1c  :  113 - 0x71
    "01110001", --   29 - 0x1d  :  113 - 0x71
    "01110001", --   30 - 0x1e  :  113 - 0x71
    "01110001", --   31 - 0x1f  :  113 - 0x71
    "00111111", --   32 - 0x20  :   63 - 0x3f -- line 0x1
    "00110000", --   33 - 0x21  :   48 - 0x30
    "00111111", --   34 - 0x22  :   63 - 0x3f
    "00110000", --   35 - 0x23  :   48 - 0x30
    "00111111", --   36 - 0x24  :   63 - 0x3f
    "00110000", --   37 - 0x25  :   48 - 0x30
    "00111111", --   38 - 0x26  :   63 - 0x3f
    "00110000", --   39 - 0x27  :   48 - 0x30
    "00111111", --   40 - 0x28  :   63 - 0x3f
    "00110000", --   41 - 0x29  :   48 - 0x30
    "00111111", --   42 - 0x2a  :   63 - 0x3f
    "00110000", --   43 - 0x2b  :   48 - 0x30
    "00111111", --   44 - 0x2c  :   63 - 0x3f
    "00110000", --   45 - 0x2d  :   48 - 0x30
    "00111111", --   46 - 0x2e  :   63 - 0x3f
    "00110000", --   47 - 0x2f  :   48 - 0x30
    "00111111", --   48 - 0x30  :   63 - 0x3f
    "00110000", --   49 - 0x31  :   48 - 0x30
    "00111111", --   50 - 0x32  :   63 - 0x3f
    "00110000", --   51 - 0x33  :   48 - 0x30
    "01100000", --   52 - 0x34  :   96 - 0x60
    "01110111", --   53 - 0x35  :  119 - 0x77
    "01110111", --   54 - 0x36  :  119 - 0x77
    "01110111", --   55 - 0x37  :  119 - 0x77
    "01110111", --   56 - 0x38  :  119 - 0x77
    "01110111", --   57 - 0x39  :  119 - 0x77
    "01110111", --   58 - 0x3a  :  119 - 0x77
    "01110111", --   59 - 0x3b  :  119 - 0x77
    "01110111", --   60 - 0x3c  :  119 - 0x77
    "01110111", --   61 - 0x3d  :  119 - 0x77
    "01110111", --   62 - 0x3e  :  119 - 0x77
    "01110111", --   63 - 0x3f  :  119 - 0x77
    "00110000", --   64 - 0x40  :   48 - 0x30 -- line 0x2
    "00111111", --   65 - 0x41  :   63 - 0x3f
    "00110000", --   66 - 0x42  :   48 - 0x30
    "00111111", --   67 - 0x43  :   63 - 0x3f
    "00110000", --   68 - 0x44  :   48 - 0x30
    "00111111", --   69 - 0x45  :   63 - 0x3f
    "00110000", --   70 - 0x46  :   48 - 0x30
    "00111111", --   71 - 0x47  :   63 - 0x3f
    "00110000", --   72 - 0x48  :   48 - 0x30
    "00111111", --   73 - 0x49  :   63 - 0x3f
    "00110000", --   74 - 0x4a  :   48 - 0x30
    "00111111", --   75 - 0x4b  :   63 - 0x3f
    "00110000", --   76 - 0x4c  :   48 - 0x30
    "00111111", --   77 - 0x4d  :   63 - 0x3f
    "00110000", --   78 - 0x4e  :   48 - 0x30
    "00111111", --   79 - 0x4f  :   63 - 0x3f
    "00110000", --   80 - 0x50  :   48 - 0x30
    "00111111", --   81 - 0x51  :   63 - 0x3f
    "00110000", --   82 - 0x52  :   48 - 0x30
    "00111111", --   83 - 0x53  :   63 - 0x3f
    "00111001", --   84 - 0x54  :   57 - 0x39
    "00111001", --   85 - 0x55  :   57 - 0x39
    "00111001", --   86 - 0x56  :   57 - 0x39
    "00111001", --   87 - 0x57  :   57 - 0x39
    "00111001", --   88 - 0x58  :   57 - 0x39
    "00111001", --   89 - 0x59  :   57 - 0x39
    "00111001", --   90 - 0x5a  :   57 - 0x39
    "00111001", --   91 - 0x5b  :   57 - 0x39
    "00111001", --   92 - 0x5c  :   57 - 0x39
    "00111001", --   93 - 0x5d  :   57 - 0x39
    "00111001", --   94 - 0x5e  :   57 - 0x39
    "00111001", --   95 - 0x5f  :   57 - 0x39
    "00111111", --   96 - 0x60  :   63 - 0x3f -- line 0x3
    "00110000", --   97 - 0x61  :   48 - 0x30
    "00111111", --   98 - 0x62  :   63 - 0x3f
    "00110000", --   99 - 0x63  :   48 - 0x30
    "00111111", --  100 - 0x64  :   63 - 0x3f
    "00110000", --  101 - 0x65  :   48 - 0x30
    "00111111", --  102 - 0x66  :   63 - 0x3f
    "00110000", --  103 - 0x67  :   48 - 0x30
    "00111111", --  104 - 0x68  :   63 - 0x3f
    "00110000", --  105 - 0x69  :   48 - 0x30
    "00111111", --  106 - 0x6a  :   63 - 0x3f
    "00110000", --  107 - 0x6b  :   48 - 0x30
    "00111111", --  108 - 0x6c  :   63 - 0x3f
    "00110000", --  109 - 0x6d  :   48 - 0x30
    "00111111", --  110 - 0x6e  :   63 - 0x3f
    "00110000", --  111 - 0x6f  :   48 - 0x30
    "00111111", --  112 - 0x70  :   63 - 0x3f
    "00110000", --  113 - 0x71  :   48 - 0x30
    "00111111", --  114 - 0x72  :   63 - 0x3f
    "00110000", --  115 - 0x73  :   48 - 0x30
    "00111111", --  116 - 0x74  :   63 - 0x3f
    "00111111", --  117 - 0x75  :   63 - 0x3f
    "00111111", --  118 - 0x76  :   63 - 0x3f
    "00111111", --  119 - 0x77  :   63 - 0x3f
    "00111111", --  120 - 0x78  :   63 - 0x3f
    "00111111", --  121 - 0x79  :   63 - 0x3f
    "00111111", --  122 - 0x7a  :   63 - 0x3f
    "00111111", --  123 - 0x7b  :   63 - 0x3f
    "00111111", --  124 - 0x7c  :   63 - 0x3f
    "00111111", --  125 - 0x7d  :   63 - 0x3f
    "00111111", --  126 - 0x7e  :   63 - 0x3f
    "00111111", --  127 - 0x7f  :   63 - 0x3f
    "00111111", --  128 - 0x80  :   63 - 0x3f -- line 0x4
    "00111111", --  129 - 0x81  :   63 - 0x3f
    "00111111", --  130 - 0x82  :   63 - 0x3f
    "00111111", --  131 - 0x83  :   63 - 0x3f
    "00111111", --  132 - 0x84  :   63 - 0x3f
    "00111111", --  133 - 0x85  :   63 - 0x3f
    "00111111", --  134 - 0x86  :   63 - 0x3f
    "00111111", --  135 - 0x87  :   63 - 0x3f
    "00111111", --  136 - 0x88  :   63 - 0x3f
    "00111111", --  137 - 0x89  :   63 - 0x3f
    "00111111", --  138 - 0x8a  :   63 - 0x3f
    "00111111", --  139 - 0x8b  :   63 - 0x3f
    "00111111", --  140 - 0x8c  :   63 - 0x3f
    "00111111", --  141 - 0x8d  :   63 - 0x3f
    "00111111", --  142 - 0x8e  :   63 - 0x3f
    "00111111", --  143 - 0x8f  :   63 - 0x3f
    "00111111", --  144 - 0x90  :   63 - 0x3f
    "00111111", --  145 - 0x91  :   63 - 0x3f
    "00111111", --  146 - 0x92  :   63 - 0x3f
    "00111111", --  147 - 0x93  :   63 - 0x3f
    "00111111", --  148 - 0x94  :   63 - 0x3f
    "00111111", --  149 - 0x95  :   63 - 0x3f
    "00111111", --  150 - 0x96  :   63 - 0x3f
    "00111111", --  151 - 0x97  :   63 - 0x3f
    "00111111", --  152 - 0x98  :   63 - 0x3f
    "00111111", --  153 - 0x99  :   63 - 0x3f
    "00000100", --  154 - 0x9a  :    4 - 0x4
    "00000110", --  155 - 0x9b  :    6 - 0x6
    "00111111", --  156 - 0x9c  :   63 - 0x3f
    "00111111", --  157 - 0x9d  :   63 - 0x3f
    "00010100", --  158 - 0x9e  :   20 - 0x14
    "00010110", --  159 - 0x9f  :   22 - 0x16
    "00111111", --  160 - 0xa0  :   63 - 0x3f -- line 0x5
    "00111111", --  161 - 0xa1  :   63 - 0x3f
    "00111111", --  162 - 0xa2  :   63 - 0x3f
    "00111111", --  163 - 0xa3  :   63 - 0x3f
    "00111111", --  164 - 0xa4  :   63 - 0x3f
    "00111111", --  165 - 0xa5  :   63 - 0x3f
    "00111111", --  166 - 0xa6  :   63 - 0x3f
    "00111111", --  167 - 0xa7  :   63 - 0x3f
    "00111111", --  168 - 0xa8  :   63 - 0x3f
    "00111111", --  169 - 0xa9  :   63 - 0x3f
    "00111111", --  170 - 0xaa  :   63 - 0x3f
    "00111111", --  171 - 0xab  :   63 - 0x3f
    "00111111", --  172 - 0xac  :   63 - 0x3f
    "00111111", --  173 - 0xad  :   63 - 0x3f
    "00111111", --  174 - 0xae  :   63 - 0x3f
    "00111111", --  175 - 0xaf  :   63 - 0x3f
    "00111111", --  176 - 0xb0  :   63 - 0x3f
    "00111111", --  177 - 0xb1  :   63 - 0x3f
    "00111111", --  178 - 0xb2  :   63 - 0x3f
    "00111111", --  179 - 0xb3  :   63 - 0x3f
    "00111111", --  180 - 0xb4  :   63 - 0x3f
    "00111111", --  181 - 0xb5  :   63 - 0x3f
    "00111111", --  182 - 0xb6  :   63 - 0x3f
    "00111111", --  183 - 0xb7  :   63 - 0x3f
    "00111111", --  184 - 0xb8  :   63 - 0x3f
    "00111111", --  185 - 0xb9  :   63 - 0x3f
    "00000101", --  186 - 0xba  :    5 - 0x5
    "00000111", --  187 - 0xbb  :    7 - 0x7
    "00111111", --  188 - 0xbc  :   63 - 0x3f
    "00111111", --  189 - 0xbd  :   63 - 0x3f
    "00010101", --  190 - 0xbe  :   21 - 0x15
    "00010111", --  191 - 0xbf  :   23 - 0x17
    "00111111", --  192 - 0xc0  :   63 - 0x3f -- line 0x6
    "00111111", --  193 - 0xc1  :   63 - 0x3f
    "00111111", --  194 - 0xc2  :   63 - 0x3f
    "00111111", --  195 - 0xc3  :   63 - 0x3f
    "00111111", --  196 - 0xc4  :   63 - 0x3f
    "00111111", --  197 - 0xc5  :   63 - 0x3f
    "00111111", --  198 - 0xc6  :   63 - 0x3f
    "00111111", --  199 - 0xc7  :   63 - 0x3f
    "00111111", --  200 - 0xc8  :   63 - 0x3f
    "00111111", --  201 - 0xc9  :   63 - 0x3f
    "00111111", --  202 - 0xca  :   63 - 0x3f
    "00111111", --  203 - 0xcb  :   63 - 0x3f
    "00111111", --  204 - 0xcc  :   63 - 0x3f
    "00111111", --  205 - 0xcd  :   63 - 0x3f
    "00111111", --  206 - 0xce  :   63 - 0x3f
    "00111111", --  207 - 0xcf  :   63 - 0x3f
    "00111111", --  208 - 0xd0  :   63 - 0x3f
    "00111111", --  209 - 0xd1  :   63 - 0x3f
    "00111111", --  210 - 0xd2  :   63 - 0x3f
    "00111111", --  211 - 0xd3  :   63 - 0x3f
    "00111111", --  212 - 0xd4  :   63 - 0x3f
    "00111111", --  213 - 0xd5  :   63 - 0x3f
    "00111111", --  214 - 0xd6  :   63 - 0x3f
    "00111111", --  215 - 0xd7  :   63 - 0x3f
    "00111111", --  216 - 0xd8  :   63 - 0x3f
    "00111111", --  217 - 0xd9  :   63 - 0x3f
    "00111111", --  218 - 0xda  :   63 - 0x3f
    "00111111", --  219 - 0xdb  :   63 - 0x3f
    "00111111", --  220 - 0xdc  :   63 - 0x3f
    "00111111", --  221 - 0xdd  :   63 - 0x3f
    "00111111", --  222 - 0xde  :   63 - 0x3f
    "00111111", --  223 - 0xdf  :   63 - 0x3f
    "00111111", --  224 - 0xe0  :   63 - 0x3f -- line 0x7
    "00111111", --  225 - 0xe1  :   63 - 0x3f
    "00111111", --  226 - 0xe2  :   63 - 0x3f
    "00111111", --  227 - 0xe3  :   63 - 0x3f
    "00111111", --  228 - 0xe4  :   63 - 0x3f
    "00111111", --  229 - 0xe5  :   63 - 0x3f
    "00111111", --  230 - 0xe6  :   63 - 0x3f
    "00111111", --  231 - 0xe7  :   63 - 0x3f
    "00111111", --  232 - 0xe8  :   63 - 0x3f
    "00111111", --  233 - 0xe9  :   63 - 0x3f
    "00111111", --  234 - 0xea  :   63 - 0x3f
    "00111111", --  235 - 0xeb  :   63 - 0x3f
    "00111111", --  236 - 0xec  :   63 - 0x3f
    "00111111", --  237 - 0xed  :   63 - 0x3f
    "00111111", --  238 - 0xee  :   63 - 0x3f
    "00111111", --  239 - 0xef  :   63 - 0x3f
    "00111111", --  240 - 0xf0  :   63 - 0x3f
    "00111111", --  241 - 0xf1  :   63 - 0x3f
    "00111111", --  242 - 0xf2  :   63 - 0x3f
    "00111111", --  243 - 0xf3  :   63 - 0x3f
    "00111111", --  244 - 0xf4  :   63 - 0x3f
    "00111111", --  245 - 0xf5  :   63 - 0x3f
    "00111111", --  246 - 0xf6  :   63 - 0x3f
    "00111111", --  247 - 0xf7  :   63 - 0x3f
    "00111111", --  248 - 0xf8  :   63 - 0x3f
    "00111111", --  249 - 0xf9  :   63 - 0x3f
    "00111111", --  250 - 0xfa  :   63 - 0x3f
    "00111111", --  251 - 0xfb  :   63 - 0x3f
    "00111111", --  252 - 0xfc  :   63 - 0x3f
    "00111111", --  253 - 0xfd  :   63 - 0x3f
    "00111111", --  254 - 0xfe  :   63 - 0x3f
    "00111111", --  255 - 0xff  :   63 - 0x3f
    "00111111", --  256 - 0x100  :   63 - 0x3f -- line 0x8
    "00111111", --  257 - 0x101  :   63 - 0x3f
    "00111111", --  258 - 0x102  :   63 - 0x3f
    "00111111", --  259 - 0x103  :   63 - 0x3f
    "00111111", --  260 - 0x104  :   63 - 0x3f
    "00111111", --  261 - 0x105  :   63 - 0x3f
    "00111111", --  262 - 0x106  :   63 - 0x3f
    "00111111", --  263 - 0x107  :   63 - 0x3f
    "00111111", --  264 - 0x108  :   63 - 0x3f
    "00111111", --  265 - 0x109  :   63 - 0x3f
    "00111111", --  266 - 0x10a  :   63 - 0x3f
    "00111111", --  267 - 0x10b  :   63 - 0x3f
    "00111111", --  268 - 0x10c  :   63 - 0x3f
    "00111111", --  269 - 0x10d  :   63 - 0x3f
    "00111111", --  270 - 0x10e  :   63 - 0x3f
    "00111111", --  271 - 0x10f  :   63 - 0x3f
    "00111111", --  272 - 0x110  :   63 - 0x3f
    "00111111", --  273 - 0x111  :   63 - 0x3f
    "00111111", --  274 - 0x112  :   63 - 0x3f
    "00111111", --  275 - 0x113  :   63 - 0x3f
    "00001100", --  276 - 0x114  :   12 - 0xc
    "00001110", --  277 - 0x115  :   14 - 0xe
    "00111111", --  278 - 0x116  :   63 - 0x3f
    "00111111", --  279 - 0x117  :   63 - 0x3f
    "00111111", --  280 - 0x118  :   63 - 0x3f
    "00111111", --  281 - 0x119  :   63 - 0x3f
    "00111111", --  282 - 0x11a  :   63 - 0x3f
    "00111111", --  283 - 0x11b  :   63 - 0x3f
    "00111111", --  284 - 0x11c  :   63 - 0x3f
    "00111111", --  285 - 0x11d  :   63 - 0x3f
    "00111111", --  286 - 0x11e  :   63 - 0x3f
    "00111111", --  287 - 0x11f  :   63 - 0x3f
    "00111111", --  288 - 0x120  :   63 - 0x3f -- line 0x9
    "00111111", --  289 - 0x121  :   63 - 0x3f
    "00111111", --  290 - 0x122  :   63 - 0x3f
    "00111111", --  291 - 0x123  :   63 - 0x3f
    "00111111", --  292 - 0x124  :   63 - 0x3f
    "00111111", --  293 - 0x125  :   63 - 0x3f
    "00111111", --  294 - 0x126  :   63 - 0x3f
    "00111111", --  295 - 0x127  :   63 - 0x3f
    "00111111", --  296 - 0x128  :   63 - 0x3f
    "00111111", --  297 - 0x129  :   63 - 0x3f
    "00111111", --  298 - 0x12a  :   63 - 0x3f
    "00111111", --  299 - 0x12b  :   63 - 0x3f
    "00111111", --  300 - 0x12c  :   63 - 0x3f
    "00111111", --  301 - 0x12d  :   63 - 0x3f
    "00111111", --  302 - 0x12e  :   63 - 0x3f
    "00111111", --  303 - 0x12f  :   63 - 0x3f
    "00111111", --  304 - 0x130  :   63 - 0x3f
    "00111111", --  305 - 0x131  :   63 - 0x3f
    "00111111", --  306 - 0x132  :   63 - 0x3f
    "00111111", --  307 - 0x133  :   63 - 0x3f
    "00001101", --  308 - 0x134  :   13 - 0xd
    "00001111", --  309 - 0x135  :   15 - 0xf
    "00111111", --  310 - 0x136  :   63 - 0x3f
    "00111111", --  311 - 0x137  :   63 - 0x3f
    "00111111", --  312 - 0x138  :   63 - 0x3f
    "00111111", --  313 - 0x139  :   63 - 0x3f
    "00111111", --  314 - 0x13a  :   63 - 0x3f
    "00111111", --  315 - 0x13b  :   63 - 0x3f
    "00111111", --  316 - 0x13c  :   63 - 0x3f
    "00111111", --  317 - 0x13d  :   63 - 0x3f
    "00111111", --  318 - 0x13e  :   63 - 0x3f
    "00111111", --  319 - 0x13f  :   63 - 0x3f
    "00111111", --  320 - 0x140  :   63 - 0x3f -- line 0xa
    "00111111", --  321 - 0x141  :   63 - 0x3f
    "00111111", --  322 - 0x142  :   63 - 0x3f
    "00111111", --  323 - 0x143  :   63 - 0x3f
    "00111111", --  324 - 0x144  :   63 - 0x3f
    "00111111", --  325 - 0x145  :   63 - 0x3f
    "00111111", --  326 - 0x146  :   63 - 0x3f
    "00111111", --  327 - 0x147  :   63 - 0x3f
    "00111111", --  328 - 0x148  :   63 - 0x3f
    "00111111", --  329 - 0x149  :   63 - 0x3f
    "00111111", --  330 - 0x14a  :   63 - 0x3f
    "00111111", --  331 - 0x14b  :   63 - 0x3f
    "00111111", --  332 - 0x14c  :   63 - 0x3f
    "00111111", --  333 - 0x14d  :   63 - 0x3f
    "00111111", --  334 - 0x14e  :   63 - 0x3f
    "00111111", --  335 - 0x14f  :   63 - 0x3f
    "00111111", --  336 - 0x150  :   63 - 0x3f
    "00111111", --  337 - 0x151  :   63 - 0x3f
    "00111111", --  338 - 0x152  :   63 - 0x3f
    "00111111", --  339 - 0x153  :   63 - 0x3f
    "01010111", --  340 - 0x154  :   87 - 0x57
    "01011000", --  341 - 0x155  :   88 - 0x58
    "01011000", --  342 - 0x156  :   88 - 0x58
    "01011000", --  343 - 0x157  :   88 - 0x58
    "01011000", --  344 - 0x158  :   88 - 0x58
    "01011000", --  345 - 0x159  :   88 - 0x58
    "01011000", --  346 - 0x15a  :   88 - 0x58
    "01011000", --  347 - 0x15b  :   88 - 0x58
    "01011000", --  348 - 0x15c  :   88 - 0x58
    "01011000", --  349 - 0x15d  :   88 - 0x58
    "01011000", --  350 - 0x15e  :   88 - 0x58
    "01011000", --  351 - 0x15f  :   88 - 0x58
    "00111111", --  352 - 0x160  :   63 - 0x3f -- line 0xb
    "00111111", --  353 - 0x161  :   63 - 0x3f
    "00111111", --  354 - 0x162  :   63 - 0x3f
    "00111111", --  355 - 0x163  :   63 - 0x3f
    "00111111", --  356 - 0x164  :   63 - 0x3f
    "00111111", --  357 - 0x165  :   63 - 0x3f
    "00111111", --  358 - 0x166  :   63 - 0x3f
    "00111111", --  359 - 0x167  :   63 - 0x3f
    "00111111", --  360 - 0x168  :   63 - 0x3f
    "00111111", --  361 - 0x169  :   63 - 0x3f
    "00111111", --  362 - 0x16a  :   63 - 0x3f
    "00111111", --  363 - 0x16b  :   63 - 0x3f
    "00111111", --  364 - 0x16c  :   63 - 0x3f
    "00111111", --  365 - 0x16d  :   63 - 0x3f
    "00111111", --  366 - 0x16e  :   63 - 0x3f
    "00111111", --  367 - 0x16f  :   63 - 0x3f
    "00111111", --  368 - 0x170  :   63 - 0x3f
    "00111111", --  369 - 0x171  :   63 - 0x3f
    "00111111", --  370 - 0x172  :   63 - 0x3f
    "00111111", --  371 - 0x173  :   63 - 0x3f
    "00111111", --  372 - 0x174  :   63 - 0x3f
    "00111111", --  373 - 0x175  :   63 - 0x3f
    "00111111", --  374 - 0x176  :   63 - 0x3f
    "00111111", --  375 - 0x177  :   63 - 0x3f
    "00111111", --  376 - 0x178  :   63 - 0x3f
    "00111111", --  377 - 0x179  :   63 - 0x3f
    "00111111", --  378 - 0x17a  :   63 - 0x3f
    "00111111", --  379 - 0x17b  :   63 - 0x3f
    "00111111", --  380 - 0x17c  :   63 - 0x3f
    "00111111", --  381 - 0x17d  :   63 - 0x3f
    "00111111", --  382 - 0x17e  :   63 - 0x3f
    "00111111", --  383 - 0x17f  :   63 - 0x3f
    "00111111", --  384 - 0x180  :   63 - 0x3f -- line 0xc
    "00111111", --  385 - 0x181  :   63 - 0x3f
    "00111111", --  386 - 0x182  :   63 - 0x3f
    "00111111", --  387 - 0x183  :   63 - 0x3f
    "00111111", --  388 - 0x184  :   63 - 0x3f
    "00111111", --  389 - 0x185  :   63 - 0x3f
    "00111111", --  390 - 0x186  :   63 - 0x3f
    "00111111", --  391 - 0x187  :   63 - 0x3f
    "00111111", --  392 - 0x188  :   63 - 0x3f
    "00111111", --  393 - 0x189  :   63 - 0x3f
    "00111111", --  394 - 0x18a  :   63 - 0x3f
    "00111111", --  395 - 0x18b  :   63 - 0x3f
    "00111111", --  396 - 0x18c  :   63 - 0x3f
    "00111111", --  397 - 0x18d  :   63 - 0x3f
    "00111111", --  398 - 0x18e  :   63 - 0x3f
    "00111111", --  399 - 0x18f  :   63 - 0x3f
    "00111111", --  400 - 0x190  :   63 - 0x3f
    "00111111", --  401 - 0x191  :   63 - 0x3f
    "00111111", --  402 - 0x192  :   63 - 0x3f
    "00111111", --  403 - 0x193  :   63 - 0x3f
    "00111111", --  404 - 0x194  :   63 - 0x3f
    "00111111", --  405 - 0x195  :   63 - 0x3f
    "00111111", --  406 - 0x196  :   63 - 0x3f
    "00111111", --  407 - 0x197  :   63 - 0x3f
    "00111111", --  408 - 0x198  :   63 - 0x3f
    "00111111", --  409 - 0x199  :   63 - 0x3f
    "00111111", --  410 - 0x19a  :   63 - 0x3f
    "00111111", --  411 - 0x19b  :   63 - 0x3f
    "00111111", --  412 - 0x19c  :   63 - 0x3f
    "00111111", --  413 - 0x19d  :   63 - 0x3f
    "00111111", --  414 - 0x19e  :   63 - 0x3f
    "00111111", --  415 - 0x19f  :   63 - 0x3f
    "00111111", --  416 - 0x1a0  :   63 - 0x3f -- line 0xd
    "00111111", --  417 - 0x1a1  :   63 - 0x3f
    "00111111", --  418 - 0x1a2  :   63 - 0x3f
    "00111111", --  419 - 0x1a3  :   63 - 0x3f
    "00111111", --  420 - 0x1a4  :   63 - 0x3f
    "00111111", --  421 - 0x1a5  :   63 - 0x3f
    "00111111", --  422 - 0x1a6  :   63 - 0x3f
    "00111111", --  423 - 0x1a7  :   63 - 0x3f
    "00111111", --  424 - 0x1a8  :   63 - 0x3f
    "00111111", --  425 - 0x1a9  :   63 - 0x3f
    "00111111", --  426 - 0x1aa  :   63 - 0x3f
    "00111111", --  427 - 0x1ab  :   63 - 0x3f
    "00111111", --  428 - 0x1ac  :   63 - 0x3f
    "00111111", --  429 - 0x1ad  :   63 - 0x3f
    "00111111", --  430 - 0x1ae  :   63 - 0x3f
    "00111111", --  431 - 0x1af  :   63 - 0x3f
    "00111111", --  432 - 0x1b0  :   63 - 0x3f
    "00111111", --  433 - 0x1b1  :   63 - 0x3f
    "00111111", --  434 - 0x1b2  :   63 - 0x3f
    "00111111", --  435 - 0x1b3  :   63 - 0x3f
    "00111111", --  436 - 0x1b4  :   63 - 0x3f
    "00111111", --  437 - 0x1b5  :   63 - 0x3f
    "00111111", --  438 - 0x1b6  :   63 - 0x3f
    "00111111", --  439 - 0x1b7  :   63 - 0x3f
    "00111111", --  440 - 0x1b8  :   63 - 0x3f
    "00111111", --  441 - 0x1b9  :   63 - 0x3f
    "00111111", --  442 - 0x1ba  :   63 - 0x3f
    "00111111", --  443 - 0x1bb  :   63 - 0x3f
    "00111111", --  444 - 0x1bc  :   63 - 0x3f
    "00111111", --  445 - 0x1bd  :   63 - 0x3f
    "00111111", --  446 - 0x1be  :   63 - 0x3f
    "00111111", --  447 - 0x1bf  :   63 - 0x3f
    "00111111", --  448 - 0x1c0  :   63 - 0x3f -- line 0xe
    "00111111", --  449 - 0x1c1  :   63 - 0x3f
    "00111111", --  450 - 0x1c2  :   63 - 0x3f
    "00111111", --  451 - 0x1c3  :   63 - 0x3f
    "00111111", --  452 - 0x1c4  :   63 - 0x3f
    "00111111", --  453 - 0x1c5  :   63 - 0x3f
    "00111111", --  454 - 0x1c6  :   63 - 0x3f
    "00111111", --  455 - 0x1c7  :   63 - 0x3f
    "00111111", --  456 - 0x1c8  :   63 - 0x3f
    "00111111", --  457 - 0x1c9  :   63 - 0x3f
    "00111111", --  458 - 0x1ca  :   63 - 0x3f
    "00111111", --  459 - 0x1cb  :   63 - 0x3f
    "00111111", --  460 - 0x1cc  :   63 - 0x3f
    "00111111", --  461 - 0x1cd  :   63 - 0x3f
    "00111111", --  462 - 0x1ce  :   63 - 0x3f
    "00111111", --  463 - 0x1cf  :   63 - 0x3f
    "00111111", --  464 - 0x1d0  :   63 - 0x3f
    "00111111", --  465 - 0x1d1  :   63 - 0x3f
    "00111111", --  466 - 0x1d2  :   63 - 0x3f
    "00111111", --  467 - 0x1d3  :   63 - 0x3f
    "00111111", --  468 - 0x1d4  :   63 - 0x3f
    "00111111", --  469 - 0x1d5  :   63 - 0x3f
    "00111111", --  470 - 0x1d6  :   63 - 0x3f
    "00111111", --  471 - 0x1d7  :   63 - 0x3f
    "00111111", --  472 - 0x1d8  :   63 - 0x3f
    "00111111", --  473 - 0x1d9  :   63 - 0x3f
    "00111111", --  474 - 0x1da  :   63 - 0x3f
    "00111111", --  475 - 0x1db  :   63 - 0x3f
    "00111111", --  476 - 0x1dc  :   63 - 0x3f
    "00111111", --  477 - 0x1dd  :   63 - 0x3f
    "00111111", --  478 - 0x1de  :   63 - 0x3f
    "00111111", --  479 - 0x1df  :   63 - 0x3f
    "00111111", --  480 - 0x1e0  :   63 - 0x3f -- line 0xf
    "00111111", --  481 - 0x1e1  :   63 - 0x3f
    "00111111", --  482 - 0x1e2  :   63 - 0x3f
    "00111111", --  483 - 0x1e3  :   63 - 0x3f
    "00111111", --  484 - 0x1e4  :   63 - 0x3f
    "00111111", --  485 - 0x1e5  :   63 - 0x3f
    "00111111", --  486 - 0x1e6  :   63 - 0x3f
    "00111111", --  487 - 0x1e7  :   63 - 0x3f
    "00111111", --  488 - 0x1e8  :   63 - 0x3f
    "00111111", --  489 - 0x1e9  :   63 - 0x3f
    "00111111", --  490 - 0x1ea  :   63 - 0x3f
    "00111111", --  491 - 0x1eb  :   63 - 0x3f
    "00111111", --  492 - 0x1ec  :   63 - 0x3f
    "00111111", --  493 - 0x1ed  :   63 - 0x3f
    "00111111", --  494 - 0x1ee  :   63 - 0x3f
    "00111111", --  495 - 0x1ef  :   63 - 0x3f
    "00111111", --  496 - 0x1f0  :   63 - 0x3f
    "00111111", --  497 - 0x1f1  :   63 - 0x3f
    "00111111", --  498 - 0x1f2  :   63 - 0x3f
    "00111111", --  499 - 0x1f3  :   63 - 0x3f
    "00111111", --  500 - 0x1f4  :   63 - 0x3f
    "00111111", --  501 - 0x1f5  :   63 - 0x3f
    "00111111", --  502 - 0x1f6  :   63 - 0x3f
    "00111111", --  503 - 0x1f7  :   63 - 0x3f
    "00111111", --  504 - 0x1f8  :   63 - 0x3f
    "00111111", --  505 - 0x1f9  :   63 - 0x3f
    "00111111", --  506 - 0x1fa  :   63 - 0x3f
    "00111111", --  507 - 0x1fb  :   63 - 0x3f
    "00111111", --  508 - 0x1fc  :   63 - 0x3f
    "00111111", --  509 - 0x1fd  :   63 - 0x3f
    "00111111", --  510 - 0x1fe  :   63 - 0x3f
    "00111111", --  511 - 0x1ff  :   63 - 0x3f
    "00111111", --  512 - 0x200  :   63 - 0x3f -- line 0x10
    "00111111", --  513 - 0x201  :   63 - 0x3f
    "00111111", --  514 - 0x202  :   63 - 0x3f
    "00111111", --  515 - 0x203  :   63 - 0x3f
    "00111111", --  516 - 0x204  :   63 - 0x3f
    "00111111", --  517 - 0x205  :   63 - 0x3f
    "00111111", --  518 - 0x206  :   63 - 0x3f
    "00111111", --  519 - 0x207  :   63 - 0x3f
    "00111111", --  520 - 0x208  :   63 - 0x3f
    "00111111", --  521 - 0x209  :   63 - 0x3f
    "00111111", --  522 - 0x20a  :   63 - 0x3f
    "00111111", --  523 - 0x20b  :   63 - 0x3f
    "00111111", --  524 - 0x20c  :   63 - 0x3f
    "00111111", --  525 - 0x20d  :   63 - 0x3f
    "00111111", --  526 - 0x20e  :   63 - 0x3f
    "00111111", --  527 - 0x20f  :   63 - 0x3f
    "00111111", --  528 - 0x210  :   63 - 0x3f
    "00111111", --  529 - 0x211  :   63 - 0x3f
    "00111111", --  530 - 0x212  :   63 - 0x3f
    "00111111", --  531 - 0x213  :   63 - 0x3f
    "00111111", --  532 - 0x214  :   63 - 0x3f
    "00111111", --  533 - 0x215  :   63 - 0x3f
    "00111111", --  534 - 0x216  :   63 - 0x3f
    "00111111", --  535 - 0x217  :   63 - 0x3f
    "00111111", --  536 - 0x218  :   63 - 0x3f
    "00111111", --  537 - 0x219  :   63 - 0x3f
    "00111111", --  538 - 0x21a  :   63 - 0x3f
    "00111111", --  539 - 0x21b  :   63 - 0x3f
    "00111111", --  540 - 0x21c  :   63 - 0x3f
    "00111111", --  541 - 0x21d  :   63 - 0x3f
    "00111111", --  542 - 0x21e  :   63 - 0x3f
    "00111111", --  543 - 0x21f  :   63 - 0x3f
    "00111111", --  544 - 0x220  :   63 - 0x3f -- line 0x11
    "00111111", --  545 - 0x221  :   63 - 0x3f
    "00111111", --  546 - 0x222  :   63 - 0x3f
    "00111111", --  547 - 0x223  :   63 - 0x3f
    "00111111", --  548 - 0x224  :   63 - 0x3f
    "00111111", --  549 - 0x225  :   63 - 0x3f
    "00111111", --  550 - 0x226  :   63 - 0x3f
    "00111111", --  551 - 0x227  :   63 - 0x3f
    "00111111", --  552 - 0x228  :   63 - 0x3f
    "00111111", --  553 - 0x229  :   63 - 0x3f
    "00111111", --  554 - 0x22a  :   63 - 0x3f
    "00111111", --  555 - 0x22b  :   63 - 0x3f
    "00111111", --  556 - 0x22c  :   63 - 0x3f
    "00111111", --  557 - 0x22d  :   63 - 0x3f
    "00111111", --  558 - 0x22e  :   63 - 0x3f
    "00111111", --  559 - 0x22f  :   63 - 0x3f
    "00111111", --  560 - 0x230  :   63 - 0x3f
    "00111111", --  561 - 0x231  :   63 - 0x3f
    "00111111", --  562 - 0x232  :   63 - 0x3f
    "00111111", --  563 - 0x233  :   63 - 0x3f
    "00111111", --  564 - 0x234  :   63 - 0x3f
    "00111111", --  565 - 0x235  :   63 - 0x3f
    "00111111", --  566 - 0x236  :   63 - 0x3f
    "00111111", --  567 - 0x237  :   63 - 0x3f
    "00111111", --  568 - 0x238  :   63 - 0x3f
    "00111111", --  569 - 0x239  :   63 - 0x3f
    "00111111", --  570 - 0x23a  :   63 - 0x3f
    "00111111", --  571 - 0x23b  :   63 - 0x3f
    "00111111", --  572 - 0x23c  :   63 - 0x3f
    "00111111", --  573 - 0x23d  :   63 - 0x3f
    "00111111", --  574 - 0x23e  :   63 - 0x3f
    "00111111", --  575 - 0x23f  :   63 - 0x3f
    "00111111", --  576 - 0x240  :   63 - 0x3f -- line 0x12
    "00111111", --  577 - 0x241  :   63 - 0x3f
    "00111111", --  578 - 0x242  :   63 - 0x3f
    "00111111", --  579 - 0x243  :   63 - 0x3f
    "00111111", --  580 - 0x244  :   63 - 0x3f
    "00111111", --  581 - 0x245  :   63 - 0x3f
    "00111111", --  582 - 0x246  :   63 - 0x3f
    "00111111", --  583 - 0x247  :   63 - 0x3f
    "00111111", --  584 - 0x248  :   63 - 0x3f
    "00111111", --  585 - 0x249  :   63 - 0x3f
    "00111111", --  586 - 0x24a  :   63 - 0x3f
    "00111111", --  587 - 0x24b  :   63 - 0x3f
    "00111111", --  588 - 0x24c  :   63 - 0x3f
    "00111111", --  589 - 0x24d  :   63 - 0x3f
    "00111111", --  590 - 0x24e  :   63 - 0x3f
    "00111111", --  591 - 0x24f  :   63 - 0x3f
    "00000000", --  592 - 0x250  :    0 - 0x0
    "00000010", --  593 - 0x251  :    2 - 0x2
    "00000000", --  594 - 0x252  :    0 - 0x0
    "00000010", --  595 - 0x253  :    2 - 0x2
    "00000000", --  596 - 0x254  :    0 - 0x0
    "00000010", --  597 - 0x255  :    2 - 0x2
    "00000100", --  598 - 0x256  :    4 - 0x4
    "00000110", --  599 - 0x257  :    6 - 0x6
    "00000000", --  600 - 0x258  :    0 - 0x0
    "00000010", --  601 - 0x259  :    2 - 0x2
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000010", --  603 - 0x25b  :    2 - 0x2
    "00000100", --  604 - 0x25c  :    4 - 0x4
    "00000110", --  605 - 0x25d  :    6 - 0x6
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000010", --  607 - 0x25f  :    2 - 0x2
    "00111111", --  608 - 0x260  :   63 - 0x3f -- line 0x13
    "00111111", --  609 - 0x261  :   63 - 0x3f
    "00111111", --  610 - 0x262  :   63 - 0x3f
    "00111111", --  611 - 0x263  :   63 - 0x3f
    "00111111", --  612 - 0x264  :   63 - 0x3f
    "00111111", --  613 - 0x265  :   63 - 0x3f
    "00111111", --  614 - 0x266  :   63 - 0x3f
    "00111111", --  615 - 0x267  :   63 - 0x3f
    "00111111", --  616 - 0x268  :   63 - 0x3f
    "00111111", --  617 - 0x269  :   63 - 0x3f
    "00111111", --  618 - 0x26a  :   63 - 0x3f
    "00111111", --  619 - 0x26b  :   63 - 0x3f
    "00111111", --  620 - 0x26c  :   63 - 0x3f
    "00111111", --  621 - 0x26d  :   63 - 0x3f
    "00111111", --  622 - 0x26e  :   63 - 0x3f
    "00111111", --  623 - 0x26f  :   63 - 0x3f
    "00000001", --  624 - 0x270  :    1 - 0x1
    "00000011", --  625 - 0x271  :    3 - 0x3
    "00000001", --  626 - 0x272  :    1 - 0x1
    "00000011", --  627 - 0x273  :    3 - 0x3
    "00000001", --  628 - 0x274  :    1 - 0x1
    "00000011", --  629 - 0x275  :    3 - 0x3
    "00000101", --  630 - 0x276  :    5 - 0x5
    "00000111", --  631 - 0x277  :    7 - 0x7
    "00000001", --  632 - 0x278  :    1 - 0x1
    "00000011", --  633 - 0x279  :    3 - 0x3
    "00000001", --  634 - 0x27a  :    1 - 0x1
    "00000011", --  635 - 0x27b  :    3 - 0x3
    "00000101", --  636 - 0x27c  :    5 - 0x5
    "00000111", --  637 - 0x27d  :    7 - 0x7
    "00000001", --  638 - 0x27e  :    1 - 0x1
    "00000011", --  639 - 0x27f  :    3 - 0x3
    "00111111", --  640 - 0x280  :   63 - 0x3f -- line 0x14
    "00111111", --  641 - 0x281  :   63 - 0x3f
    "00111111", --  642 - 0x282  :   63 - 0x3f
    "00111111", --  643 - 0x283  :   63 - 0x3f
    "00111111", --  644 - 0x284  :   63 - 0x3f
    "00111111", --  645 - 0x285  :   63 - 0x3f
    "00111111", --  646 - 0x286  :   63 - 0x3f
    "00111111", --  647 - 0x287  :   63 - 0x3f
    "00111111", --  648 - 0x288  :   63 - 0x3f
    "00111111", --  649 - 0x289  :   63 - 0x3f
    "00111111", --  650 - 0x28a  :   63 - 0x3f
    "00111111", --  651 - 0x28b  :   63 - 0x3f
    "00111111", --  652 - 0x28c  :   63 - 0x3f
    "00111111", --  653 - 0x28d  :   63 - 0x3f
    "00111111", --  654 - 0x28e  :   63 - 0x3f
    "00111111", --  655 - 0x28f  :   63 - 0x3f
    "00111111", --  656 - 0x290  :   63 - 0x3f
    "00111111", --  657 - 0x291  :   63 - 0x3f
    "00111111", --  658 - 0x292  :   63 - 0x3f
    "00111111", --  659 - 0x293  :   63 - 0x3f
    "00111111", --  660 - 0x294  :   63 - 0x3f
    "00111111", --  661 - 0x295  :   63 - 0x3f
    "00111111", --  662 - 0x296  :   63 - 0x3f
    "00111111", --  663 - 0x297  :   63 - 0x3f
    "00111111", --  664 - 0x298  :   63 - 0x3f
    "00111111", --  665 - 0x299  :   63 - 0x3f
    "00111111", --  666 - 0x29a  :   63 - 0x3f
    "00111111", --  667 - 0x29b  :   63 - 0x3f
    "00111111", --  668 - 0x29c  :   63 - 0x3f
    "00111111", --  669 - 0x29d  :   63 - 0x3f
    "00111111", --  670 - 0x29e  :   63 - 0x3f
    "00111111", --  671 - 0x29f  :   63 - 0x3f
    "00111111", --  672 - 0x2a0  :   63 - 0x3f -- line 0x15
    "00111111", --  673 - 0x2a1  :   63 - 0x3f
    "00111111", --  674 - 0x2a2  :   63 - 0x3f
    "00111111", --  675 - 0x2a3  :   63 - 0x3f
    "00111111", --  676 - 0x2a4  :   63 - 0x3f
    "00111111", --  677 - 0x2a5  :   63 - 0x3f
    "00111111", --  678 - 0x2a6  :   63 - 0x3f
    "00111111", --  679 - 0x2a7  :   63 - 0x3f
    "00111111", --  680 - 0x2a8  :   63 - 0x3f
    "00111111", --  681 - 0x2a9  :   63 - 0x3f
    "00111111", --  682 - 0x2aa  :   63 - 0x3f
    "00111111", --  683 - 0x2ab  :   63 - 0x3f
    "00111111", --  684 - 0x2ac  :   63 - 0x3f
    "00111111", --  685 - 0x2ad  :   63 - 0x3f
    "00111111", --  686 - 0x2ae  :   63 - 0x3f
    "00111111", --  687 - 0x2af  :   63 - 0x3f
    "00111111", --  688 - 0x2b0  :   63 - 0x3f
    "00111111", --  689 - 0x2b1  :   63 - 0x3f
    "00111111", --  690 - 0x2b2  :   63 - 0x3f
    "00111111", --  691 - 0x2b3  :   63 - 0x3f
    "00111111", --  692 - 0x2b4  :   63 - 0x3f
    "00111111", --  693 - 0x2b5  :   63 - 0x3f
    "00111111", --  694 - 0x2b6  :   63 - 0x3f
    "00111111", --  695 - 0x2b7  :   63 - 0x3f
    "00111111", --  696 - 0x2b8  :   63 - 0x3f
    "00111111", --  697 - 0x2b9  :   63 - 0x3f
    "00111111", --  698 - 0x2ba  :   63 - 0x3f
    "00111111", --  699 - 0x2bb  :   63 - 0x3f
    "00111111", --  700 - 0x2bc  :   63 - 0x3f
    "00111111", --  701 - 0x2bd  :   63 - 0x3f
    "00111111", --  702 - 0x2be  :   63 - 0x3f
    "00111111", --  703 - 0x2bf  :   63 - 0x3f
    "00111111", --  704 - 0x2c0  :   63 - 0x3f -- line 0x16
    "00111111", --  705 - 0x2c1  :   63 - 0x3f
    "00111111", --  706 - 0x2c2  :   63 - 0x3f
    "00111111", --  707 - 0x2c3  :   63 - 0x3f
    "00111111", --  708 - 0x2c4  :   63 - 0x3f
    "00111111", --  709 - 0x2c5  :   63 - 0x3f
    "00111111", --  710 - 0x2c6  :   63 - 0x3f
    "00111111", --  711 - 0x2c7  :   63 - 0x3f
    "00111111", --  712 - 0x2c8  :   63 - 0x3f
    "00111111", --  713 - 0x2c9  :   63 - 0x3f
    "00111111", --  714 - 0x2ca  :   63 - 0x3f
    "00111111", --  715 - 0x2cb  :   63 - 0x3f
    "00111111", --  716 - 0x2cc  :   63 - 0x3f
    "00111111", --  717 - 0x2cd  :   63 - 0x3f
    "00111111", --  718 - 0x2ce  :   63 - 0x3f
    "00111111", --  719 - 0x2cf  :   63 - 0x3f
    "00111111", --  720 - 0x2d0  :   63 - 0x3f
    "00111111", --  721 - 0x2d1  :   63 - 0x3f
    "00111111", --  722 - 0x2d2  :   63 - 0x3f
    "00111111", --  723 - 0x2d3  :   63 - 0x3f
    "00111111", --  724 - 0x2d4  :   63 - 0x3f
    "00111111", --  725 - 0x2d5  :   63 - 0x3f
    "00111111", --  726 - 0x2d6  :   63 - 0x3f
    "00111111", --  727 - 0x2d7  :   63 - 0x3f
    "00111111", --  728 - 0x2d8  :   63 - 0x3f
    "00111111", --  729 - 0x2d9  :   63 - 0x3f
    "00111111", --  730 - 0x2da  :   63 - 0x3f
    "00111111", --  731 - 0x2db  :   63 - 0x3f
    "00111111", --  732 - 0x2dc  :   63 - 0x3f
    "00111111", --  733 - 0x2dd  :   63 - 0x3f
    "00111111", --  734 - 0x2de  :   63 - 0x3f
    "00111111", --  735 - 0x2df  :   63 - 0x3f
    "00111111", --  736 - 0x2e0  :   63 - 0x3f -- line 0x17
    "00111111", --  737 - 0x2e1  :   63 - 0x3f
    "00111111", --  738 - 0x2e2  :   63 - 0x3f
    "00111111", --  739 - 0x2e3  :   63 - 0x3f
    "00111111", --  740 - 0x2e4  :   63 - 0x3f
    "00111111", --  741 - 0x2e5  :   63 - 0x3f
    "00111111", --  742 - 0x2e6  :   63 - 0x3f
    "00111111", --  743 - 0x2e7  :   63 - 0x3f
    "00111111", --  744 - 0x2e8  :   63 - 0x3f
    "00111111", --  745 - 0x2e9  :   63 - 0x3f
    "00111111", --  746 - 0x2ea  :   63 - 0x3f
    "00111111", --  747 - 0x2eb  :   63 - 0x3f
    "00111111", --  748 - 0x2ec  :   63 - 0x3f
    "00111111", --  749 - 0x2ed  :   63 - 0x3f
    "00111111", --  750 - 0x2ee  :   63 - 0x3f
    "00111111", --  751 - 0x2ef  :   63 - 0x3f
    "11000101", --  752 - 0x2f0  :  197 - 0xc5
    "11010110", --  753 - 0x2f1  :  214 - 0xd6
    "11000101", --  754 - 0x2f2  :  197 - 0xc5
    "11010110", --  755 - 0x2f3  :  214 - 0xd6
    "11000101", --  756 - 0x2f4  :  197 - 0xc5
    "11010110", --  757 - 0x2f5  :  214 - 0xd6
    "11000101", --  758 - 0x2f6  :  197 - 0xc5
    "11010110", --  759 - 0x2f7  :  214 - 0xd6
    "11000101", --  760 - 0x2f8  :  197 - 0xc5
    "11010110", --  761 - 0x2f9  :  214 - 0xd6
    "11000101", --  762 - 0x2fa  :  197 - 0xc5
    "11010110", --  763 - 0x2fb  :  214 - 0xd6
    "11000101", --  764 - 0x2fc  :  197 - 0xc5
    "11010110", --  765 - 0x2fd  :  214 - 0xd6
    "11000101", --  766 - 0x2fe  :  197 - 0xc5
    "11010110", --  767 - 0x2ff  :  214 - 0xd6
    "00111111", --  768 - 0x300  :   63 - 0x3f -- line 0x18
    "00111111", --  769 - 0x301  :   63 - 0x3f
    "00111111", --  770 - 0x302  :   63 - 0x3f
    "00111111", --  771 - 0x303  :   63 - 0x3f
    "00011100", --  772 - 0x304  :   28 - 0x1c
    "00011110", --  773 - 0x305  :   30 - 0x1e
    "00111111", --  774 - 0x306  :   63 - 0x3f
    "00111111", --  775 - 0x307  :   63 - 0x3f
    "00111111", --  776 - 0x308  :   63 - 0x3f
    "00111111", --  777 - 0x309  :   63 - 0x3f
    "00111111", --  778 - 0x30a  :   63 - 0x3f
    "00111111", --  779 - 0x30b  :   63 - 0x3f
    "00111111", --  780 - 0x30c  :   63 - 0x3f
    "00111111", --  781 - 0x30d  :   63 - 0x3f
    "00111111", --  782 - 0x30e  :   63 - 0x3f
    "00111111", --  783 - 0x30f  :   63 - 0x3f
    "11000111", --  784 - 0x310  :  199 - 0xc7
    "11001001", --  785 - 0x311  :  201 - 0xc9
    "11000111", --  786 - 0x312  :  199 - 0xc7
    "11001001", --  787 - 0x313  :  201 - 0xc9
    "11000111", --  788 - 0x314  :  199 - 0xc7
    "11001001", --  789 - 0x315  :  201 - 0xc9
    "11000111", --  790 - 0x316  :  199 - 0xc7
    "11001001", --  791 - 0x317  :  201 - 0xc9
    "11000111", --  792 - 0x318  :  199 - 0xc7
    "11001001", --  793 - 0x319  :  201 - 0xc9
    "11000111", --  794 - 0x31a  :  199 - 0xc7
    "11001001", --  795 - 0x31b  :  201 - 0xc9
    "11000111", --  796 - 0x31c  :  199 - 0xc7
    "11001001", --  797 - 0x31d  :  201 - 0xc9
    "11000111", --  798 - 0x31e  :  199 - 0xc7
    "11001001", --  799 - 0x31f  :  201 - 0xc9
    "00111111", --  800 - 0x320  :   63 - 0x3f -- line 0x19
    "00111111", --  801 - 0x321  :   63 - 0x3f
    "00111111", --  802 - 0x322  :   63 - 0x3f
    "00111111", --  803 - 0x323  :   63 - 0x3f
    "00011101", --  804 - 0x324  :   29 - 0x1d
    "00011111", --  805 - 0x325  :   31 - 0x1f
    "00111111", --  806 - 0x326  :   63 - 0x3f
    "00111111", --  807 - 0x327  :   63 - 0x3f
    "00111111", --  808 - 0x328  :   63 - 0x3f
    "00111111", --  809 - 0x329  :   63 - 0x3f
    "00111111", --  810 - 0x32a  :   63 - 0x3f
    "00111111", --  811 - 0x32b  :   63 - 0x3f
    "00111111", --  812 - 0x32c  :   63 - 0x3f
    "00111111", --  813 - 0x32d  :   63 - 0x3f
    "00111111", --  814 - 0x32e  :   63 - 0x3f
    "00111111", --  815 - 0x32f  :   63 - 0x3f
    "11010111", --  816 - 0x330  :  215 - 0xd7
    "11011001", --  817 - 0x331  :  217 - 0xd9
    "11010111", --  818 - 0x332  :  215 - 0xd7
    "11011001", --  819 - 0x333  :  217 - 0xd9
    "11010111", --  820 - 0x334  :  215 - 0xd7
    "11011001", --  821 - 0x335  :  217 - 0xd9
    "11010111", --  822 - 0x336  :  215 - 0xd7
    "11011001", --  823 - 0x337  :  217 - 0xd9
    "11010111", --  824 - 0x338  :  215 - 0xd7
    "11011001", --  825 - 0x339  :  217 - 0xd9
    "11010111", --  826 - 0x33a  :  215 - 0xd7
    "11011001", --  827 - 0x33b  :  217 - 0xd9
    "11010111", --  828 - 0x33c  :  215 - 0xd7
    "11011001", --  829 - 0x33d  :  217 - 0xd9
    "11010111", --  830 - 0x33e  :  215 - 0xd7
    "11011001", --  831 - 0x33f  :  217 - 0xd9
    "01110000", --  832 - 0x340  :  112 - 0x70 -- line 0x1a
    "01110001", --  833 - 0x341  :  113 - 0x71
    "01110001", --  834 - 0x342  :  113 - 0x71
    "01110001", --  835 - 0x343  :  113 - 0x71
    "01110001", --  836 - 0x344  :  113 - 0x71
    "01110001", --  837 - 0x345  :  113 - 0x71
    "01110001", --  838 - 0x346  :  113 - 0x71
    "01110001", --  839 - 0x347  :  113 - 0x71
    "01110001", --  840 - 0x348  :  113 - 0x71
    "01110001", --  841 - 0x349  :  113 - 0x71
    "01110001", --  842 - 0x34a  :  113 - 0x71
    "01110001", --  843 - 0x34b  :  113 - 0x71
    "01110001", --  844 - 0x34c  :  113 - 0x71
    "01110001", --  845 - 0x34d  :  113 - 0x71
    "01110001", --  846 - 0x34e  :  113 - 0x71
    "01110001", --  847 - 0x34f  :  113 - 0x71
    "01110001", --  848 - 0x350  :  113 - 0x71
    "01110001", --  849 - 0x351  :  113 - 0x71
    "01110001", --  850 - 0x352  :  113 - 0x71
    "01110001", --  851 - 0x353  :  113 - 0x71
    "01110001", --  852 - 0x354  :  113 - 0x71
    "01110001", --  853 - 0x355  :  113 - 0x71
    "01110001", --  854 - 0x356  :  113 - 0x71
    "01110001", --  855 - 0x357  :  113 - 0x71
    "01110001", --  856 - 0x358  :  113 - 0x71
    "01110001", --  857 - 0x359  :  113 - 0x71
    "01110001", --  858 - 0x35a  :  113 - 0x71
    "01110001", --  859 - 0x35b  :  113 - 0x71
    "01110001", --  860 - 0x35c  :  113 - 0x71
    "01110001", --  861 - 0x35d  :  113 - 0x71
    "01110001", --  862 - 0x35e  :  113 - 0x71
    "01110001", --  863 - 0x35f  :  113 - 0x71
    "01100000", --  864 - 0x360  :   96 - 0x60 -- line 0x1b
    "01110111", --  865 - 0x361  :  119 - 0x77
    "01110111", --  866 - 0x362  :  119 - 0x77
    "01110111", --  867 - 0x363  :  119 - 0x77
    "01110111", --  868 - 0x364  :  119 - 0x77
    "01110111", --  869 - 0x365  :  119 - 0x77
    "01110111", --  870 - 0x366  :  119 - 0x77
    "01110111", --  871 - 0x367  :  119 - 0x77
    "01110111", --  872 - 0x368  :  119 - 0x77
    "01110111", --  873 - 0x369  :  119 - 0x77
    "01110111", --  874 - 0x36a  :  119 - 0x77
    "01110111", --  875 - 0x36b  :  119 - 0x77
    "01110111", --  876 - 0x36c  :  119 - 0x77
    "01110111", --  877 - 0x36d  :  119 - 0x77
    "01110111", --  878 - 0x36e  :  119 - 0x77
    "01110111", --  879 - 0x36f  :  119 - 0x77
    "01110111", --  880 - 0x370  :  119 - 0x77
    "01110111", --  881 - 0x371  :  119 - 0x77
    "01110111", --  882 - 0x372  :  119 - 0x77
    "01110111", --  883 - 0x373  :  119 - 0x77
    "01110111", --  884 - 0x374  :  119 - 0x77
    "01110111", --  885 - 0x375  :  119 - 0x77
    "01110111", --  886 - 0x376  :  119 - 0x77
    "01110111", --  887 - 0x377  :  119 - 0x77
    "01110111", --  888 - 0x378  :  119 - 0x77
    "01110111", --  889 - 0x379  :  119 - 0x77
    "01110111", --  890 - 0x37a  :  119 - 0x77
    "01110111", --  891 - 0x37b  :  119 - 0x77
    "01110111", --  892 - 0x37c  :  119 - 0x77
    "01110111", --  893 - 0x37d  :  119 - 0x77
    "01110111", --  894 - 0x37e  :  119 - 0x77
    "01110111", --  895 - 0x37f  :  119 - 0x77
    "01100000", --  896 - 0x380  :   96 - 0x60 -- line 0x1c
    "01110011", --  897 - 0x381  :  115 - 0x73
    "01110011", --  898 - 0x382  :  115 - 0x73
    "01110011", --  899 - 0x383  :  115 - 0x73
    "01110011", --  900 - 0x384  :  115 - 0x73
    "01110011", --  901 - 0x385  :  115 - 0x73
    "01110011", --  902 - 0x386  :  115 - 0x73
    "01110011", --  903 - 0x387  :  115 - 0x73
    "01110011", --  904 - 0x388  :  115 - 0x73
    "01110011", --  905 - 0x389  :  115 - 0x73
    "01110011", --  906 - 0x38a  :  115 - 0x73
    "01110011", --  907 - 0x38b  :  115 - 0x73
    "01110011", --  908 - 0x38c  :  115 - 0x73
    "01110011", --  909 - 0x38d  :  115 - 0x73
    "01110011", --  910 - 0x38e  :  115 - 0x73
    "01110011", --  911 - 0x38f  :  115 - 0x73
    "01110011", --  912 - 0x390  :  115 - 0x73
    "01110011", --  913 - 0x391  :  115 - 0x73
    "01110011", --  914 - 0x392  :  115 - 0x73
    "01110011", --  915 - 0x393  :  115 - 0x73
    "01110011", --  916 - 0x394  :  115 - 0x73
    "01110011", --  917 - 0x395  :  115 - 0x73
    "01110011", --  918 - 0x396  :  115 - 0x73
    "01110011", --  919 - 0x397  :  115 - 0x73
    "01110011", --  920 - 0x398  :  115 - 0x73
    "01110011", --  921 - 0x399  :  115 - 0x73
    "01110011", --  922 - 0x39a  :  115 - 0x73
    "01110011", --  923 - 0x39b  :  115 - 0x73
    "01110011", --  924 - 0x39c  :  115 - 0x73
    "01110011", --  925 - 0x39d  :  115 - 0x73
    "01110011", --  926 - 0x39e  :  115 - 0x73
    "01110011", --  927 - 0x39f  :  115 - 0x73
    "01100000", --  928 - 0x3a0  :   96 - 0x60 -- line 0x1d
    "01110011", --  929 - 0x3a1  :  115 - 0x73
    "01110011", --  930 - 0x3a2  :  115 - 0x73
    "01110011", --  931 - 0x3a3  :  115 - 0x73
    "01110011", --  932 - 0x3a4  :  115 - 0x73
    "01110011", --  933 - 0x3a5  :  115 - 0x73
    "01110011", --  934 - 0x3a6  :  115 - 0x73
    "01110011", --  935 - 0x3a7  :  115 - 0x73
    "01110011", --  936 - 0x3a8  :  115 - 0x73
    "01110011", --  937 - 0x3a9  :  115 - 0x73
    "01110011", --  938 - 0x3aa  :  115 - 0x73
    "01110011", --  939 - 0x3ab  :  115 - 0x73
    "01110011", --  940 - 0x3ac  :  115 - 0x73
    "01110011", --  941 - 0x3ad  :  115 - 0x73
    "01110011", --  942 - 0x3ae  :  115 - 0x73
    "01110011", --  943 - 0x3af  :  115 - 0x73
    "01110011", --  944 - 0x3b0  :  115 - 0x73
    "01110011", --  945 - 0x3b1  :  115 - 0x73
    "01110011", --  946 - 0x3b2  :  115 - 0x73
    "01110011", --  947 - 0x3b3  :  115 - 0x73
    "01110011", --  948 - 0x3b4  :  115 - 0x73
    "01110011", --  949 - 0x3b5  :  115 - 0x73
    "01110011", --  950 - 0x3b6  :  115 - 0x73
    "01110011", --  951 - 0x3b7  :  115 - 0x73
    "01110011", --  952 - 0x3b8  :  115 - 0x73
    "01110011", --  953 - 0x3b9  :  115 - 0x73
    "01110011", --  954 - 0x3ba  :  115 - 0x73
    "01110011", --  955 - 0x3bb  :  115 - 0x73
    "01110011", --  956 - 0x3bc  :  115 - 0x73
    "01110011", --  957 - 0x3bd  :  115 - 0x73
    "01110011", --  958 - 0x3be  :  115 - 0x73
    "01110011", --  959 - 0x3bf  :  115 - 0x73
        ---- Attribute Table 0----
    "00000000", --  960 - 0x3c0  :    0 - 0x0
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00001000", --  974 - 0x3ce  :    8 - 0x8
    "00001000", --  975 - 0x3cf  :    8 - 0x8
    "00000000", --  976 - 0x3d0  :    0 - 0x0
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "01010001", --  981 - 0x3d5  :   81 - 0x51
    "01010000", --  982 - 0x3d6  :   80 - 0x50
    "01010000", --  983 - 0x3d7  :   80 - 0x50
    "00000000", --  984 - 0x3d8  :    0 - 0x0
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "10100000", --  996 - 0x3e4  :  160 - 0xa0
    "10100000", --  997 - 0x3e5  :  160 - 0xa0
    "10100000", --  998 - 0x3e6  :  160 - 0xa0
    "10100000", --  999 - 0x3e7  :  160 - 0xa0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0
    "00000010", -- 1009 - 0x3f1  :    2 - 0x2
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
     ------- Name Table 1---------
    "01110001", -- 1024 - 0x400  :  113 - 0x71 -- line 0x0
    "01110001", -- 1025 - 0x401  :  113 - 0x71
    "01110001", -- 1026 - 0x402  :  113 - 0x71
    "01110001", -- 1027 - 0x403  :  113 - 0x71
    "01110001", -- 1028 - 0x404  :  113 - 0x71
    "01110001", -- 1029 - 0x405  :  113 - 0x71
    "01110001", -- 1030 - 0x406  :  113 - 0x71
    "01110001", -- 1031 - 0x407  :  113 - 0x71
    "01110001", -- 1032 - 0x408  :  113 - 0x71
    "01110010", -- 1033 - 0x409  :  114 - 0x72
    "00010000", -- 1034 - 0x40a  :   16 - 0x10
    "00010001", -- 1035 - 0x40b  :   17 - 0x11
    "00001100", -- 1036 - 0x40c  :   12 - 0xc
    "00001110", -- 1037 - 0x40d  :   14 - 0xe
    "00110000", -- 1038 - 0x40e  :   48 - 0x30
    "00111111", -- 1039 - 0x40f  :   63 - 0x3f
    "00110000", -- 1040 - 0x410  :   48 - 0x30
    "00111111", -- 1041 - 0x411  :   63 - 0x3f
    "00110000", -- 1042 - 0x412  :   48 - 0x30
    "00111111", -- 1043 - 0x413  :   63 - 0x3f
    "00110000", -- 1044 - 0x414  :   48 - 0x30
    "00111111", -- 1045 - 0x415  :   63 - 0x3f
    "00110000", -- 1046 - 0x416  :   48 - 0x30
    "00111111", -- 1047 - 0x417  :   63 - 0x3f
    "00110000", -- 1048 - 0x418  :   48 - 0x30
    "00111111", -- 1049 - 0x419  :   63 - 0x3f
    "00110000", -- 1050 - 0x41a  :   48 - 0x30
    "00111111", -- 1051 - 0x41b  :   63 - 0x3f
    "00110000", -- 1052 - 0x41c  :   48 - 0x30
    "00111111", -- 1053 - 0x41d  :   63 - 0x3f
    "00110000", -- 1054 - 0x41e  :   48 - 0x30
    "00111111", -- 1055 - 0x41f  :   63 - 0x3f
    "01110111", -- 1056 - 0x420  :  119 - 0x77 -- line 0x1
    "01110111", -- 1057 - 0x421  :  119 - 0x77
    "01110111", -- 1058 - 0x422  :  119 - 0x77
    "01110111", -- 1059 - 0x423  :  119 - 0x77
    "01110111", -- 1060 - 0x424  :  119 - 0x77
    "01110111", -- 1061 - 0x425  :  119 - 0x77
    "01110111", -- 1062 - 0x426  :  119 - 0x77
    "01110111", -- 1063 - 0x427  :  119 - 0x77
    "01110111", -- 1064 - 0x428  :  119 - 0x77
    "01100001", -- 1065 - 0x429  :   97 - 0x61
    "00010000", -- 1066 - 0x42a  :   16 - 0x10
    "00010001", -- 1067 - 0x42b  :   17 - 0x11
    "00001101", -- 1068 - 0x42c  :   13 - 0xd
    "00001111", -- 1069 - 0x42d  :   15 - 0xf
    "00111111", -- 1070 - 0x42e  :   63 - 0x3f
    "00110000", -- 1071 - 0x42f  :   48 - 0x30
    "00111111", -- 1072 - 0x430  :   63 - 0x3f
    "00110000", -- 1073 - 0x431  :   48 - 0x30
    "00111111", -- 1074 - 0x432  :   63 - 0x3f
    "00110000", -- 1075 - 0x433  :   48 - 0x30
    "00111111", -- 1076 - 0x434  :   63 - 0x3f
    "00110000", -- 1077 - 0x435  :   48 - 0x30
    "00111111", -- 1078 - 0x436  :   63 - 0x3f
    "00110000", -- 1079 - 0x437  :   48 - 0x30
    "00111111", -- 1080 - 0x438  :   63 - 0x3f
    "00110000", -- 1081 - 0x439  :   48 - 0x30
    "00111111", -- 1082 - 0x43a  :   63 - 0x3f
    "00110000", -- 1083 - 0x43b  :   48 - 0x30
    "00111111", -- 1084 - 0x43c  :   63 - 0x3f
    "00110000", -- 1085 - 0x43d  :   48 - 0x30
    "00111111", -- 1086 - 0x43e  :   63 - 0x3f
    "00110000", -- 1087 - 0x43f  :   48 - 0x30
    "00111001", -- 1088 - 0x440  :   57 - 0x39 -- line 0x2
    "00111001", -- 1089 - 0x441  :   57 - 0x39
    "00111001", -- 1090 - 0x442  :   57 - 0x39
    "00111001", -- 1091 - 0x443  :   57 - 0x39
    "00111001", -- 1092 - 0x444  :   57 - 0x39
    "00111001", -- 1093 - 0x445  :   57 - 0x39
    "00111001", -- 1094 - 0x446  :   57 - 0x39
    "00111001", -- 1095 - 0x447  :   57 - 0x39
    "00111001", -- 1096 - 0x448  :   57 - 0x39
    "00111001", -- 1097 - 0x449  :   57 - 0x39
    "00010000", -- 1098 - 0x44a  :   16 - 0x10
    "00010001", -- 1099 - 0x44b  :   17 - 0x11
    "00001100", -- 1100 - 0x44c  :   12 - 0xc
    "00001110", -- 1101 - 0x44d  :   14 - 0xe
    "00110000", -- 1102 - 0x44e  :   48 - 0x30
    "00111111", -- 1103 - 0x44f  :   63 - 0x3f
    "00110000", -- 1104 - 0x450  :   48 - 0x30
    "00111111", -- 1105 - 0x451  :   63 - 0x3f
    "00110000", -- 1106 - 0x452  :   48 - 0x30
    "00111111", -- 1107 - 0x453  :   63 - 0x3f
    "00110000", -- 1108 - 0x454  :   48 - 0x30
    "00111111", -- 1109 - 0x455  :   63 - 0x3f
    "00110000", -- 1110 - 0x456  :   48 - 0x30
    "00111111", -- 1111 - 0x457  :   63 - 0x3f
    "00110000", -- 1112 - 0x458  :   48 - 0x30
    "00111111", -- 1113 - 0x459  :   63 - 0x3f
    "00110000", -- 1114 - 0x45a  :   48 - 0x30
    "00111111", -- 1115 - 0x45b  :   63 - 0x3f
    "00110000", -- 1116 - 0x45c  :   48 - 0x30
    "00111111", -- 1117 - 0x45d  :   63 - 0x3f
    "00110000", -- 1118 - 0x45e  :   48 - 0x30
    "00111111", -- 1119 - 0x45f  :   63 - 0x3f
    "00111111", -- 1120 - 0x460  :   63 - 0x3f -- line 0x3
    "00111111", -- 1121 - 0x461  :   63 - 0x3f
    "00111111", -- 1122 - 0x462  :   63 - 0x3f
    "00111111", -- 1123 - 0x463  :   63 - 0x3f
    "00111111", -- 1124 - 0x464  :   63 - 0x3f
    "00111111", -- 1125 - 0x465  :   63 - 0x3f
    "00111111", -- 1126 - 0x466  :   63 - 0x3f
    "00111111", -- 1127 - 0x467  :   63 - 0x3f
    "00111111", -- 1128 - 0x468  :   63 - 0x3f
    "00111111", -- 1129 - 0x469  :   63 - 0x3f
    "00010000", -- 1130 - 0x46a  :   16 - 0x10
    "00010001", -- 1131 - 0x46b  :   17 - 0x11
    "00001101", -- 1132 - 0x46c  :   13 - 0xd
    "00001111", -- 1133 - 0x46d  :   15 - 0xf
    "00111111", -- 1134 - 0x46e  :   63 - 0x3f
    "00110000", -- 1135 - 0x46f  :   48 - 0x30
    "00111111", -- 1136 - 0x470  :   63 - 0x3f
    "00110000", -- 1137 - 0x471  :   48 - 0x30
    "00111111", -- 1138 - 0x472  :   63 - 0x3f
    "00110000", -- 1139 - 0x473  :   48 - 0x30
    "00111111", -- 1140 - 0x474  :   63 - 0x3f
    "00110000", -- 1141 - 0x475  :   48 - 0x30
    "00111111", -- 1142 - 0x476  :   63 - 0x3f
    "00110000", -- 1143 - 0x477  :   48 - 0x30
    "00111111", -- 1144 - 0x478  :   63 - 0x3f
    "00110000", -- 1145 - 0x479  :   48 - 0x30
    "00111111", -- 1146 - 0x47a  :   63 - 0x3f
    "00110000", -- 1147 - 0x47b  :   48 - 0x30
    "00111111", -- 1148 - 0x47c  :   63 - 0x3f
    "00110000", -- 1149 - 0x47d  :   48 - 0x30
    "00111111", -- 1150 - 0x47e  :   63 - 0x3f
    "00110000", -- 1151 - 0x47f  :   48 - 0x30
    "00010100", -- 1152 - 0x480  :   20 - 0x14 -- line 0x4
    "00010110", -- 1153 - 0x481  :   22 - 0x16
    "00010100", -- 1154 - 0x482  :   20 - 0x14
    "00010110", -- 1155 - 0x483  :   22 - 0x16
    "00010100", -- 1156 - 0x484  :   20 - 0x14
    "00010110", -- 1157 - 0x485  :   22 - 0x16
    "00111111", -- 1158 - 0x486  :   63 - 0x3f
    "00111111", -- 1159 - 0x487  :   63 - 0x3f
    "00111111", -- 1160 - 0x488  :   63 - 0x3f
    "00111111", -- 1161 - 0x489  :   63 - 0x3f
    "00010000", -- 1162 - 0x48a  :   16 - 0x10
    "00010001", -- 1163 - 0x48b  :   17 - 0x11
    "00001100", -- 1164 - 0x48c  :   12 - 0xc
    "00001110", -- 1165 - 0x48d  :   14 - 0xe
    "00111111", -- 1166 - 0x48e  :   63 - 0x3f
    "00111111", -- 1167 - 0x48f  :   63 - 0x3f
    "00111111", -- 1168 - 0x490  :   63 - 0x3f
    "00111111", -- 1169 - 0x491  :   63 - 0x3f
    "00111111", -- 1170 - 0x492  :   63 - 0x3f
    "00111111", -- 1171 - 0x493  :   63 - 0x3f
    "00111111", -- 1172 - 0x494  :   63 - 0x3f
    "00111111", -- 1173 - 0x495  :   63 - 0x3f
    "00111111", -- 1174 - 0x496  :   63 - 0x3f
    "00111111", -- 1175 - 0x497  :   63 - 0x3f
    "00111111", -- 1176 - 0x498  :   63 - 0x3f
    "00111111", -- 1177 - 0x499  :   63 - 0x3f
    "00111111", -- 1178 - 0x49a  :   63 - 0x3f
    "00111111", -- 1179 - 0x49b  :   63 - 0x3f
    "00111111", -- 1180 - 0x49c  :   63 - 0x3f
    "00111111", -- 1181 - 0x49d  :   63 - 0x3f
    "00111111", -- 1182 - 0x49e  :   63 - 0x3f
    "00111111", -- 1183 - 0x49f  :   63 - 0x3f
    "00010101", -- 1184 - 0x4a0  :   21 - 0x15 -- line 0x5
    "00010111", -- 1185 - 0x4a1  :   23 - 0x17
    "00010101", -- 1186 - 0x4a2  :   21 - 0x15
    "00010111", -- 1187 - 0x4a3  :   23 - 0x17
    "00010101", -- 1188 - 0x4a4  :   21 - 0x15
    "00010111", -- 1189 - 0x4a5  :   23 - 0x17
    "00111111", -- 1190 - 0x4a6  :   63 - 0x3f
    "00111111", -- 1191 - 0x4a7  :   63 - 0x3f
    "00111111", -- 1192 - 0x4a8  :   63 - 0x3f
    "00111111", -- 1193 - 0x4a9  :   63 - 0x3f
    "00010000", -- 1194 - 0x4aa  :   16 - 0x10
    "00010001", -- 1195 - 0x4ab  :   17 - 0x11
    "00001101", -- 1196 - 0x4ac  :   13 - 0xd
    "00001111", -- 1197 - 0x4ad  :   15 - 0xf
    "00111111", -- 1198 - 0x4ae  :   63 - 0x3f
    "00111111", -- 1199 - 0x4af  :   63 - 0x3f
    "00111111", -- 1200 - 0x4b0  :   63 - 0x3f
    "00111111", -- 1201 - 0x4b1  :   63 - 0x3f
    "00111111", -- 1202 - 0x4b2  :   63 - 0x3f
    "00111111", -- 1203 - 0x4b3  :   63 - 0x3f
    "00111111", -- 1204 - 0x4b4  :   63 - 0x3f
    "00111111", -- 1205 - 0x4b5  :   63 - 0x3f
    "00111111", -- 1206 - 0x4b6  :   63 - 0x3f
    "00111111", -- 1207 - 0x4b7  :   63 - 0x3f
    "00111111", -- 1208 - 0x4b8  :   63 - 0x3f
    "00111111", -- 1209 - 0x4b9  :   63 - 0x3f
    "00111111", -- 1210 - 0x4ba  :   63 - 0x3f
    "00111111", -- 1211 - 0x4bb  :   63 - 0x3f
    "00111111", -- 1212 - 0x4bc  :   63 - 0x3f
    "00111111", -- 1213 - 0x4bd  :   63 - 0x3f
    "00111111", -- 1214 - 0x4be  :   63 - 0x3f
    "00111111", -- 1215 - 0x4bf  :   63 - 0x3f
    "00111111", -- 1216 - 0x4c0  :   63 - 0x3f -- line 0x6
    "00111111", -- 1217 - 0x4c1  :   63 - 0x3f
    "00111111", -- 1218 - 0x4c2  :   63 - 0x3f
    "00111111", -- 1219 - 0x4c3  :   63 - 0x3f
    "00111111", -- 1220 - 0x4c4  :   63 - 0x3f
    "00111111", -- 1221 - 0x4c5  :   63 - 0x3f
    "00111111", -- 1222 - 0x4c6  :   63 - 0x3f
    "00111111", -- 1223 - 0x4c7  :   63 - 0x3f
    "00111111", -- 1224 - 0x4c8  :   63 - 0x3f
    "00111111", -- 1225 - 0x4c9  :   63 - 0x3f
    "00010000", -- 1226 - 0x4ca  :   16 - 0x10
    "00010001", -- 1227 - 0x4cb  :   17 - 0x11
    "00001100", -- 1228 - 0x4cc  :   12 - 0xc
    "00001110", -- 1229 - 0x4cd  :   14 - 0xe
    "00111111", -- 1230 - 0x4ce  :   63 - 0x3f
    "00111111", -- 1231 - 0x4cf  :   63 - 0x3f
    "00111111", -- 1232 - 0x4d0  :   63 - 0x3f
    "00111111", -- 1233 - 0x4d1  :   63 - 0x3f
    "00111111", -- 1234 - 0x4d2  :   63 - 0x3f
    "00111111", -- 1235 - 0x4d3  :   63 - 0x3f
    "00111111", -- 1236 - 0x4d4  :   63 - 0x3f
    "00111111", -- 1237 - 0x4d5  :   63 - 0x3f
    "00111111", -- 1238 - 0x4d6  :   63 - 0x3f
    "00111111", -- 1239 - 0x4d7  :   63 - 0x3f
    "00111111", -- 1240 - 0x4d8  :   63 - 0x3f
    "00111111", -- 1241 - 0x4d9  :   63 - 0x3f
    "00111111", -- 1242 - 0x4da  :   63 - 0x3f
    "00111111", -- 1243 - 0x4db  :   63 - 0x3f
    "00111111", -- 1244 - 0x4dc  :   63 - 0x3f
    "00111111", -- 1245 - 0x4dd  :   63 - 0x3f
    "00111111", -- 1246 - 0x4de  :   63 - 0x3f
    "00111111", -- 1247 - 0x4df  :   63 - 0x3f
    "00111111", -- 1248 - 0x4e0  :   63 - 0x3f -- line 0x7
    "00111111", -- 1249 - 0x4e1  :   63 - 0x3f
    "00111111", -- 1250 - 0x4e2  :   63 - 0x3f
    "00111111", -- 1251 - 0x4e3  :   63 - 0x3f
    "00111111", -- 1252 - 0x4e4  :   63 - 0x3f
    "00111111", -- 1253 - 0x4e5  :   63 - 0x3f
    "00111111", -- 1254 - 0x4e6  :   63 - 0x3f
    "00111111", -- 1255 - 0x4e7  :   63 - 0x3f
    "00111111", -- 1256 - 0x4e8  :   63 - 0x3f
    "00111111", -- 1257 - 0x4e9  :   63 - 0x3f
    "00010000", -- 1258 - 0x4ea  :   16 - 0x10
    "00010001", -- 1259 - 0x4eb  :   17 - 0x11
    "00001101", -- 1260 - 0x4ec  :   13 - 0xd
    "00001111", -- 1261 - 0x4ed  :   15 - 0xf
    "00111111", -- 1262 - 0x4ee  :   63 - 0x3f
    "00111111", -- 1263 - 0x4ef  :   63 - 0x3f
    "00111111", -- 1264 - 0x4f0  :   63 - 0x3f
    "00111111", -- 1265 - 0x4f1  :   63 - 0x3f
    "00111111", -- 1266 - 0x4f2  :   63 - 0x3f
    "00111111", -- 1267 - 0x4f3  :   63 - 0x3f
    "00111111", -- 1268 - 0x4f4  :   63 - 0x3f
    "00111111", -- 1269 - 0x4f5  :   63 - 0x3f
    "00111111", -- 1270 - 0x4f6  :   63 - 0x3f
    "00111111", -- 1271 - 0x4f7  :   63 - 0x3f
    "00111111", -- 1272 - 0x4f8  :   63 - 0x3f
    "00111111", -- 1273 - 0x4f9  :   63 - 0x3f
    "00111111", -- 1274 - 0x4fa  :   63 - 0x3f
    "00111111", -- 1275 - 0x4fb  :   63 - 0x3f
    "00111111", -- 1276 - 0x4fc  :   63 - 0x3f
    "00111111", -- 1277 - 0x4fd  :   63 - 0x3f
    "00111111", -- 1278 - 0x4fe  :   63 - 0x3f
    "00111111", -- 1279 - 0x4ff  :   63 - 0x3f
    "00111111", -- 1280 - 0x500  :   63 - 0x3f -- line 0x8
    "00111111", -- 1281 - 0x501  :   63 - 0x3f
    "00001100", -- 1282 - 0x502  :   12 - 0xc
    "00001110", -- 1283 - 0x503  :   14 - 0xe
    "00001100", -- 1284 - 0x504  :   12 - 0xc
    "00001110", -- 1285 - 0x505  :   14 - 0xe
    "00001100", -- 1286 - 0x506  :   12 - 0xc
    "00001110", -- 1287 - 0x507  :   14 - 0xe
    "00001100", -- 1288 - 0x508  :   12 - 0xc
    "00001110", -- 1289 - 0x509  :   14 - 0xe
    "00001100", -- 1290 - 0x50a  :   12 - 0xc
    "00001110", -- 1291 - 0x50b  :   14 - 0xe
    "00001100", -- 1292 - 0x50c  :   12 - 0xc
    "00001110", -- 1293 - 0x50d  :   14 - 0xe
    "00111111", -- 1294 - 0x50e  :   63 - 0x3f
    "00111111", -- 1295 - 0x50f  :   63 - 0x3f
    "00111111", -- 1296 - 0x510  :   63 - 0x3f
    "00111111", -- 1297 - 0x511  :   63 - 0x3f
    "00111111", -- 1298 - 0x512  :   63 - 0x3f
    "00111111", -- 1299 - 0x513  :   63 - 0x3f
    "00111111", -- 1300 - 0x514  :   63 - 0x3f
    "00111111", -- 1301 - 0x515  :   63 - 0x3f
    "00111111", -- 1302 - 0x516  :   63 - 0x3f
    "00111111", -- 1303 - 0x517  :   63 - 0x3f
    "00111111", -- 1304 - 0x518  :   63 - 0x3f
    "00111111", -- 1305 - 0x519  :   63 - 0x3f
    "00111111", -- 1306 - 0x51a  :   63 - 0x3f
    "00111111", -- 1307 - 0x51b  :   63 - 0x3f
    "00111111", -- 1308 - 0x51c  :   63 - 0x3f
    "00111111", -- 1309 - 0x51d  :   63 - 0x3f
    "00111111", -- 1310 - 0x51e  :   63 - 0x3f
    "00111111", -- 1311 - 0x51f  :   63 - 0x3f
    "00111111", -- 1312 - 0x520  :   63 - 0x3f -- line 0x9
    "00111111", -- 1313 - 0x521  :   63 - 0x3f
    "00001101", -- 1314 - 0x522  :   13 - 0xd
    "00001111", -- 1315 - 0x523  :   15 - 0xf
    "00001101", -- 1316 - 0x524  :   13 - 0xd
    "00001111", -- 1317 - 0x525  :   15 - 0xf
    "00001101", -- 1318 - 0x526  :   13 - 0xd
    "00001111", -- 1319 - 0x527  :   15 - 0xf
    "00001101", -- 1320 - 0x528  :   13 - 0xd
    "00001111", -- 1321 - 0x529  :   15 - 0xf
    "00001101", -- 1322 - 0x52a  :   13 - 0xd
    "00001111", -- 1323 - 0x52b  :   15 - 0xf
    "00001101", -- 1324 - 0x52c  :   13 - 0xd
    "00001111", -- 1325 - 0x52d  :   15 - 0xf
    "00111111", -- 1326 - 0x52e  :   63 - 0x3f
    "00111111", -- 1327 - 0x52f  :   63 - 0x3f
    "00111111", -- 1328 - 0x530  :   63 - 0x3f
    "00111111", -- 1329 - 0x531  :   63 - 0x3f
    "00111111", -- 1330 - 0x532  :   63 - 0x3f
    "00111111", -- 1331 - 0x533  :   63 - 0x3f
    "00111111", -- 1332 - 0x534  :   63 - 0x3f
    "00111111", -- 1333 - 0x535  :   63 - 0x3f
    "00111111", -- 1334 - 0x536  :   63 - 0x3f
    "00111111", -- 1335 - 0x537  :   63 - 0x3f
    "00111111", -- 1336 - 0x538  :   63 - 0x3f
    "00111111", -- 1337 - 0x539  :   63 - 0x3f
    "00111111", -- 1338 - 0x53a  :   63 - 0x3f
    "00111111", -- 1339 - 0x53b  :   63 - 0x3f
    "00111111", -- 1340 - 0x53c  :   63 - 0x3f
    "00111111", -- 1341 - 0x53d  :   63 - 0x3f
    "00111111", -- 1342 - 0x53e  :   63 - 0x3f
    "00111111", -- 1343 - 0x53f  :   63 - 0x3f
    "01011000", -- 1344 - 0x540  :   88 - 0x58 -- line 0xa
    "01011000", -- 1345 - 0x541  :   88 - 0x58
    "01011000", -- 1346 - 0x542  :   88 - 0x58
    "01011001", -- 1347 - 0x543  :   89 - 0x59
    "00111111", -- 1348 - 0x544  :   63 - 0x3f
    "00111111", -- 1349 - 0x545  :   63 - 0x3f
    "00111111", -- 1350 - 0x546  :   63 - 0x3f
    "00111111", -- 1351 - 0x547  :   63 - 0x3f
    "00111111", -- 1352 - 0x548  :   63 - 0x3f
    "00111111", -- 1353 - 0x549  :   63 - 0x3f
    "00111111", -- 1354 - 0x54a  :   63 - 0x3f
    "00111111", -- 1355 - 0x54b  :   63 - 0x3f
    "00111111", -- 1356 - 0x54c  :   63 - 0x3f
    "00111111", -- 1357 - 0x54d  :   63 - 0x3f
    "00111111", -- 1358 - 0x54e  :   63 - 0x3f
    "00111111", -- 1359 - 0x54f  :   63 - 0x3f
    "00111111", -- 1360 - 0x550  :   63 - 0x3f
    "00111111", -- 1361 - 0x551  :   63 - 0x3f
    "00111111", -- 1362 - 0x552  :   63 - 0x3f
    "00111111", -- 1363 - 0x553  :   63 - 0x3f
    "00111111", -- 1364 - 0x554  :   63 - 0x3f
    "00111111", -- 1365 - 0x555  :   63 - 0x3f
    "00111111", -- 1366 - 0x556  :   63 - 0x3f
    "00111111", -- 1367 - 0x557  :   63 - 0x3f
    "00111111", -- 1368 - 0x558  :   63 - 0x3f
    "00111111", -- 1369 - 0x559  :   63 - 0x3f
    "00010100", -- 1370 - 0x55a  :   20 - 0x14
    "00010110", -- 1371 - 0x55b  :   22 - 0x16
    "00010100", -- 1372 - 0x55c  :   20 - 0x14
    "00010110", -- 1373 - 0x55d  :   22 - 0x16
    "00010100", -- 1374 - 0x55e  :   20 - 0x14
    "00010110", -- 1375 - 0x55f  :   22 - 0x16
    "00111111", -- 1376 - 0x560  :   63 - 0x3f -- line 0xb
    "00111111", -- 1377 - 0x561  :   63 - 0x3f
    "00111111", -- 1378 - 0x562  :   63 - 0x3f
    "00111111", -- 1379 - 0x563  :   63 - 0x3f
    "00111111", -- 1380 - 0x564  :   63 - 0x3f
    "00111111", -- 1381 - 0x565  :   63 - 0x3f
    "00111111", -- 1382 - 0x566  :   63 - 0x3f
    "00111111", -- 1383 - 0x567  :   63 - 0x3f
    "00111111", -- 1384 - 0x568  :   63 - 0x3f
    "00111111", -- 1385 - 0x569  :   63 - 0x3f
    "00111111", -- 1386 - 0x56a  :   63 - 0x3f
    "00111111", -- 1387 - 0x56b  :   63 - 0x3f
    "00111111", -- 1388 - 0x56c  :   63 - 0x3f
    "00111111", -- 1389 - 0x56d  :   63 - 0x3f
    "00111111", -- 1390 - 0x56e  :   63 - 0x3f
    "00111111", -- 1391 - 0x56f  :   63 - 0x3f
    "00111111", -- 1392 - 0x570  :   63 - 0x3f
    "00111111", -- 1393 - 0x571  :   63 - 0x3f
    "00111111", -- 1394 - 0x572  :   63 - 0x3f
    "00111111", -- 1395 - 0x573  :   63 - 0x3f
    "00111111", -- 1396 - 0x574  :   63 - 0x3f
    "00111111", -- 1397 - 0x575  :   63 - 0x3f
    "00111111", -- 1398 - 0x576  :   63 - 0x3f
    "00111111", -- 1399 - 0x577  :   63 - 0x3f
    "00111111", -- 1400 - 0x578  :   63 - 0x3f
    "00111111", -- 1401 - 0x579  :   63 - 0x3f
    "00010101", -- 1402 - 0x57a  :   21 - 0x15
    "00010111", -- 1403 - 0x57b  :   23 - 0x17
    "00010101", -- 1404 - 0x57c  :   21 - 0x15
    "00010111", -- 1405 - 0x57d  :   23 - 0x17
    "00010101", -- 1406 - 0x57e  :   21 - 0x15
    "00010111", -- 1407 - 0x57f  :   23 - 0x17
    "00111111", -- 1408 - 0x580  :   63 - 0x3f -- line 0xc
    "00111111", -- 1409 - 0x581  :   63 - 0x3f
    "00111111", -- 1410 - 0x582  :   63 - 0x3f
    "00111111", -- 1411 - 0x583  :   63 - 0x3f
    "00111111", -- 1412 - 0x584  :   63 - 0x3f
    "00111111", -- 1413 - 0x585  :   63 - 0x3f
    "00111111", -- 1414 - 0x586  :   63 - 0x3f
    "00111111", -- 1415 - 0x587  :   63 - 0x3f
    "00111111", -- 1416 - 0x588  :   63 - 0x3f
    "00111111", -- 1417 - 0x589  :   63 - 0x3f
    "00111111", -- 1418 - 0x58a  :   63 - 0x3f
    "00111111", -- 1419 - 0x58b  :   63 - 0x3f
    "00111111", -- 1420 - 0x58c  :   63 - 0x3f
    "00111111", -- 1421 - 0x58d  :   63 - 0x3f
    "00111111", -- 1422 - 0x58e  :   63 - 0x3f
    "00111111", -- 1423 - 0x58f  :   63 - 0x3f
    "00111111", -- 1424 - 0x590  :   63 - 0x3f
    "00111111", -- 1425 - 0x591  :   63 - 0x3f
    "00111111", -- 1426 - 0x592  :   63 - 0x3f
    "00111111", -- 1427 - 0x593  :   63 - 0x3f
    "00111111", -- 1428 - 0x594  :   63 - 0x3f
    "00111111", -- 1429 - 0x595  :   63 - 0x3f
    "00111111", -- 1430 - 0x596  :   63 - 0x3f
    "00111111", -- 1431 - 0x597  :   63 - 0x3f
    "00111111", -- 1432 - 0x598  :   63 - 0x3f
    "00111111", -- 1433 - 0x599  :   63 - 0x3f
    "00111111", -- 1434 - 0x59a  :   63 - 0x3f
    "00111111", -- 1435 - 0x59b  :   63 - 0x3f
    "00111111", -- 1436 - 0x59c  :   63 - 0x3f
    "00111111", -- 1437 - 0x59d  :   63 - 0x3f
    "00111111", -- 1438 - 0x59e  :   63 - 0x3f
    "00111111", -- 1439 - 0x59f  :   63 - 0x3f
    "00111111", -- 1440 - 0x5a0  :   63 - 0x3f -- line 0xd
    "00111111", -- 1441 - 0x5a1  :   63 - 0x3f
    "00111111", -- 1442 - 0x5a2  :   63 - 0x3f
    "00111111", -- 1443 - 0x5a3  :   63 - 0x3f
    "00111111", -- 1444 - 0x5a4  :   63 - 0x3f
    "00111111", -- 1445 - 0x5a5  :   63 - 0x3f
    "00111111", -- 1446 - 0x5a6  :   63 - 0x3f
    "00111111", -- 1447 - 0x5a7  :   63 - 0x3f
    "00111111", -- 1448 - 0x5a8  :   63 - 0x3f
    "00111111", -- 1449 - 0x5a9  :   63 - 0x3f
    "00111111", -- 1450 - 0x5aa  :   63 - 0x3f
    "00111111", -- 1451 - 0x5ab  :   63 - 0x3f
    "00111111", -- 1452 - 0x5ac  :   63 - 0x3f
    "00111111", -- 1453 - 0x5ad  :   63 - 0x3f
    "00111111", -- 1454 - 0x5ae  :   63 - 0x3f
    "00111111", -- 1455 - 0x5af  :   63 - 0x3f
    "00111111", -- 1456 - 0x5b0  :   63 - 0x3f
    "00111111", -- 1457 - 0x5b1  :   63 - 0x3f
    "00111111", -- 1458 - 0x5b2  :   63 - 0x3f
    "00111111", -- 1459 - 0x5b3  :   63 - 0x3f
    "00111111", -- 1460 - 0x5b4  :   63 - 0x3f
    "00111111", -- 1461 - 0x5b5  :   63 - 0x3f
    "00111111", -- 1462 - 0x5b6  :   63 - 0x3f
    "00111111", -- 1463 - 0x5b7  :   63 - 0x3f
    "00111111", -- 1464 - 0x5b8  :   63 - 0x3f
    "00111111", -- 1465 - 0x5b9  :   63 - 0x3f
    "00111111", -- 1466 - 0x5ba  :   63 - 0x3f
    "00111111", -- 1467 - 0x5bb  :   63 - 0x3f
    "00111111", -- 1468 - 0x5bc  :   63 - 0x3f
    "00111111", -- 1469 - 0x5bd  :   63 - 0x3f
    "00111111", -- 1470 - 0x5be  :   63 - 0x3f
    "00111111", -- 1471 - 0x5bf  :   63 - 0x3f
    "00111111", -- 1472 - 0x5c0  :   63 - 0x3f -- line 0xe
    "00111111", -- 1473 - 0x5c1  :   63 - 0x3f
    "00111111", -- 1474 - 0x5c2  :   63 - 0x3f
    "00111111", -- 1475 - 0x5c3  :   63 - 0x3f
    "00111111", -- 1476 - 0x5c4  :   63 - 0x3f
    "00111111", -- 1477 - 0x5c5  :   63 - 0x3f
    "00111111", -- 1478 - 0x5c6  :   63 - 0x3f
    "00111111", -- 1479 - 0x5c7  :   63 - 0x3f
    "00111111", -- 1480 - 0x5c8  :   63 - 0x3f
    "00111111", -- 1481 - 0x5c9  :   63 - 0x3f
    "00111111", -- 1482 - 0x5ca  :   63 - 0x3f
    "00111111", -- 1483 - 0x5cb  :   63 - 0x3f
    "00111111", -- 1484 - 0x5cc  :   63 - 0x3f
    "00111111", -- 1485 - 0x5cd  :   63 - 0x3f
    "00111111", -- 1486 - 0x5ce  :   63 - 0x3f
    "00111111", -- 1487 - 0x5cf  :   63 - 0x3f
    "00111111", -- 1488 - 0x5d0  :   63 - 0x3f
    "00111111", -- 1489 - 0x5d1  :   63 - 0x3f
    "00111111", -- 1490 - 0x5d2  :   63 - 0x3f
    "00111111", -- 1491 - 0x5d3  :   63 - 0x3f
    "00111111", -- 1492 - 0x5d4  :   63 - 0x3f
    "00111111", -- 1493 - 0x5d5  :   63 - 0x3f
    "00111111", -- 1494 - 0x5d6  :   63 - 0x3f
    "00111111", -- 1495 - 0x5d7  :   63 - 0x3f
    "01010111", -- 1496 - 0x5d8  :   87 - 0x57
    "01011000", -- 1497 - 0x5d9  :   88 - 0x58
    "01011000", -- 1498 - 0x5da  :   88 - 0x58
    "01011000", -- 1499 - 0x5db  :   88 - 0x58
    "01011000", -- 1500 - 0x5dc  :   88 - 0x58
    "01011000", -- 1501 - 0x5dd  :   88 - 0x58
    "01011000", -- 1502 - 0x5de  :   88 - 0x58
    "01011000", -- 1503 - 0x5df  :   88 - 0x58
    "00111111", -- 1504 - 0x5e0  :   63 - 0x3f -- line 0xf
    "00111111", -- 1505 - 0x5e1  :   63 - 0x3f
    "00111111", -- 1506 - 0x5e2  :   63 - 0x3f
    "00111111", -- 1507 - 0x5e3  :   63 - 0x3f
    "00111111", -- 1508 - 0x5e4  :   63 - 0x3f
    "00111111", -- 1509 - 0x5e5  :   63 - 0x3f
    "00111111", -- 1510 - 0x5e6  :   63 - 0x3f
    "00111111", -- 1511 - 0x5e7  :   63 - 0x3f
    "00111111", -- 1512 - 0x5e8  :   63 - 0x3f
    "00111111", -- 1513 - 0x5e9  :   63 - 0x3f
    "00111111", -- 1514 - 0x5ea  :   63 - 0x3f
    "00111111", -- 1515 - 0x5eb  :   63 - 0x3f
    "00111111", -- 1516 - 0x5ec  :   63 - 0x3f
    "00111111", -- 1517 - 0x5ed  :   63 - 0x3f
    "00111111", -- 1518 - 0x5ee  :   63 - 0x3f
    "00111111", -- 1519 - 0x5ef  :   63 - 0x3f
    "00111111", -- 1520 - 0x5f0  :   63 - 0x3f
    "00111111", -- 1521 - 0x5f1  :   63 - 0x3f
    "00111111", -- 1522 - 0x5f2  :   63 - 0x3f
    "00111111", -- 1523 - 0x5f3  :   63 - 0x3f
    "00111111", -- 1524 - 0x5f4  :   63 - 0x3f
    "00111111", -- 1525 - 0x5f5  :   63 - 0x3f
    "00111111", -- 1526 - 0x5f6  :   63 - 0x3f
    "00111111", -- 1527 - 0x5f7  :   63 - 0x3f
    "00111111", -- 1528 - 0x5f8  :   63 - 0x3f
    "00111111", -- 1529 - 0x5f9  :   63 - 0x3f
    "00111111", -- 1530 - 0x5fa  :   63 - 0x3f
    "00111111", -- 1531 - 0x5fb  :   63 - 0x3f
    "00111111", -- 1532 - 0x5fc  :   63 - 0x3f
    "00111111", -- 1533 - 0x5fd  :   63 - 0x3f
    "00111111", -- 1534 - 0x5fe  :   63 - 0x3f
    "00111111", -- 1535 - 0x5ff  :   63 - 0x3f
    "00111111", -- 1536 - 0x600  :   63 - 0x3f -- line 0x10
    "00111111", -- 1537 - 0x601  :   63 - 0x3f
    "00111111", -- 1538 - 0x602  :   63 - 0x3f
    "00111111", -- 1539 - 0x603  :   63 - 0x3f
    "00111111", -- 1540 - 0x604  :   63 - 0x3f
    "00111111", -- 1541 - 0x605  :   63 - 0x3f
    "00111111", -- 1542 - 0x606  :   63 - 0x3f
    "00111111", -- 1543 - 0x607  :   63 - 0x3f
    "00111111", -- 1544 - 0x608  :   63 - 0x3f
    "00111111", -- 1545 - 0x609  :   63 - 0x3f
    "00111111", -- 1546 - 0x60a  :   63 - 0x3f
    "00111111", -- 1547 - 0x60b  :   63 - 0x3f
    "00111111", -- 1548 - 0x60c  :   63 - 0x3f
    "00111111", -- 1549 - 0x60d  :   63 - 0x3f
    "00111111", -- 1550 - 0x60e  :   63 - 0x3f
    "00111111", -- 1551 - 0x60f  :   63 - 0x3f
    "00111111", -- 1552 - 0x610  :   63 - 0x3f
    "00111111", -- 1553 - 0x611  :   63 - 0x3f
    "00111111", -- 1554 - 0x612  :   63 - 0x3f
    "00111111", -- 1555 - 0x613  :   63 - 0x3f
    "00111111", -- 1556 - 0x614  :   63 - 0x3f
    "00111111", -- 1557 - 0x615  :   63 - 0x3f
    "00111111", -- 1558 - 0x616  :   63 - 0x3f
    "00111111", -- 1559 - 0x617  :   63 - 0x3f
    "00111111", -- 1560 - 0x618  :   63 - 0x3f
    "00111111", -- 1561 - 0x619  :   63 - 0x3f
    "00111111", -- 1562 - 0x61a  :   63 - 0x3f
    "00111111", -- 1563 - 0x61b  :   63 - 0x3f
    "00111111", -- 1564 - 0x61c  :   63 - 0x3f
    "00111111", -- 1565 - 0x61d  :   63 - 0x3f
    "00111111", -- 1566 - 0x61e  :   63 - 0x3f
    "00111111", -- 1567 - 0x61f  :   63 - 0x3f
    "00111111", -- 1568 - 0x620  :   63 - 0x3f -- line 0x11
    "00111111", -- 1569 - 0x621  :   63 - 0x3f
    "00111111", -- 1570 - 0x622  :   63 - 0x3f
    "00111111", -- 1571 - 0x623  :   63 - 0x3f
    "00111111", -- 1572 - 0x624  :   63 - 0x3f
    "00111111", -- 1573 - 0x625  :   63 - 0x3f
    "00111111", -- 1574 - 0x626  :   63 - 0x3f
    "00111111", -- 1575 - 0x627  :   63 - 0x3f
    "00111111", -- 1576 - 0x628  :   63 - 0x3f
    "00111111", -- 1577 - 0x629  :   63 - 0x3f
    "00111111", -- 1578 - 0x62a  :   63 - 0x3f
    "00111111", -- 1579 - 0x62b  :   63 - 0x3f
    "00111111", -- 1580 - 0x62c  :   63 - 0x3f
    "00111111", -- 1581 - 0x62d  :   63 - 0x3f
    "00111111", -- 1582 - 0x62e  :   63 - 0x3f
    "00111111", -- 1583 - 0x62f  :   63 - 0x3f
    "00111111", -- 1584 - 0x630  :   63 - 0x3f
    "00111111", -- 1585 - 0x631  :   63 - 0x3f
    "00111111", -- 1586 - 0x632  :   63 - 0x3f
    "00111111", -- 1587 - 0x633  :   63 - 0x3f
    "00111111", -- 1588 - 0x634  :   63 - 0x3f
    "00111111", -- 1589 - 0x635  :   63 - 0x3f
    "00111111", -- 1590 - 0x636  :   63 - 0x3f
    "00111111", -- 1591 - 0x637  :   63 - 0x3f
    "00111111", -- 1592 - 0x638  :   63 - 0x3f
    "00111111", -- 1593 - 0x639  :   63 - 0x3f
    "00111111", -- 1594 - 0x63a  :   63 - 0x3f
    "00111111", -- 1595 - 0x63b  :   63 - 0x3f
    "00111111", -- 1596 - 0x63c  :   63 - 0x3f
    "00111111", -- 1597 - 0x63d  :   63 - 0x3f
    "00111111", -- 1598 - 0x63e  :   63 - 0x3f
    "00111111", -- 1599 - 0x63f  :   63 - 0x3f
    "00111111", -- 1600 - 0x640  :   63 - 0x3f -- line 0x12
    "00111111", -- 1601 - 0x641  :   63 - 0x3f
    "00111111", -- 1602 - 0x642  :   63 - 0x3f
    "00111111", -- 1603 - 0x643  :   63 - 0x3f
    "00111111", -- 1604 - 0x644  :   63 - 0x3f
    "00111111", -- 1605 - 0x645  :   63 - 0x3f
    "00111111", -- 1606 - 0x646  :   63 - 0x3f
    "00111111", -- 1607 - 0x647  :   63 - 0x3f
    "00111111", -- 1608 - 0x648  :   63 - 0x3f
    "00111111", -- 1609 - 0x649  :   63 - 0x3f
    "00111111", -- 1610 - 0x64a  :   63 - 0x3f
    "00111111", -- 1611 - 0x64b  :   63 - 0x3f
    "11011100", -- 1612 - 0x64c  :  220 - 0xdc
    "11011101", -- 1613 - 0x64d  :  221 - 0xdd
    "11001100", -- 1614 - 0x64e  :  204 - 0xcc
    "11001101", -- 1615 - 0x64f  :  205 - 0xcd
    "00111111", -- 1616 - 0x650  :   63 - 0x3f
    "00111111", -- 1617 - 0x651  :   63 - 0x3f
    "00111111", -- 1618 - 0x652  :   63 - 0x3f
    "00111111", -- 1619 - 0x653  :   63 - 0x3f
    "00111111", -- 1620 - 0x654  :   63 - 0x3f
    "00111111", -- 1621 - 0x655  :   63 - 0x3f
    "00111111", -- 1622 - 0x656  :   63 - 0x3f
    "00111111", -- 1623 - 0x657  :   63 - 0x3f
    "00111111", -- 1624 - 0x658  :   63 - 0x3f
    "00111111", -- 1625 - 0x659  :   63 - 0x3f
    "00111111", -- 1626 - 0x65a  :   63 - 0x3f
    "00111111", -- 1627 - 0x65b  :   63 - 0x3f
    "00111111", -- 1628 - 0x65c  :   63 - 0x3f
    "00111111", -- 1629 - 0x65d  :   63 - 0x3f
    "00111111", -- 1630 - 0x65e  :   63 - 0x3f
    "00111111", -- 1631 - 0x65f  :   63 - 0x3f
    "00111111", -- 1632 - 0x660  :   63 - 0x3f -- line 0x13
    "00111111", -- 1633 - 0x661  :   63 - 0x3f
    "00111111", -- 1634 - 0x662  :   63 - 0x3f
    "00111111", -- 1635 - 0x663  :   63 - 0x3f
    "00111111", -- 1636 - 0x664  :   63 - 0x3f
    "00111111", -- 1637 - 0x665  :   63 - 0x3f
    "00111111", -- 1638 - 0x666  :   63 - 0x3f
    "00111111", -- 1639 - 0x667  :   63 - 0x3f
    "00111111", -- 1640 - 0x668  :   63 - 0x3f
    "00111111", -- 1641 - 0x669  :   63 - 0x3f
    "00111111", -- 1642 - 0x66a  :   63 - 0x3f
    "00111111", -- 1643 - 0x66b  :   63 - 0x3f
    "11011010", -- 1644 - 0x66c  :  218 - 0xda
    "11011011", -- 1645 - 0x66d  :  219 - 0xdb
    "11011010", -- 1646 - 0x66e  :  218 - 0xda
    "11011011", -- 1647 - 0x66f  :  219 - 0xdb
    "00111111", -- 1648 - 0x670  :   63 - 0x3f
    "00111111", -- 1649 - 0x671  :   63 - 0x3f
    "00011000", -- 1650 - 0x672  :   24 - 0x18
    "00011001", -- 1651 - 0x673  :   25 - 0x19
    "00111111", -- 1652 - 0x674  :   63 - 0x3f
    "00111111", -- 1653 - 0x675  :   63 - 0x3f
    "00111111", -- 1654 - 0x676  :   63 - 0x3f
    "00111111", -- 1655 - 0x677  :   63 - 0x3f
    "00111111", -- 1656 - 0x678  :   63 - 0x3f
    "00111111", -- 1657 - 0x679  :   63 - 0x3f
    "00111111", -- 1658 - 0x67a  :   63 - 0x3f
    "00111111", -- 1659 - 0x67b  :   63 - 0x3f
    "00111111", -- 1660 - 0x67c  :   63 - 0x3f
    "00111111", -- 1661 - 0x67d  :   63 - 0x3f
    "00111111", -- 1662 - 0x67e  :   63 - 0x3f
    "00111111", -- 1663 - 0x67f  :   63 - 0x3f
    "00111111", -- 1664 - 0x680  :   63 - 0x3f -- line 0x14
    "00111111", -- 1665 - 0x681  :   63 - 0x3f
    "00111111", -- 1666 - 0x682  :   63 - 0x3f
    "00111111", -- 1667 - 0x683  :   63 - 0x3f
    "00111111", -- 1668 - 0x684  :   63 - 0x3f
    "00111111", -- 1669 - 0x685  :   63 - 0x3f
    "00111111", -- 1670 - 0x686  :   63 - 0x3f
    "00111111", -- 1671 - 0x687  :   63 - 0x3f
    "00111111", -- 1672 - 0x688  :   63 - 0x3f
    "00111111", -- 1673 - 0x689  :   63 - 0x3f
    "01110000", -- 1674 - 0x68a  :  112 - 0x70
    "01110001", -- 1675 - 0x68b  :  113 - 0x71
    "01110001", -- 1676 - 0x68c  :  113 - 0x71
    "01110001", -- 1677 - 0x68d  :  113 - 0x71
    "01110001", -- 1678 - 0x68e  :  113 - 0x71
    "01110001", -- 1679 - 0x68f  :  113 - 0x71
    "01110001", -- 1680 - 0x690  :  113 - 0x71
    "01110001", -- 1681 - 0x691  :  113 - 0x71
    "01110001", -- 1682 - 0x692  :  113 - 0x71
    "01110001", -- 1683 - 0x693  :  113 - 0x71
    "01110001", -- 1684 - 0x694  :  113 - 0x71
    "01110010", -- 1685 - 0x695  :  114 - 0x72
    "00111111", -- 1686 - 0x696  :   63 - 0x3f
    "00111111", -- 1687 - 0x697  :   63 - 0x3f
    "00111111", -- 1688 - 0x698  :   63 - 0x3f
    "00111111", -- 1689 - 0x699  :   63 - 0x3f
    "00111111", -- 1690 - 0x69a  :   63 - 0x3f
    "00111111", -- 1691 - 0x69b  :   63 - 0x3f
    "00111111", -- 1692 - 0x69c  :   63 - 0x3f
    "00111111", -- 1693 - 0x69d  :   63 - 0x3f
    "00111111", -- 1694 - 0x69e  :   63 - 0x3f
    "00111111", -- 1695 - 0x69f  :   63 - 0x3f
    "00111111", -- 1696 - 0x6a0  :   63 - 0x3f -- line 0x15
    "00111111", -- 1697 - 0x6a1  :   63 - 0x3f
    "00111111", -- 1698 - 0x6a2  :   63 - 0x3f
    "00111111", -- 1699 - 0x6a3  :   63 - 0x3f
    "00111111", -- 1700 - 0x6a4  :   63 - 0x3f
    "00111111", -- 1701 - 0x6a5  :   63 - 0x3f
    "00111111", -- 1702 - 0x6a6  :   63 - 0x3f
    "00111111", -- 1703 - 0x6a7  :   63 - 0x3f
    "00111111", -- 1704 - 0x6a8  :   63 - 0x3f
    "00111111", -- 1705 - 0x6a9  :   63 - 0x3f
    "01100000", -- 1706 - 0x6aa  :   96 - 0x60
    "01110111", -- 1707 - 0x6ab  :  119 - 0x77
    "01110111", -- 1708 - 0x6ac  :  119 - 0x77
    "01110111", -- 1709 - 0x6ad  :  119 - 0x77
    "01110111", -- 1710 - 0x6ae  :  119 - 0x77
    "01110111", -- 1711 - 0x6af  :  119 - 0x77
    "01110111", -- 1712 - 0x6b0  :  119 - 0x77
    "01110111", -- 1713 - 0x6b1  :  119 - 0x77
    "01110111", -- 1714 - 0x6b2  :  119 - 0x77
    "01110111", -- 1715 - 0x6b3  :  119 - 0x77
    "01110111", -- 1716 - 0x6b4  :  119 - 0x77
    "01100001", -- 1717 - 0x6b5  :   97 - 0x61
    "00111111", -- 1718 - 0x6b6  :   63 - 0x3f
    "00111111", -- 1719 - 0x6b7  :   63 - 0x3f
    "00111111", -- 1720 - 0x6b8  :   63 - 0x3f
    "00111111", -- 1721 - 0x6b9  :   63 - 0x3f
    "00111111", -- 1722 - 0x6ba  :   63 - 0x3f
    "00111111", -- 1723 - 0x6bb  :   63 - 0x3f
    "00111111", -- 1724 - 0x6bc  :   63 - 0x3f
    "00111111", -- 1725 - 0x6bd  :   63 - 0x3f
    "00111111", -- 1726 - 0x6be  :   63 - 0x3f
    "00111111", -- 1727 - 0x6bf  :   63 - 0x3f
    "00111111", -- 1728 - 0x6c0  :   63 - 0x3f -- line 0x16
    "00111111", -- 1729 - 0x6c1  :   63 - 0x3f
    "00111111", -- 1730 - 0x6c2  :   63 - 0x3f
    "00111111", -- 1731 - 0x6c3  :   63 - 0x3f
    "00111111", -- 1732 - 0x6c4  :   63 - 0x3f
    "00111111", -- 1733 - 0x6c5  :   63 - 0x3f
    "00111111", -- 1734 - 0x6c6  :   63 - 0x3f
    "00111111", -- 1735 - 0x6c7  :   63 - 0x3f
    "00111111", -- 1736 - 0x6c8  :   63 - 0x3f
    "00111111", -- 1737 - 0x6c9  :   63 - 0x3f
    "01100000", -- 1738 - 0x6ca  :   96 - 0x60
    "01110011", -- 1739 - 0x6cb  :  115 - 0x73
    "01110011", -- 1740 - 0x6cc  :  115 - 0x73
    "01110011", -- 1741 - 0x6cd  :  115 - 0x73
    "01110011", -- 1742 - 0x6ce  :  115 - 0x73
    "01110011", -- 1743 - 0x6cf  :  115 - 0x73
    "01110011", -- 1744 - 0x6d0  :  115 - 0x73
    "01110011", -- 1745 - 0x6d1  :  115 - 0x73
    "01110011", -- 1746 - 0x6d2  :  115 - 0x73
    "01110011", -- 1747 - 0x6d3  :  115 - 0x73
    "01110011", -- 1748 - 0x6d4  :  115 - 0x73
    "01100001", -- 1749 - 0x6d5  :   97 - 0x61
    "00111111", -- 1750 - 0x6d6  :   63 - 0x3f
    "00111111", -- 1751 - 0x6d7  :   63 - 0x3f
    "00111111", -- 1752 - 0x6d8  :   63 - 0x3f
    "00111111", -- 1753 - 0x6d9  :   63 - 0x3f
    "00111111", -- 1754 - 0x6da  :   63 - 0x3f
    "00111111", -- 1755 - 0x6db  :   63 - 0x3f
    "00111111", -- 1756 - 0x6dc  :   63 - 0x3f
    "00111111", -- 1757 - 0x6dd  :   63 - 0x3f
    "00111111", -- 1758 - 0x6de  :   63 - 0x3f
    "00111111", -- 1759 - 0x6df  :   63 - 0x3f
    "11000101", -- 1760 - 0x6e0  :  197 - 0xc5 -- line 0x17
    "11010110", -- 1761 - 0x6e1  :  214 - 0xd6
    "00111111", -- 1762 - 0x6e2  :   63 - 0x3f
    "00111111", -- 1763 - 0x6e3  :   63 - 0x3f
    "00111111", -- 1764 - 0x6e4  :   63 - 0x3f
    "00111111", -- 1765 - 0x6e5  :   63 - 0x3f
    "00111111", -- 1766 - 0x6e6  :   63 - 0x3f
    "00111111", -- 1767 - 0x6e7  :   63 - 0x3f
    "00111111", -- 1768 - 0x6e8  :   63 - 0x3f
    "00111111", -- 1769 - 0x6e9  :   63 - 0x3f
    "01100000", -- 1770 - 0x6ea  :   96 - 0x60
    "01110011", -- 1771 - 0x6eb  :  115 - 0x73
    "01110011", -- 1772 - 0x6ec  :  115 - 0x73
    "01110011", -- 1773 - 0x6ed  :  115 - 0x73
    "01110011", -- 1774 - 0x6ee  :  115 - 0x73
    "01110011", -- 1775 - 0x6ef  :  115 - 0x73
    "01110011", -- 1776 - 0x6f0  :  115 - 0x73
    "01110011", -- 1777 - 0x6f1  :  115 - 0x73
    "01110011", -- 1778 - 0x6f2  :  115 - 0x73
    "01110011", -- 1779 - 0x6f3  :  115 - 0x73
    "01110011", -- 1780 - 0x6f4  :  115 - 0x73
    "01100001", -- 1781 - 0x6f5  :   97 - 0x61
    "00111111", -- 1782 - 0x6f6  :   63 - 0x3f
    "00111111", -- 1783 - 0x6f7  :   63 - 0x3f
    "00111111", -- 1784 - 0x6f8  :   63 - 0x3f
    "00111111", -- 1785 - 0x6f9  :   63 - 0x3f
    "00111111", -- 1786 - 0x6fa  :   63 - 0x3f
    "00111111", -- 1787 - 0x6fb  :   63 - 0x3f
    "00111111", -- 1788 - 0x6fc  :   63 - 0x3f
    "00111111", -- 1789 - 0x6fd  :   63 - 0x3f
    "00111111", -- 1790 - 0x6fe  :   63 - 0x3f
    "00111111", -- 1791 - 0x6ff  :   63 - 0x3f
    "11000111", -- 1792 - 0x700  :  199 - 0xc7 -- line 0x18
    "11001001", -- 1793 - 0x701  :  201 - 0xc9
    "00111111", -- 1794 - 0x702  :   63 - 0x3f
    "00111111", -- 1795 - 0x703  :   63 - 0x3f
    "00111111", -- 1796 - 0x704  :   63 - 0x3f
    "00111111", -- 1797 - 0x705  :   63 - 0x3f
    "00111111", -- 1798 - 0x706  :   63 - 0x3f
    "00111111", -- 1799 - 0x707  :   63 - 0x3f
    "00111111", -- 1800 - 0x708  :   63 - 0x3f
    "00111111", -- 1801 - 0x709  :   63 - 0x3f
    "01100000", -- 1802 - 0x70a  :   96 - 0x60
    "01110011", -- 1803 - 0x70b  :  115 - 0x73
    "01110011", -- 1804 - 0x70c  :  115 - 0x73
    "01110011", -- 1805 - 0x70d  :  115 - 0x73
    "01110011", -- 1806 - 0x70e  :  115 - 0x73
    "01110011", -- 1807 - 0x70f  :  115 - 0x73
    "01110011", -- 1808 - 0x710  :  115 - 0x73
    "01110011", -- 1809 - 0x711  :  115 - 0x73
    "01110011", -- 1810 - 0x712  :  115 - 0x73
    "01110011", -- 1811 - 0x713  :  115 - 0x73
    "01110011", -- 1812 - 0x714  :  115 - 0x73
    "01100001", -- 1813 - 0x715  :   97 - 0x61
    "00111111", -- 1814 - 0x716  :   63 - 0x3f
    "00111111", -- 1815 - 0x717  :   63 - 0x3f
    "00111111", -- 1816 - 0x718  :   63 - 0x3f
    "00111111", -- 1817 - 0x719  :   63 - 0x3f
    "00111111", -- 1818 - 0x71a  :   63 - 0x3f
    "00111111", -- 1819 - 0x71b  :   63 - 0x3f
    "00111111", -- 1820 - 0x71c  :   63 - 0x3f
    "00111111", -- 1821 - 0x71d  :   63 - 0x3f
    "00111111", -- 1822 - 0x71e  :   63 - 0x3f
    "00111111", -- 1823 - 0x71f  :   63 - 0x3f
    "11010111", -- 1824 - 0x720  :  215 - 0xd7 -- line 0x19
    "11011001", -- 1825 - 0x721  :  217 - 0xd9
    "00111111", -- 1826 - 0x722  :   63 - 0x3f
    "00111111", -- 1827 - 0x723  :   63 - 0x3f
    "00111111", -- 1828 - 0x724  :   63 - 0x3f
    "00111111", -- 1829 - 0x725  :   63 - 0x3f
    "00111111", -- 1830 - 0x726  :   63 - 0x3f
    "00111111", -- 1831 - 0x727  :   63 - 0x3f
    "00011000", -- 1832 - 0x728  :   24 - 0x18
    "00011001", -- 1833 - 0x729  :   25 - 0x19
    "01100000", -- 1834 - 0x72a  :   96 - 0x60
    "01110011", -- 1835 - 0x72b  :  115 - 0x73
    "01110011", -- 1836 - 0x72c  :  115 - 0x73
    "01110011", -- 1837 - 0x72d  :  115 - 0x73
    "01110011", -- 1838 - 0x72e  :  115 - 0x73
    "01110011", -- 1839 - 0x72f  :  115 - 0x73
    "01110011", -- 1840 - 0x730  :  115 - 0x73
    "01110011", -- 1841 - 0x731  :  115 - 0x73
    "01110011", -- 1842 - 0x732  :  115 - 0x73
    "01110011", -- 1843 - 0x733  :  115 - 0x73
    "01110011", -- 1844 - 0x734  :  115 - 0x73
    "01100001", -- 1845 - 0x735  :   97 - 0x61
    "00111111", -- 1846 - 0x736  :   63 - 0x3f
    "00111111", -- 1847 - 0x737  :   63 - 0x3f
    "00111111", -- 1848 - 0x738  :   63 - 0x3f
    "00111111", -- 1849 - 0x739  :   63 - 0x3f
    "00111111", -- 1850 - 0x73a  :   63 - 0x3f
    "00111111", -- 1851 - 0x73b  :   63 - 0x3f
    "00111111", -- 1852 - 0x73c  :   63 - 0x3f
    "00111111", -- 1853 - 0x73d  :   63 - 0x3f
    "00111111", -- 1854 - 0x73e  :   63 - 0x3f
    "00111111", -- 1855 - 0x73f  :   63 - 0x3f
    "01110001", -- 1856 - 0x740  :  113 - 0x71 -- line 0x1a
    "01110001", -- 1857 - 0x741  :  113 - 0x71
    "01110001", -- 1858 - 0x742  :  113 - 0x71
    "01110001", -- 1859 - 0x743  :  113 - 0x71
    "01110001", -- 1860 - 0x744  :  113 - 0x71
    "01110001", -- 1861 - 0x745  :  113 - 0x71
    "01110001", -- 1862 - 0x746  :  113 - 0x71
    "01110001", -- 1863 - 0x747  :  113 - 0x71
    "01110001", -- 1864 - 0x748  :  113 - 0x71
    "01110001", -- 1865 - 0x749  :  113 - 0x71
    "01100000", -- 1866 - 0x74a  :   96 - 0x60
    "01110011", -- 1867 - 0x74b  :  115 - 0x73
    "01110011", -- 1868 - 0x74c  :  115 - 0x73
    "01110011", -- 1869 - 0x74d  :  115 - 0x73
    "01110011", -- 1870 - 0x74e  :  115 - 0x73
    "01110011", -- 1871 - 0x74f  :  115 - 0x73
    "01110011", -- 1872 - 0x750  :  115 - 0x73
    "01110011", -- 1873 - 0x751  :  115 - 0x73
    "01110011", -- 1874 - 0x752  :  115 - 0x73
    "01110011", -- 1875 - 0x753  :  115 - 0x73
    "01110011", -- 1876 - 0x754  :  115 - 0x73
    "01100001", -- 1877 - 0x755  :   97 - 0x61
    "00111111", -- 1878 - 0x756  :   63 - 0x3f
    "00111111", -- 1879 - 0x757  :   63 - 0x3f
    "00111111", -- 1880 - 0x758  :   63 - 0x3f
    "00111111", -- 1881 - 0x759  :   63 - 0x3f
    "00111111", -- 1882 - 0x75a  :   63 - 0x3f
    "00111111", -- 1883 - 0x75b  :   63 - 0x3f
    "00111111", -- 1884 - 0x75c  :   63 - 0x3f
    "00111111", -- 1885 - 0x75d  :   63 - 0x3f
    "00111111", -- 1886 - 0x75e  :   63 - 0x3f
    "00111111", -- 1887 - 0x75f  :   63 - 0x3f
    "01110111", -- 1888 - 0x760  :  119 - 0x77 -- line 0x1b
    "01110111", -- 1889 - 0x761  :  119 - 0x77
    "01110111", -- 1890 - 0x762  :  119 - 0x77
    "01110111", -- 1891 - 0x763  :  119 - 0x77
    "01110111", -- 1892 - 0x764  :  119 - 0x77
    "01110111", -- 1893 - 0x765  :  119 - 0x77
    "01110111", -- 1894 - 0x766  :  119 - 0x77
    "01110111", -- 1895 - 0x767  :  119 - 0x77
    "01110111", -- 1896 - 0x768  :  119 - 0x77
    "01110111", -- 1897 - 0x769  :  119 - 0x77
    "01110011", -- 1898 - 0x76a  :  115 - 0x73
    "01110011", -- 1899 - 0x76b  :  115 - 0x73
    "01110011", -- 1900 - 0x76c  :  115 - 0x73
    "01110011", -- 1901 - 0x76d  :  115 - 0x73
    "01110011", -- 1902 - 0x76e  :  115 - 0x73
    "01110011", -- 1903 - 0x76f  :  115 - 0x73
    "01110011", -- 1904 - 0x770  :  115 - 0x73
    "01110011", -- 1905 - 0x771  :  115 - 0x73
    "01110011", -- 1906 - 0x772  :  115 - 0x73
    "01110011", -- 1907 - 0x773  :  115 - 0x73
    "01110011", -- 1908 - 0x774  :  115 - 0x73
    "01100001", -- 1909 - 0x775  :   97 - 0x61
    "00111111", -- 1910 - 0x776  :   63 - 0x3f
    "00111111", -- 1911 - 0x777  :   63 - 0x3f
    "00111111", -- 1912 - 0x778  :   63 - 0x3f
    "00111111", -- 1913 - 0x779  :   63 - 0x3f
    "00111111", -- 1914 - 0x77a  :   63 - 0x3f
    "00111111", -- 1915 - 0x77b  :   63 - 0x3f
    "00111111", -- 1916 - 0x77c  :   63 - 0x3f
    "00111111", -- 1917 - 0x77d  :   63 - 0x3f
    "00111111", -- 1918 - 0x77e  :   63 - 0x3f
    "00111111", -- 1919 - 0x77f  :   63 - 0x3f
    "01110011", -- 1920 - 0x780  :  115 - 0x73 -- line 0x1c
    "01110011", -- 1921 - 0x781  :  115 - 0x73
    "01110011", -- 1922 - 0x782  :  115 - 0x73
    "01110011", -- 1923 - 0x783  :  115 - 0x73
    "01110011", -- 1924 - 0x784  :  115 - 0x73
    "01110011", -- 1925 - 0x785  :  115 - 0x73
    "01110011", -- 1926 - 0x786  :  115 - 0x73
    "01110011", -- 1927 - 0x787  :  115 - 0x73
    "01110011", -- 1928 - 0x788  :  115 - 0x73
    "01110011", -- 1929 - 0x789  :  115 - 0x73
    "01110011", -- 1930 - 0x78a  :  115 - 0x73
    "01110011", -- 1931 - 0x78b  :  115 - 0x73
    "01110011", -- 1932 - 0x78c  :  115 - 0x73
    "01110011", -- 1933 - 0x78d  :  115 - 0x73
    "01110011", -- 1934 - 0x78e  :  115 - 0x73
    "01110011", -- 1935 - 0x78f  :  115 - 0x73
    "01110011", -- 1936 - 0x790  :  115 - 0x73
    "01110011", -- 1937 - 0x791  :  115 - 0x73
    "01110011", -- 1938 - 0x792  :  115 - 0x73
    "01110011", -- 1939 - 0x793  :  115 - 0x73
    "01110011", -- 1940 - 0x794  :  115 - 0x73
    "01100001", -- 1941 - 0x795  :   97 - 0x61
    "00111111", -- 1942 - 0x796  :   63 - 0x3f
    "00111111", -- 1943 - 0x797  :   63 - 0x3f
    "00111111", -- 1944 - 0x798  :   63 - 0x3f
    "00111111", -- 1945 - 0x799  :   63 - 0x3f
    "00111111", -- 1946 - 0x79a  :   63 - 0x3f
    "00111111", -- 1947 - 0x79b  :   63 - 0x3f
    "00111111", -- 1948 - 0x79c  :   63 - 0x3f
    "00111111", -- 1949 - 0x79d  :   63 - 0x3f
    "00111111", -- 1950 - 0x79e  :   63 - 0x3f
    "00111111", -- 1951 - 0x79f  :   63 - 0x3f
    "01110011", -- 1952 - 0x7a0  :  115 - 0x73 -- line 0x1d
    "01110011", -- 1953 - 0x7a1  :  115 - 0x73
    "01110011", -- 1954 - 0x7a2  :  115 - 0x73
    "01110011", -- 1955 - 0x7a3  :  115 - 0x73
    "01110011", -- 1956 - 0x7a4  :  115 - 0x73
    "01110011", -- 1957 - 0x7a5  :  115 - 0x73
    "01110011", -- 1958 - 0x7a6  :  115 - 0x73
    "01110011", -- 1959 - 0x7a7  :  115 - 0x73
    "01110011", -- 1960 - 0x7a8  :  115 - 0x73
    "01110011", -- 1961 - 0x7a9  :  115 - 0x73
    "01110011", -- 1962 - 0x7aa  :  115 - 0x73
    "01110011", -- 1963 - 0x7ab  :  115 - 0x73
    "01110011", -- 1964 - 0x7ac  :  115 - 0x73
    "01110011", -- 1965 - 0x7ad  :  115 - 0x73
    "01110011", -- 1966 - 0x7ae  :  115 - 0x73
    "01110011", -- 1967 - 0x7af  :  115 - 0x73
    "01110011", -- 1968 - 0x7b0  :  115 - 0x73
    "01110011", -- 1969 - 0x7b1  :  115 - 0x73
    "01110011", -- 1970 - 0x7b2  :  115 - 0x73
    "01110011", -- 1971 - 0x7b3  :  115 - 0x73
    "01110011", -- 1972 - 0x7b4  :  115 - 0x73
    "01100001", -- 1973 - 0x7b5  :   97 - 0x61
    "00111111", -- 1974 - 0x7b6  :   63 - 0x3f
    "00111111", -- 1975 - 0x7b7  :   63 - 0x3f
    "00111111", -- 1976 - 0x7b8  :   63 - 0x3f
    "00111111", -- 1977 - 0x7b9  :   63 - 0x3f
    "00111111", -- 1978 - 0x7ba  :   63 - 0x3f
    "00111111", -- 1979 - 0x7bb  :   63 - 0x3f
    "00111111", -- 1980 - 0x7bc  :   63 - 0x3f
    "00111111", -- 1981 - 0x7bd  :   63 - 0x3f
    "00111111", -- 1982 - 0x7be  :   63 - 0x3f
    "00111111", -- 1983 - 0x7bf  :   63 - 0x3f
        ---- Attribute Table 1----
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "10001000", -- 1986 - 0x7c2  :  136 - 0x88
    "00010001", -- 1987 - 0x7c3  :   17 - 0x11
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00001010", -- 1992 - 0x7c8  :   10 - 0xa
    "00000010", -- 1993 - 0x7c9  :    2 - 0x2
    "10001000", -- 1994 - 0x7ca  :  136 - 0x88
    "00010001", -- 1995 - 0x7cb  :   17 - 0x11
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "01010100", -- 2000 - 0x7d0  :   84 - 0x54
    "00000101", -- 2001 - 0x7d1  :    5 - 0x5
    "00000101", -- 2002 - 0x7d2  :    5 - 0x5
    "00000001", -- 2003 - 0x7d3  :    1 - 0x1
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "10000000", -- 2006 - 0x7d6  :  128 - 0x80
    "10100000", -- 2007 - 0x7d7  :  160 - 0xa0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "01010000", -- 2014 - 0x7de  :   80 - 0x50
    "01010000", -- 2015 - 0x7df  :   80 - 0x50
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "10000000", -- 2020 - 0x7e4  :  128 - 0x80
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000010", -- 2034 - 0x7f2  :    2 - 0x2
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
