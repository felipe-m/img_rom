//-   Sprites Pattern table COLOR PLANE 0
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: donkeykong_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_DONKEYKONG_SPR_PLN0
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table COLOR PLANE 0
      11'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      11'h1: dout  = 8'b00000011; //    1 :   3 - 0x3
      11'h2: dout  = 8'b00000111; //    2 :   7 - 0x7
      11'h3: dout  = 8'b00000111; //    3 :   7 - 0x7
      11'h4: dout  = 8'b00001001; //    4 :   9 - 0x9
      11'h5: dout  = 8'b00001001; //    5 :   9 - 0x9
      11'h6: dout  = 8'b00011100; //    6 :  28 - 0x1c
      11'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      11'h8: dout  = 8'b00001111; //    8 :  15 - 0xf -- Sprite 0x1
      11'h9: dout  = 8'b00001111; //    9 :  15 - 0xf
      11'hA: dout  = 8'b00001111; //   10 :  15 - 0xf
      11'hB: dout  = 8'b11111111; //   11 : 255 - 0xff
      11'hC: dout  = 8'b11111111; //   12 : 255 - 0xff
      11'hD: dout  = 8'b11111100; //   13 : 252 - 0xfc
      11'hE: dout  = 8'b10000001; //   14 : 129 - 0x81
      11'hF: dout  = 8'b00000001; //   15 :   1 - 0x1
      11'h10: dout  = 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x2
      11'h11: dout  = 8'b11000000; //   17 : 192 - 0xc0
      11'h12: dout  = 8'b11111000; //   18 : 248 - 0xf8
      11'h13: dout  = 8'b10000000; //   19 : 128 - 0x80
      11'h14: dout  = 8'b00100000; //   20 :  32 - 0x20
      11'h15: dout  = 8'b10010000; //   21 : 144 - 0x90
      11'h16: dout  = 8'b00111100; //   22 :  60 - 0x3c
      11'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      11'h18: dout  = 8'b11000000; //   24 : 192 - 0xc0 -- Sprite 0x3
      11'h19: dout  = 8'b11000000; //   25 : 192 - 0xc0
      11'h1A: dout  = 8'b11000000; //   26 : 192 - 0xc0
      11'h1B: dout  = 8'b11110000; //   27 : 240 - 0xf0
      11'h1C: dout  = 8'b11110000; //   28 : 240 - 0xf0
      11'h1D: dout  = 8'b11100000; //   29 : 224 - 0xe0
      11'h1E: dout  = 8'b11000000; //   30 : 192 - 0xc0
      11'h1F: dout  = 8'b11100000; //   31 : 224 - 0xe0
      11'h20: dout  = 8'b00000111; //   32 :   7 - 0x7 -- Sprite 0x4
      11'h21: dout  = 8'b00001111; //   33 :  15 - 0xf
      11'h22: dout  = 8'b00001111; //   34 :  15 - 0xf
      11'h23: dout  = 8'b00010010; //   35 :  18 - 0x12
      11'h24: dout  = 8'b00010011; //   36 :  19 - 0x13
      11'h25: dout  = 8'b00111000; //   37 :  56 - 0x38
      11'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      11'h27: dout  = 8'b00001111; //   39 :  15 - 0xf
      11'h28: dout  = 8'b00011111; //   40 :  31 - 0x1f -- Sprite 0x5
      11'h29: dout  = 8'b00011111; //   41 :  31 - 0x1f
      11'h2A: dout  = 8'b00011111; //   42 :  31 - 0x1f
      11'h2B: dout  = 8'b00011000; //   43 :  24 - 0x18
      11'h2C: dout  = 8'b00011001; //   44 :  25 - 0x19
      11'h2D: dout  = 8'b00011110; //   45 :  30 - 0x1e
      11'h2E: dout  = 8'b00011100; //   46 :  28 - 0x1c
      11'h2F: dout  = 8'b00011110; //   47 :  30 - 0x1e
      11'h30: dout  = 8'b10000000; //   48 : 128 - 0x80 -- Sprite 0x6
      11'h31: dout  = 8'b11110000; //   49 : 240 - 0xf0
      11'h32: dout  = 8'b00000000; //   50 :   0 - 0x0
      11'h33: dout  = 8'b01000000; //   51 :  64 - 0x40
      11'h34: dout  = 8'b00100000; //   52 :  32 - 0x20
      11'h35: dout  = 8'b01111000; //   53 : 120 - 0x78
      11'h36: dout  = 8'b00000000; //   54 :   0 - 0x0
      11'h37: dout  = 8'b11000000; //   55 : 192 - 0xc0
      11'h38: dout  = 8'b11100000; //   56 : 224 - 0xe0 -- Sprite 0x7
      11'h39: dout  = 8'b01100000; //   57 :  96 - 0x60
      11'h3A: dout  = 8'b11110000; //   58 : 240 - 0xf0
      11'h3B: dout  = 8'b11110000; //   59 : 240 - 0xf0
      11'h3C: dout  = 8'b11110000; //   60 : 240 - 0xf0
      11'h3D: dout  = 8'b11100000; //   61 : 224 - 0xe0
      11'h3E: dout  = 8'b11100000; //   62 : 224 - 0xe0
      11'h3F: dout  = 8'b11110000; //   63 : 240 - 0xf0
      11'h40: dout  = 8'b00000111; //   64 :   7 - 0x7 -- Sprite 0x8
      11'h41: dout  = 8'b00001111; //   65 :  15 - 0xf
      11'h42: dout  = 8'b00001111; //   66 :  15 - 0xf
      11'h43: dout  = 8'b00010010; //   67 :  18 - 0x12
      11'h44: dout  = 8'b00010011; //   68 :  19 - 0x13
      11'h45: dout  = 8'b00111000; //   69 :  56 - 0x38
      11'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      11'h47: dout  = 8'b00111111; //   71 :  63 - 0x3f
      11'h48: dout  = 8'b00111111; //   72 :  63 - 0x3f -- Sprite 0x9
      11'h49: dout  = 8'b00001110; //   73 :  14 - 0xe
      11'h4A: dout  = 8'b00001111; //   74 :  15 - 0xf
      11'h4B: dout  = 8'b00011111; //   75 :  31 - 0x1f
      11'h4C: dout  = 8'b00111111; //   76 :  63 - 0x3f
      11'h4D: dout  = 8'b01111100; //   77 : 124 - 0x7c
      11'h4E: dout  = 8'b01110000; //   78 : 112 - 0x70
      11'h4F: dout  = 8'b00111000; //   79 :  56 - 0x38
      11'h50: dout  = 8'b10000000; //   80 : 128 - 0x80 -- Sprite 0xa
      11'h51: dout  = 8'b11110000; //   81 : 240 - 0xf0
      11'h52: dout  = 8'b00000000; //   82 :   0 - 0x0
      11'h53: dout  = 8'b01000000; //   83 :  64 - 0x40
      11'h54: dout  = 8'b00100000; //   84 :  32 - 0x20
      11'h55: dout  = 8'b01111000; //   85 : 120 - 0x78
      11'h56: dout  = 8'b00000000; //   86 :   0 - 0x0
      11'h57: dout  = 8'b11000000; //   87 : 192 - 0xc0
      11'h58: dout  = 8'b11110000; //   88 : 240 - 0xf0 -- Sprite 0xb
      11'h59: dout  = 8'b11111000; //   89 : 248 - 0xf8
      11'h5A: dout  = 8'b11100100; //   90 : 228 - 0xe4
      11'h5B: dout  = 8'b11111100; //   91 : 252 - 0xfc
      11'h5C: dout  = 8'b11111100; //   92 : 252 - 0xfc
      11'h5D: dout  = 8'b01111100; //   93 : 124 - 0x7c
      11'h5E: dout  = 8'b00000000; //   94 :   0 - 0x0
      11'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      11'h60: dout  = 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0xc
      11'h61: dout  = 8'b00000010; //   97 :   2 - 0x2
      11'h62: dout  = 8'b00000110; //   98 :   6 - 0x6
      11'h63: dout  = 8'b00000111; //   99 :   7 - 0x7
      11'h64: dout  = 8'b00001001; //  100 :   9 - 0x9
      11'h65: dout  = 8'b00001001; //  101 :   9 - 0x9
      11'h66: dout  = 8'b00011101; //  102 :  29 - 0x1d
      11'h67: dout  = 8'b00000011; //  103 :   3 - 0x3
      11'h68: dout  = 8'b00001111; //  104 :  15 - 0xf -- Sprite 0xd
      11'h69: dout  = 8'b00001111; //  105 :  15 - 0xf
      11'h6A: dout  = 8'b00001111; //  106 :  15 - 0xf
      11'h6B: dout  = 8'b11111111; //  107 : 255 - 0xff
      11'h6C: dout  = 8'b11111111; //  108 : 255 - 0xff
      11'h6D: dout  = 8'b11111100; //  109 : 252 - 0xfc
      11'h6E: dout  = 8'b10000001; //  110 : 129 - 0x81
      11'h6F: dout  = 8'b00000001; //  111 :   1 - 0x1
      11'h70: dout  = 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0xe
      11'h71: dout  = 8'b00000000; //  113 :   0 - 0x0
      11'h72: dout  = 8'b00111000; //  114 :  56 - 0x38
      11'h73: dout  = 8'b11000000; //  115 : 192 - 0xc0
      11'h74: dout  = 8'b11100000; //  116 : 224 - 0xe0
      11'h75: dout  = 8'b11010000; //  117 : 208 - 0xd0
      11'h76: dout  = 8'b11111100; //  118 : 252 - 0xfc
      11'h77: dout  = 8'b11000000; //  119 : 192 - 0xc0
      11'h78: dout  = 8'b11100000; //  120 : 224 - 0xe0 -- Sprite 0xf
      11'h79: dout  = 8'b11100000; //  121 : 224 - 0xe0
      11'h7A: dout  = 8'b10110000; //  122 : 176 - 0xb0
      11'h7B: dout  = 8'b11110000; //  123 : 240 - 0xf0
      11'h7C: dout  = 8'b11110000; //  124 : 240 - 0xf0
      11'h7D: dout  = 8'b11100000; //  125 : 224 - 0xe0
      11'h7E: dout  = 8'b11000000; //  126 : 192 - 0xc0
      11'h7F: dout  = 8'b11100000; //  127 : 224 - 0xe0
      11'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      11'h81: dout  = 8'b00000011; //  129 :   3 - 0x3
      11'h82: dout  = 8'b00000111; //  130 :   7 - 0x7
      11'h83: dout  = 8'b00000111; //  131 :   7 - 0x7
      11'h84: dout  = 8'b00001001; //  132 :   9 - 0x9
      11'h85: dout  = 8'b00001001; //  133 :   9 - 0x9
      11'h86: dout  = 8'b00011100; //  134 :  28 - 0x1c
      11'h87: dout  = 8'b00000000; //  135 :   0 - 0x0
      11'h88: dout  = 8'b00001111; //  136 :  15 - 0xf -- Sprite 0x11
      11'h89: dout  = 8'b00001111; //  137 :  15 - 0xf
      11'h8A: dout  = 8'b00001111; //  138 :  15 - 0xf
      11'h8B: dout  = 8'b11111111; //  139 : 255 - 0xff
      11'h8C: dout  = 8'b11111111; //  140 : 255 - 0xff
      11'h8D: dout  = 8'b11111100; //  141 : 252 - 0xfc
      11'h8E: dout  = 8'b10000001; //  142 : 129 - 0x81
      11'h8F: dout  = 8'b00000001; //  143 :   1 - 0x1
      11'h90: dout  = 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x12
      11'h91: dout  = 8'b11000000; //  145 : 192 - 0xc0
      11'h92: dout  = 8'b11111000; //  146 : 248 - 0xf8
      11'h93: dout  = 8'b10000000; //  147 : 128 - 0x80
      11'h94: dout  = 8'b00100000; //  148 :  32 - 0x20
      11'h95: dout  = 8'b10010000; //  149 : 144 - 0x90
      11'h96: dout  = 8'b00111100; //  150 :  60 - 0x3c
      11'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      11'h98: dout  = 8'b11100000; //  152 : 224 - 0xe0 -- Sprite 0x13
      11'h99: dout  = 8'b11110000; //  153 : 240 - 0xf0
      11'h9A: dout  = 8'b11110000; //  154 : 240 - 0xf0
      11'h9B: dout  = 8'b11110000; //  155 : 240 - 0xf0
      11'h9C: dout  = 8'b11110000; //  156 : 240 - 0xf0
      11'h9D: dout  = 8'b11100000; //  157 : 224 - 0xe0
      11'h9E: dout  = 8'b11000000; //  158 : 192 - 0xc0
      11'h9F: dout  = 8'b11100000; //  159 : 224 - 0xe0
      11'hA0: dout  = 8'b00000100; //  160 :   4 - 0x4 -- Sprite 0x14
      11'hA1: dout  = 8'b00001100; //  161 :  12 - 0xc
      11'hA2: dout  = 8'b00001100; //  162 :  12 - 0xc
      11'hA3: dout  = 8'b00010011; //  163 :  19 - 0x13
      11'hA4: dout  = 8'b00010011; //  164 :  19 - 0x13
      11'hA5: dout  = 8'b00111011; //  165 :  59 - 0x3b
      11'hA6: dout  = 8'b00000111; //  166 :   7 - 0x7
      11'hA7: dout  = 8'b00001111; //  167 :  15 - 0xf
      11'hA8: dout  = 8'b00001111; //  168 :  15 - 0xf -- Sprite 0x15
      11'hA9: dout  = 8'b00001111; //  169 :  15 - 0xf
      11'hAA: dout  = 8'b00001111; //  170 :  15 - 0xf
      11'hAB: dout  = 8'b00011111; //  171 :  31 - 0x1f
      11'hAC: dout  = 8'b00011111; //  172 :  31 - 0x1f
      11'hAD: dout  = 8'b00011110; //  173 :  30 - 0x1e
      11'hAE: dout  = 8'b00011100; //  174 :  28 - 0x1c
      11'hAF: dout  = 8'b00011110; //  175 :  30 - 0x1e
      11'hB0: dout  = 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0x16
      11'hB1: dout  = 8'b01110000; //  177 : 112 - 0x70
      11'hB2: dout  = 8'b00000000; //  178 :   0 - 0x0
      11'hB3: dout  = 8'b11000000; //  179 : 192 - 0xc0
      11'hB4: dout  = 8'b10100000; //  180 : 160 - 0xa0
      11'hB5: dout  = 8'b11111000; //  181 : 248 - 0xf8
      11'hB6: dout  = 8'b10000000; //  182 : 128 - 0x80
      11'hB7: dout  = 8'b11000000; //  183 : 192 - 0xc0
      11'hB8: dout  = 8'b11100000; //  184 : 224 - 0xe0 -- Sprite 0x17
      11'hB9: dout  = 8'b01100000; //  185 :  96 - 0x60
      11'hBA: dout  = 8'b11110000; //  186 : 240 - 0xf0
      11'hBB: dout  = 8'b11110000; //  187 : 240 - 0xf0
      11'hBC: dout  = 8'b11110000; //  188 : 240 - 0xf0
      11'hBD: dout  = 8'b11100000; //  189 : 224 - 0xe0
      11'hBE: dout  = 8'b11100000; //  190 : 224 - 0xe0
      11'hBF: dout  = 8'b11110000; //  191 : 240 - 0xf0
      11'hC0: dout  = 8'b00000111; //  192 :   7 - 0x7 -- Sprite 0x18
      11'hC1: dout  = 8'b00001111; //  193 :  15 - 0xf
      11'hC2: dout  = 8'b00001111; //  194 :  15 - 0xf
      11'hC3: dout  = 8'b00010010; //  195 :  18 - 0x12
      11'hC4: dout  = 8'b00010011; //  196 :  19 - 0x13
      11'hC5: dout  = 8'b00111000; //  197 :  56 - 0x38
      11'hC6: dout  = 8'b00000000; //  198 :   0 - 0x0
      11'hC7: dout  = 8'b00001111; //  199 :  15 - 0xf
      11'hC8: dout  = 8'b00011111; //  200 :  31 - 0x1f -- Sprite 0x19
      11'hC9: dout  = 8'b00011111; //  201 :  31 - 0x1f
      11'hCA: dout  = 8'b00011111; //  202 :  31 - 0x1f
      11'hCB: dout  = 8'b00011111; //  203 :  31 - 0x1f
      11'hCC: dout  = 8'b00011111; //  204 :  31 - 0x1f
      11'hCD: dout  = 8'b00011110; //  205 :  30 - 0x1e
      11'hCE: dout  = 8'b00011100; //  206 :  28 - 0x1c
      11'hCF: dout  = 8'b00011110; //  207 :  30 - 0x1e
      11'hD0: dout  = 8'b10000000; //  208 : 128 - 0x80 -- Sprite 0x1a
      11'hD1: dout  = 8'b11110000; //  209 : 240 - 0xf0
      11'hD2: dout  = 8'b00000000; //  210 :   0 - 0x0
      11'hD3: dout  = 8'b01000000; //  211 :  64 - 0x40
      11'hD4: dout  = 8'b00100000; //  212 :  32 - 0x20
      11'hD5: dout  = 8'b01111000; //  213 : 120 - 0x78
      11'hD6: dout  = 8'b00000000; //  214 :   0 - 0x0
      11'hD7: dout  = 8'b11000000; //  215 : 192 - 0xc0
      11'hD8: dout  = 8'b11111000; //  216 : 248 - 0xf8 -- Sprite 0x1b
      11'hD9: dout  = 8'b11111000; //  217 : 248 - 0xf8
      11'hDA: dout  = 8'b11110000; //  218 : 240 - 0xf0
      11'hDB: dout  = 8'b11110000; //  219 : 240 - 0xf0
      11'hDC: dout  = 8'b11110000; //  220 : 240 - 0xf0
      11'hDD: dout  = 8'b11100000; //  221 : 224 - 0xe0
      11'hDE: dout  = 8'b11100000; //  222 : 224 - 0xe0
      11'hDF: dout  = 8'b11110000; //  223 : 240 - 0xf0
      11'hE0: dout  = 8'b00000100; //  224 :   4 - 0x4 -- Sprite 0x1c
      11'hE1: dout  = 8'b00001100; //  225 :  12 - 0xc
      11'hE2: dout  = 8'b00001100; //  226 :  12 - 0xc
      11'hE3: dout  = 8'b00010011; //  227 :  19 - 0x13
      11'hE4: dout  = 8'b00010011; //  228 :  19 - 0x13
      11'hE5: dout  = 8'b00111111; //  229 :  63 - 0x3f
      11'hE6: dout  = 8'b00000111; //  230 :   7 - 0x7
      11'hE7: dout  = 8'b00001111; //  231 :  15 - 0xf
      11'hE8: dout  = 8'b00001111; //  232 :  15 - 0xf -- Sprite 0x1d
      11'hE9: dout  = 8'b00001111; //  233 :  15 - 0xf
      11'hEA: dout  = 8'b00001111; //  234 :  15 - 0xf
      11'hEB: dout  = 8'b00011111; //  235 :  31 - 0x1f
      11'hEC: dout  = 8'b00111111; //  236 :  63 - 0x3f
      11'hED: dout  = 8'b01111100; //  237 : 124 - 0x7c
      11'hEE: dout  = 8'b01110000; //  238 : 112 - 0x70
      11'hEF: dout  = 8'b00111000; //  239 :  56 - 0x38
      11'hF0: dout  = 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0x1e
      11'hF1: dout  = 8'b01110000; //  241 : 112 - 0x70
      11'hF2: dout  = 8'b00000000; //  242 :   0 - 0x0
      11'hF3: dout  = 8'b11000000; //  243 : 192 - 0xc0
      11'hF4: dout  = 8'b10100000; //  244 : 160 - 0xa0
      11'hF5: dout  = 8'b11111000; //  245 : 248 - 0xf8
      11'hF6: dout  = 8'b10000000; //  246 : 128 - 0x80
      11'hF7: dout  = 8'b11000000; //  247 : 192 - 0xc0
      11'hF8: dout  = 8'b11000000; //  248 : 192 - 0xc0 -- Sprite 0x1f
      11'hF9: dout  = 8'b01100000; //  249 :  96 - 0x60
      11'hFA: dout  = 8'b11100100; //  250 : 228 - 0xe4
      11'hFB: dout  = 8'b11111100; //  251 : 252 - 0xfc
      11'hFC: dout  = 8'b11111100; //  252 : 252 - 0xfc
      11'hFD: dout  = 8'b01111100; //  253 : 124 - 0x7c
      11'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      11'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout  = 8'b00000111; //  256 :   7 - 0x7 -- Sprite 0x20
      11'h101: dout  = 8'b00001111; //  257 :  15 - 0xf
      11'h102: dout  = 8'b00001111; //  258 :  15 - 0xf
      11'h103: dout  = 8'b00010010; //  259 :  18 - 0x12
      11'h104: dout  = 8'b00010011; //  260 :  19 - 0x13
      11'h105: dout  = 8'b00111000; //  261 :  56 - 0x38
      11'h106: dout  = 8'b00000000; //  262 :   0 - 0x0
      11'h107: dout  = 8'b00000111; //  263 :   7 - 0x7
      11'h108: dout  = 8'b00001111; //  264 :  15 - 0xf -- Sprite 0x21
      11'h109: dout  = 8'b00001111; //  265 :  15 - 0xf
      11'h10A: dout  = 8'b00001111; //  266 :  15 - 0xf
      11'h10B: dout  = 8'b00011111; //  267 :  31 - 0x1f
      11'h10C: dout  = 8'b00111111; //  268 :  63 - 0x3f
      11'h10D: dout  = 8'b01111100; //  269 : 124 - 0x7c
      11'h10E: dout  = 8'b01110000; //  270 : 112 - 0x70
      11'h10F: dout  = 8'b00111000; //  271 :  56 - 0x38
      11'h110: dout  = 8'b10000000; //  272 : 128 - 0x80 -- Sprite 0x22
      11'h111: dout  = 8'b11110000; //  273 : 240 - 0xf0
      11'h112: dout  = 8'b00000000; //  274 :   0 - 0x0
      11'h113: dout  = 8'b01000000; //  275 :  64 - 0x40
      11'h114: dout  = 8'b00100000; //  276 :  32 - 0x20
      11'h115: dout  = 8'b01111000; //  277 : 120 - 0x78
      11'h116: dout  = 8'b00000000; //  278 :   0 - 0x0
      11'h117: dout  = 8'b11000000; //  279 : 192 - 0xc0
      11'h118: dout  = 8'b11111000; //  280 : 248 - 0xf8 -- Sprite 0x23
      11'h119: dout  = 8'b11111000; //  281 : 248 - 0xf8
      11'h11A: dout  = 8'b11100000; //  282 : 224 - 0xe0
      11'h11B: dout  = 8'b11111100; //  283 : 252 - 0xfc
      11'h11C: dout  = 8'b11111100; //  284 : 252 - 0xfc
      11'h11D: dout  = 8'b01111100; //  285 : 124 - 0x7c
      11'h11E: dout  = 8'b00000000; //  286 :   0 - 0x0
      11'h11F: dout  = 8'b00000000; //  287 :   0 - 0x0
      11'h120: dout  = 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x24
      11'h121: dout  = 8'b00000111; //  289 :   7 - 0x7
      11'h122: dout  = 8'b00000111; //  290 :   7 - 0x7
      11'h123: dout  = 8'b00001111; //  291 :  15 - 0xf
      11'h124: dout  = 8'b00001111; //  292 :  15 - 0xf
      11'h125: dout  = 8'b00111000; //  293 :  56 - 0x38
      11'h126: dout  = 8'b01111111; //  294 : 127 - 0x7f
      11'h127: dout  = 8'b01111111; //  295 : 127 - 0x7f
      11'h128: dout  = 8'b00011111; //  296 :  31 - 0x1f -- Sprite 0x25
      11'h129: dout  = 8'b00011111; //  297 :  31 - 0x1f
      11'h12A: dout  = 8'b00011111; //  298 :  31 - 0x1f
      11'h12B: dout  = 8'b00011111; //  299 :  31 - 0x1f
      11'h12C: dout  = 8'b00001111; //  300 :  15 - 0xf
      11'h12D: dout  = 8'b00001111; //  301 :  15 - 0xf
      11'h12E: dout  = 8'b00001111; //  302 :  15 - 0xf
      11'h12F: dout  = 8'b00000111; //  303 :   7 - 0x7
      11'h130: dout  = 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      11'h131: dout  = 8'b11100000; //  305 : 224 - 0xe0
      11'h132: dout  = 8'b11111000; //  306 : 248 - 0xf8
      11'h133: dout  = 8'b11111100; //  307 : 252 - 0xfc
      11'h134: dout  = 8'b11111100; //  308 : 252 - 0xfc
      11'h135: dout  = 8'b00011100; //  309 :  28 - 0x1c
      11'h136: dout  = 8'b11111000; //  310 : 248 - 0xf8
      11'h137: dout  = 8'b11111000; //  311 : 248 - 0xf8
      11'h138: dout  = 8'b11111000; //  312 : 248 - 0xf8 -- Sprite 0x27
      11'h139: dout  = 8'b11111100; //  313 : 252 - 0xfc
      11'h13A: dout  = 8'b11111100; //  314 : 252 - 0xfc
      11'h13B: dout  = 8'b11111000; //  315 : 248 - 0xf8
      11'h13C: dout  = 8'b01111000; //  316 : 120 - 0x78
      11'h13D: dout  = 8'b10000000; //  317 : 128 - 0x80
      11'h13E: dout  = 8'b11000000; //  318 : 192 - 0xc0
      11'h13F: dout  = 8'b11000000; //  319 : 192 - 0xc0
      11'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      11'h141: dout  = 8'b00000011; //  321 :   3 - 0x3
      11'h142: dout  = 8'b00000111; //  322 :   7 - 0x7
      11'h143: dout  = 8'b00000111; //  323 :   7 - 0x7
      11'h144: dout  = 8'b00001001; //  324 :   9 - 0x9
      11'h145: dout  = 8'b00001001; //  325 :   9 - 0x9
      11'h146: dout  = 8'b00011100; //  326 :  28 - 0x1c
      11'h147: dout  = 8'b00000000; //  327 :   0 - 0x0
      11'h148: dout  = 8'b00011111; //  328 :  31 - 0x1f -- Sprite 0x29
      11'h149: dout  = 8'b00001111; //  329 :  15 - 0xf
      11'h14A: dout  = 8'b00000111; //  330 :   7 - 0x7
      11'h14B: dout  = 8'b00110111; //  331 :  55 - 0x37
      11'h14C: dout  = 8'b01111111; //  332 : 127 - 0x7f
      11'h14D: dout  = 8'b11011111; //  333 : 223 - 0xdf
      11'h14E: dout  = 8'b00001111; //  334 :  15 - 0xf
      11'h14F: dout  = 8'b00000110; //  335 :   6 - 0x6
      11'h150: dout  = 8'b00000000; //  336 :   0 - 0x0 -- Sprite 0x2a
      11'h151: dout  = 8'b11000000; //  337 : 192 - 0xc0
      11'h152: dout  = 8'b11111000; //  338 : 248 - 0xf8
      11'h153: dout  = 8'b10000000; //  339 : 128 - 0x80
      11'h154: dout  = 8'b00100000; //  340 :  32 - 0x20
      11'h155: dout  = 8'b10010000; //  341 : 144 - 0x90
      11'h156: dout  = 8'b00111100; //  342 :  60 - 0x3c
      11'h157: dout  = 8'b00000000; //  343 :   0 - 0x0
      11'h158: dout  = 8'b11100100; //  344 : 228 - 0xe4 -- Sprite 0x2b
      11'h159: dout  = 8'b11111110; //  345 : 254 - 0xfe
      11'h15A: dout  = 8'b01110000; //  346 : 112 - 0x70
      11'h15B: dout  = 8'b11110001; //  347 : 241 - 0xf1
      11'h15C: dout  = 8'b11111111; //  348 : 255 - 0xff
      11'h15D: dout  = 8'b11111111; //  349 : 255 - 0xff
      11'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      11'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      11'h160: dout  = 8'b00000111; //  352 :   7 - 0x7 -- Sprite 0x2c
      11'h161: dout  = 8'b00001111; //  353 :  15 - 0xf
      11'h162: dout  = 8'b00001111; //  354 :  15 - 0xf
      11'h163: dout  = 8'b00010010; //  355 :  18 - 0x12
      11'h164: dout  = 8'b00010011; //  356 :  19 - 0x13
      11'h165: dout  = 8'b00111000; //  357 :  56 - 0x38
      11'h166: dout  = 8'b01110000; //  358 : 112 - 0x70
      11'h167: dout  = 8'b11111111; //  359 : 255 - 0xff
      11'h168: dout  = 8'b11011111; //  360 : 223 - 0xdf -- Sprite 0x2d
      11'h169: dout  = 8'b00011110; //  361 :  30 - 0x1e
      11'h16A: dout  = 8'b00011111; //  362 :  31 - 0x1f
      11'h16B: dout  = 8'b00011111; //  363 :  31 - 0x1f
      11'h16C: dout  = 8'b00011111; //  364 :  31 - 0x1f
      11'h16D: dout  = 8'b00001111; //  365 :  15 - 0xf
      11'h16E: dout  = 8'b00000111; //  366 :   7 - 0x7
      11'h16F: dout  = 8'b00000001; //  367 :   1 - 0x1
      11'h170: dout  = 8'b10000000; //  368 : 128 - 0x80 -- Sprite 0x2e
      11'h171: dout  = 8'b11110000; //  369 : 240 - 0xf0
      11'h172: dout  = 8'b00000000; //  370 :   0 - 0x0
      11'h173: dout  = 8'b01000000; //  371 :  64 - 0x40
      11'h174: dout  = 8'b00100000; //  372 :  32 - 0x20
      11'h175: dout  = 8'b01111000; //  373 : 120 - 0x78
      11'h176: dout  = 8'b00000000; //  374 :   0 - 0x0
      11'h177: dout  = 8'b11111100; //  375 : 252 - 0xfc
      11'h178: dout  = 8'b11110000; //  376 : 240 - 0xf0 -- Sprite 0x2f
      11'h179: dout  = 8'b11100000; //  377 : 224 - 0xe0
      11'h17A: dout  = 8'b11100000; //  378 : 224 - 0xe0
      11'h17B: dout  = 8'b11110000; //  379 : 240 - 0xf0
      11'h17C: dout  = 8'b11111010; //  380 : 250 - 0xfa
      11'h17D: dout  = 8'b11111110; //  381 : 254 - 0xfe
      11'h17E: dout  = 8'b11111100; //  382 : 252 - 0xfc
      11'h17F: dout  = 8'b11011000; //  383 : 216 - 0xd8
      11'h180: dout  = 8'b00000000; //  384 :   0 - 0x0 -- Sprite 0x30
      11'h181: dout  = 8'b00000000; //  385 :   0 - 0x0
      11'h182: dout  = 8'b00000111; //  386 :   7 - 0x7
      11'h183: dout  = 8'b00001000; //  387 :   8 - 0x8
      11'h184: dout  = 8'b00010000; //  388 :  16 - 0x10
      11'h185: dout  = 8'b00100000; //  389 :  32 - 0x20
      11'h186: dout  = 8'b01000000; //  390 :  64 - 0x40
      11'h187: dout  = 8'b01000000; //  391 :  64 - 0x40
      11'h188: dout  = 8'b01000000; //  392 :  64 - 0x40 -- Sprite 0x31
      11'h189: dout  = 8'b01000000; //  393 :  64 - 0x40
      11'h18A: dout  = 8'b00100000; //  394 :  32 - 0x20
      11'h18B: dout  = 8'b00010000; //  395 :  16 - 0x10
      11'h18C: dout  = 8'b00001000; //  396 :   8 - 0x8
      11'h18D: dout  = 8'b00000111; //  397 :   7 - 0x7
      11'h18E: dout  = 8'b00000000; //  398 :   0 - 0x0
      11'h18F: dout  = 8'b00000000; //  399 :   0 - 0x0
      11'h190: dout  = 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      11'h191: dout  = 8'b00000000; //  401 :   0 - 0x0
      11'h192: dout  = 8'b11100000; //  402 : 224 - 0xe0
      11'h193: dout  = 8'b00010000; //  403 :  16 - 0x10
      11'h194: dout  = 8'b00001000; //  404 :   8 - 0x8
      11'h195: dout  = 8'b00000100; //  405 :   4 - 0x4
      11'h196: dout  = 8'b00000010; //  406 :   2 - 0x2
      11'h197: dout  = 8'b00000010; //  407 :   2 - 0x2
      11'h198: dout  = 8'b00000010; //  408 :   2 - 0x2 -- Sprite 0x33
      11'h199: dout  = 8'b00000010; //  409 :   2 - 0x2
      11'h19A: dout  = 8'b00000100; //  410 :   4 - 0x4
      11'h19B: dout  = 8'b00001000; //  411 :   8 - 0x8
      11'h19C: dout  = 8'b00010000; //  412 :  16 - 0x10
      11'h19D: dout  = 8'b11100000; //  413 : 224 - 0xe0
      11'h19E: dout  = 8'b00000000; //  414 :   0 - 0x0
      11'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      11'h1A0: dout  = 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x34
      11'h1A1: dout  = 8'b00000000; //  417 :   0 - 0x0
      11'h1A2: dout  = 8'b00000000; //  418 :   0 - 0x0
      11'h1A3: dout  = 8'b00000000; //  419 :   0 - 0x0
      11'h1A4: dout  = 8'b00000011; //  420 :   3 - 0x3
      11'h1A5: dout  = 8'b00000100; //  421 :   4 - 0x4
      11'h1A6: dout  = 8'b00001000; //  422 :   8 - 0x8
      11'h1A7: dout  = 8'b00010000; //  423 :  16 - 0x10
      11'h1A8: dout  = 8'b00010000; //  424 :  16 - 0x10 -- Sprite 0x35
      11'h1A9: dout  = 8'b00001000; //  425 :   8 - 0x8
      11'h1AA: dout  = 8'b00000100; //  426 :   4 - 0x4
      11'h1AB: dout  = 8'b00000011; //  427 :   3 - 0x3
      11'h1AC: dout  = 8'b00000000; //  428 :   0 - 0x0
      11'h1AD: dout  = 8'b00000000; //  429 :   0 - 0x0
      11'h1AE: dout  = 8'b00000000; //  430 :   0 - 0x0
      11'h1AF: dout  = 8'b00000000; //  431 :   0 - 0x0
      11'h1B0: dout  = 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x36
      11'h1B1: dout  = 8'b00000000; //  433 :   0 - 0x0
      11'h1B2: dout  = 8'b00000000; //  434 :   0 - 0x0
      11'h1B3: dout  = 8'b00000000; //  435 :   0 - 0x0
      11'h1B4: dout  = 8'b11000000; //  436 : 192 - 0xc0
      11'h1B5: dout  = 8'b00100000; //  437 :  32 - 0x20
      11'h1B6: dout  = 8'b00010000; //  438 :  16 - 0x10
      11'h1B7: dout  = 8'b00001000; //  439 :   8 - 0x8
      11'h1B8: dout  = 8'b00001000; //  440 :   8 - 0x8 -- Sprite 0x37
      11'h1B9: dout  = 8'b00010000; //  441 :  16 - 0x10
      11'h1BA: dout  = 8'b00100000; //  442 :  32 - 0x20
      11'h1BB: dout  = 8'b11000000; //  443 : 192 - 0xc0
      11'h1BC: dout  = 8'b00000000; //  444 :   0 - 0x0
      11'h1BD: dout  = 8'b00000000; //  445 :   0 - 0x0
      11'h1BE: dout  = 8'b00000000; //  446 :   0 - 0x0
      11'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      11'h1C0: dout  = 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      11'h1C1: dout  = 8'b00000000; //  449 :   0 - 0x0
      11'h1C2: dout  = 8'b00000000; //  450 :   0 - 0x0
      11'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      11'h1C4: dout  = 8'b00000000; //  452 :   0 - 0x0
      11'h1C5: dout  = 8'b00000000; //  453 :   0 - 0x0
      11'h1C6: dout  = 8'b00000000; //  454 :   0 - 0x0
      11'h1C7: dout  = 8'b00000001; //  455 :   1 - 0x1
      11'h1C8: dout  = 8'b00000010; //  456 :   2 - 0x2 -- Sprite 0x39
      11'h1C9: dout  = 8'b00000001; //  457 :   1 - 0x1
      11'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      11'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      11'h1CC: dout  = 8'b00000000; //  460 :   0 - 0x0
      11'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      11'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      11'h1D2: dout  = 8'b00000000; //  466 :   0 - 0x0
      11'h1D3: dout  = 8'b00000000; //  467 :   0 - 0x0
      11'h1D4: dout  = 8'b00000000; //  468 :   0 - 0x0
      11'h1D5: dout  = 8'b00000000; //  469 :   0 - 0x0
      11'h1D6: dout  = 8'b00000000; //  470 :   0 - 0x0
      11'h1D7: dout  = 8'b00000000; //  471 :   0 - 0x0
      11'h1D8: dout  = 8'b10000000; //  472 : 128 - 0x80 -- Sprite 0x3b
      11'h1D9: dout  = 8'b00000000; //  473 :   0 - 0x0
      11'h1DA: dout  = 8'b00000000; //  474 :   0 - 0x0
      11'h1DB: dout  = 8'b00000000; //  475 :   0 - 0x0
      11'h1DC: dout  = 8'b00000000; //  476 :   0 - 0x0
      11'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      11'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      11'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      11'h1E1: dout  = 8'b00000000; //  481 :   0 - 0x0
      11'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      11'h1E3: dout  = 8'b00000001; //  483 :   1 - 0x1
      11'h1E4: dout  = 8'b00100001; //  484 :  33 - 0x21
      11'h1E5: dout  = 8'b00010000; //  485 :  16 - 0x10
      11'h1E6: dout  = 8'b00000000; //  486 :   0 - 0x0
      11'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout  = 8'b01100000; //  488 :  96 - 0x60 -- Sprite 0x3d
      11'h1E9: dout  = 8'b00000000; //  489 :   0 - 0x0
      11'h1EA: dout  = 8'b00000000; //  490 :   0 - 0x0
      11'h1EB: dout  = 8'b00010000; //  491 :  16 - 0x10
      11'h1EC: dout  = 8'b00100001; //  492 :  33 - 0x21
      11'h1ED: dout  = 8'b00000001; //  493 :   1 - 0x1
      11'h1EE: dout  = 8'b00000000; //  494 :   0 - 0x0
      11'h1EF: dout  = 8'b00000000; //  495 :   0 - 0x0
      11'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      11'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      11'h1F2: dout  = 8'b00000000; //  498 :   0 - 0x0
      11'h1F3: dout  = 8'b00000000; //  499 :   0 - 0x0
      11'h1F4: dout  = 8'b00001000; //  500 :   8 - 0x8
      11'h1F5: dout  = 8'b00010000; //  501 :  16 - 0x10
      11'h1F6: dout  = 8'b00000000; //  502 :   0 - 0x0
      11'h1F7: dout  = 8'b00000000; //  503 :   0 - 0x0
      11'h1F8: dout  = 8'b00001100; //  504 :  12 - 0xc -- Sprite 0x3f
      11'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      11'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      11'h1FB: dout  = 8'b00010000; //  507 :  16 - 0x10
      11'h1FC: dout  = 8'b00001000; //  508 :   8 - 0x8
      11'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      11'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      11'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      11'h200: dout  = 8'b00000100; //  512 :   4 - 0x4 -- Sprite 0x40
      11'h201: dout  = 8'b00000010; //  513 :   2 - 0x2
      11'h202: dout  = 8'b00000001; //  514 :   1 - 0x1
      11'h203: dout  = 8'b00000000; //  515 :   0 - 0x0
      11'h204: dout  = 8'b00000000; //  516 :   0 - 0x0
      11'h205: dout  = 8'b00000000; //  517 :   0 - 0x0
      11'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      11'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      11'h208: dout  = 8'b00000000; //  520 :   0 - 0x0 -- Sprite 0x41
      11'h209: dout  = 8'b00000000; //  521 :   0 - 0x0
      11'h20A: dout  = 8'b00000000; //  522 :   0 - 0x0
      11'h20B: dout  = 8'b00000000; //  523 :   0 - 0x0
      11'h20C: dout  = 8'b00000000; //  524 :   0 - 0x0
      11'h20D: dout  = 8'b00000000; //  525 :   0 - 0x0
      11'h20E: dout  = 8'b00000001; //  526 :   1 - 0x1
      11'h20F: dout  = 8'b00000011; //  527 :   3 - 0x3
      11'h210: dout  = 8'b00000111; //  528 :   7 - 0x7 -- Sprite 0x42
      11'h211: dout  = 8'b00000111; //  529 :   7 - 0x7
      11'h212: dout  = 8'b00000111; //  530 :   7 - 0x7
      11'h213: dout  = 8'b00000011; //  531 :   3 - 0x3
      11'h214: dout  = 8'b00000001; //  532 :   1 - 0x1
      11'h215: dout  = 8'b00000000; //  533 :   0 - 0x0
      11'h216: dout  = 8'b00000000; //  534 :   0 - 0x0
      11'h217: dout  = 8'b00000000; //  535 :   0 - 0x0
      11'h218: dout  = 8'b00000000; //  536 :   0 - 0x0 -- Sprite 0x43
      11'h219: dout  = 8'b00000000; //  537 :   0 - 0x0
      11'h21A: dout  = 8'b00000000; //  538 :   0 - 0x0
      11'h21B: dout  = 8'b00000000; //  539 :   0 - 0x0
      11'h21C: dout  = 8'b00000000; //  540 :   0 - 0x0
      11'h21D: dout  = 8'b00000000; //  541 :   0 - 0x0
      11'h21E: dout  = 8'b00000000; //  542 :   0 - 0x0
      11'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      11'h220: dout  = 8'b00000000; //  544 :   0 - 0x0 -- Sprite 0x44
      11'h221: dout  = 8'b01000010; //  545 :  66 - 0x42
      11'h222: dout  = 8'b00111001; //  546 :  57 - 0x39
      11'h223: dout  = 8'b11111111; //  547 : 255 - 0xff
      11'h224: dout  = 8'b11111111; //  548 : 255 - 0xff
      11'h225: dout  = 8'b11111111; //  549 : 255 - 0xff
      11'h226: dout  = 8'b11111111; //  550 : 255 - 0xff
      11'h227: dout  = 8'b11111111; //  551 : 255 - 0xff
      11'h228: dout  = 8'b01111111; //  552 : 127 - 0x7f -- Sprite 0x45
      11'h229: dout  = 8'b00111111; //  553 :  63 - 0x3f
      11'h22A: dout  = 8'b00011111; //  554 :  31 - 0x1f
      11'h22B: dout  = 8'b00001111; //  555 :  15 - 0xf
      11'h22C: dout  = 8'b00011111; //  556 :  31 - 0x1f
      11'h22D: dout  = 8'b11111111; //  557 : 255 - 0xff
      11'h22E: dout  = 8'b11111111; //  558 : 255 - 0xff
      11'h22F: dout  = 8'b11111111; //  559 : 255 - 0xff
      11'h230: dout  = 8'b11111000; //  560 : 248 - 0xf8 -- Sprite 0x46
      11'h231: dout  = 8'b11110111; //  561 : 247 - 0xf7
      11'h232: dout  = 8'b11101111; //  562 : 239 - 0xef
      11'h233: dout  = 8'b11111111; //  563 : 255 - 0xff
      11'h234: dout  = 8'b11111111; //  564 : 255 - 0xff
      11'h235: dout  = 8'b11111110; //  565 : 254 - 0xfe
      11'h236: dout  = 8'b01111110; //  566 : 126 - 0x7e
      11'h237: dout  = 8'b00111110; //  567 :  62 - 0x3e
      11'h238: dout  = 8'b00000111; //  568 :   7 - 0x7 -- Sprite 0x47
      11'h239: dout  = 8'b00000000; //  569 :   0 - 0x0
      11'h23A: dout  = 8'b00000000; //  570 :   0 - 0x0
      11'h23B: dout  = 8'b00000000; //  571 :   0 - 0x0
      11'h23C: dout  = 8'b00000000; //  572 :   0 - 0x0
      11'h23D: dout  = 8'b00000000; //  573 :   0 - 0x0
      11'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      11'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout  = 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x48
      11'h241: dout  = 8'b00000000; //  577 :   0 - 0x0
      11'h242: dout  = 8'b00000000; //  578 :   0 - 0x0
      11'h243: dout  = 8'b11000000; //  579 : 192 - 0xc0
      11'h244: dout  = 8'b11100000; //  580 : 224 - 0xe0
      11'h245: dout  = 8'b11110000; //  581 : 240 - 0xf0
      11'h246: dout  = 8'b11011011; //  582 : 219 - 0xdb
      11'h247: dout  = 8'b11110110; //  583 : 246 - 0xf6
      11'h248: dout  = 8'b11001011; //  584 : 203 - 0xcb -- Sprite 0x49
      11'h249: dout  = 8'b11100000; //  585 : 224 - 0xe0
      11'h24A: dout  = 8'b11000100; //  586 : 196 - 0xc4
      11'h24B: dout  = 8'b00000010; //  587 :   2 - 0x2
      11'h24C: dout  = 8'b11010001; //  588 : 209 - 0xd1
      11'h24D: dout  = 8'b11100001; //  589 : 225 - 0xe1
      11'h24E: dout  = 8'b11010001; //  590 : 209 - 0xd1
      11'h24F: dout  = 8'b10000011; //  591 : 131 - 0x83
      11'h250: dout  = 8'b00001111; //  592 :  15 - 0xf -- Sprite 0x4a
      11'h251: dout  = 8'b11111111; //  593 : 255 - 0xff
      11'h252: dout  = 8'b11100000; //  594 : 224 - 0xe0
      11'h253: dout  = 8'b10001111; //  595 : 143 - 0x8f
      11'h254: dout  = 8'b01101110; //  596 : 110 - 0x6e
      11'h255: dout  = 8'b01000100; //  597 :  68 - 0x44
      11'h256: dout  = 8'b11101110; //  598 : 238 - 0xee
      11'h257: dout  = 8'b01100000; //  599 :  96 - 0x60
      11'h258: dout  = 8'b10000011; //  600 : 131 - 0x83 -- Sprite 0x4b
      11'h259: dout  = 8'b11100000; //  601 : 224 - 0xe0
      11'h25A: dout  = 8'b11100100; //  602 : 228 - 0xe4
      11'h25B: dout  = 8'b11000110; //  603 : 198 - 0xc6
      11'h25C: dout  = 8'b01100001; //  604 :  97 - 0x61
      11'h25D: dout  = 8'b00110011; //  605 :  51 - 0x33
      11'h25E: dout  = 8'b00011111; //  606 :  31 - 0x1f
      11'h25F: dout  = 8'b00001111; //  607 :  15 - 0xf
      11'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x4c
      11'h261: dout  = 8'b00000000; //  609 :   0 - 0x0
      11'h262: dout  = 8'b00000000; //  610 :   0 - 0x0
      11'h263: dout  = 8'b00000011; //  611 :   3 - 0x3
      11'h264: dout  = 8'b00000111; //  612 :   7 - 0x7
      11'h265: dout  = 8'b00001111; //  613 :  15 - 0xf
      11'h266: dout  = 8'b01011011; //  614 :  91 - 0x5b
      11'h267: dout  = 8'b10100111; //  615 : 167 - 0xa7
      11'h268: dout  = 8'b01110011; //  616 : 115 - 0x73 -- Sprite 0x4d
      11'h269: dout  = 8'b00000111; //  617 :   7 - 0x7
      11'h26A: dout  = 8'b00100111; //  618 :  39 - 0x27
      11'h26B: dout  = 8'b01000000; //  619 :  64 - 0x40
      11'h26C: dout  = 8'b10001011; //  620 : 139 - 0x8b
      11'h26D: dout  = 8'b10000111; //  621 : 135 - 0x87
      11'h26E: dout  = 8'b10001011; //  622 : 139 - 0x8b
      11'h26F: dout  = 8'b11000001; //  623 : 193 - 0xc1
      11'h270: dout  = 8'b11110000; //  624 : 240 - 0xf0 -- Sprite 0x4e
      11'h271: dout  = 8'b11111111; //  625 : 255 - 0xff
      11'h272: dout  = 8'b00001111; //  626 :  15 - 0xf
      11'h273: dout  = 8'b11100001; //  627 : 225 - 0xe1
      11'h274: dout  = 8'b11101100; //  628 : 236 - 0xec
      11'h275: dout  = 8'b01000100; //  629 :  68 - 0x44
      11'h276: dout  = 8'b11101110; //  630 : 238 - 0xee
      11'h277: dout  = 8'b00001100; //  631 :  12 - 0xc
      11'h278: dout  = 8'b10000000; //  632 : 128 - 0x80 -- Sprite 0x4f
      11'h279: dout  = 8'b00001110; //  633 :  14 - 0xe
      11'h27A: dout  = 8'b01001110; //  634 :  78 - 0x4e
      11'h27B: dout  = 8'b11000110; //  635 : 198 - 0xc6
      11'h27C: dout  = 8'b00001100; //  636 :  12 - 0xc
      11'h27D: dout  = 8'b10011000; //  637 : 152 - 0x98
      11'h27E: dout  = 8'b11110000; //  638 : 240 - 0xf0
      11'h27F: dout  = 8'b11100000; //  639 : 224 - 0xe0
      11'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x50
      11'h281: dout  = 8'b01000010; //  641 :  66 - 0x42
      11'h282: dout  = 8'b10011100; //  642 : 156 - 0x9c
      11'h283: dout  = 8'b11111111; //  643 : 255 - 0xff
      11'h284: dout  = 8'b11111111; //  644 : 255 - 0xff
      11'h285: dout  = 8'b11111111; //  645 : 255 - 0xff
      11'h286: dout  = 8'b11111111; //  646 : 255 - 0xff
      11'h287: dout  = 8'b11111111; //  647 : 255 - 0xff
      11'h288: dout  = 8'b11111110; //  648 : 254 - 0xfe -- Sprite 0x51
      11'h289: dout  = 8'b11111100; //  649 : 252 - 0xfc
      11'h28A: dout  = 8'b11111000; //  650 : 248 - 0xf8
      11'h28B: dout  = 8'b11110000; //  651 : 240 - 0xf0
      11'h28C: dout  = 8'b11111000; //  652 : 248 - 0xf8
      11'h28D: dout  = 8'b11111111; //  653 : 255 - 0xff
      11'h28E: dout  = 8'b11111111; //  654 : 255 - 0xff
      11'h28F: dout  = 8'b11111111; //  655 : 255 - 0xff
      11'h290: dout  = 8'b00011111; //  656 :  31 - 0x1f -- Sprite 0x52
      11'h291: dout  = 8'b11101111; //  657 : 239 - 0xef
      11'h292: dout  = 8'b11110111; //  658 : 247 - 0xf7
      11'h293: dout  = 8'b11111111; //  659 : 255 - 0xff
      11'h294: dout  = 8'b11111111; //  660 : 255 - 0xff
      11'h295: dout  = 8'b11111110; //  661 : 254 - 0xfe
      11'h296: dout  = 8'b01111100; //  662 : 124 - 0x7c
      11'h297: dout  = 8'b01110000; //  663 : 112 - 0x70
      11'h298: dout  = 8'b11100000; //  664 : 224 - 0xe0 -- Sprite 0x53
      11'h299: dout  = 8'b00000000; //  665 :   0 - 0x0
      11'h29A: dout  = 8'b00000000; //  666 :   0 - 0x0
      11'h29B: dout  = 8'b00000000; //  667 :   0 - 0x0
      11'h29C: dout  = 8'b00000000; //  668 :   0 - 0x0
      11'h29D: dout  = 8'b00000000; //  669 :   0 - 0x0
      11'h29E: dout  = 8'b00000000; //  670 :   0 - 0x0
      11'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      11'h2A0: dout  = 8'b00100000; //  672 :  32 - 0x20 -- Sprite 0x54
      11'h2A1: dout  = 8'b01000000; //  673 :  64 - 0x40
      11'h2A2: dout  = 8'b10000000; //  674 : 128 - 0x80
      11'h2A3: dout  = 8'b00000000; //  675 :   0 - 0x0
      11'h2A4: dout  = 8'b00000000; //  676 :   0 - 0x0
      11'h2A5: dout  = 8'b00000000; //  677 :   0 - 0x0
      11'h2A6: dout  = 8'b00000000; //  678 :   0 - 0x0
      11'h2A7: dout  = 8'b00000000; //  679 :   0 - 0x0
      11'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      11'h2A9: dout  = 8'b00000000; //  681 :   0 - 0x0
      11'h2AA: dout  = 8'b00000000; //  682 :   0 - 0x0
      11'h2AB: dout  = 8'b00000000; //  683 :   0 - 0x0
      11'h2AC: dout  = 8'b00000000; //  684 :   0 - 0x0
      11'h2AD: dout  = 8'b00000000; //  685 :   0 - 0x0
      11'h2AE: dout  = 8'b10000000; //  686 : 128 - 0x80
      11'h2AF: dout  = 8'b11000000; //  687 : 192 - 0xc0
      11'h2B0: dout  = 8'b11100000; //  688 : 224 - 0xe0 -- Sprite 0x56
      11'h2B1: dout  = 8'b11100000; //  689 : 224 - 0xe0
      11'h2B2: dout  = 8'b11100000; //  690 : 224 - 0xe0
      11'h2B3: dout  = 8'b11000000; //  691 : 192 - 0xc0
      11'h2B4: dout  = 8'b10000000; //  692 : 128 - 0x80
      11'h2B5: dout  = 8'b00000000; //  693 :   0 - 0x0
      11'h2B6: dout  = 8'b00000000; //  694 :   0 - 0x0
      11'h2B7: dout  = 8'b00000000; //  695 :   0 - 0x0
      11'h2B8: dout  = 8'b00000000; //  696 :   0 - 0x0 -- Sprite 0x57
      11'h2B9: dout  = 8'b00000000; //  697 :   0 - 0x0
      11'h2BA: dout  = 8'b00000000; //  698 :   0 - 0x0
      11'h2BB: dout  = 8'b00000000; //  699 :   0 - 0x0
      11'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      11'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      11'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      11'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      11'h2C0: dout  = 8'b11111111; //  704 : 255 - 0xff -- Sprite 0x58
      11'h2C1: dout  = 8'b11111111; //  705 : 255 - 0xff
      11'h2C2: dout  = 8'b11111111; //  706 : 255 - 0xff
      11'h2C3: dout  = 8'b11111111; //  707 : 255 - 0xff
      11'h2C4: dout  = 8'b11111111; //  708 : 255 - 0xff
      11'h2C5: dout  = 8'b11111111; //  709 : 255 - 0xff
      11'h2C6: dout  = 8'b11111111; //  710 : 255 - 0xff
      11'h2C7: dout  = 8'b11111111; //  711 : 255 - 0xff
      11'h2C8: dout  = 8'b11111111; //  712 : 255 - 0xff -- Sprite 0x59
      11'h2C9: dout  = 8'b11111111; //  713 : 255 - 0xff
      11'h2CA: dout  = 8'b11111111; //  714 : 255 - 0xff
      11'h2CB: dout  = 8'b11111111; //  715 : 255 - 0xff
      11'h2CC: dout  = 8'b11111111; //  716 : 255 - 0xff
      11'h2CD: dout  = 8'b11111111; //  717 : 255 - 0xff
      11'h2CE: dout  = 8'b11111111; //  718 : 255 - 0xff
      11'h2CF: dout  = 8'b11111111; //  719 : 255 - 0xff
      11'h2D0: dout  = 8'b11111111; //  720 : 255 - 0xff -- Sprite 0x5a
      11'h2D1: dout  = 8'b11111111; //  721 : 255 - 0xff
      11'h2D2: dout  = 8'b11111111; //  722 : 255 - 0xff
      11'h2D3: dout  = 8'b11111111; //  723 : 255 - 0xff
      11'h2D4: dout  = 8'b11111111; //  724 : 255 - 0xff
      11'h2D5: dout  = 8'b11111111; //  725 : 255 - 0xff
      11'h2D6: dout  = 8'b11111111; //  726 : 255 - 0xff
      11'h2D7: dout  = 8'b11111111; //  727 : 255 - 0xff
      11'h2D8: dout  = 8'b11111111; //  728 : 255 - 0xff -- Sprite 0x5b
      11'h2D9: dout  = 8'b11111111; //  729 : 255 - 0xff
      11'h2DA: dout  = 8'b11111111; //  730 : 255 - 0xff
      11'h2DB: dout  = 8'b11111111; //  731 : 255 - 0xff
      11'h2DC: dout  = 8'b11111111; //  732 : 255 - 0xff
      11'h2DD: dout  = 8'b11111111; //  733 : 255 - 0xff
      11'h2DE: dout  = 8'b11111111; //  734 : 255 - 0xff
      11'h2DF: dout  = 8'b11111111; //  735 : 255 - 0xff
      11'h2E0: dout  = 8'b11111111; //  736 : 255 - 0xff -- Sprite 0x5c
      11'h2E1: dout  = 8'b11111111; //  737 : 255 - 0xff
      11'h2E2: dout  = 8'b11111111; //  738 : 255 - 0xff
      11'h2E3: dout  = 8'b11111111; //  739 : 255 - 0xff
      11'h2E4: dout  = 8'b11111111; //  740 : 255 - 0xff
      11'h2E5: dout  = 8'b11111111; //  741 : 255 - 0xff
      11'h2E6: dout  = 8'b11111111; //  742 : 255 - 0xff
      11'h2E7: dout  = 8'b11111111; //  743 : 255 - 0xff
      11'h2E8: dout  = 8'b11111111; //  744 : 255 - 0xff -- Sprite 0x5d
      11'h2E9: dout  = 8'b11111111; //  745 : 255 - 0xff
      11'h2EA: dout  = 8'b11111111; //  746 : 255 - 0xff
      11'h2EB: dout  = 8'b11111111; //  747 : 255 - 0xff
      11'h2EC: dout  = 8'b11111111; //  748 : 255 - 0xff
      11'h2ED: dout  = 8'b11111111; //  749 : 255 - 0xff
      11'h2EE: dout  = 8'b11111111; //  750 : 255 - 0xff
      11'h2EF: dout  = 8'b11111111; //  751 : 255 - 0xff
      11'h2F0: dout  = 8'b11111111; //  752 : 255 - 0xff -- Sprite 0x5e
      11'h2F1: dout  = 8'b11111111; //  753 : 255 - 0xff
      11'h2F2: dout  = 8'b11111111; //  754 : 255 - 0xff
      11'h2F3: dout  = 8'b11111111; //  755 : 255 - 0xff
      11'h2F4: dout  = 8'b11111111; //  756 : 255 - 0xff
      11'h2F5: dout  = 8'b11111111; //  757 : 255 - 0xff
      11'h2F6: dout  = 8'b11111111; //  758 : 255 - 0xff
      11'h2F7: dout  = 8'b11111111; //  759 : 255 - 0xff
      11'h2F8: dout  = 8'b11111111; //  760 : 255 - 0xff -- Sprite 0x5f
      11'h2F9: dout  = 8'b11111111; //  761 : 255 - 0xff
      11'h2FA: dout  = 8'b11111111; //  762 : 255 - 0xff
      11'h2FB: dout  = 8'b11111111; //  763 : 255 - 0xff
      11'h2FC: dout  = 8'b11111111; //  764 : 255 - 0xff
      11'h2FD: dout  = 8'b11111111; //  765 : 255 - 0xff
      11'h2FE: dout  = 8'b11111111; //  766 : 255 - 0xff
      11'h2FF: dout  = 8'b11111111; //  767 : 255 - 0xff
      11'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      11'h301: dout  = 8'b00000000; //  769 :   0 - 0x0
      11'h302: dout  = 8'b00011111; //  770 :  31 - 0x1f
      11'h303: dout  = 8'b00111111; //  771 :  63 - 0x3f
      11'h304: dout  = 8'b00111111; //  772 :  63 - 0x3f
      11'h305: dout  = 8'b01111111; //  773 : 127 - 0x7f
      11'h306: dout  = 8'b01111111; //  774 : 127 - 0x7f
      11'h307: dout  = 8'b01111111; //  775 : 127 - 0x7f
      11'h308: dout  = 8'b01111111; //  776 : 127 - 0x7f -- Sprite 0x61
      11'h309: dout  = 8'b00111110; //  777 :  62 - 0x3e
      11'h30A: dout  = 8'b00011111; //  778 :  31 - 0x1f
      11'h30B: dout  = 8'b00011111; //  779 :  31 - 0x1f
      11'h30C: dout  = 8'b00001111; //  780 :  15 - 0xf
      11'h30D: dout  = 8'b00001111; //  781 :  15 - 0xf
      11'h30E: dout  = 8'b00001111; //  782 :  15 - 0xf
      11'h30F: dout  = 8'b00000111; //  783 :   7 - 0x7
      11'h310: dout  = 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x62
      11'h311: dout  = 8'b01100000; //  785 :  96 - 0x60
      11'h312: dout  = 8'b11110000; //  786 : 240 - 0xf0
      11'h313: dout  = 8'b11111000; //  787 : 248 - 0xf8
      11'h314: dout  = 8'b11111000; //  788 : 248 - 0xf8
      11'h315: dout  = 8'b11111000; //  789 : 248 - 0xf8
      11'h316: dout  = 8'b11111100; //  790 : 252 - 0xfc
      11'h317: dout  = 8'b11111100; //  791 : 252 - 0xfc
      11'h318: dout  = 8'b11111000; //  792 : 248 - 0xf8 -- Sprite 0x63
      11'h319: dout  = 8'b11110000; //  793 : 240 - 0xf0
      11'h31A: dout  = 8'b11110000; //  794 : 240 - 0xf0
      11'h31B: dout  = 8'b11100000; //  795 : 224 - 0xe0
      11'h31C: dout  = 8'b10000000; //  796 : 128 - 0x80
      11'h31D: dout  = 8'b10000000; //  797 : 128 - 0x80
      11'h31E: dout  = 8'b11000000; //  798 : 192 - 0xc0
      11'h31F: dout  = 8'b11000000; //  799 : 192 - 0xc0
      11'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x64
      11'h321: dout  = 8'b00011111; //  801 :  31 - 0x1f
      11'h322: dout  = 8'b00111111; //  802 :  63 - 0x3f
      11'h323: dout  = 8'b01111111; //  803 : 127 - 0x7f
      11'h324: dout  = 8'b11111111; //  804 : 255 - 0xff
      11'h325: dout  = 8'b11111111; //  805 : 255 - 0xff
      11'h326: dout  = 8'b00111110; //  806 :  62 - 0x3e
      11'h327: dout  = 8'b00001111; //  807 :  15 - 0xf
      11'h328: dout  = 8'b00000000; //  808 :   0 - 0x0 -- Sprite 0x65
      11'h329: dout  = 8'b00000000; //  809 :   0 - 0x0
      11'h32A: dout  = 8'b00000000; //  810 :   0 - 0x0
      11'h32B: dout  = 8'b00000001; //  811 :   1 - 0x1
      11'h32C: dout  = 8'b00000000; //  812 :   0 - 0x0
      11'h32D: dout  = 8'b00000000; //  813 :   0 - 0x0
      11'h32E: dout  = 8'b00000000; //  814 :   0 - 0x0
      11'h32F: dout  = 8'b00000000; //  815 :   0 - 0x0
      11'h330: dout  = 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x66
      11'h331: dout  = 8'b11100000; //  817 : 224 - 0xe0
      11'h332: dout  = 8'b11110000; //  818 : 240 - 0xf0
      11'h333: dout  = 8'b11111100; //  819 : 252 - 0xfc
      11'h334: dout  = 8'b11111110; //  820 : 254 - 0xfe
      11'h335: dout  = 8'b11111110; //  821 : 254 - 0xfe
      11'h336: dout  = 8'b11111111; //  822 : 255 - 0xff
      11'h337: dout  = 8'b11111100; //  823 : 252 - 0xfc
      11'h338: dout  = 8'b01111100; //  824 : 124 - 0x7c -- Sprite 0x67
      11'h339: dout  = 8'b11111100; //  825 : 252 - 0xfc
      11'h33A: dout  = 8'b11111000; //  826 : 248 - 0xf8
      11'h33B: dout  = 8'b11110000; //  827 : 240 - 0xf0
      11'h33C: dout  = 8'b11100000; //  828 : 224 - 0xe0
      11'h33D: dout  = 8'b00000000; //  829 :   0 - 0x0
      11'h33E: dout  = 8'b00000000; //  830 :   0 - 0x0
      11'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      11'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      11'h341: dout  = 8'b00000111; //  833 :   7 - 0x7
      11'h342: dout  = 8'b00000111; //  834 :   7 - 0x7
      11'h343: dout  = 8'b00001111; //  835 :  15 - 0xf
      11'h344: dout  = 8'b00001111; //  836 :  15 - 0xf
      11'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      11'h346: dout  = 8'b00011111; //  838 :  31 - 0x1f
      11'h347: dout  = 8'b00111111; //  839 :  63 - 0x3f
      11'h348: dout  = 8'b01111111; //  840 : 127 - 0x7f -- Sprite 0x69
      11'h349: dout  = 8'b01111111; //  841 : 127 - 0x7f
      11'h34A: dout  = 8'b00011111; //  842 :  31 - 0x1f
      11'h34B: dout  = 8'b00011111; //  843 :  31 - 0x1f
      11'h34C: dout  = 8'b00011111; //  844 :  31 - 0x1f
      11'h34D: dout  = 8'b00011110; //  845 :  30 - 0x1e
      11'h34E: dout  = 8'b00001111; //  846 :  15 - 0xf
      11'h34F: dout  = 8'b00011111; //  847 :  31 - 0x1f
      11'h350: dout  = 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      11'h351: dout  = 8'b11100000; //  849 : 224 - 0xe0
      11'h352: dout  = 8'b11100000; //  850 : 224 - 0xe0
      11'h353: dout  = 8'b11110000; //  851 : 240 - 0xf0
      11'h354: dout  = 8'b11110000; //  852 : 240 - 0xf0
      11'h355: dout  = 8'b00000000; //  853 :   0 - 0x0
      11'h356: dout  = 8'b11111000; //  854 : 248 - 0xf8
      11'h357: dout  = 8'b11111100; //  855 : 252 - 0xfc
      11'h358: dout  = 8'b11111110; //  856 : 254 - 0xfe -- Sprite 0x6b
      11'h359: dout  = 8'b11111110; //  857 : 254 - 0xfe
      11'h35A: dout  = 8'b11111000; //  858 : 248 - 0xf8
      11'h35B: dout  = 8'b11111000; //  859 : 248 - 0xf8
      11'h35C: dout  = 8'b11111000; //  860 : 248 - 0xf8
      11'h35D: dout  = 8'b01111000; //  861 : 120 - 0x78
      11'h35E: dout  = 8'b11110000; //  862 : 240 - 0xf0
      11'h35F: dout  = 8'b11111000; //  863 : 248 - 0xf8
      11'h360: dout  = 8'b00000011; //  864 :   3 - 0x3 -- Sprite 0x6c
      11'h361: dout  = 8'b00000111; //  865 :   7 - 0x7
      11'h362: dout  = 8'b00000101; //  866 :   5 - 0x5
      11'h363: dout  = 8'b00001000; //  867 :   8 - 0x8
      11'h364: dout  = 8'b00011011; //  868 :  27 - 0x1b
      11'h365: dout  = 8'b00011001; //  869 :  25 - 0x19
      11'h366: dout  = 8'b00000101; //  870 :   5 - 0x5
      11'h367: dout  = 8'b00111111; //  871 :  63 - 0x3f
      11'h368: dout  = 8'b00111111; //  872 :  63 - 0x3f -- Sprite 0x6d
      11'h369: dout  = 8'b00001111; //  873 :  15 - 0xf
      11'h36A: dout  = 8'b00000101; //  874 :   5 - 0x5
      11'h36B: dout  = 8'b00110111; //  875 :  55 - 0x37
      11'h36C: dout  = 8'b00111111; //  876 :  63 - 0x3f
      11'h36D: dout  = 8'b00111111; //  877 :  63 - 0x3f
      11'h36E: dout  = 8'b00111110; //  878 :  62 - 0x3e
      11'h36F: dout  = 8'b00011100; //  879 :  28 - 0x1c
      11'h370: dout  = 8'b11100000; //  880 : 224 - 0xe0 -- Sprite 0x6e
      11'h371: dout  = 8'b11110000; //  881 : 240 - 0xf0
      11'h372: dout  = 8'b01010000; //  882 :  80 - 0x50
      11'h373: dout  = 8'b00001000; //  883 :   8 - 0x8
      11'h374: dout  = 8'b01101100; //  884 : 108 - 0x6c
      11'h375: dout  = 8'b11001100; //  885 : 204 - 0xcc
      11'h376: dout  = 8'b11010000; //  886 : 208 - 0xd0
      11'h377: dout  = 8'b11111110; //  887 : 254 - 0xfe
      11'h378: dout  = 8'b11111110; //  888 : 254 - 0xfe -- Sprite 0x6f
      11'h379: dout  = 8'b11111000; //  889 : 248 - 0xf8
      11'h37A: dout  = 8'b11010000; //  890 : 208 - 0xd0
      11'h37B: dout  = 8'b11111011; //  891 : 251 - 0xfb
      11'h37C: dout  = 8'b11111111; //  892 : 255 - 0xff
      11'h37D: dout  = 8'b11111111; //  893 : 255 - 0xff
      11'h37E: dout  = 8'b00111110; //  894 :  62 - 0x3e
      11'h37F: dout  = 8'b00001100; //  895 :  12 - 0xc
      11'h380: dout  = 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x70
      11'h381: dout  = 8'b00000000; //  897 :   0 - 0x0
      11'h382: dout  = 8'b01111001; //  898 : 121 - 0x79
      11'h383: dout  = 8'b11111001; //  899 : 249 - 0xf9
      11'h384: dout  = 8'b11110011; //  900 : 243 - 0xf3
      11'h385: dout  = 8'b11111111; //  901 : 255 - 0xff
      11'h386: dout  = 8'b01111011; //  902 : 123 - 0x7b
      11'h387: dout  = 8'b00111111; //  903 :  63 - 0x3f
      11'h388: dout  = 8'b00111111; //  904 :  63 - 0x3f -- Sprite 0x71
      11'h389: dout  = 8'b00111111; //  905 :  63 - 0x3f
      11'h38A: dout  = 8'b01111011; //  906 : 123 - 0x7b
      11'h38B: dout  = 8'b01111111; //  907 : 127 - 0x7f
      11'h38C: dout  = 8'b11111011; //  908 : 251 - 0xfb
      11'h38D: dout  = 8'b11110001; //  909 : 241 - 0xf1
      11'h38E: dout  = 8'b01111001; //  910 : 121 - 0x79
      11'h38F: dout  = 8'b00111000; //  911 :  56 - 0x38
      11'h390: dout  = 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x72
      11'h391: dout  = 8'b00000000; //  913 :   0 - 0x0
      11'h392: dout  = 8'b10000000; //  914 : 128 - 0x80
      11'h393: dout  = 8'b10110000; //  915 : 176 - 0xb0
      11'h394: dout  = 8'b10111000; //  916 : 184 - 0xb8
      11'h395: dout  = 8'b11000110; //  917 : 198 - 0xc6
      11'h396: dout  = 8'b10010011; //  918 : 147 - 0x93
      11'h397: dout  = 8'b11110111; //  919 : 247 - 0xf7
      11'h398: dout  = 8'b11100011; //  920 : 227 - 0xe3 -- Sprite 0x73
      11'h399: dout  = 8'b11110111; //  921 : 247 - 0xf7
      11'h39A: dout  = 8'b10010011; //  922 : 147 - 0x93
      11'h39B: dout  = 8'b11000110; //  923 : 198 - 0xc6
      11'h39C: dout  = 8'b10111000; //  924 : 184 - 0xb8
      11'h39D: dout  = 8'b10110000; //  925 : 176 - 0xb0
      11'h39E: dout  = 8'b10000000; //  926 : 128 - 0x80
      11'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      11'h3A0: dout  = 8'b00110000; //  928 :  48 - 0x30 -- Sprite 0x74
      11'h3A1: dout  = 8'b01111100; //  929 : 124 - 0x7c
      11'h3A2: dout  = 8'b11111111; //  930 : 255 - 0xff
      11'h3A3: dout  = 8'b11111111; //  931 : 255 - 0xff
      11'h3A4: dout  = 8'b11011111; //  932 : 223 - 0xdf
      11'h3A5: dout  = 8'b00001011; //  933 :  11 - 0xb
      11'h3A6: dout  = 8'b00011111; //  934 :  31 - 0x1f
      11'h3A7: dout  = 8'b01111111; //  935 : 127 - 0x7f
      11'h3A8: dout  = 8'b01111111; //  936 : 127 - 0x7f -- Sprite 0x75
      11'h3A9: dout  = 8'b00001011; //  937 :  11 - 0xb
      11'h3AA: dout  = 8'b00110011; //  938 :  51 - 0x33
      11'h3AB: dout  = 8'b00110110; //  939 :  54 - 0x36
      11'h3AC: dout  = 8'b00010000; //  940 :  16 - 0x10
      11'h3AD: dout  = 8'b00001010; //  941 :  10 - 0xa
      11'h3AE: dout  = 8'b00001111; //  942 :  15 - 0xf
      11'h3AF: dout  = 8'b00000111; //  943 :   7 - 0x7
      11'h3B0: dout  = 8'b00111000; //  944 :  56 - 0x38 -- Sprite 0x76
      11'h3B1: dout  = 8'b01111100; //  945 : 124 - 0x7c
      11'h3B2: dout  = 8'b11111100; //  946 : 252 - 0xfc
      11'h3B3: dout  = 8'b11111100; //  947 : 252 - 0xfc
      11'h3B4: dout  = 8'b11101100; //  948 : 236 - 0xec
      11'h3B5: dout  = 8'b10100000; //  949 : 160 - 0xa0
      11'h3B6: dout  = 8'b11110000; //  950 : 240 - 0xf0
      11'h3B7: dout  = 8'b11111100; //  951 : 252 - 0xfc
      11'h3B8: dout  = 8'b11111100; //  952 : 252 - 0xfc -- Sprite 0x77
      11'h3B9: dout  = 8'b10100000; //  953 : 160 - 0xa0
      11'h3BA: dout  = 8'b10011000; //  954 : 152 - 0x98
      11'h3BB: dout  = 8'b11011000; //  955 : 216 - 0xd8
      11'h3BC: dout  = 8'b00010000; //  956 :  16 - 0x10
      11'h3BD: dout  = 8'b10100000; //  957 : 160 - 0xa0
      11'h3BE: dout  = 8'b11100000; //  958 : 224 - 0xe0
      11'h3BF: dout  = 8'b11000000; //  959 : 192 - 0xc0
      11'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x78
      11'h3C1: dout  = 8'b00000001; //  961 :   1 - 0x1
      11'h3C2: dout  = 8'b00001101; //  962 :  13 - 0xd
      11'h3C3: dout  = 8'b00011101; //  963 :  29 - 0x1d
      11'h3C4: dout  = 8'b01100011; //  964 :  99 - 0x63
      11'h3C5: dout  = 8'b11001001; //  965 : 201 - 0xc9
      11'h3C6: dout  = 8'b11101111; //  966 : 239 - 0xef
      11'h3C7: dout  = 8'b11000111; //  967 : 199 - 0xc7
      11'h3C8: dout  = 8'b11101111; //  968 : 239 - 0xef -- Sprite 0x79
      11'h3C9: dout  = 8'b11001001; //  969 : 201 - 0xc9
      11'h3CA: dout  = 8'b01100011; //  970 :  99 - 0x63
      11'h3CB: dout  = 8'b00011101; //  971 :  29 - 0x1d
      11'h3CC: dout  = 8'b00001101; //  972 :  13 - 0xd
      11'h3CD: dout  = 8'b00000001; //  973 :   1 - 0x1
      11'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      11'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      11'h3D0: dout  = 8'b00011100; //  976 :  28 - 0x1c -- Sprite 0x7a
      11'h3D1: dout  = 8'b10011110; //  977 : 158 - 0x9e
      11'h3D2: dout  = 8'b10001111; //  978 : 143 - 0x8f
      11'h3D3: dout  = 8'b11011111; //  979 : 223 - 0xdf
      11'h3D4: dout  = 8'b11111110; //  980 : 254 - 0xfe
      11'h3D5: dout  = 8'b11011110; //  981 : 222 - 0xde
      11'h3D6: dout  = 8'b11111100; //  982 : 252 - 0xfc
      11'h3D7: dout  = 8'b11111100; //  983 : 252 - 0xfc
      11'h3D8: dout  = 8'b11111100; //  984 : 252 - 0xfc -- Sprite 0x7b
      11'h3D9: dout  = 8'b11011110; //  985 : 222 - 0xde
      11'h3DA: dout  = 8'b11111111; //  986 : 255 - 0xff
      11'h3DB: dout  = 8'b11001111; //  987 : 207 - 0xcf
      11'h3DC: dout  = 8'b10011111; //  988 : 159 - 0x9f
      11'h3DD: dout  = 8'b10011110; //  989 : 158 - 0x9e
      11'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      11'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      11'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      11'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      11'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      11'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      11'h3E4: dout  = 8'b00011110; //  996 :  30 - 0x1e
      11'h3E5: dout  = 8'b00111111; //  997 :  63 - 0x3f
      11'h3E6: dout  = 8'b01111101; //  998 : 125 - 0x7d
      11'h3E7: dout  = 8'b01111000; //  999 : 120 - 0x78
      11'h3E8: dout  = 8'b01111100; // 1000 : 124 - 0x7c -- Sprite 0x7d
      11'h3E9: dout  = 8'b11111011; // 1001 : 251 - 0xfb
      11'h3EA: dout  = 8'b11111111; // 1002 : 255 - 0xff
      11'h3EB: dout  = 8'b11111111; // 1003 : 255 - 0xff
      11'h3EC: dout  = 8'b01011111; // 1004 :  95 - 0x5f
      11'h3ED: dout  = 8'b00011111; // 1005 :  31 - 0x1f
      11'h3EE: dout  = 8'b00011111; // 1006 :  31 - 0x1f
      11'h3EF: dout  = 8'b00011111; // 1007 :  31 - 0x1f
      11'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x7e
      11'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      11'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      11'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      11'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      11'h3F5: dout  = 8'b10000000; // 1013 : 128 - 0x80
      11'h3F6: dout  = 8'b10000000; // 1014 : 128 - 0x80
      11'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      11'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0 -- Sprite 0x7f
      11'h3F9: dout  = 8'b00100001; // 1017 :  33 - 0x21
      11'h3FA: dout  = 8'b10100010; // 1018 : 162 - 0xa2
      11'h3FB: dout  = 8'b10100011; // 1019 : 163 - 0xa3
      11'h3FC: dout  = 8'b10110011; // 1020 : 179 - 0xb3
      11'h3FD: dout  = 8'b10001111; // 1021 : 143 - 0x8f
      11'h3FE: dout  = 8'b00100111; // 1022 :  39 - 0x27
      11'h3FF: dout  = 8'b11111110; // 1023 : 254 - 0xfe
      11'h400: dout  = 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x80
      11'h401: dout  = 8'b00000000; // 1025 :   0 - 0x0
      11'h402: dout  = 8'b00000000; // 1026 :   0 - 0x0
      11'h403: dout  = 8'b00000000; // 1027 :   0 - 0x0
      11'h404: dout  = 8'b00000011; // 1028 :   3 - 0x3
      11'h405: dout  = 8'b00001111; // 1029 :  15 - 0xf
      11'h406: dout  = 8'b00011111; // 1030 :  31 - 0x1f
      11'h407: dout  = 8'b00011111; // 1031 :  31 - 0x1f
      11'h408: dout  = 8'b00011111; // 1032 :  31 - 0x1f -- Sprite 0x81
      11'h409: dout  = 8'b00011111; // 1033 :  31 - 0x1f
      11'h40A: dout  = 8'b00001111; // 1034 :  15 - 0xf
      11'h40B: dout  = 8'b00000011; // 1035 :   3 - 0x3
      11'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      11'h40D: dout  = 8'b00000000; // 1037 :   0 - 0x0
      11'h40E: dout  = 8'b00000000; // 1038 :   0 - 0x0
      11'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      11'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x82
      11'h411: dout  = 8'b00000000; // 1041 :   0 - 0x0
      11'h412: dout  = 8'b00000000; // 1042 :   0 - 0x0
      11'h413: dout  = 8'b00000000; // 1043 :   0 - 0x0
      11'h414: dout  = 8'b11000000; // 1044 : 192 - 0xc0
      11'h415: dout  = 8'b11110000; // 1045 : 240 - 0xf0
      11'h416: dout  = 8'b11111000; // 1046 : 248 - 0xf8
      11'h417: dout  = 8'b11111000; // 1047 : 248 - 0xf8
      11'h418: dout  = 8'b11111000; // 1048 : 248 - 0xf8 -- Sprite 0x83
      11'h419: dout  = 8'b11111000; // 1049 : 248 - 0xf8
      11'h41A: dout  = 8'b11110000; // 1050 : 240 - 0xf0
      11'h41B: dout  = 8'b11000000; // 1051 : 192 - 0xc0
      11'h41C: dout  = 8'b00000000; // 1052 :   0 - 0x0
      11'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      11'h41E: dout  = 8'b00000000; // 1054 :   0 - 0x0
      11'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      11'h420: dout  = 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x84
      11'h421: dout  = 8'b00000000; // 1057 :   0 - 0x0
      11'h422: dout  = 8'b00000000; // 1058 :   0 - 0x0
      11'h423: dout  = 8'b00000000; // 1059 :   0 - 0x0
      11'h424: dout  = 8'b00000011; // 1060 :   3 - 0x3
      11'h425: dout  = 8'b00001111; // 1061 :  15 - 0xf
      11'h426: dout  = 8'b00011111; // 1062 :  31 - 0x1f
      11'h427: dout  = 8'b00011111; // 1063 :  31 - 0x1f
      11'h428: dout  = 8'b00011111; // 1064 :  31 - 0x1f -- Sprite 0x85
      11'h429: dout  = 8'b00011111; // 1065 :  31 - 0x1f
      11'h42A: dout  = 8'b00001111; // 1066 :  15 - 0xf
      11'h42B: dout  = 8'b00000011; // 1067 :   3 - 0x3
      11'h42C: dout  = 8'b00000000; // 1068 :   0 - 0x0
      11'h42D: dout  = 8'b00000000; // 1069 :   0 - 0x0
      11'h42E: dout  = 8'b00000000; // 1070 :   0 - 0x0
      11'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      11'h430: dout  = 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x86
      11'h431: dout  = 8'b00000000; // 1073 :   0 - 0x0
      11'h432: dout  = 8'b00000000; // 1074 :   0 - 0x0
      11'h433: dout  = 8'b00000000; // 1075 :   0 - 0x0
      11'h434: dout  = 8'b11000000; // 1076 : 192 - 0xc0
      11'h435: dout  = 8'b11110000; // 1077 : 240 - 0xf0
      11'h436: dout  = 8'b11111000; // 1078 : 248 - 0xf8
      11'h437: dout  = 8'b11111000; // 1079 : 248 - 0xf8
      11'h438: dout  = 8'b11111000; // 1080 : 248 - 0xf8 -- Sprite 0x87
      11'h439: dout  = 8'b11111000; // 1081 : 248 - 0xf8
      11'h43A: dout  = 8'b11110000; // 1082 : 240 - 0xf0
      11'h43B: dout  = 8'b11000000; // 1083 : 192 - 0xc0
      11'h43C: dout  = 8'b00000000; // 1084 :   0 - 0x0
      11'h43D: dout  = 8'b00000000; // 1085 :   0 - 0x0
      11'h43E: dout  = 8'b00000000; // 1086 :   0 - 0x0
      11'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      11'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x88
      11'h441: dout  = 8'b00000000; // 1089 :   0 - 0x0
      11'h442: dout  = 8'b00000000; // 1090 :   0 - 0x0
      11'h443: dout  = 8'b00000000; // 1091 :   0 - 0x0
      11'h444: dout  = 8'b00000011; // 1092 :   3 - 0x3
      11'h445: dout  = 8'b00001111; // 1093 :  15 - 0xf
      11'h446: dout  = 8'b00011111; // 1094 :  31 - 0x1f
      11'h447: dout  = 8'b00011111; // 1095 :  31 - 0x1f
      11'h448: dout  = 8'b00011111; // 1096 :  31 - 0x1f -- Sprite 0x89
      11'h449: dout  = 8'b00011111; // 1097 :  31 - 0x1f
      11'h44A: dout  = 8'b00001111; // 1098 :  15 - 0xf
      11'h44B: dout  = 8'b00000011; // 1099 :   3 - 0x3
      11'h44C: dout  = 8'b00000000; // 1100 :   0 - 0x0
      11'h44D: dout  = 8'b00000000; // 1101 :   0 - 0x0
      11'h44E: dout  = 8'b00000000; // 1102 :   0 - 0x0
      11'h44F: dout  = 8'b00000000; // 1103 :   0 - 0x0
      11'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x8a
      11'h451: dout  = 8'b00000000; // 1105 :   0 - 0x0
      11'h452: dout  = 8'b00000000; // 1106 :   0 - 0x0
      11'h453: dout  = 8'b00000000; // 1107 :   0 - 0x0
      11'h454: dout  = 8'b11000000; // 1108 : 192 - 0xc0
      11'h455: dout  = 8'b11110000; // 1109 : 240 - 0xf0
      11'h456: dout  = 8'b11111000; // 1110 : 248 - 0xf8
      11'h457: dout  = 8'b11111000; // 1111 : 248 - 0xf8
      11'h458: dout  = 8'b11111000; // 1112 : 248 - 0xf8 -- Sprite 0x8b
      11'h459: dout  = 8'b11111000; // 1113 : 248 - 0xf8
      11'h45A: dout  = 8'b11110000; // 1114 : 240 - 0xf0
      11'h45B: dout  = 8'b11000000; // 1115 : 192 - 0xc0
      11'h45C: dout  = 8'b00000000; // 1116 :   0 - 0x0
      11'h45D: dout  = 8'b00000000; // 1117 :   0 - 0x0
      11'h45E: dout  = 8'b00000000; // 1118 :   0 - 0x0
      11'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      11'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x8c
      11'h461: dout  = 8'b00000000; // 1121 :   0 - 0x0
      11'h462: dout  = 8'b00000000; // 1122 :   0 - 0x0
      11'h463: dout  = 8'b00000000; // 1123 :   0 - 0x0
      11'h464: dout  = 8'b00000011; // 1124 :   3 - 0x3
      11'h465: dout  = 8'b00001111; // 1125 :  15 - 0xf
      11'h466: dout  = 8'b00011111; // 1126 :  31 - 0x1f
      11'h467: dout  = 8'b00011111; // 1127 :  31 - 0x1f
      11'h468: dout  = 8'b00011111; // 1128 :  31 - 0x1f -- Sprite 0x8d
      11'h469: dout  = 8'b00011111; // 1129 :  31 - 0x1f
      11'h46A: dout  = 8'b00001111; // 1130 :  15 - 0xf
      11'h46B: dout  = 8'b00000011; // 1131 :   3 - 0x3
      11'h46C: dout  = 8'b00000000; // 1132 :   0 - 0x0
      11'h46D: dout  = 8'b00000000; // 1133 :   0 - 0x0
      11'h46E: dout  = 8'b00000000; // 1134 :   0 - 0x0
      11'h46F: dout  = 8'b00000000; // 1135 :   0 - 0x0
      11'h470: dout  = 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x8e
      11'h471: dout  = 8'b00000000; // 1137 :   0 - 0x0
      11'h472: dout  = 8'b00000000; // 1138 :   0 - 0x0
      11'h473: dout  = 8'b00000000; // 1139 :   0 - 0x0
      11'h474: dout  = 8'b11000000; // 1140 : 192 - 0xc0
      11'h475: dout  = 8'b11110000; // 1141 : 240 - 0xf0
      11'h476: dout  = 8'b11111000; // 1142 : 248 - 0xf8
      11'h477: dout  = 8'b11111000; // 1143 : 248 - 0xf8
      11'h478: dout  = 8'b11111000; // 1144 : 248 - 0xf8 -- Sprite 0x8f
      11'h479: dout  = 8'b11111000; // 1145 : 248 - 0xf8
      11'h47A: dout  = 8'b11110000; // 1146 : 240 - 0xf0
      11'h47B: dout  = 8'b11000000; // 1147 : 192 - 0xc0
      11'h47C: dout  = 8'b00000000; // 1148 :   0 - 0x0
      11'h47D: dout  = 8'b00000000; // 1149 :   0 - 0x0
      11'h47E: dout  = 8'b00000000; // 1150 :   0 - 0x0
      11'h47F: dout  = 8'b00000000; // 1151 :   0 - 0x0
      11'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      11'h481: dout  = 8'b00000000; // 1153 :   0 - 0x0
      11'h482: dout  = 8'b00000000; // 1154 :   0 - 0x0
      11'h483: dout  = 8'b00001111; // 1155 :  15 - 0xf
      11'h484: dout  = 8'b00110000; // 1156 :  48 - 0x30
      11'h485: dout  = 8'b01100000; // 1157 :  96 - 0x60
      11'h486: dout  = 8'b00111111; // 1158 :  63 - 0x3f
      11'h487: dout  = 8'b01111111; // 1159 : 127 - 0x7f
      11'h488: dout  = 8'b01111111; // 1160 : 127 - 0x7f -- Sprite 0x91
      11'h489: dout  = 8'b00111111; // 1161 :  63 - 0x3f
      11'h48A: dout  = 8'b01100000; // 1162 :  96 - 0x60
      11'h48B: dout  = 8'b00110000; // 1163 :  48 - 0x30
      11'h48C: dout  = 8'b00001111; // 1164 :  15 - 0xf
      11'h48D: dout  = 8'b00000000; // 1165 :   0 - 0x0
      11'h48E: dout  = 8'b00000000; // 1166 :   0 - 0x0
      11'h48F: dout  = 8'b00000000; // 1167 :   0 - 0x0
      11'h490: dout  = 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x92
      11'h491: dout  = 8'b00000000; // 1169 :   0 - 0x0
      11'h492: dout  = 8'b00000000; // 1170 :   0 - 0x0
      11'h493: dout  = 8'b11111000; // 1171 : 248 - 0xf8
      11'h494: dout  = 8'b00000110; // 1172 :   6 - 0x6
      11'h495: dout  = 8'b00000011; // 1173 :   3 - 0x3
      11'h496: dout  = 8'b11111110; // 1174 : 254 - 0xfe
      11'h497: dout  = 8'b11111111; // 1175 : 255 - 0xff
      11'h498: dout  = 8'b11111111; // 1176 : 255 - 0xff -- Sprite 0x93
      11'h499: dout  = 8'b11111110; // 1177 : 254 - 0xfe
      11'h49A: dout  = 8'b00000011; // 1178 :   3 - 0x3
      11'h49B: dout  = 8'b00000110; // 1179 :   6 - 0x6
      11'h49C: dout  = 8'b11111000; // 1180 : 248 - 0xf8
      11'h49D: dout  = 8'b00000000; // 1181 :   0 - 0x0
      11'h49E: dout  = 8'b00000000; // 1182 :   0 - 0x0
      11'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      11'h4A0: dout  = 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x94
      11'h4A1: dout  = 8'b00000000; // 1185 :   0 - 0x0
      11'h4A2: dout  = 8'b00000000; // 1186 :   0 - 0x0
      11'h4A3: dout  = 8'b00000000; // 1187 :   0 - 0x0
      11'h4A4: dout  = 8'b00101111; // 1188 :  47 - 0x2f
      11'h4A5: dout  = 8'b00111111; // 1189 :  63 - 0x3f
      11'h4A6: dout  = 8'b01100000; // 1190 :  96 - 0x60
      11'h4A7: dout  = 8'b00100000; // 1191 :  32 - 0x20
      11'h4A8: dout  = 8'b00100000; // 1192 :  32 - 0x20 -- Sprite 0x95
      11'h4A9: dout  = 8'b01100000; // 1193 :  96 - 0x60
      11'h4AA: dout  = 8'b00111111; // 1194 :  63 - 0x3f
      11'h4AB: dout  = 8'b00101111; // 1195 :  47 - 0x2f
      11'h4AC: dout  = 8'b00000000; // 1196 :   0 - 0x0
      11'h4AD: dout  = 8'b00000000; // 1197 :   0 - 0x0
      11'h4AE: dout  = 8'b00000000; // 1198 :   0 - 0x0
      11'h4AF: dout  = 8'b00000000; // 1199 :   0 - 0x0
      11'h4B0: dout  = 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x96
      11'h4B1: dout  = 8'b00000000; // 1201 :   0 - 0x0
      11'h4B2: dout  = 8'b00000000; // 1202 :   0 - 0x0
      11'h4B3: dout  = 8'b00000000; // 1203 :   0 - 0x0
      11'h4B4: dout  = 8'b11111010; // 1204 : 250 - 0xfa
      11'h4B5: dout  = 8'b11111110; // 1205 : 254 - 0xfe
      11'h4B6: dout  = 8'b00000011; // 1206 :   3 - 0x3
      11'h4B7: dout  = 8'b00000010; // 1207 :   2 - 0x2
      11'h4B8: dout  = 8'b00000010; // 1208 :   2 - 0x2 -- Sprite 0x97
      11'h4B9: dout  = 8'b00000011; // 1209 :   3 - 0x3
      11'h4BA: dout  = 8'b11111110; // 1210 : 254 - 0xfe
      11'h4BB: dout  = 8'b11111010; // 1211 : 250 - 0xfa
      11'h4BC: dout  = 8'b00000000; // 1212 :   0 - 0x0
      11'h4BD: dout  = 8'b00000000; // 1213 :   0 - 0x0
      11'h4BE: dout  = 8'b00000000; // 1214 :   0 - 0x0
      11'h4BF: dout  = 8'b00000000; // 1215 :   0 - 0x0
      11'h4C0: dout  = 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x98
      11'h4C1: dout  = 8'b01000100; // 1217 :  68 - 0x44
      11'h4C2: dout  = 8'b00000000; // 1218 :   0 - 0x0
      11'h4C3: dout  = 8'b01000001; // 1219 :  65 - 0x41
      11'h4C4: dout  = 8'b00100000; // 1220 :  32 - 0x20
      11'h4C5: dout  = 8'b01001011; // 1221 :  75 - 0x4b
      11'h4C6: dout  = 8'b00100111; // 1222 :  39 - 0x27
      11'h4C7: dout  = 8'b00011111; // 1223 :  31 - 0x1f
      11'h4C8: dout  = 8'b00001111; // 1224 :  15 - 0xf -- Sprite 0x99
      11'h4C9: dout  = 8'b00011110; // 1225 :  30 - 0x1e
      11'h4CA: dout  = 8'b00011111; // 1226 :  31 - 0x1f
      11'h4CB: dout  = 8'b00011111; // 1227 :  31 - 0x1f
      11'h4CC: dout  = 8'b00011111; // 1228 :  31 - 0x1f
      11'h4CD: dout  = 8'b00001111; // 1229 :  15 - 0xf
      11'h4CE: dout  = 8'b00001111; // 1230 :  15 - 0xf
      11'h4CF: dout  = 8'b00000011; // 1231 :   3 - 0x3
      11'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      11'h4D1: dout  = 8'b00100000; // 1233 :  32 - 0x20
      11'h4D2: dout  = 8'b01010000; // 1234 :  80 - 0x50
      11'h4D3: dout  = 8'b00100000; // 1235 :  32 - 0x20
      11'h4D4: dout  = 8'b01100000; // 1236 :  96 - 0x60
      11'h4D5: dout  = 8'b01001000; // 1237 :  72 - 0x48
      11'h4D6: dout  = 8'b11100000; // 1238 : 224 - 0xe0
      11'h4D7: dout  = 8'b11110000; // 1239 : 240 - 0xf0
      11'h4D8: dout  = 8'b11111000; // 1240 : 248 - 0xf8 -- Sprite 0x9b
      11'h4D9: dout  = 8'b01111000; // 1241 : 120 - 0x78
      11'h4DA: dout  = 8'b00111100; // 1242 :  60 - 0x3c
      11'h4DB: dout  = 8'b00111100; // 1243 :  60 - 0x3c
      11'h4DC: dout  = 8'b00111100; // 1244 :  60 - 0x3c
      11'h4DD: dout  = 8'b11111100; // 1245 : 252 - 0xfc
      11'h4DE: dout  = 8'b11111000; // 1246 : 248 - 0xf8
      11'h4DF: dout  = 8'b11100000; // 1247 : 224 - 0xe0
      11'h4E0: dout  = 8'b00010000; // 1248 :  16 - 0x10 -- Sprite 0x9c
      11'h4E1: dout  = 8'b00000001; // 1249 :   1 - 0x1
      11'h4E2: dout  = 8'b00101010; // 1250 :  42 - 0x2a
      11'h4E3: dout  = 8'b00001100; // 1251 :  12 - 0xc
      11'h4E4: dout  = 8'b10100110; // 1252 : 166 - 0xa6
      11'h4E5: dout  = 8'b00010111; // 1253 :  23 - 0x17
      11'h4E6: dout  = 8'b00011111; // 1254 :  31 - 0x1f
      11'h4E7: dout  = 8'b00011111; // 1255 :  31 - 0x1f
      11'h4E8: dout  = 8'b01011110; // 1256 :  94 - 0x5e -- Sprite 0x9d
      11'h4E9: dout  = 8'b00111100; // 1257 :  60 - 0x3c
      11'h4EA: dout  = 8'b00111101; // 1258 :  61 - 0x3d
      11'h4EB: dout  = 8'b00111101; // 1259 :  61 - 0x3d
      11'h4EC: dout  = 8'b00111110; // 1260 :  62 - 0x3e
      11'h4ED: dout  = 8'b00011111; // 1261 :  31 - 0x1f
      11'h4EE: dout  = 8'b00001111; // 1262 :  15 - 0xf
      11'h4EF: dout  = 8'b00000111; // 1263 :   7 - 0x7
      11'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Sprite 0x9e
      11'h4F1: dout  = 8'b00000000; // 1265 :   0 - 0x0
      11'h4F2: dout  = 8'b10000000; // 1266 : 128 - 0x80
      11'h4F3: dout  = 8'b11001000; // 1267 : 200 - 0xc8
      11'h4F4: dout  = 8'b01100000; // 1268 :  96 - 0x60
      11'h4F5: dout  = 8'b11100000; // 1269 : 224 - 0xe0
      11'h4F6: dout  = 8'b11110100; // 1270 : 244 - 0xf4
      11'h4F7: dout  = 8'b11111000; // 1271 : 248 - 0xf8
      11'h4F8: dout  = 8'b01111100; // 1272 : 124 - 0x7c -- Sprite 0x9f
      11'h4F9: dout  = 8'b00011100; // 1273 :  28 - 0x1c
      11'h4FA: dout  = 8'b00101110; // 1274 :  46 - 0x2e
      11'h4FB: dout  = 8'b00101110; // 1275 :  46 - 0x2e
      11'h4FC: dout  = 8'b00011110; // 1276 :  30 - 0x1e
      11'h4FD: dout  = 8'b11111100; // 1277 : 252 - 0xfc
      11'h4FE: dout  = 8'b11111000; // 1278 : 248 - 0xf8
      11'h4FF: dout  = 8'b11100000; // 1279 : 224 - 0xe0
      11'h500: dout  = 8'b11111111; // 1280 : 255 - 0xff -- Sprite 0xa0
      11'h501: dout  = 8'b11111111; // 1281 : 255 - 0xff
      11'h502: dout  = 8'b00111000; // 1282 :  56 - 0x38
      11'h503: dout  = 8'b01101100; // 1283 : 108 - 0x6c
      11'h504: dout  = 8'b11000110; // 1284 : 198 - 0xc6
      11'h505: dout  = 8'b10000011; // 1285 : 131 - 0x83
      11'h506: dout  = 8'b11111111; // 1286 : 255 - 0xff
      11'h507: dout  = 8'b11111111; // 1287 : 255 - 0xff
      11'h508: dout  = 8'b11111111; // 1288 : 255 - 0xff -- Sprite 0xa1
      11'h509: dout  = 8'b11111111; // 1289 : 255 - 0xff
      11'h50A: dout  = 8'b00111000; // 1290 :  56 - 0x38
      11'h50B: dout  = 8'b01101100; // 1291 : 108 - 0x6c
      11'h50C: dout  = 8'b11000110; // 1292 : 198 - 0xc6
      11'h50D: dout  = 8'b10000011; // 1293 : 131 - 0x83
      11'h50E: dout  = 8'b11111111; // 1294 : 255 - 0xff
      11'h50F: dout  = 8'b11111111; // 1295 : 255 - 0xff
      11'h510: dout  = 8'b10010010; // 1296 : 146 - 0x92 -- Sprite 0xa2
      11'h511: dout  = 8'b01010100; // 1297 :  84 - 0x54
      11'h512: dout  = 8'b00111000; // 1298 :  56 - 0x38
      11'h513: dout  = 8'b11111110; // 1299 : 254 - 0xfe
      11'h514: dout  = 8'b00111000; // 1300 :  56 - 0x38
      11'h515: dout  = 8'b01010100; // 1301 :  84 - 0x54
      11'h516: dout  = 8'b10010010; // 1302 : 146 - 0x92
      11'h517: dout  = 8'b00000000; // 1303 :   0 - 0x0
      11'h518: dout  = 8'b11111111; // 1304 : 255 - 0xff -- Sprite 0xa3
      11'h519: dout  = 8'b11111111; // 1305 : 255 - 0xff
      11'h51A: dout  = 8'b11111111; // 1306 : 255 - 0xff
      11'h51B: dout  = 8'b11111111; // 1307 : 255 - 0xff
      11'h51C: dout  = 8'b11111111; // 1308 : 255 - 0xff
      11'h51D: dout  = 8'b11111111; // 1309 : 255 - 0xff
      11'h51E: dout  = 8'b11111111; // 1310 : 255 - 0xff
      11'h51F: dout  = 8'b11111111; // 1311 : 255 - 0xff
      11'h520: dout  = 8'b11111111; // 1312 : 255 - 0xff -- Sprite 0xa4
      11'h521: dout  = 8'b11111111; // 1313 : 255 - 0xff
      11'h522: dout  = 8'b11111111; // 1314 : 255 - 0xff
      11'h523: dout  = 8'b11111111; // 1315 : 255 - 0xff
      11'h524: dout  = 8'b11111111; // 1316 : 255 - 0xff
      11'h525: dout  = 8'b11111111; // 1317 : 255 - 0xff
      11'h526: dout  = 8'b11111111; // 1318 : 255 - 0xff
      11'h527: dout  = 8'b11111111; // 1319 : 255 - 0xff
      11'h528: dout  = 8'b11111111; // 1320 : 255 - 0xff -- Sprite 0xa5
      11'h529: dout  = 8'b11111111; // 1321 : 255 - 0xff
      11'h52A: dout  = 8'b11111111; // 1322 : 255 - 0xff
      11'h52B: dout  = 8'b11111111; // 1323 : 255 - 0xff
      11'h52C: dout  = 8'b11111111; // 1324 : 255 - 0xff
      11'h52D: dout  = 8'b11111111; // 1325 : 255 - 0xff
      11'h52E: dout  = 8'b11111111; // 1326 : 255 - 0xff
      11'h52F: dout  = 8'b11111111; // 1327 : 255 - 0xff
      11'h530: dout  = 8'b11111111; // 1328 : 255 - 0xff -- Sprite 0xa6
      11'h531: dout  = 8'b11111111; // 1329 : 255 - 0xff
      11'h532: dout  = 8'b11111111; // 1330 : 255 - 0xff
      11'h533: dout  = 8'b11111111; // 1331 : 255 - 0xff
      11'h534: dout  = 8'b11111111; // 1332 : 255 - 0xff
      11'h535: dout  = 8'b11111111; // 1333 : 255 - 0xff
      11'h536: dout  = 8'b11111111; // 1334 : 255 - 0xff
      11'h537: dout  = 8'b11111111; // 1335 : 255 - 0xff
      11'h538: dout  = 8'b11111111; // 1336 : 255 - 0xff -- Sprite 0xa7
      11'h539: dout  = 8'b11111111; // 1337 : 255 - 0xff
      11'h53A: dout  = 8'b11111111; // 1338 : 255 - 0xff
      11'h53B: dout  = 8'b11111111; // 1339 : 255 - 0xff
      11'h53C: dout  = 8'b11111111; // 1340 : 255 - 0xff
      11'h53D: dout  = 8'b11111111; // 1341 : 255 - 0xff
      11'h53E: dout  = 8'b11111111; // 1342 : 255 - 0xff
      11'h53F: dout  = 8'b11111111; // 1343 : 255 - 0xff
      11'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0xa8
      11'h541: dout  = 8'b00000000; // 1345 :   0 - 0x0
      11'h542: dout  = 8'b00000000; // 1346 :   0 - 0x0
      11'h543: dout  = 8'b00000000; // 1347 :   0 - 0x0
      11'h544: dout  = 8'b00000000; // 1348 :   0 - 0x0
      11'h545: dout  = 8'b00100011; // 1349 :  35 - 0x23
      11'h546: dout  = 8'b10010111; // 1350 : 151 - 0x97
      11'h547: dout  = 8'b00101111; // 1351 :  47 - 0x2f
      11'h548: dout  = 8'b01101110; // 1352 : 110 - 0x6e -- Sprite 0xa9
      11'h549: dout  = 8'b11101111; // 1353 : 239 - 0xef
      11'h54A: dout  = 8'b11110111; // 1354 : 247 - 0xf7
      11'h54B: dout  = 8'b11111111; // 1355 : 255 - 0xff
      11'h54C: dout  = 8'b01111111; // 1356 : 127 - 0x7f
      11'h54D: dout  = 8'b00111111; // 1357 :  63 - 0x3f
      11'h54E: dout  = 8'b01011111; // 1358 :  95 - 0x5f
      11'h54F: dout  = 8'b00001111; // 1359 :  15 - 0xf
      11'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      11'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      11'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      11'h553: dout  = 8'b00000000; // 1363 :   0 - 0x0
      11'h554: dout  = 8'b11111000; // 1364 : 248 - 0xf8
      11'h555: dout  = 8'b11111100; // 1365 : 252 - 0xfc
      11'h556: dout  = 8'b11111110; // 1366 : 254 - 0xfe
      11'h557: dout  = 8'b01011110; // 1367 :  94 - 0x5e
      11'h558: dout  = 8'b01011110; // 1368 :  94 - 0x5e -- Sprite 0xab
      11'h559: dout  = 8'b00001100; // 1369 :  12 - 0xc
      11'h55A: dout  = 8'b10011110; // 1370 : 158 - 0x9e
      11'h55B: dout  = 8'b11111110; // 1371 : 254 - 0xfe
      11'h55C: dout  = 8'b11111110; // 1372 : 254 - 0xfe
      11'h55D: dout  = 8'b11111110; // 1373 : 254 - 0xfe
      11'h55E: dout  = 8'b11111000; // 1374 : 248 - 0xf8
      11'h55F: dout  = 8'b11000000; // 1375 : 192 - 0xc0
      11'h560: dout  = 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      11'h561: dout  = 8'b00000000; // 1377 :   0 - 0x0
      11'h562: dout  = 8'b00000000; // 1378 :   0 - 0x0
      11'h563: dout  = 8'b00000000; // 1379 :   0 - 0x0
      11'h564: dout  = 8'b00000000; // 1380 :   0 - 0x0
      11'h565: dout  = 8'b00000011; // 1381 :   3 - 0x3
      11'h566: dout  = 8'b00000111; // 1382 :   7 - 0x7
      11'h567: dout  = 8'b00101111; // 1383 :  47 - 0x2f
      11'h568: dout  = 8'b01001110; // 1384 :  78 - 0x4e -- Sprite 0xad
      11'h569: dout  = 8'b01101110; // 1385 : 110 - 0x6e
      11'h56A: dout  = 8'b11111110; // 1386 : 254 - 0xfe
      11'h56B: dout  = 8'b01111111; // 1387 : 127 - 0x7f
      11'h56C: dout  = 8'b00111111; // 1388 :  63 - 0x3f
      11'h56D: dout  = 8'b00011111; // 1389 :  31 - 0x1f
      11'h56E: dout  = 8'b00001111; // 1390 :  15 - 0xf
      11'h56F: dout  = 8'b00000011; // 1391 :   3 - 0x3
      11'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      11'h571: dout  = 8'b00000000; // 1393 :   0 - 0x0
      11'h572: dout  = 8'b00000000; // 1394 :   0 - 0x0
      11'h573: dout  = 8'b00000000; // 1395 :   0 - 0x0
      11'h574: dout  = 8'b11111000; // 1396 : 248 - 0xf8
      11'h575: dout  = 8'b11111100; // 1397 : 252 - 0xfc
      11'h576: dout  = 8'b11111110; // 1398 : 254 - 0xfe
      11'h577: dout  = 8'b01010110; // 1399 :  86 - 0x56
      11'h578: dout  = 8'b01010110; // 1400 :  86 - 0x56 -- Sprite 0xaf
      11'h579: dout  = 8'b00001100; // 1401 :  12 - 0xc
      11'h57A: dout  = 8'b00001110; // 1402 :  14 - 0xe
      11'h57B: dout  = 8'b00011111; // 1403 :  31 - 0x1f
      11'h57C: dout  = 8'b11111111; // 1404 : 255 - 0xff
      11'h57D: dout  = 8'b11111111; // 1405 : 255 - 0xff
      11'h57E: dout  = 8'b11111110; // 1406 : 254 - 0xfe
      11'h57F: dout  = 8'b11111000; // 1407 : 248 - 0xf8
      11'h580: dout  = 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0xb0
      11'h581: dout  = 8'b11111111; // 1409 : 255 - 0xff
      11'h582: dout  = 8'b11111111; // 1410 : 255 - 0xff
      11'h583: dout  = 8'b11111111; // 1411 : 255 - 0xff
      11'h584: dout  = 8'b11111111; // 1412 : 255 - 0xff
      11'h585: dout  = 8'b11111111; // 1413 : 255 - 0xff
      11'h586: dout  = 8'b11111111; // 1414 : 255 - 0xff
      11'h587: dout  = 8'b11111111; // 1415 : 255 - 0xff
      11'h588: dout  = 8'b11111111; // 1416 : 255 - 0xff -- Sprite 0xb1
      11'h589: dout  = 8'b11111111; // 1417 : 255 - 0xff
      11'h58A: dout  = 8'b11111111; // 1418 : 255 - 0xff
      11'h58B: dout  = 8'b11111111; // 1419 : 255 - 0xff
      11'h58C: dout  = 8'b11111111; // 1420 : 255 - 0xff
      11'h58D: dout  = 8'b11111111; // 1421 : 255 - 0xff
      11'h58E: dout  = 8'b11111111; // 1422 : 255 - 0xff
      11'h58F: dout  = 8'b11111111; // 1423 : 255 - 0xff
      11'h590: dout  = 8'b11111111; // 1424 : 255 - 0xff -- Sprite 0xb2
      11'h591: dout  = 8'b11111111; // 1425 : 255 - 0xff
      11'h592: dout  = 8'b11111111; // 1426 : 255 - 0xff
      11'h593: dout  = 8'b11111111; // 1427 : 255 - 0xff
      11'h594: dout  = 8'b11111111; // 1428 : 255 - 0xff
      11'h595: dout  = 8'b11111111; // 1429 : 255 - 0xff
      11'h596: dout  = 8'b11111111; // 1430 : 255 - 0xff
      11'h597: dout  = 8'b11111111; // 1431 : 255 - 0xff
      11'h598: dout  = 8'b11111111; // 1432 : 255 - 0xff -- Sprite 0xb3
      11'h599: dout  = 8'b11111111; // 1433 : 255 - 0xff
      11'h59A: dout  = 8'b11111111; // 1434 : 255 - 0xff
      11'h59B: dout  = 8'b11111111; // 1435 : 255 - 0xff
      11'h59C: dout  = 8'b11111111; // 1436 : 255 - 0xff
      11'h59D: dout  = 8'b11111111; // 1437 : 255 - 0xff
      11'h59E: dout  = 8'b11111111; // 1438 : 255 - 0xff
      11'h59F: dout  = 8'b11111111; // 1439 : 255 - 0xff
      11'h5A0: dout  = 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0xb4
      11'h5A1: dout  = 8'b11111111; // 1441 : 255 - 0xff
      11'h5A2: dout  = 8'b11111111; // 1442 : 255 - 0xff
      11'h5A3: dout  = 8'b11111111; // 1443 : 255 - 0xff
      11'h5A4: dout  = 8'b11111111; // 1444 : 255 - 0xff
      11'h5A5: dout  = 8'b11111111; // 1445 : 255 - 0xff
      11'h5A6: dout  = 8'b11111111; // 1446 : 255 - 0xff
      11'h5A7: dout  = 8'b11111111; // 1447 : 255 - 0xff
      11'h5A8: dout  = 8'b11111111; // 1448 : 255 - 0xff -- Sprite 0xb5
      11'h5A9: dout  = 8'b11111111; // 1449 : 255 - 0xff
      11'h5AA: dout  = 8'b11111111; // 1450 : 255 - 0xff
      11'h5AB: dout  = 8'b11111111; // 1451 : 255 - 0xff
      11'h5AC: dout  = 8'b11111111; // 1452 : 255 - 0xff
      11'h5AD: dout  = 8'b11111111; // 1453 : 255 - 0xff
      11'h5AE: dout  = 8'b11111111; // 1454 : 255 - 0xff
      11'h5AF: dout  = 8'b11111111; // 1455 : 255 - 0xff
      11'h5B0: dout  = 8'b11111111; // 1456 : 255 - 0xff -- Sprite 0xb6
      11'h5B1: dout  = 8'b11111111; // 1457 : 255 - 0xff
      11'h5B2: dout  = 8'b11111111; // 1458 : 255 - 0xff
      11'h5B3: dout  = 8'b11111111; // 1459 : 255 - 0xff
      11'h5B4: dout  = 8'b11111111; // 1460 : 255 - 0xff
      11'h5B5: dout  = 8'b11111111; // 1461 : 255 - 0xff
      11'h5B6: dout  = 8'b11111111; // 1462 : 255 - 0xff
      11'h5B7: dout  = 8'b11111111; // 1463 : 255 - 0xff
      11'h5B8: dout  = 8'b11111111; // 1464 : 255 - 0xff -- Sprite 0xb7
      11'h5B9: dout  = 8'b11111111; // 1465 : 255 - 0xff
      11'h5BA: dout  = 8'b11111111; // 1466 : 255 - 0xff
      11'h5BB: dout  = 8'b11111111; // 1467 : 255 - 0xff
      11'h5BC: dout  = 8'b11111111; // 1468 : 255 - 0xff
      11'h5BD: dout  = 8'b11111111; // 1469 : 255 - 0xff
      11'h5BE: dout  = 8'b11111111; // 1470 : 255 - 0xff
      11'h5BF: dout  = 8'b11111111; // 1471 : 255 - 0xff
      11'h5C0: dout  = 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0xb8
      11'h5C1: dout  = 8'b00000111; // 1473 :   7 - 0x7
      11'h5C2: dout  = 8'b00001000; // 1474 :   8 - 0x8
      11'h5C3: dout  = 8'b00010000; // 1475 :  16 - 0x10
      11'h5C4: dout  = 8'b00010000; // 1476 :  16 - 0x10
      11'h5C5: dout  = 8'b00100000; // 1477 :  32 - 0x20
      11'h5C6: dout  = 8'b00100000; // 1478 :  32 - 0x20
      11'h5C7: dout  = 8'b00100000; // 1479 :  32 - 0x20
      11'h5C8: dout  = 8'b00011111; // 1480 :  31 - 0x1f -- Sprite 0xb9
      11'h5C9: dout  = 8'b00101111; // 1481 :  47 - 0x2f
      11'h5CA: dout  = 8'b00110111; // 1482 :  55 - 0x37
      11'h5CB: dout  = 8'b00111010; // 1483 :  58 - 0x3a
      11'h5CC: dout  = 8'b00111101; // 1484 :  61 - 0x3d
      11'h5CD: dout  = 8'b00111110; // 1485 :  62 - 0x3e
      11'h5CE: dout  = 8'b00111111; // 1486 :  63 - 0x3f
      11'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      11'h5D0: dout  = 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0xba
      11'h5D1: dout  = 8'b00000101; // 1489 :   5 - 0x5
      11'h5D2: dout  = 8'b00011001; // 1490 :  25 - 0x19
      11'h5D3: dout  = 8'b00110011; // 1491 :  51 - 0x33
      11'h5D4: dout  = 8'b01100011; // 1492 :  99 - 0x63
      11'h5D5: dout  = 8'b11000111; // 1493 : 199 - 0xc7
      11'h5D6: dout  = 8'b11000111; // 1494 : 199 - 0xc7
      11'h5D7: dout  = 8'b11000100; // 1495 : 196 - 0xc4
      11'h5D8: dout  = 8'b10000000; // 1496 : 128 - 0x80 -- Sprite 0xbb
      11'h5D9: dout  = 8'b00000000; // 1497 :   0 - 0x0
      11'h5DA: dout  = 8'b00000000; // 1498 :   0 - 0x0
      11'h5DB: dout  = 8'b00000000; // 1499 :   0 - 0x0
      11'h5DC: dout  = 8'b00000000; // 1500 :   0 - 0x0
      11'h5DD: dout  = 8'b00000011; // 1501 :   3 - 0x3
      11'h5DE: dout  = 8'b00000011; // 1502 :   3 - 0x3
      11'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      11'h5E0: dout  = 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0xbc
      11'h5E1: dout  = 8'b00000000; // 1505 :   0 - 0x0
      11'h5E2: dout  = 8'b00000000; // 1506 :   0 - 0x0
      11'h5E3: dout  = 8'b00000000; // 1507 :   0 - 0x0
      11'h5E4: dout  = 8'b00000000; // 1508 :   0 - 0x0
      11'h5E5: dout  = 8'b00000000; // 1509 :   0 - 0x0
      11'h5E6: dout  = 8'b00000000; // 1510 :   0 - 0x0
      11'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      11'h5E8: dout  = 8'b00000000; // 1512 :   0 - 0x0 -- Sprite 0xbd
      11'h5E9: dout  = 8'b00000000; // 1513 :   0 - 0x0
      11'h5EA: dout  = 8'b00001111; // 1514 :  15 - 0xf
      11'h5EB: dout  = 8'b00000000; // 1515 :   0 - 0x0
      11'h5EC: dout  = 8'b10000000; // 1516 : 128 - 0x80
      11'h5ED: dout  = 8'b01100011; // 1517 :  99 - 0x63
      11'h5EE: dout  = 8'b00011110; // 1518 :  30 - 0x1e
      11'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      11'h5F0: dout  = 8'b00000001; // 1520 :   1 - 0x1 -- Sprite 0xbe
      11'h5F1: dout  = 8'b00000011; // 1521 :   3 - 0x3
      11'h5F2: dout  = 8'b00011001; // 1522 :  25 - 0x19
      11'h5F3: dout  = 8'b00111100; // 1523 :  60 - 0x3c
      11'h5F4: dout  = 8'b00011001; // 1524 :  25 - 0x19
      11'h5F5: dout  = 8'b00100011; // 1525 :  35 - 0x23
      11'h5F6: dout  = 8'b01010001; // 1526 :  81 - 0x51
      11'h5F7: dout  = 8'b00100000; // 1527 :  32 - 0x20
      11'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      11'h5F9: dout  = 8'b00000000; // 1529 :   0 - 0x0
      11'h5FA: dout  = 8'b00000000; // 1530 :   0 - 0x0
      11'h5FB: dout  = 8'b00000000; // 1531 :   0 - 0x0
      11'h5FC: dout  = 8'b00000000; // 1532 :   0 - 0x0
      11'h5FD: dout  = 8'b00000000; // 1533 :   0 - 0x0
      11'h5FE: dout  = 8'b00000000; // 1534 :   0 - 0x0
      11'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      11'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      11'h601: dout  = 8'b00111111; // 1537 :  63 - 0x3f
      11'h602: dout  = 8'b00011111; // 1538 :  31 - 0x1f
      11'h603: dout  = 8'b00000000; // 1539 :   0 - 0x0
      11'h604: dout  = 8'b00000001; // 1540 :   1 - 0x1
      11'h605: dout  = 8'b00000000; // 1541 :   0 - 0x0
      11'h606: dout  = 8'b00000001; // 1542 :   1 - 0x1
      11'h607: dout  = 8'b00000000; // 1543 :   0 - 0x0
      11'h608: dout  = 8'b00010001; // 1544 :  17 - 0x11 -- Sprite 0xc1
      11'h609: dout  = 8'b00000000; // 1545 :   0 - 0x0
      11'h60A: dout  = 8'b00000001; // 1546 :   1 - 0x1
      11'h60B: dout  = 8'b00000000; // 1547 :   0 - 0x0
      11'h60C: dout  = 8'b00000001; // 1548 :   1 - 0x1
      11'h60D: dout  = 8'b00000000; // 1549 :   0 - 0x0
      11'h60E: dout  = 8'b00011111; // 1550 :  31 - 0x1f
      11'h60F: dout  = 8'b00111111; // 1551 :  63 - 0x3f
      11'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      11'h611: dout  = 8'b11111100; // 1553 : 252 - 0xfc
      11'h612: dout  = 8'b11111000; // 1554 : 248 - 0xf8
      11'h613: dout  = 8'b00000000; // 1555 :   0 - 0x0
      11'h614: dout  = 8'b10000000; // 1556 : 128 - 0x80
      11'h615: dout  = 8'b00000000; // 1557 :   0 - 0x0
      11'h616: dout  = 8'b10000000; // 1558 : 128 - 0x80
      11'h617: dout  = 8'b00000000; // 1559 :   0 - 0x0
      11'h618: dout  = 8'b10001000; // 1560 : 136 - 0x88 -- Sprite 0xc3
      11'h619: dout  = 8'b00000000; // 1561 :   0 - 0x0
      11'h61A: dout  = 8'b10000000; // 1562 : 128 - 0x80
      11'h61B: dout  = 8'b00000000; // 1563 :   0 - 0x0
      11'h61C: dout  = 8'b10000000; // 1564 : 128 - 0x80
      11'h61D: dout  = 8'b00000000; // 1565 :   0 - 0x0
      11'h61E: dout  = 8'b11111000; // 1566 : 248 - 0xf8
      11'h61F: dout  = 8'b11111100; // 1567 : 252 - 0xfc
      11'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      11'h621: dout  = 8'b00000000; // 1569 :   0 - 0x0
      11'h622: dout  = 8'b00000000; // 1570 :   0 - 0x0
      11'h623: dout  = 8'b00000000; // 1571 :   0 - 0x0
      11'h624: dout  = 8'b00000000; // 1572 :   0 - 0x0
      11'h625: dout  = 8'b00111111; // 1573 :  63 - 0x3f
      11'h626: dout  = 8'b00011111; // 1574 :  31 - 0x1f
      11'h627: dout  = 8'b00000000; // 1575 :   0 - 0x0
      11'h628: dout  = 8'b00000001; // 1576 :   1 - 0x1 -- Sprite 0xc5
      11'h629: dout  = 8'b00000001; // 1577 :   1 - 0x1
      11'h62A: dout  = 8'b01000001; // 1578 :  65 - 0x41
      11'h62B: dout  = 8'b00000001; // 1579 :   1 - 0x1
      11'h62C: dout  = 8'b00000001; // 1580 :   1 - 0x1
      11'h62D: dout  = 8'b00000000; // 1581 :   0 - 0x0
      11'h62E: dout  = 8'b00011111; // 1582 :  31 - 0x1f
      11'h62F: dout  = 8'b00111111; // 1583 :  63 - 0x3f
      11'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0xc6
      11'h631: dout  = 8'b00000000; // 1585 :   0 - 0x0
      11'h632: dout  = 8'b00000000; // 1586 :   0 - 0x0
      11'h633: dout  = 8'b00000000; // 1587 :   0 - 0x0
      11'h634: dout  = 8'b00000000; // 1588 :   0 - 0x0
      11'h635: dout  = 8'b11111100; // 1589 : 252 - 0xfc
      11'h636: dout  = 8'b11111000; // 1590 : 248 - 0xf8
      11'h637: dout  = 8'b00000000; // 1591 :   0 - 0x0
      11'h638: dout  = 8'b10000000; // 1592 : 128 - 0x80 -- Sprite 0xc7
      11'h639: dout  = 8'b10000000; // 1593 : 128 - 0x80
      11'h63A: dout  = 8'b10000010; // 1594 : 130 - 0x82
      11'h63B: dout  = 8'b10000000; // 1595 : 128 - 0x80
      11'h63C: dout  = 8'b10000000; // 1596 : 128 - 0x80
      11'h63D: dout  = 8'b00000000; // 1597 :   0 - 0x0
      11'h63E: dout  = 8'b11111000; // 1598 : 248 - 0xf8
      11'h63F: dout  = 8'b11111100; // 1599 : 252 - 0xfc
      11'h640: dout  = 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      11'h641: dout  = 8'b00000000; // 1601 :   0 - 0x0
      11'h642: dout  = 8'b00000000; // 1602 :   0 - 0x0
      11'h643: dout  = 8'b00011110; // 1603 :  30 - 0x1e
      11'h644: dout  = 8'b00111111; // 1604 :  63 - 0x3f
      11'h645: dout  = 8'b00111111; // 1605 :  63 - 0x3f
      11'h646: dout  = 8'b00111111; // 1606 :  63 - 0x3f
      11'h647: dout  = 8'b00111111; // 1607 :  63 - 0x3f
      11'h648: dout  = 8'b00011111; // 1608 :  31 - 0x1f -- Sprite 0xc9
      11'h649: dout  = 8'b00001111; // 1609 :  15 - 0xf
      11'h64A: dout  = 8'b00000111; // 1610 :   7 - 0x7
      11'h64B: dout  = 8'b00000011; // 1611 :   3 - 0x3
      11'h64C: dout  = 8'b00000001; // 1612 :   1 - 0x1
      11'h64D: dout  = 8'b00000000; // 1613 :   0 - 0x0
      11'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      11'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      11'h650: dout  = 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      11'h651: dout  = 8'b00000000; // 1617 :   0 - 0x0
      11'h652: dout  = 8'b00000000; // 1618 :   0 - 0x0
      11'h653: dout  = 8'b00111100; // 1619 :  60 - 0x3c
      11'h654: dout  = 8'b01111110; // 1620 : 126 - 0x7e
      11'h655: dout  = 8'b11111110; // 1621 : 254 - 0xfe
      11'h656: dout  = 8'b11111110; // 1622 : 254 - 0xfe
      11'h657: dout  = 8'b11111110; // 1623 : 254 - 0xfe
      11'h658: dout  = 8'b11111100; // 1624 : 252 - 0xfc -- Sprite 0xcb
      11'h659: dout  = 8'b11111000; // 1625 : 248 - 0xf8
      11'h65A: dout  = 8'b11110000; // 1626 : 240 - 0xf0
      11'h65B: dout  = 8'b11100000; // 1627 : 224 - 0xe0
      11'h65C: dout  = 8'b11000000; // 1628 : 192 - 0xc0
      11'h65D: dout  = 8'b10000000; // 1629 : 128 - 0x80
      11'h65E: dout  = 8'b00000000; // 1630 :   0 - 0x0
      11'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      11'h660: dout  = 8'b11111111; // 1632 : 255 - 0xff -- Sprite 0xcc
      11'h661: dout  = 8'b11111111; // 1633 : 255 - 0xff
      11'h662: dout  = 8'b11111111; // 1634 : 255 - 0xff
      11'h663: dout  = 8'b11111111; // 1635 : 255 - 0xff
      11'h664: dout  = 8'b11111111; // 1636 : 255 - 0xff
      11'h665: dout  = 8'b11111111; // 1637 : 255 - 0xff
      11'h666: dout  = 8'b11111111; // 1638 : 255 - 0xff
      11'h667: dout  = 8'b11111111; // 1639 : 255 - 0xff
      11'h668: dout  = 8'b11111111; // 1640 : 255 - 0xff -- Sprite 0xcd
      11'h669: dout  = 8'b11111111; // 1641 : 255 - 0xff
      11'h66A: dout  = 8'b11111111; // 1642 : 255 - 0xff
      11'h66B: dout  = 8'b11111111; // 1643 : 255 - 0xff
      11'h66C: dout  = 8'b11111111; // 1644 : 255 - 0xff
      11'h66D: dout  = 8'b11111111; // 1645 : 255 - 0xff
      11'h66E: dout  = 8'b11111111; // 1646 : 255 - 0xff
      11'h66F: dout  = 8'b11111111; // 1647 : 255 - 0xff
      11'h670: dout  = 8'b11111111; // 1648 : 255 - 0xff -- Sprite 0xce
      11'h671: dout  = 8'b11111111; // 1649 : 255 - 0xff
      11'h672: dout  = 8'b11111111; // 1650 : 255 - 0xff
      11'h673: dout  = 8'b11111111; // 1651 : 255 - 0xff
      11'h674: dout  = 8'b11111111; // 1652 : 255 - 0xff
      11'h675: dout  = 8'b11111111; // 1653 : 255 - 0xff
      11'h676: dout  = 8'b11111111; // 1654 : 255 - 0xff
      11'h677: dout  = 8'b11111111; // 1655 : 255 - 0xff
      11'h678: dout  = 8'b11111111; // 1656 : 255 - 0xff -- Sprite 0xcf
      11'h679: dout  = 8'b11111111; // 1657 : 255 - 0xff
      11'h67A: dout  = 8'b11111111; // 1658 : 255 - 0xff
      11'h67B: dout  = 8'b11111111; // 1659 : 255 - 0xff
      11'h67C: dout  = 8'b11111111; // 1660 : 255 - 0xff
      11'h67D: dout  = 8'b11111111; // 1661 : 255 - 0xff
      11'h67E: dout  = 8'b11111111; // 1662 : 255 - 0xff
      11'h67F: dout  = 8'b11111111; // 1663 : 255 - 0xff
      11'h680: dout  = 8'b00001000; // 1664 :   8 - 0x8 -- Sprite 0xd0
      11'h681: dout  = 8'b00011001; // 1665 :  25 - 0x19
      11'h682: dout  = 8'b00001001; // 1666 :   9 - 0x9
      11'h683: dout  = 8'b00001001; // 1667 :   9 - 0x9
      11'h684: dout  = 8'b00001001; // 1668 :   9 - 0x9
      11'h685: dout  = 8'b00001001; // 1669 :   9 - 0x9
      11'h686: dout  = 8'b00011100; // 1670 :  28 - 0x1c
      11'h687: dout  = 8'b00000000; // 1671 :   0 - 0x0
      11'h688: dout  = 8'b00111000; // 1672 :  56 - 0x38 -- Sprite 0xd1
      11'h689: dout  = 8'b00000101; // 1673 :   5 - 0x5
      11'h68A: dout  = 8'b00000101; // 1674 :   5 - 0x5
      11'h68B: dout  = 8'b00011001; // 1675 :  25 - 0x19
      11'h68C: dout  = 8'b00000101; // 1676 :   5 - 0x5
      11'h68D: dout  = 8'b00000101; // 1677 :   5 - 0x5
      11'h68E: dout  = 8'b00111000; // 1678 :  56 - 0x38
      11'h68F: dout  = 8'b00000000; // 1679 :   0 - 0x0
      11'h690: dout  = 8'b00111100; // 1680 :  60 - 0x3c -- Sprite 0xd2
      11'h691: dout  = 8'b00100001; // 1681 :  33 - 0x21
      11'h692: dout  = 8'b00100001; // 1682 :  33 - 0x21
      11'h693: dout  = 8'b00111101; // 1683 :  61 - 0x3d
      11'h694: dout  = 8'b00000101; // 1684 :   5 - 0x5
      11'h695: dout  = 8'b00000101; // 1685 :   5 - 0x5
      11'h696: dout  = 8'b00111000; // 1686 :  56 - 0x38
      11'h697: dout  = 8'b00000000; // 1687 :   0 - 0x0
      11'h698: dout  = 8'b00011000; // 1688 :  24 - 0x18 -- Sprite 0xd3
      11'h699: dout  = 8'b00100101; // 1689 :  37 - 0x25
      11'h69A: dout  = 8'b00100101; // 1690 :  37 - 0x25
      11'h69B: dout  = 8'b00011001; // 1691 :  25 - 0x19
      11'h69C: dout  = 8'b00100101; // 1692 :  37 - 0x25
      11'h69D: dout  = 8'b00100101; // 1693 :  37 - 0x25
      11'h69E: dout  = 8'b00011000; // 1694 :  24 - 0x18
      11'h69F: dout  = 8'b00000000; // 1695 :   0 - 0x0
      11'h6A0: dout  = 8'b11000110; // 1696 : 198 - 0xc6 -- Sprite 0xd4
      11'h6A1: dout  = 8'b00101001; // 1697 :  41 - 0x29
      11'h6A2: dout  = 8'b00101001; // 1698 :  41 - 0x29
      11'h6A3: dout  = 8'b00101001; // 1699 :  41 - 0x29
      11'h6A4: dout  = 8'b00101001; // 1700 :  41 - 0x29
      11'h6A5: dout  = 8'b00101001; // 1701 :  41 - 0x29
      11'h6A6: dout  = 8'b11000110; // 1702 : 198 - 0xc6
      11'h6A7: dout  = 8'b00000000; // 1703 :   0 - 0x0
      11'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0 -- Sprite 0xd5
      11'h6A9: dout  = 8'b00000000; // 1705 :   0 - 0x0
      11'h6AA: dout  = 8'b00000000; // 1706 :   0 - 0x0
      11'h6AB: dout  = 8'b00000000; // 1707 :   0 - 0x0
      11'h6AC: dout  = 8'b00000000; // 1708 :   0 - 0x0
      11'h6AD: dout  = 8'b00000000; // 1709 :   0 - 0x0
      11'h6AE: dout  = 8'b00000000; // 1710 :   0 - 0x0
      11'h6AF: dout  = 8'b00000000; // 1711 :   0 - 0x0
      11'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      11'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      11'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      11'h6B3: dout  = 8'b00000000; // 1715 :   0 - 0x0
      11'h6B4: dout  = 8'b00111100; // 1716 :  60 - 0x3c
      11'h6B5: dout  = 8'b10110110; // 1717 : 182 - 0xb6
      11'h6B6: dout  = 8'b01111100; // 1718 : 124 - 0x7c
      11'h6B7: dout  = 8'b11111000; // 1719 : 248 - 0xf8
      11'h6B8: dout  = 8'b00000011; // 1720 :   3 - 0x3 -- Sprite 0xd7
      11'h6B9: dout  = 8'b00000011; // 1721 :   3 - 0x3
      11'h6BA: dout  = 8'b00000011; // 1722 :   3 - 0x3
      11'h6BB: dout  = 8'b00000111; // 1723 :   7 - 0x7
      11'h6BC: dout  = 8'b00001100; // 1724 :  12 - 0xc
      11'h6BD: dout  = 8'b00011011; // 1725 :  27 - 0x1b
      11'h6BE: dout  = 8'b01110111; // 1726 : 119 - 0x77
      11'h6BF: dout  = 8'b00000111; // 1727 :   7 - 0x7
      11'h6C0: dout  = 8'b00001111; // 1728 :  15 - 0xf -- Sprite 0xd8
      11'h6C1: dout  = 8'b00001111; // 1729 :  15 - 0xf
      11'h6C2: dout  = 8'b00011111; // 1730 :  31 - 0x1f
      11'h6C3: dout  = 8'b00111111; // 1731 :  63 - 0x3f
      11'h6C4: dout  = 8'b01111111; // 1732 : 127 - 0x7f
      11'h6C5: dout  = 8'b00111111; // 1733 :  63 - 0x3f
      11'h6C6: dout  = 8'b00000000; // 1734 :   0 - 0x0
      11'h6C7: dout  = 8'b00000000; // 1735 :   0 - 0x0
      11'h6C8: dout  = 8'b11100000; // 1736 : 224 - 0xe0 -- Sprite 0xd9
      11'h6C9: dout  = 8'b11110000; // 1737 : 240 - 0xf0
      11'h6CA: dout  = 8'b11110000; // 1738 : 240 - 0xf0
      11'h6CB: dout  = 8'b11110000; // 1739 : 240 - 0xf0
      11'h6CC: dout  = 8'b00011000; // 1740 :  24 - 0x18
      11'h6CD: dout  = 8'b11111100; // 1741 : 252 - 0xfc
      11'h6CE: dout  = 8'b11111100; // 1742 : 252 - 0xfc
      11'h6CF: dout  = 8'b11111100; // 1743 : 252 - 0xfc
      11'h6D0: dout  = 8'b11111000; // 1744 : 248 - 0xf8 -- Sprite 0xda
      11'h6D1: dout  = 8'b11111100; // 1745 : 252 - 0xfc
      11'h6D2: dout  = 8'b11111111; // 1746 : 255 - 0xff
      11'h6D3: dout  = 8'b11111111; // 1747 : 255 - 0xff
      11'h6D4: dout  = 8'b11111110; // 1748 : 254 - 0xfe
      11'h6D5: dout  = 8'b11110000; // 1749 : 240 - 0xf0
      11'h6D6: dout  = 8'b00000000; // 1750 :   0 - 0x0
      11'h6D7: dout  = 8'b00000000; // 1751 :   0 - 0x0
      11'h6D8: dout  = 8'b00000011; // 1752 :   3 - 0x3 -- Sprite 0xdb
      11'h6D9: dout  = 8'b00000011; // 1753 :   3 - 0x3
      11'h6DA: dout  = 8'b00000011; // 1754 :   3 - 0x3
      11'h6DB: dout  = 8'b00000011; // 1755 :   3 - 0x3
      11'h6DC: dout  = 8'b00000001; // 1756 :   1 - 0x1
      11'h6DD: dout  = 8'b00000000; // 1757 :   0 - 0x0
      11'h6DE: dout  = 8'b00000111; // 1758 :   7 - 0x7
      11'h6DF: dout  = 8'b00011111; // 1759 :  31 - 0x1f
      11'h6E0: dout  = 8'b11111111; // 1760 : 255 - 0xff -- Sprite 0xdc
      11'h6E1: dout  = 8'b11111111; // 1761 : 255 - 0xff
      11'h6E2: dout  = 8'b01111111; // 1762 : 127 - 0x7f
      11'h6E3: dout  = 8'b00111111; // 1763 :  63 - 0x3f
      11'h6E4: dout  = 8'b00001111; // 1764 :  15 - 0xf
      11'h6E5: dout  = 8'b00000011; // 1765 :   3 - 0x3
      11'h6E6: dout  = 8'b00000000; // 1766 :   0 - 0x0
      11'h6E7: dout  = 8'b00000000; // 1767 :   0 - 0x0
      11'h6E8: dout  = 8'b11100000; // 1768 : 224 - 0xe0 -- Sprite 0xdd
      11'h6E9: dout  = 8'b11110000; // 1769 : 240 - 0xf0
      11'h6EA: dout  = 8'b11110000; // 1770 : 240 - 0xf0
      11'h6EB: dout  = 8'b11100000; // 1771 : 224 - 0xe0
      11'h6EC: dout  = 8'b11111110; // 1772 : 254 - 0xfe
      11'h6ED: dout  = 8'b00111100; // 1773 :  60 - 0x3c
      11'h6EE: dout  = 8'b11110000; // 1774 : 240 - 0xf0
      11'h6EF: dout  = 8'b11111100; // 1775 : 252 - 0xfc
      11'h6F0: dout  = 8'b11111100; // 1776 : 252 - 0xfc -- Sprite 0xde
      11'h6F1: dout  = 8'b11111000; // 1777 : 248 - 0xf8
      11'h6F2: dout  = 8'b11111000; // 1778 : 248 - 0xf8
      11'h6F3: dout  = 8'b11111000; // 1779 : 248 - 0xf8
      11'h6F4: dout  = 8'b11111000; // 1780 : 248 - 0xf8
      11'h6F5: dout  = 8'b11111000; // 1781 : 248 - 0xf8
      11'h6F6: dout  = 8'b11111000; // 1782 : 248 - 0xf8
      11'h6F7: dout  = 8'b00000000; // 1783 :   0 - 0x0
      11'h6F8: dout  = 8'b11111111; // 1784 : 255 - 0xff -- Sprite 0xdf
      11'h6F9: dout  = 8'b11111111; // 1785 : 255 - 0xff
      11'h6FA: dout  = 8'b11111111; // 1786 : 255 - 0xff
      11'h6FB: dout  = 8'b11111111; // 1787 : 255 - 0xff
      11'h6FC: dout  = 8'b11111111; // 1788 : 255 - 0xff
      11'h6FD: dout  = 8'b11111111; // 1789 : 255 - 0xff
      11'h6FE: dout  = 8'b11111111; // 1790 : 255 - 0xff
      11'h6FF: dout  = 8'b11111111; // 1791 : 255 - 0xff
      11'h700: dout  = 8'b11111111; // 1792 : 255 - 0xff -- Sprite 0xe0
      11'h701: dout  = 8'b11111111; // 1793 : 255 - 0xff
      11'h702: dout  = 8'b11111111; // 1794 : 255 - 0xff
      11'h703: dout  = 8'b11111111; // 1795 : 255 - 0xff
      11'h704: dout  = 8'b11111111; // 1796 : 255 - 0xff
      11'h705: dout  = 8'b11111111; // 1797 : 255 - 0xff
      11'h706: dout  = 8'b11111111; // 1798 : 255 - 0xff
      11'h707: dout  = 8'b11111111; // 1799 : 255 - 0xff
      11'h708: dout  = 8'b11111111; // 1800 : 255 - 0xff -- Sprite 0xe1
      11'h709: dout  = 8'b11111111; // 1801 : 255 - 0xff
      11'h70A: dout  = 8'b11111111; // 1802 : 255 - 0xff
      11'h70B: dout  = 8'b11111111; // 1803 : 255 - 0xff
      11'h70C: dout  = 8'b11111111; // 1804 : 255 - 0xff
      11'h70D: dout  = 8'b11111111; // 1805 : 255 - 0xff
      11'h70E: dout  = 8'b11111111; // 1806 : 255 - 0xff
      11'h70F: dout  = 8'b11111111; // 1807 : 255 - 0xff
      11'h710: dout  = 8'b11111111; // 1808 : 255 - 0xff -- Sprite 0xe2
      11'h711: dout  = 8'b11111111; // 1809 : 255 - 0xff
      11'h712: dout  = 8'b11111111; // 1810 : 255 - 0xff
      11'h713: dout  = 8'b11111111; // 1811 : 255 - 0xff
      11'h714: dout  = 8'b11111111; // 1812 : 255 - 0xff
      11'h715: dout  = 8'b11111111; // 1813 : 255 - 0xff
      11'h716: dout  = 8'b11111111; // 1814 : 255 - 0xff
      11'h717: dout  = 8'b11111111; // 1815 : 255 - 0xff
      11'h718: dout  = 8'b11111111; // 1816 : 255 - 0xff -- Sprite 0xe3
      11'h719: dout  = 8'b11111111; // 1817 : 255 - 0xff
      11'h71A: dout  = 8'b11111111; // 1818 : 255 - 0xff
      11'h71B: dout  = 8'b11111111; // 1819 : 255 - 0xff
      11'h71C: dout  = 8'b11111111; // 1820 : 255 - 0xff
      11'h71D: dout  = 8'b11111111; // 1821 : 255 - 0xff
      11'h71E: dout  = 8'b11111111; // 1822 : 255 - 0xff
      11'h71F: dout  = 8'b11111111; // 1823 : 255 - 0xff
      11'h720: dout  = 8'b11111111; // 1824 : 255 - 0xff -- Sprite 0xe4
      11'h721: dout  = 8'b11111111; // 1825 : 255 - 0xff
      11'h722: dout  = 8'b11111111; // 1826 : 255 - 0xff
      11'h723: dout  = 8'b11111111; // 1827 : 255 - 0xff
      11'h724: dout  = 8'b11111111; // 1828 : 255 - 0xff
      11'h725: dout  = 8'b11111111; // 1829 : 255 - 0xff
      11'h726: dout  = 8'b11111111; // 1830 : 255 - 0xff
      11'h727: dout  = 8'b11111111; // 1831 : 255 - 0xff
      11'h728: dout  = 8'b11111111; // 1832 : 255 - 0xff -- Sprite 0xe5
      11'h729: dout  = 8'b11111111; // 1833 : 255 - 0xff
      11'h72A: dout  = 8'b11111111; // 1834 : 255 - 0xff
      11'h72B: dout  = 8'b11111111; // 1835 : 255 - 0xff
      11'h72C: dout  = 8'b11111111; // 1836 : 255 - 0xff
      11'h72D: dout  = 8'b11111111; // 1837 : 255 - 0xff
      11'h72E: dout  = 8'b11111111; // 1838 : 255 - 0xff
      11'h72F: dout  = 8'b11111111; // 1839 : 255 - 0xff
      11'h730: dout  = 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0xe6
      11'h731: dout  = 8'b11111111; // 1841 : 255 - 0xff
      11'h732: dout  = 8'b11111111; // 1842 : 255 - 0xff
      11'h733: dout  = 8'b11111111; // 1843 : 255 - 0xff
      11'h734: dout  = 8'b11111111; // 1844 : 255 - 0xff
      11'h735: dout  = 8'b11111111; // 1845 : 255 - 0xff
      11'h736: dout  = 8'b11111111; // 1846 : 255 - 0xff
      11'h737: dout  = 8'b11111111; // 1847 : 255 - 0xff
      11'h738: dout  = 8'b11111111; // 1848 : 255 - 0xff -- Sprite 0xe7
      11'h739: dout  = 8'b11111111; // 1849 : 255 - 0xff
      11'h73A: dout  = 8'b11111111; // 1850 : 255 - 0xff
      11'h73B: dout  = 8'b11111111; // 1851 : 255 - 0xff
      11'h73C: dout  = 8'b11111111; // 1852 : 255 - 0xff
      11'h73D: dout  = 8'b11111111; // 1853 : 255 - 0xff
      11'h73E: dout  = 8'b11111111; // 1854 : 255 - 0xff
      11'h73F: dout  = 8'b11111111; // 1855 : 255 - 0xff
      11'h740: dout  = 8'b11111111; // 1856 : 255 - 0xff -- Sprite 0xe8
      11'h741: dout  = 8'b11111111; // 1857 : 255 - 0xff
      11'h742: dout  = 8'b11111111; // 1858 : 255 - 0xff
      11'h743: dout  = 8'b11111111; // 1859 : 255 - 0xff
      11'h744: dout  = 8'b11111111; // 1860 : 255 - 0xff
      11'h745: dout  = 8'b11111111; // 1861 : 255 - 0xff
      11'h746: dout  = 8'b11111111; // 1862 : 255 - 0xff
      11'h747: dout  = 8'b11111111; // 1863 : 255 - 0xff
      11'h748: dout  = 8'b11111111; // 1864 : 255 - 0xff -- Sprite 0xe9
      11'h749: dout  = 8'b11111111; // 1865 : 255 - 0xff
      11'h74A: dout  = 8'b11111111; // 1866 : 255 - 0xff
      11'h74B: dout  = 8'b11111111; // 1867 : 255 - 0xff
      11'h74C: dout  = 8'b11111111; // 1868 : 255 - 0xff
      11'h74D: dout  = 8'b11111111; // 1869 : 255 - 0xff
      11'h74E: dout  = 8'b11111111; // 1870 : 255 - 0xff
      11'h74F: dout  = 8'b11111111; // 1871 : 255 - 0xff
      11'h750: dout  = 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0xea
      11'h751: dout  = 8'b11111111; // 1873 : 255 - 0xff
      11'h752: dout  = 8'b11111111; // 1874 : 255 - 0xff
      11'h753: dout  = 8'b11111111; // 1875 : 255 - 0xff
      11'h754: dout  = 8'b11111111; // 1876 : 255 - 0xff
      11'h755: dout  = 8'b11111111; // 1877 : 255 - 0xff
      11'h756: dout  = 8'b11111111; // 1878 : 255 - 0xff
      11'h757: dout  = 8'b11111111; // 1879 : 255 - 0xff
      11'h758: dout  = 8'b11111111; // 1880 : 255 - 0xff -- Sprite 0xeb
      11'h759: dout  = 8'b11111111; // 1881 : 255 - 0xff
      11'h75A: dout  = 8'b11111111; // 1882 : 255 - 0xff
      11'h75B: dout  = 8'b11111111; // 1883 : 255 - 0xff
      11'h75C: dout  = 8'b11111111; // 1884 : 255 - 0xff
      11'h75D: dout  = 8'b11111111; // 1885 : 255 - 0xff
      11'h75E: dout  = 8'b11111111; // 1886 : 255 - 0xff
      11'h75F: dout  = 8'b11111111; // 1887 : 255 - 0xff
      11'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      11'h761: dout  = 8'b00000001; // 1889 :   1 - 0x1
      11'h762: dout  = 8'b00000011; // 1890 :   3 - 0x3
      11'h763: dout  = 8'b00110011; // 1891 :  51 - 0x33
      11'h764: dout  = 8'b00011001; // 1892 :  25 - 0x19
      11'h765: dout  = 8'b00001111; // 1893 :  15 - 0xf
      11'h766: dout  = 8'b00111111; // 1894 :  63 - 0x3f
      11'h767: dout  = 8'b00011111; // 1895 :  31 - 0x1f
      11'h768: dout  = 8'b00101011; // 1896 :  43 - 0x2b -- Sprite 0xed
      11'h769: dout  = 8'b00000111; // 1897 :   7 - 0x7
      11'h76A: dout  = 8'b00000101; // 1898 :   5 - 0x5
      11'h76B: dout  = 8'b00001101; // 1899 :  13 - 0xd
      11'h76C: dout  = 8'b00001011; // 1900 :  11 - 0xb
      11'h76D: dout  = 8'b00011011; // 1901 :  27 - 0x1b
      11'h76E: dout  = 8'b00011011; // 1902 :  27 - 0x1b
      11'h76F: dout  = 8'b00111011; // 1903 :  59 - 0x3b
      11'h770: dout  = 8'b00001001; // 1904 :   9 - 0x9 -- Sprite 0xee
      11'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      11'h772: dout  = 8'b00000111; // 1906 :   7 - 0x7
      11'h773: dout  = 8'b00000111; // 1907 :   7 - 0x7
      11'h774: dout  = 8'b00001111; // 1908 :  15 - 0xf
      11'h775: dout  = 8'b00001101; // 1909 :  13 - 0xd
      11'h776: dout  = 8'b00000001; // 1910 :   1 - 0x1
      11'h777: dout  = 8'b00000000; // 1911 :   0 - 0x0
      11'h778: dout  = 8'b11111000; // 1912 : 248 - 0xf8 -- Sprite 0xef
      11'h779: dout  = 8'b11111100; // 1913 : 252 - 0xfc
      11'h77A: dout  = 8'b11111000; // 1914 : 248 - 0xf8
      11'h77B: dout  = 8'b11101100; // 1915 : 236 - 0xec
      11'h77C: dout  = 8'b11111000; // 1916 : 248 - 0xf8
      11'h77D: dout  = 8'b11110000; // 1917 : 240 - 0xf0
      11'h77E: dout  = 8'b11000000; // 1918 : 192 - 0xc0
      11'h77F: dout  = 8'b11000000; // 1919 : 192 - 0xc0
      11'h780: dout  = 8'b11110000; // 1920 : 240 - 0xf0 -- Sprite 0xf0
      11'h781: dout  = 8'b11111000; // 1921 : 248 - 0xf8
      11'h782: dout  = 8'b11111000; // 1922 : 248 - 0xf8
      11'h783: dout  = 8'b11101000; // 1923 : 232 - 0xe8
      11'h784: dout  = 8'b11001100; // 1924 : 204 - 0xcc
      11'h785: dout  = 8'b11100110; // 1925 : 230 - 0xe6
      11'h786: dout  = 8'b11111011; // 1926 : 251 - 0xfb
      11'h787: dout  = 8'b11111111; // 1927 : 255 - 0xff
      11'h788: dout  = 8'b11111111; // 1928 : 255 - 0xff -- Sprite 0xf1
      11'h789: dout  = 8'b11111110; // 1929 : 254 - 0xfe
      11'h78A: dout  = 8'b11111110; // 1930 : 254 - 0xfe
      11'h78B: dout  = 8'b11111110; // 1931 : 254 - 0xfe
      11'h78C: dout  = 8'b11111110; // 1932 : 254 - 0xfe
      11'h78D: dout  = 8'b10001111; // 1933 : 143 - 0x8f
      11'h78E: dout  = 8'b00000000; // 1934 :   0 - 0x0
      11'h78F: dout  = 8'b00000000; // 1935 :   0 - 0x0
      11'h790: dout  = 8'b00000001; // 1936 :   1 - 0x1 -- Sprite 0xf2
      11'h791: dout  = 8'b00001111; // 1937 :  15 - 0xf
      11'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      11'h793: dout  = 8'b00000000; // 1939 :   0 - 0x0
      11'h794: dout  = 8'b00000100; // 1940 :   4 - 0x4
      11'h795: dout  = 8'b00011110; // 1941 :  30 - 0x1e
      11'h796: dout  = 8'b00000000; // 1942 :   0 - 0x0
      11'h797: dout  = 8'b00000011; // 1943 :   3 - 0x3
      11'h798: dout  = 8'b00000111; // 1944 :   7 - 0x7 -- Sprite 0xf3
      11'h799: dout  = 8'b00001111; // 1945 :  15 - 0xf
      11'h79A: dout  = 8'b00011111; // 1946 :  31 - 0x1f
      11'h79B: dout  = 8'b00001111; // 1947 :  15 - 0xf
      11'h79C: dout  = 8'b00000111; // 1948 :   7 - 0x7
      11'h79D: dout  = 8'b00001111; // 1949 :  15 - 0xf
      11'h79E: dout  = 8'b00001111; // 1950 :  15 - 0xf
      11'h79F: dout  = 8'b00000011; // 1951 :   3 - 0x3
      11'h7A0: dout  = 8'b11100000; // 1952 : 224 - 0xe0 -- Sprite 0xf4
      11'h7A1: dout  = 8'b11110000; // 1953 : 240 - 0xf0
      11'h7A2: dout  = 8'b11110000; // 1954 : 240 - 0xf0
      11'h7A3: dout  = 8'b01001000; // 1955 :  72 - 0x48
      11'h7A4: dout  = 8'b11001000; // 1956 : 200 - 0xc8
      11'h7A5: dout  = 8'b10011100; // 1957 : 156 - 0x9c
      11'h7A6: dout  = 8'b00000000; // 1958 :   0 - 0x0
      11'h7A7: dout  = 8'b11110000; // 1959 : 240 - 0xf0
      11'h7A8: dout  = 8'b11111000; // 1960 : 248 - 0xf8 -- Sprite 0xf5
      11'h7A9: dout  = 8'b11111100; // 1961 : 252 - 0xfc
      11'h7AA: dout  = 8'b11111100; // 1962 : 252 - 0xfc
      11'h7AB: dout  = 8'b11111000; // 1963 : 248 - 0xf8
      11'h7AC: dout  = 8'b11111000; // 1964 : 248 - 0xf8
      11'h7AD: dout  = 8'b01111000; // 1965 : 120 - 0x78
      11'h7AE: dout  = 8'b01110000; // 1966 : 112 - 0x70
      11'h7AF: dout  = 8'b01100000; // 1967 :  96 - 0x60
      11'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      11'h7B1: dout  = 8'b00000000; // 1969 :   0 - 0x0
      11'h7B2: dout  = 8'b01111100; // 1970 : 124 - 0x7c
      11'h7B3: dout  = 8'b10001010; // 1971 : 138 - 0x8a
      11'h7B4: dout  = 8'b11111110; // 1972 : 254 - 0xfe
      11'h7B5: dout  = 8'b11111110; // 1973 : 254 - 0xfe
      11'h7B6: dout  = 8'b11111110; // 1974 : 254 - 0xfe
      11'h7B7: dout  = 8'b11111110; // 1975 : 254 - 0xfe
      11'h7B8: dout  = 8'b11111110; // 1976 : 254 - 0xfe -- Sprite 0xf7
      11'h7B9: dout  = 8'b01111100; // 1977 : 124 - 0x7c
      11'h7BA: dout  = 8'b00000000; // 1978 :   0 - 0x0
      11'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      11'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      11'h7BD: dout  = 8'b00000000; // 1981 :   0 - 0x0
      11'h7BE: dout  = 8'b00000000; // 1982 :   0 - 0x0
      11'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      11'h7C0: dout  = 8'b00000111; // 1984 :   7 - 0x7 -- Sprite 0xf8
      11'h7C1: dout  = 8'b00001011; // 1985 :  11 - 0xb
      11'h7C2: dout  = 8'b00001111; // 1986 :  15 - 0xf
      11'h7C3: dout  = 8'b00001011; // 1987 :  11 - 0xb
      11'h7C4: dout  = 8'b00001011; // 1988 :  11 - 0xb
      11'h7C5: dout  = 8'b00001011; // 1989 :  11 - 0xb
      11'h7C6: dout  = 8'b00001011; // 1990 :  11 - 0xb
      11'h7C7: dout  = 8'b00000111; // 1991 :   7 - 0x7
      11'h7C8: dout  = 8'b11000000; // 1992 : 192 - 0xc0 -- Sprite 0xf9
      11'h7C9: dout  = 8'b11100000; // 1993 : 224 - 0xe0
      11'h7CA: dout  = 8'b11100000; // 1994 : 224 - 0xe0
      11'h7CB: dout  = 8'b11100000; // 1995 : 224 - 0xe0
      11'h7CC: dout  = 8'b11100000; // 1996 : 224 - 0xe0
      11'h7CD: dout  = 8'b11100000; // 1997 : 224 - 0xe0
      11'h7CE: dout  = 8'b11100000; // 1998 : 224 - 0xe0
      11'h7CF: dout  = 8'b11000000; // 1999 : 192 - 0xc0
      11'h7D0: dout  = 8'b00000011; // 2000 :   3 - 0x3 -- Sprite 0xfa
      11'h7D1: dout  = 8'b00000111; // 2001 :   7 - 0x7
      11'h7D2: dout  = 8'b00000111; // 2002 :   7 - 0x7
      11'h7D3: dout  = 8'b00000111; // 2003 :   7 - 0x7
      11'h7D4: dout  = 8'b00000111; // 2004 :   7 - 0x7
      11'h7D5: dout  = 8'b00000111; // 2005 :   7 - 0x7
      11'h7D6: dout  = 8'b00000111; // 2006 :   7 - 0x7
      11'h7D7: dout  = 8'b00000011; // 2007 :   3 - 0x3
      11'h7D8: dout  = 8'b11100000; // 2008 : 224 - 0xe0 -- Sprite 0xfb
      11'h7D9: dout  = 8'b11010000; // 2009 : 208 - 0xd0
      11'h7DA: dout  = 8'b11010000; // 2010 : 208 - 0xd0
      11'h7DB: dout  = 8'b11010000; // 2011 : 208 - 0xd0
      11'h7DC: dout  = 8'b11010000; // 2012 : 208 - 0xd0
      11'h7DD: dout  = 8'b11110000; // 2013 : 240 - 0xf0
      11'h7DE: dout  = 8'b11010000; // 2014 : 208 - 0xd0
      11'h7DF: dout  = 8'b11100000; // 2015 : 224 - 0xe0
      11'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      11'h7E1: dout  = 8'b00000001; // 2017 :   1 - 0x1
      11'h7E2: dout  = 8'b00010011; // 2018 :  19 - 0x13
      11'h7E3: dout  = 8'b00110111; // 2019 :  55 - 0x37
      11'h7E4: dout  = 8'b00111011; // 2020 :  59 - 0x3b
      11'h7E5: dout  = 8'b01110100; // 2021 : 116 - 0x74
      11'h7E6: dout  = 8'b01111010; // 2022 : 122 - 0x7a
      11'h7E7: dout  = 8'b00111110; // 2023 :  62 - 0x3e
      11'h7E8: dout  = 8'b11011000; // 2024 : 216 - 0xd8 -- Sprite 0xfd
      11'h7E9: dout  = 8'b10011000; // 2025 : 152 - 0x98
      11'h7EA: dout  = 8'b10101000; // 2026 : 168 - 0xa8
      11'h7EB: dout  = 8'b11011000; // 2027 : 216 - 0xd8
      11'h7EC: dout  = 8'b11011010; // 2028 : 218 - 0xda
      11'h7ED: dout  = 8'b01110100; // 2029 : 116 - 0x74
      11'h7EE: dout  = 8'b00101000; // 2030 :  40 - 0x28
      11'h7EF: dout  = 8'b11001000; // 2031 : 200 - 0xc8
      11'h7F0: dout  = 8'b00001000; // 2032 :   8 - 0x8 -- Sprite 0xfe
      11'h7F1: dout  = 8'b01011001; // 2033 :  89 - 0x59
      11'h7F2: dout  = 8'b00110000; // 2034 :  48 - 0x30
      11'h7F3: dout  = 8'b01110001; // 2035 : 113 - 0x71
      11'h7F4: dout  = 8'b01111001; // 2036 : 121 - 0x79
      11'h7F5: dout  = 8'b00101011; // 2037 :  43 - 0x2b
      11'h7F6: dout  = 8'b00110110; // 2038 :  54 - 0x36
      11'h7F7: dout  = 8'b00010110; // 2039 :  22 - 0x16
      11'h7F8: dout  = 8'b11000110; // 2040 : 198 - 0xc6 -- Sprite 0xff
      11'h7F9: dout  = 8'b11000100; // 2041 : 196 - 0xc4
      11'h7FA: dout  = 8'b11001100; // 2042 : 204 - 0xcc
      11'h7FB: dout  = 8'b11001100; // 2043 : 204 - 0xcc
      11'h7FC: dout  = 8'b10111000; // 2044 : 184 - 0xb8
      11'h7FD: dout  = 8'b01111100; // 2045 : 124 - 0x7c
      11'h7FE: dout  = 8'b11101100; // 2046 : 236 - 0xec
      11'h7FF: dout  = 8'b11001000; // 2047 : 200 - 0xc8
    endcase
  end

endmodule
