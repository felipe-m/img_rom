//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: lawnmower_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_LAWN_color1
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout <= 8'b00000000; //    1 :   0 - 0x0
      12'h2: dout <= 8'b00000000; //    2 :   0 - 0x0
      12'h3: dout <= 8'b00000000; //    3 :   0 - 0x0
      12'h4: dout <= 8'b00000000; //    4 :   0 - 0x0
      12'h5: dout <= 8'b00000000; //    5 :   0 - 0x0
      12'h6: dout <= 8'b00000000; //    6 :   0 - 0x0
      12'h7: dout <= 8'b00000000; //    7 :   0 - 0x0
      12'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      12'h9: dout <= 8'b00000000; //    9 :   0 - 0x0
      12'hA: dout <= 8'b00000000; //   10 :   0 - 0x0
      12'hB: dout <= 8'b00000000; //   11 :   0 - 0x0
      12'hC: dout <= 8'b00000000; //   12 :   0 - 0x0
      12'hD: dout <= 8'b00000111; //   13 :   7 - 0x7
      12'hE: dout <= 8'b00000111; //   14 :   7 - 0x7
      12'hF: dout <= 8'b00000110; //   15 :   6 - 0x6
      12'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x2
      12'h11: dout <= 8'b00000000; //   17 :   0 - 0x0
      12'h12: dout <= 8'b00000000; //   18 :   0 - 0x0
      12'h13: dout <= 8'b00000000; //   19 :   0 - 0x0
      12'h14: dout <= 8'b00000000; //   20 :   0 - 0x0
      12'h15: dout <= 8'b11111111; //   21 : 255 - 0xff
      12'h16: dout <= 8'b11111111; //   22 : 255 - 0xff
      12'h17: dout <= 8'b00000000; //   23 :   0 - 0x0
      12'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- Sprite 0x3
      12'h19: dout <= 8'b00000000; //   25 :   0 - 0x0
      12'h1A: dout <= 8'b00000000; //   26 :   0 - 0x0
      12'h1B: dout <= 8'b00000000; //   27 :   0 - 0x0
      12'h1C: dout <= 8'b00000000; //   28 :   0 - 0x0
      12'h1D: dout <= 8'b11100000; //   29 : 224 - 0xe0
      12'h1E: dout <= 8'b11100000; //   30 : 224 - 0xe0
      12'h1F: dout <= 8'b01100000; //   31 :  96 - 0x60
      12'h20: dout <= 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x4
      12'h21: dout <= 8'b00000000; //   33 :   0 - 0x0
      12'h22: dout <= 8'b00000000; //   34 :   0 - 0x0
      12'h23: dout <= 8'b00000000; //   35 :   0 - 0x0
      12'h24: dout <= 8'b00000000; //   36 :   0 - 0x0
      12'h25: dout <= 8'b00011111; //   37 :  31 - 0x1f
      12'h26: dout <= 8'b01111111; //   38 : 127 - 0x7f
      12'h27: dout <= 8'b11110000; //   39 : 240 - 0xf0
      12'h28: dout <= 8'b00000000; //   40 :   0 - 0x0 -- Sprite 0x5
      12'h29: dout <= 8'b00000000; //   41 :   0 - 0x0
      12'h2A: dout <= 8'b00000000; //   42 :   0 - 0x0
      12'h2B: dout <= 8'b00000000; //   43 :   0 - 0x0
      12'h2C: dout <= 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout <= 8'b11111000; //   45 : 248 - 0xf8
      12'h2E: dout <= 8'b11111110; //   46 : 254 - 0xfe
      12'h2F: dout <= 8'b00001111; //   47 :  15 - 0xf
      12'h30: dout <= 8'b00000000; //   48 :   0 - 0x0 -- Sprite 0x6
      12'h31: dout <= 8'b00000000; //   49 :   0 - 0x0
      12'h32: dout <= 8'b00000000; //   50 :   0 - 0x0
      12'h33: dout <= 8'b00000000; //   51 :   0 - 0x0
      12'h34: dout <= 8'b00000000; //   52 :   0 - 0x0
      12'h35: dout <= 8'b11100111; //   53 : 231 - 0xe7
      12'h36: dout <= 8'b11100111; //   54 : 231 - 0xe7
      12'h37: dout <= 8'b01100110; //   55 : 102 - 0x66
      12'h38: dout <= 8'b00000000; //   56 :   0 - 0x0 -- Sprite 0x7
      12'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      12'h3A: dout <= 8'b00000000; //   58 :   0 - 0x0
      12'h3B: dout <= 8'b00000000; //   59 :   0 - 0x0
      12'h3C: dout <= 8'b00000000; //   60 :   0 - 0x0
      12'h3D: dout <= 8'b11000111; //   61 : 199 - 0xc7
      12'h3E: dout <= 8'b11000111; //   62 : 199 - 0xc7
      12'h3F: dout <= 8'b01100110; //   63 : 102 - 0x66
      12'h40: dout <= 8'b00000110; //   64 :   6 - 0x6 -- Sprite 0x8
      12'h41: dout <= 8'b00000110; //   65 :   6 - 0x6
      12'h42: dout <= 8'b00000110; //   66 :   6 - 0x6
      12'h43: dout <= 8'b00000110; //   67 :   6 - 0x6
      12'h44: dout <= 8'b00000110; //   68 :   6 - 0x6
      12'h45: dout <= 8'b00000110; //   69 :   6 - 0x6
      12'h46: dout <= 8'b00000110; //   70 :   6 - 0x6
      12'h47: dout <= 8'b00000110; //   71 :   6 - 0x6
      12'h48: dout <= 8'b11111111; //   72 : 255 - 0xff -- Sprite 0x9
      12'h49: dout <= 8'b11111111; //   73 : 255 - 0xff
      12'h4A: dout <= 8'b11111111; //   74 : 255 - 0xff
      12'h4B: dout <= 8'b11111111; //   75 : 255 - 0xff
      12'h4C: dout <= 8'b11111111; //   76 : 255 - 0xff
      12'h4D: dout <= 8'b11111111; //   77 : 255 - 0xff
      12'h4E: dout <= 8'b11111111; //   78 : 255 - 0xff
      12'h4F: dout <= 8'b11111111; //   79 : 255 - 0xff
      12'h50: dout <= 8'b01100000; //   80 :  96 - 0x60 -- Sprite 0xa
      12'h51: dout <= 8'b01100000; //   81 :  96 - 0x60
      12'h52: dout <= 8'b01100000; //   82 :  96 - 0x60
      12'h53: dout <= 8'b01100000; //   83 :  96 - 0x60
      12'h54: dout <= 8'b01100000; //   84 :  96 - 0x60
      12'h55: dout <= 8'b01100000; //   85 :  96 - 0x60
      12'h56: dout <= 8'b01100000; //   86 :  96 - 0x60
      12'h57: dout <= 8'b01100000; //   87 :  96 - 0x60
      12'h58: dout <= 8'b00000001; //   88 :   1 - 0x1 -- Sprite 0xb
      12'h59: dout <= 8'b00000011; //   89 :   3 - 0x3
      12'h5A: dout <= 8'b00000011; //   90 :   3 - 0x3
      12'h5B: dout <= 8'b00000111; //   91 :   7 - 0x7
      12'h5C: dout <= 8'b00000110; //   92 :   6 - 0x6
      12'h5D: dout <= 8'b00000110; //   93 :   6 - 0x6
      12'h5E: dout <= 8'b00000110; //   94 :   6 - 0x6
      12'h5F: dout <= 8'b00000110; //   95 :   6 - 0x6
      12'h60: dout <= 8'b11000111; //   96 : 199 - 0xc7 -- Sprite 0xc
      12'h61: dout <= 8'b10011111; //   97 : 159 - 0x9f
      12'h62: dout <= 8'b00111111; //   98 :  63 - 0x3f
      12'h63: dout <= 8'b01111111; //   99 : 127 - 0x7f
      12'h64: dout <= 8'b01111111; //  100 : 127 - 0x7f
      12'h65: dout <= 8'b11111111; //  101 : 255 - 0xff
      12'h66: dout <= 8'b11111111; //  102 : 255 - 0xff
      12'h67: dout <= 8'b11111111; //  103 : 255 - 0xff
      12'h68: dout <= 8'b11100011; //  104 : 227 - 0xe3 -- Sprite 0xd
      12'h69: dout <= 8'b11111001; //  105 : 249 - 0xf9
      12'h6A: dout <= 8'b11111100; //  106 : 252 - 0xfc
      12'h6B: dout <= 8'b11111110; //  107 : 254 - 0xfe
      12'h6C: dout <= 8'b11111110; //  108 : 254 - 0xfe
      12'h6D: dout <= 8'b11111111; //  109 : 255 - 0xff
      12'h6E: dout <= 8'b11111111; //  110 : 255 - 0xff
      12'h6F: dout <= 8'b11111111; //  111 : 255 - 0xff
      12'h70: dout <= 8'b10000110; //  112 : 134 - 0x86 -- Sprite 0xe
      12'h71: dout <= 8'b11000110; //  113 : 198 - 0xc6
      12'h72: dout <= 8'b11000110; //  114 : 198 - 0xc6
      12'h73: dout <= 8'b11100110; //  115 : 230 - 0xe6
      12'h74: dout <= 8'b01100110; //  116 : 102 - 0x66
      12'h75: dout <= 8'b01100110; //  117 : 102 - 0x66
      12'h76: dout <= 8'b01100110; //  118 : 102 - 0x66
      12'h77: dout <= 8'b01100110; //  119 : 102 - 0x66
      12'h78: dout <= 8'b01100110; //  120 : 102 - 0x66 -- Sprite 0xf
      12'h79: dout <= 8'b01100110; //  121 : 102 - 0x66
      12'h7A: dout <= 8'b01100110; //  122 : 102 - 0x66
      12'h7B: dout <= 8'b01100110; //  123 : 102 - 0x66
      12'h7C: dout <= 8'b01100110; //  124 : 102 - 0x66
      12'h7D: dout <= 8'b01100110; //  125 : 102 - 0x66
      12'h7E: dout <= 8'b01100110; //  126 : 102 - 0x66
      12'h7F: dout <= 8'b01100110; //  127 : 102 - 0x66
      12'h80: dout <= 8'b01100110; //  128 : 102 - 0x66 -- Sprite 0x10
      12'h81: dout <= 8'b00110110; //  129 :  54 - 0x36
      12'h82: dout <= 8'b10110110; //  130 : 182 - 0xb6
      12'h83: dout <= 8'b10011110; //  131 : 158 - 0x9e
      12'h84: dout <= 8'b11011110; //  132 : 222 - 0xde
      12'h85: dout <= 8'b11001110; //  133 : 206 - 0xce
      12'h86: dout <= 8'b11101110; //  134 : 238 - 0xee
      12'h87: dout <= 8'b11100110; //  135 : 230 - 0xe6
      12'h88: dout <= 8'b10000001; //  136 : 129 - 0x81 -- Sprite 0x11
      12'h89: dout <= 8'b00111100; //  137 :  60 - 0x3c
      12'h8A: dout <= 8'b01111110; //  138 : 126 - 0x7e
      12'h8B: dout <= 8'b01100110; //  139 : 102 - 0x66
      12'h8C: dout <= 8'b01100110; //  140 : 102 - 0x66
      12'h8D: dout <= 8'b01100110; //  141 : 102 - 0x66
      12'h8E: dout <= 8'b01100110; //  142 : 102 - 0x66
      12'h8F: dout <= 8'b01100110; //  143 : 102 - 0x66
      12'h90: dout <= 8'b11110110; //  144 : 246 - 0xf6 -- Sprite 0x12
      12'h91: dout <= 8'b11110010; //  145 : 242 - 0xf2
      12'h92: dout <= 8'b11111010; //  146 : 250 - 0xfa
      12'h93: dout <= 8'b11111000; //  147 : 248 - 0xf8
      12'h94: dout <= 8'b11111100; //  148 : 252 - 0xfc
      12'h95: dout <= 8'b11111100; //  149 : 252 - 0xfc
      12'h96: dout <= 8'b11111110; //  150 : 254 - 0xfe
      12'h97: dout <= 8'b11111110; //  151 : 254 - 0xfe
      12'h98: dout <= 8'b01100110; //  152 : 102 - 0x66 -- Sprite 0x13
      12'h99: dout <= 8'b01100110; //  153 : 102 - 0x66
      12'h9A: dout <= 8'b01100110; //  154 : 102 - 0x66
      12'h9B: dout <= 8'b01100110; //  155 : 102 - 0x66
      12'h9C: dout <= 8'b01100110; //  156 : 102 - 0x66
      12'h9D: dout <= 8'b01100110; //  157 : 102 - 0x66
      12'h9E: dout <= 8'b01100110; //  158 : 102 - 0x66
      12'h9F: dout <= 8'b01111110; //  159 : 126 - 0x7e
      12'hA0: dout <= 8'b11111111; //  160 : 255 - 0xff -- Sprite 0x14
      12'hA1: dout <= 8'b01111111; //  161 : 127 - 0x7f
      12'hA2: dout <= 8'b01111111; //  162 : 127 - 0x7f
      12'hA3: dout <= 8'b00111111; //  163 :  63 - 0x3f
      12'hA4: dout <= 8'b00111111; //  164 :  63 - 0x3f
      12'hA5: dout <= 8'b00011111; //  165 :  31 - 0x1f
      12'hA6: dout <= 8'b01011111; //  166 :  95 - 0x5f
      12'hA7: dout <= 8'b01001111; //  167 :  79 - 0x4f
      12'hA8: dout <= 8'b01100110; //  168 : 102 - 0x66 -- Sprite 0x15
      12'hA9: dout <= 8'b01100110; //  169 : 102 - 0x66
      12'hAA: dout <= 8'b01100110; //  170 : 102 - 0x66
      12'hAB: dout <= 8'b01100110; //  171 : 102 - 0x66
      12'hAC: dout <= 8'b01100110; //  172 : 102 - 0x66
      12'hAD: dout <= 8'b01111110; //  173 : 126 - 0x7e
      12'hAE: dout <= 8'b01111110; //  174 : 126 - 0x7e
      12'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      12'hB0: dout <= 8'b01111110; //  176 : 126 - 0x7e -- Sprite 0x16
      12'hB1: dout <= 8'b01100110; //  177 : 102 - 0x66
      12'hB2: dout <= 8'b01000010; //  178 :  66 - 0x42
      12'hB3: dout <= 8'b00011000; //  179 :  24 - 0x18
      12'hB4: dout <= 8'b00111100; //  180 :  60 - 0x3c
      12'hB5: dout <= 8'b01111110; //  181 : 126 - 0x7e
      12'hB6: dout <= 8'b11111111; //  182 : 255 - 0xff
      12'hB7: dout <= 8'b11111111; //  183 : 255 - 0xff
      12'hB8: dout <= 8'b01101111; //  184 : 111 - 0x6f -- Sprite 0x17
      12'hB9: dout <= 8'b01100111; //  185 : 103 - 0x67
      12'hBA: dout <= 8'b01110111; //  186 : 119 - 0x77
      12'hBB: dout <= 8'b01110011; //  187 : 115 - 0x73
      12'hBC: dout <= 8'b01111011; //  188 : 123 - 0x7b
      12'hBD: dout <= 8'b01111001; //  189 : 121 - 0x79
      12'hBE: dout <= 8'b01101101; //  190 : 109 - 0x6d
      12'hBF: dout <= 8'b01101100; //  191 : 108 - 0x6c
      12'hC0: dout <= 8'b01100000; //  192 :  96 - 0x60 -- Sprite 0x18
      12'hC1: dout <= 8'b01100000; //  193 :  96 - 0x60
      12'hC2: dout <= 8'b01100000; //  194 :  96 - 0x60
      12'hC3: dout <= 8'b01100000; //  195 :  96 - 0x60
      12'hC4: dout <= 8'b01100000; //  196 :  96 - 0x60
      12'hC5: dout <= 8'b01111111; //  197 : 127 - 0x7f
      12'hC6: dout <= 8'b01111111; //  198 : 127 - 0x7f
      12'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      12'hC8: dout <= 8'b00000110; //  200 :   6 - 0x6 -- Sprite 0x19
      12'hC9: dout <= 8'b00000110; //  201 :   6 - 0x6
      12'hCA: dout <= 8'b00000110; //  202 :   6 - 0x6
      12'hCB: dout <= 8'b00000110; //  203 :   6 - 0x6
      12'hCC: dout <= 8'b00000110; //  204 :   6 - 0x6
      12'hCD: dout <= 8'b11100110; //  205 : 230 - 0xe6
      12'hCE: dout <= 8'b11100110; //  206 : 230 - 0xe6
      12'hCF: dout <= 8'b01100110; //  207 : 102 - 0x66
      12'hD0: dout <= 8'b11111111; //  208 : 255 - 0xff -- Sprite 0x1a
      12'hD1: dout <= 8'b11111111; //  209 : 255 - 0xff
      12'hD2: dout <= 8'b11111111; //  210 : 255 - 0xff
      12'hD3: dout <= 8'b11111111; //  211 : 255 - 0xff
      12'hD4: dout <= 8'b11100111; //  212 : 231 - 0xe7
      12'hD5: dout <= 8'b11000011; //  213 : 195 - 0xc3
      12'hD6: dout <= 8'b10011001; //  214 : 153 - 0x99
      12'hD7: dout <= 8'b00111100; //  215 :  60 - 0x3c
      12'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x1b
      12'hD9: dout <= 8'b01111110; //  217 : 126 - 0x7e
      12'hDA: dout <= 8'b01111110; //  218 : 126 - 0x7e
      12'hDB: dout <= 8'b01100110; //  219 : 102 - 0x66
      12'hDC: dout <= 8'b01100110; //  220 : 102 - 0x66
      12'hDD: dout <= 8'b01100110; //  221 : 102 - 0x66
      12'hDE: dout <= 8'b01100110; //  222 : 102 - 0x66
      12'hDF: dout <= 8'b01100110; //  223 : 102 - 0x66
      12'hE0: dout <= 8'b11111110; //  224 : 254 - 0xfe -- Sprite 0x1c
      12'hE1: dout <= 8'b11111100; //  225 : 252 - 0xfc
      12'hE2: dout <= 8'b11111001; //  226 : 249 - 0xf9
      12'hE3: dout <= 8'b11110011; //  227 : 243 - 0xf3
      12'hE4: dout <= 8'b11100111; //  228 : 231 - 0xe7
      12'hE5: dout <= 8'b11001110; //  229 : 206 - 0xce
      12'hE6: dout <= 8'b10011100; //  230 : 156 - 0x9c
      12'hE7: dout <= 8'b00111000; //  231 :  56 - 0x38
      12'hE8: dout <= 8'b01111110; //  232 : 126 - 0x7e -- Sprite 0x1d
      12'hE9: dout <= 8'b11100111; //  233 : 231 - 0xe7
      12'hEA: dout <= 8'b11000011; //  234 : 195 - 0xc3
      12'hEB: dout <= 8'b10000001; //  235 : 129 - 0x81
      12'hEC: dout <= 8'b00000000; //  236 :   0 - 0x0
      12'hED: dout <= 8'b00000000; //  237 :   0 - 0x0
      12'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      12'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      12'hF0: dout <= 8'b01111111; //  240 : 127 - 0x7f -- Sprite 0x1e
      12'hF1: dout <= 8'b00111111; //  241 :  63 - 0x3f
      12'hF2: dout <= 8'b10011111; //  242 : 159 - 0x9f
      12'hF3: dout <= 8'b11001111; //  243 : 207 - 0xcf
      12'hF4: dout <= 8'b11100111; //  244 : 231 - 0xe7
      12'hF5: dout <= 8'b01110011; //  245 : 115 - 0x73
      12'hF6: dout <= 8'b00111001; //  246 :  57 - 0x39
      12'hF7: dout <= 8'b00011100; //  247 :  28 - 0x1c
      12'hF8: dout <= 8'b00000110; //  248 :   6 - 0x6 -- Sprite 0x1f
      12'hF9: dout <= 8'b00000111; //  249 :   7 - 0x7
      12'hFA: dout <= 8'b00000111; //  250 :   7 - 0x7
      12'hFB: dout <= 8'b00000000; //  251 :   0 - 0x0
      12'hFC: dout <= 8'b00000000; //  252 :   0 - 0x0
      12'hFD: dout <= 8'b00000000; //  253 :   0 - 0x0
      12'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      12'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      12'h101: dout <= 8'b11111111; //  257 : 255 - 0xff
      12'h102: dout <= 8'b11111111; //  258 : 255 - 0xff
      12'h103: dout <= 8'b00000000; //  259 :   0 - 0x0
      12'h104: dout <= 8'b00000000; //  260 :   0 - 0x0
      12'h105: dout <= 8'b00000000; //  261 :   0 - 0x0
      12'h106: dout <= 8'b00000000; //  262 :   0 - 0x0
      12'h107: dout <= 8'b00000000; //  263 :   0 - 0x0
      12'h108: dout <= 8'b01100110; //  264 : 102 - 0x66 -- Sprite 0x21
      12'h109: dout <= 8'b11100111; //  265 : 231 - 0xe7
      12'h10A: dout <= 8'b11100111; //  266 : 231 - 0xe7
      12'h10B: dout <= 8'b00000000; //  267 :   0 - 0x0
      12'h10C: dout <= 8'b00000000; //  268 :   0 - 0x0
      12'h10D: dout <= 8'b00000000; //  269 :   0 - 0x0
      12'h10E: dout <= 8'b00000000; //  270 :   0 - 0x0
      12'h10F: dout <= 8'b00000000; //  271 :   0 - 0x0
      12'h110: dout <= 8'b01110000; //  272 : 112 - 0x70 -- Sprite 0x22
      12'h111: dout <= 8'b11100000; //  273 : 224 - 0xe0
      12'h112: dout <= 8'b11000000; //  274 : 192 - 0xc0
      12'h113: dout <= 8'b00000000; //  275 :   0 - 0x0
      12'h114: dout <= 8'b00000000; //  276 :   0 - 0x0
      12'h115: dout <= 8'b00000000; //  277 :   0 - 0x0
      12'h116: dout <= 8'b00000000; //  278 :   0 - 0x0
      12'h117: dout <= 8'b00000000; //  279 :   0 - 0x0
      12'h118: dout <= 8'b00001110; //  280 :  14 - 0xe -- Sprite 0x23
      12'h119: dout <= 8'b00000111; //  281 :   7 - 0x7
      12'h11A: dout <= 8'b00000011; //  282 :   3 - 0x3
      12'h11B: dout <= 8'b00000000; //  283 :   0 - 0x0
      12'h11C: dout <= 8'b00000000; //  284 :   0 - 0x0
      12'h11D: dout <= 8'b00000000; //  285 :   0 - 0x0
      12'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      12'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      12'h120: dout <= 8'b01100000; //  288 :  96 - 0x60 -- Sprite 0x24
      12'h121: dout <= 8'b11100000; //  289 : 224 - 0xe0
      12'h122: dout <= 8'b11100000; //  290 : 224 - 0xe0
      12'h123: dout <= 8'b00000000; //  291 :   0 - 0x0
      12'h124: dout <= 8'b00000000; //  292 :   0 - 0x0
      12'h125: dout <= 8'b00000000; //  293 :   0 - 0x0
      12'h126: dout <= 8'b00000000; //  294 :   0 - 0x0
      12'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout <= 8'b00000000; //  296 :   0 - 0x0 -- Sprite 0x25
      12'h129: dout <= 8'b00000000; //  297 :   0 - 0x0
      12'h12A: dout <= 8'b00000000; //  298 :   0 - 0x0
      12'h12B: dout <= 8'b00000000; //  299 :   0 - 0x0
      12'h12C: dout <= 8'b00000000; //  300 :   0 - 0x0
      12'h12D: dout <= 8'b11000000; //  301 : 192 - 0xc0
      12'h12E: dout <= 8'b11100000; //  302 : 224 - 0xe0
      12'h12F: dout <= 8'b01110000; //  303 : 112 - 0x70
      12'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      12'h131: dout <= 8'b00000000; //  305 :   0 - 0x0
      12'h132: dout <= 8'b00000000; //  306 :   0 - 0x0
      12'h133: dout <= 8'b00000000; //  307 :   0 - 0x0
      12'h134: dout <= 8'b00000000; //  308 :   0 - 0x0
      12'h135: dout <= 8'b00000011; //  309 :   3 - 0x3
      12'h136: dout <= 8'b00000111; //  310 :   7 - 0x7
      12'h137: dout <= 8'b00001110; //  311 :  14 - 0xe
      12'h138: dout <= 8'b00111000; //  312 :  56 - 0x38 -- Sprite 0x27
      12'h139: dout <= 8'b10011100; //  313 : 156 - 0x9c
      12'h13A: dout <= 8'b11001110; //  314 : 206 - 0xce
      12'h13B: dout <= 8'b11100111; //  315 : 231 - 0xe7
      12'h13C: dout <= 8'b11110011; //  316 : 243 - 0xf3
      12'h13D: dout <= 8'b11111001; //  317 : 249 - 0xf9
      12'h13E: dout <= 8'b11111100; //  318 : 252 - 0xfc
      12'h13F: dout <= 8'b11111110; //  319 : 254 - 0xfe
      12'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      12'h141: dout <= 8'b00000000; //  321 :   0 - 0x0
      12'h142: dout <= 8'b00000000; //  322 :   0 - 0x0
      12'h143: dout <= 8'b00000000; //  323 :   0 - 0x0
      12'h144: dout <= 8'b10000001; //  324 : 129 - 0x81
      12'h145: dout <= 8'b11000011; //  325 : 195 - 0xc3
      12'h146: dout <= 8'b11100111; //  326 : 231 - 0xe7
      12'h147: dout <= 8'b01111110; //  327 : 126 - 0x7e
      12'h148: dout <= 8'b00011100; //  328 :  28 - 0x1c -- Sprite 0x29
      12'h149: dout <= 8'b00111001; //  329 :  57 - 0x39
      12'h14A: dout <= 8'b01110011; //  330 : 115 - 0x73
      12'h14B: dout <= 8'b11100111; //  331 : 231 - 0xe7
      12'h14C: dout <= 8'b11001111; //  332 : 207 - 0xcf
      12'h14D: dout <= 8'b10011111; //  333 : 159 - 0x9f
      12'h14E: dout <= 8'b00111111; //  334 :  63 - 0x3f
      12'h14F: dout <= 8'b01111111; //  335 : 127 - 0x7f
      12'h150: dout <= 8'b01100001; //  336 :  97 - 0x61 -- Sprite 0x2a
      12'h151: dout <= 8'b01100011; //  337 :  99 - 0x63
      12'h152: dout <= 8'b01100011; //  338 :  99 - 0x63
      12'h153: dout <= 8'b01100111; //  339 : 103 - 0x67
      12'h154: dout <= 8'b01100110; //  340 : 102 - 0x66
      12'h155: dout <= 8'b01100110; //  341 : 102 - 0x66
      12'h156: dout <= 8'b01100110; //  342 : 102 - 0x66
      12'h157: dout <= 8'b01100110; //  343 : 102 - 0x66
      12'h158: dout <= 8'b10000000; //  344 : 128 - 0x80 -- Sprite 0x2b
      12'h159: dout <= 8'b11000000; //  345 : 192 - 0xc0
      12'h15A: dout <= 8'b11000000; //  346 : 192 - 0xc0
      12'h15B: dout <= 8'b11100000; //  347 : 224 - 0xe0
      12'h15C: dout <= 8'b01100000; //  348 :  96 - 0x60
      12'h15D: dout <= 8'b01100000; //  349 :  96 - 0x60
      12'h15E: dout <= 8'b01100000; //  350 :  96 - 0x60
      12'h15F: dout <= 8'b01100000; //  351 :  96 - 0x60
      12'h160: dout <= 8'b00111100; //  352 :  60 - 0x3c -- Sprite 0x2c
      12'h161: dout <= 8'b10011001; //  353 : 153 - 0x99
      12'h162: dout <= 8'b11000011; //  354 : 195 - 0xc3
      12'h163: dout <= 8'b11100111; //  355 : 231 - 0xe7
      12'h164: dout <= 8'b11111111; //  356 : 255 - 0xff
      12'h165: dout <= 8'b11111111; //  357 : 255 - 0xff
      12'h166: dout <= 8'b11111111; //  358 : 255 - 0xff
      12'h167: dout <= 8'b11111111; //  359 : 255 - 0xff
      12'h168: dout <= 8'b00000000; //  360 :   0 - 0x0 -- Sprite 0x2d
      12'h169: dout <= 8'b01111111; //  361 : 127 - 0x7f
      12'h16A: dout <= 8'b01111111; //  362 : 127 - 0x7f
      12'h16B: dout <= 8'b01100000; //  363 :  96 - 0x60
      12'h16C: dout <= 8'b01100000; //  364 :  96 - 0x60
      12'h16D: dout <= 8'b01100000; //  365 :  96 - 0x60
      12'h16E: dout <= 8'b01100000; //  366 :  96 - 0x60
      12'h16F: dout <= 8'b01100000; //  367 :  96 - 0x60
      12'h170: dout <= 8'b01100110; //  368 : 102 - 0x66 -- Sprite 0x2e
      12'h171: dout <= 8'b11100110; //  369 : 230 - 0xe6
      12'h172: dout <= 8'b11100110; //  370 : 230 - 0xe6
      12'h173: dout <= 8'b00000110; //  371 :   6 - 0x6
      12'h174: dout <= 8'b00000110; //  372 :   6 - 0x6
      12'h175: dout <= 8'b00000110; //  373 :   6 - 0x6
      12'h176: dout <= 8'b00000110; //  374 :   6 - 0x6
      12'h177: dout <= 8'b00000110; //  375 :   6 - 0x6
      12'h178: dout <= 8'b00000001; //  376 :   1 - 0x1 -- Sprite 0x2f
      12'h179: dout <= 8'b01111100; //  377 : 124 - 0x7c
      12'h17A: dout <= 8'b01111110; //  378 : 126 - 0x7e
      12'h17B: dout <= 8'b01100110; //  379 : 102 - 0x66
      12'h17C: dout <= 8'b01100110; //  380 : 102 - 0x66
      12'h17D: dout <= 8'b01100110; //  381 : 102 - 0x66
      12'h17E: dout <= 8'b01100110; //  382 : 102 - 0x66
      12'h17F: dout <= 8'b01100110; //  383 : 102 - 0x66
      12'h180: dout <= 8'b11111111; //  384 : 255 - 0xff -- Sprite 0x30
      12'h181: dout <= 8'b11111111; //  385 : 255 - 0xff
      12'h182: dout <= 8'b01111110; //  386 : 126 - 0x7e
      12'h183: dout <= 8'b00111100; //  387 :  60 - 0x3c
      12'h184: dout <= 8'b00011000; //  388 :  24 - 0x18
      12'h185: dout <= 8'b01000010; //  389 :  66 - 0x42
      12'h186: dout <= 8'b01100110; //  390 : 102 - 0x66
      12'h187: dout <= 8'b01111110; //  391 : 126 - 0x7e
      12'h188: dout <= 8'b01100000; //  392 :  96 - 0x60 -- Sprite 0x31
      12'h189: dout <= 8'b01111111; //  393 : 127 - 0x7f
      12'h18A: dout <= 8'b01111111; //  394 : 127 - 0x7f
      12'h18B: dout <= 8'b00000000; //  395 :   0 - 0x0
      12'h18C: dout <= 8'b11111111; //  396 : 255 - 0xff
      12'h18D: dout <= 8'b11111111; //  397 : 255 - 0xff
      12'h18E: dout <= 8'b11111111; //  398 : 255 - 0xff
      12'h18F: dout <= 8'b11111111; //  399 : 255 - 0xff
      12'h190: dout <= 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      12'h191: dout <= 8'b11111111; //  401 : 255 - 0xff
      12'h192: dout <= 8'b11111111; //  402 : 255 - 0xff
      12'h193: dout <= 8'b00000000; //  403 :   0 - 0x0
      12'h194: dout <= 8'b11111111; //  404 : 255 - 0xff
      12'h195: dout <= 8'b11111111; //  405 : 255 - 0xff
      12'h196: dout <= 8'b11111111; //  406 : 255 - 0xff
      12'h197: dout <= 8'b11111111; //  407 : 255 - 0xff
      12'h198: dout <= 8'b00000000; //  408 :   0 - 0x0 -- Sprite 0x33
      12'h199: dout <= 8'b11100000; //  409 : 224 - 0xe0
      12'h19A: dout <= 8'b11100000; //  410 : 224 - 0xe0
      12'h19B: dout <= 8'b01100000; //  411 :  96 - 0x60
      12'h19C: dout <= 8'b01100000; //  412 :  96 - 0x60
      12'h19D: dout <= 8'b01100000; //  413 :  96 - 0x60
      12'h19E: dout <= 8'b01100000; //  414 :  96 - 0x60
      12'h19F: dout <= 8'b01100000; //  415 :  96 - 0x60
      12'h1A0: dout <= 8'b01111110; //  416 : 126 - 0x7e -- Sprite 0x34
      12'h1A1: dout <= 8'b01100110; //  417 : 102 - 0x66
      12'h1A2: dout <= 8'b01100110; //  418 : 102 - 0x66
      12'h1A3: dout <= 8'b01100110; //  419 : 102 - 0x66
      12'h1A4: dout <= 8'b01100110; //  420 : 102 - 0x66
      12'h1A5: dout <= 8'b01100110; //  421 : 102 - 0x66
      12'h1A6: dout <= 8'b01100110; //  422 : 102 - 0x66
      12'h1A7: dout <= 8'b01100110; //  423 : 102 - 0x66
      12'h1A8: dout <= 8'b11111111; //  424 : 255 - 0xff -- Sprite 0x35
      12'h1A9: dout <= 8'b11111111; //  425 : 255 - 0xff
      12'h1AA: dout <= 8'b11111111; //  426 : 255 - 0xff
      12'h1AB: dout <= 8'b11111111; //  427 : 255 - 0xff
      12'h1AC: dout <= 8'b00000000; //  428 :   0 - 0x0
      12'h1AD: dout <= 8'b01111111; //  429 : 127 - 0x7f
      12'h1AE: dout <= 8'b01111111; //  430 : 127 - 0x7f
      12'h1AF: dout <= 8'b01100000; //  431 :  96 - 0x60
      12'h1B0: dout <= 8'b11111111; //  432 : 255 - 0xff -- Sprite 0x36
      12'h1B1: dout <= 8'b11111111; //  433 : 255 - 0xff
      12'h1B2: dout <= 8'b11111111; //  434 : 255 - 0xff
      12'h1B3: dout <= 8'b11111111; //  435 : 255 - 0xff
      12'h1B4: dout <= 8'b00000000; //  436 :   0 - 0x0
      12'h1B5: dout <= 8'b11111111; //  437 : 255 - 0xff
      12'h1B6: dout <= 8'b11111111; //  438 : 255 - 0xff
      12'h1B7: dout <= 8'b00000000; //  439 :   0 - 0x0
      12'h1B8: dout <= 8'b01100000; //  440 :  96 - 0x60 -- Sprite 0x37
      12'h1B9: dout <= 8'b01100000; //  441 :  96 - 0x60
      12'h1BA: dout <= 8'b01100000; //  442 :  96 - 0x60
      12'h1BB: dout <= 8'b01100000; //  443 :  96 - 0x60
      12'h1BC: dout <= 8'b01100000; //  444 :  96 - 0x60
      12'h1BD: dout <= 8'b11100000; //  445 : 224 - 0xe0
      12'h1BE: dout <= 8'b11100000; //  446 : 224 - 0xe0
      12'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout <= 8'b01100110; //  448 : 102 - 0x66 -- Sprite 0x38
      12'h1C1: dout <= 8'b01100110; //  449 : 102 - 0x66
      12'h1C2: dout <= 8'b01100110; //  450 : 102 - 0x66
      12'h1C3: dout <= 8'b01100110; //  451 : 102 - 0x66
      12'h1C4: dout <= 8'b01100110; //  452 : 102 - 0x66
      12'h1C5: dout <= 8'b01111110; //  453 : 126 - 0x7e
      12'h1C6: dout <= 8'b01111100; //  454 : 124 - 0x7c
      12'h1C7: dout <= 8'b00000001; //  455 :   1 - 0x1
      12'h1C8: dout <= 8'b11111111; //  456 : 255 - 0xff -- Sprite 0x39
      12'h1C9: dout <= 8'b11111111; //  457 : 255 - 0xff
      12'h1CA: dout <= 8'b11111111; //  458 : 255 - 0xff
      12'h1CB: dout <= 8'b11111111; //  459 : 255 - 0xff
      12'h1CC: dout <= 8'b11111111; //  460 : 255 - 0xff
      12'h1CD: dout <= 8'b11111111; //  461 : 255 - 0xff
      12'h1CE: dout <= 8'b11111111; //  462 : 255 - 0xff
      12'h1CF: dout <= 8'b11111110; //  463 : 254 - 0xfe
      12'h1D0: dout <= 8'b01100110; //  464 : 102 - 0x66 -- Sprite 0x3a
      12'h1D1: dout <= 8'b01100110; //  465 : 102 - 0x66
      12'h1D2: dout <= 8'b01100110; //  466 : 102 - 0x66
      12'h1D3: dout <= 8'b01100110; //  467 : 102 - 0x66
      12'h1D4: dout <= 8'b01100110; //  468 : 102 - 0x66
      12'h1D5: dout <= 8'b01111110; //  469 : 126 - 0x7e
      12'h1D6: dout <= 8'b00111100; //  470 :  60 - 0x3c
      12'h1D7: dout <= 8'b10000001; //  471 : 129 - 0x81
      12'h1D8: dout <= 8'b01100000; //  472 :  96 - 0x60 -- Sprite 0x3b
      12'h1D9: dout <= 8'b01100000; //  473 :  96 - 0x60
      12'h1DA: dout <= 8'b01100000; //  474 :  96 - 0x60
      12'h1DB: dout <= 8'b01100000; //  475 :  96 - 0x60
      12'h1DC: dout <= 8'b01100000; //  476 :  96 - 0x60
      12'h1DD: dout <= 8'b01111111; //  477 : 127 - 0x7f
      12'h1DE: dout <= 8'b01111111; //  478 : 127 - 0x7f
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      12'h1E1: dout <= 8'b00000000; //  481 :   0 - 0x0
      12'h1E2: dout <= 8'b00000000; //  482 :   0 - 0x0
      12'h1E3: dout <= 8'b00000000; //  483 :   0 - 0x0
      12'h1E4: dout <= 8'b00000000; //  484 :   0 - 0x0
      12'h1E5: dout <= 8'b11111111; //  485 : 255 - 0xff
      12'h1E6: dout <= 8'b11111111; //  486 : 255 - 0xff
      12'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      12'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      12'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      12'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      12'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      12'h1ED: dout <= 8'b11111111; //  493 : 255 - 0xff
      12'h1EE: dout <= 8'b11111111; //  494 : 255 - 0xff
      12'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout <= 8'b11111110; //  496 : 254 - 0xfe -- Sprite 0x3e
      12'h1F1: dout <= 8'b11111100; //  497 : 252 - 0xfc
      12'h1F2: dout <= 8'b11111001; //  498 : 249 - 0xf9
      12'h1F3: dout <= 8'b11110011; //  499 : 243 - 0xf3
      12'h1F4: dout <= 8'b11110011; //  500 : 243 - 0xf3
      12'h1F5: dout <= 8'b11111001; //  501 : 249 - 0xf9
      12'h1F6: dout <= 8'b11111100; //  502 : 252 - 0xfc
      12'h1F7: dout <= 8'b11111110; //  503 : 254 - 0xfe
      12'h1F8: dout <= 8'b11100000; //  504 : 224 - 0xe0 -- Sprite 0x3f
      12'h1F9: dout <= 8'b11000000; //  505 : 192 - 0xc0
      12'h1FA: dout <= 8'b11000000; //  506 : 192 - 0xc0
      12'h1FB: dout <= 8'b10000000; //  507 : 128 - 0x80
      12'h1FC: dout <= 8'b10000000; //  508 : 128 - 0x80
      12'h1FD: dout <= 8'b11000000; //  509 : 192 - 0xc0
      12'h1FE: dout <= 8'b11000000; //  510 : 192 - 0xc0
      12'h1FF: dout <= 8'b11100000; //  511 : 224 - 0xe0
      12'h200: dout <= 8'b01100110; //  512 : 102 - 0x66 -- Sprite 0x40
      12'h201: dout <= 8'b01100110; //  513 : 102 - 0x66
      12'h202: dout <= 8'b01100110; //  514 : 102 - 0x66
      12'h203: dout <= 8'b01100110; //  515 : 102 - 0x66
      12'h204: dout <= 8'b01100111; //  516 : 103 - 0x67
      12'h205: dout <= 8'b01100011; //  517 :  99 - 0x63
      12'h206: dout <= 8'b01100011; //  518 :  99 - 0x63
      12'h207: dout <= 8'b01100001; //  519 :  97 - 0x61
      12'h208: dout <= 8'b11111111; //  520 : 255 - 0xff -- Sprite 0x41
      12'h209: dout <= 8'b11111111; //  521 : 255 - 0xff
      12'h20A: dout <= 8'b11111111; //  522 : 255 - 0xff
      12'h20B: dout <= 8'b01111111; //  523 : 127 - 0x7f
      12'h20C: dout <= 8'b01111111; //  524 : 127 - 0x7f
      12'h20D: dout <= 8'b00111111; //  525 :  63 - 0x3f
      12'h20E: dout <= 8'b10011111; //  526 : 159 - 0x9f
      12'h20F: dout <= 8'b11000111; //  527 : 199 - 0xc7
      12'h210: dout <= 8'b11111111; //  528 : 255 - 0xff -- Sprite 0x42
      12'h211: dout <= 8'b11111111; //  529 : 255 - 0xff
      12'h212: dout <= 8'b11111111; //  530 : 255 - 0xff
      12'h213: dout <= 8'b11111110; //  531 : 254 - 0xfe
      12'h214: dout <= 8'b11111110; //  532 : 254 - 0xfe
      12'h215: dout <= 8'b11111100; //  533 : 252 - 0xfc
      12'h216: dout <= 8'b11111001; //  534 : 249 - 0xf9
      12'h217: dout <= 8'b11100011; //  535 : 227 - 0xe3
      12'h218: dout <= 8'b01100110; //  536 : 102 - 0x66 -- Sprite 0x43
      12'h219: dout <= 8'b01100110; //  537 : 102 - 0x66
      12'h21A: dout <= 8'b01100110; //  538 : 102 - 0x66
      12'h21B: dout <= 8'b01100110; //  539 : 102 - 0x66
      12'h21C: dout <= 8'b11100110; //  540 : 230 - 0xe6
      12'h21D: dout <= 8'b11000110; //  541 : 198 - 0xc6
      12'h21E: dout <= 8'b11000110; //  542 : 198 - 0xc6
      12'h21F: dout <= 8'b10000110; //  543 : 134 - 0x86
      12'h220: dout <= 8'b11111110; //  544 : 254 - 0xfe -- Sprite 0x44
      12'h221: dout <= 8'b11111111; //  545 : 255 - 0xff
      12'h222: dout <= 8'b11111111; //  546 : 255 - 0xff
      12'h223: dout <= 8'b11111111; //  547 : 255 - 0xff
      12'h224: dout <= 8'b11111111; //  548 : 255 - 0xff
      12'h225: dout <= 8'b11111111; //  549 : 255 - 0xff
      12'h226: dout <= 8'b11111111; //  550 : 255 - 0xff
      12'h227: dout <= 8'b11111111; //  551 : 255 - 0xff
      12'h228: dout <= 8'b01100000; //  552 :  96 - 0x60 -- Sprite 0x45
      12'h229: dout <= 8'b01100000; //  553 :  96 - 0x60
      12'h22A: dout <= 8'b01100000; //  554 :  96 - 0x60
      12'h22B: dout <= 8'b01100000; //  555 :  96 - 0x60
      12'h22C: dout <= 8'b01100000; //  556 :  96 - 0x60
      12'h22D: dout <= 8'b01100000; //  557 :  96 - 0x60
      12'h22E: dout <= 8'b01100000; //  558 :  96 - 0x60
      12'h22F: dout <= 8'b01100000; //  559 :  96 - 0x60
      12'h230: dout <= 8'b11110000; //  560 : 240 - 0xf0 -- Sprite 0x46
      12'h231: dout <= 8'b01111111; //  561 : 127 - 0x7f
      12'h232: dout <= 8'b00011111; //  562 :  31 - 0x1f
      12'h233: dout <= 8'b00000000; //  563 :   0 - 0x0
      12'h234: dout <= 8'b00000000; //  564 :   0 - 0x0
      12'h235: dout <= 8'b00000000; //  565 :   0 - 0x0
      12'h236: dout <= 8'b00000000; //  566 :   0 - 0x0
      12'h237: dout <= 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout <= 8'b00001111; //  568 :  15 - 0xf -- Sprite 0x47
      12'h239: dout <= 8'b11111110; //  569 : 254 - 0xfe
      12'h23A: dout <= 8'b11111000; //  570 : 248 - 0xf8
      12'h23B: dout <= 8'b00000000; //  571 :   0 - 0x0
      12'h23C: dout <= 8'b00000000; //  572 :   0 - 0x0
      12'h23D: dout <= 8'b00000000; //  573 :   0 - 0x0
      12'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout <= 8'b00000110; //  576 :   6 - 0x6 -- Sprite 0x48
      12'h241: dout <= 8'b00000111; //  577 :   7 - 0x7
      12'h242: dout <= 8'b00000111; //  578 :   7 - 0x7
      12'h243: dout <= 8'b00000000; //  579 :   0 - 0x0
      12'h244: dout <= 8'b00000000; //  580 :   0 - 0x0
      12'h245: dout <= 8'b00000000; //  581 :   0 - 0x0
      12'h246: dout <= 8'b00000000; //  582 :   0 - 0x0
      12'h247: dout <= 8'b00000000; //  583 :   0 - 0x0
      12'h248: dout <= 8'b00000000; //  584 :   0 - 0x0 -- Sprite 0x49
      12'h249: dout <= 8'b00000000; //  585 :   0 - 0x0
      12'h24A: dout <= 8'b00000000; //  586 :   0 - 0x0
      12'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      12'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      12'h24D: dout <= 8'b00000000; //  589 :   0 - 0x0
      12'h24E: dout <= 8'b00000000; //  590 :   0 - 0x0
      12'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout <= 8'b00000000; //  592 :   0 - 0x0 -- Sprite 0x4a
      12'h251: dout <= 8'b01110110; //  593 : 118 - 0x76
      12'h252: dout <= 8'b01010111; //  594 :  87 - 0x57
      12'h253: dout <= 8'b01010101; //  595 :  85 - 0x55
      12'h254: dout <= 8'b01010101; //  596 :  85 - 0x55
      12'h255: dout <= 8'b01110101; //  597 : 117 - 0x75
      12'h256: dout <= 8'b01000111; //  598 :  71 - 0x47
      12'h257: dout <= 8'b00000000; //  599 :   0 - 0x0
      12'h258: dout <= 8'b00000000; //  600 :   0 - 0x0 -- Sprite 0x4b
      12'h259: dout <= 8'b01110111; //  601 : 119 - 0x77
      12'h25A: dout <= 8'b00010101; //  602 :  21 - 0x15
      12'h25B: dout <= 8'b01110101; //  603 : 117 - 0x75
      12'h25C: dout <= 8'b01000101; //  604 :  69 - 0x45
      12'h25D: dout <= 8'b01000101; //  605 :  69 - 0x45
      12'h25E: dout <= 8'b01110111; //  606 : 119 - 0x77
      12'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout <= 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x4c
      12'h261: dout <= 8'b00100100; //  609 :  36 - 0x24
      12'h262: dout <= 8'b01101100; //  610 : 108 - 0x6c
      12'h263: dout <= 8'b00100100; //  611 :  36 - 0x24
      12'h264: dout <= 8'b00100100; //  612 :  36 - 0x24
      12'h265: dout <= 8'b00100100; //  613 :  36 - 0x24
      12'h266: dout <= 8'b00100101; //  614 :  37 - 0x25
      12'h267: dout <= 8'b00000000; //  615 :   0 - 0x0
      12'h268: dout <= 8'b00000000; //  616 :   0 - 0x0 -- Sprite 0x4d
      12'h269: dout <= 8'b01110100; //  617 : 116 - 0x74
      12'h26A: dout <= 8'b01000111; //  618 :  71 - 0x47
      12'h26B: dout <= 8'b01110101; //  619 : 117 - 0x75
      12'h26C: dout <= 8'b00010101; //  620 :  21 - 0x15
      12'h26D: dout <= 8'b00010101; //  621 :  21 - 0x15
      12'h26E: dout <= 8'b01110101; //  622 : 117 - 0x75
      12'h26F: dout <= 8'b00000000; //  623 :   0 - 0x0
      12'h270: dout <= 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x4e
      12'h271: dout <= 8'b01000000; //  625 :  64 - 0x40
      12'h272: dout <= 8'b00011101; //  626 :  29 - 0x1d
      12'h273: dout <= 8'b01010101; //  627 :  85 - 0x55
      12'h274: dout <= 8'b01010001; //  628 :  81 - 0x51
      12'h275: dout <= 8'b01010001; //  629 :  81 - 0x51
      12'h276: dout <= 8'b01010001; //  630 :  81 - 0x51
      12'h277: dout <= 8'b00000000; //  631 :   0 - 0x0
      12'h278: dout <= 8'b00000000; //  632 :   0 - 0x0 -- Sprite 0x4f
      12'h279: dout <= 8'b00000000; //  633 :   0 - 0x0
      12'h27A: dout <= 8'b01001000; //  634 :  72 - 0x48
      12'h27B: dout <= 8'b01000001; //  635 :  65 - 0x41
      12'h27C: dout <= 8'b01000100; //  636 :  68 - 0x44
      12'h27D: dout <= 8'b01000000; //  637 :  64 - 0x40
      12'h27E: dout <= 8'b11010000; //  638 : 208 - 0xd0
      12'h27F: dout <= 8'b00000010; //  639 :   2 - 0x2
      12'h280: dout <= 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x50
      12'h281: dout <= 8'b00000000; //  641 :   0 - 0x0
      12'h282: dout <= 8'b11111100; //  642 : 252 - 0xfc
      12'h283: dout <= 8'b11111110; //  643 : 254 - 0xfe
      12'h284: dout <= 8'b11101110; //  644 : 238 - 0xee
      12'h285: dout <= 8'b11101110; //  645 : 238 - 0xee
      12'h286: dout <= 8'b11101110; //  646 : 238 - 0xee
      12'h287: dout <= 8'b11101110; //  647 : 238 - 0xee
      12'h288: dout <= 8'b00000000; //  648 :   0 - 0x0 -- Sprite 0x51
      12'h289: dout <= 8'b00000000; //  649 :   0 - 0x0
      12'h28A: dout <= 8'b11111100; //  650 : 252 - 0xfc
      12'h28B: dout <= 8'b11111110; //  651 : 254 - 0xfe
      12'h28C: dout <= 8'b11101110; //  652 : 238 - 0xee
      12'h28D: dout <= 8'b11101110; //  653 : 238 - 0xee
      12'h28E: dout <= 8'b11101110; //  654 : 238 - 0xee
      12'h28F: dout <= 8'b11101110; //  655 : 238 - 0xee
      12'h290: dout <= 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      12'h291: dout <= 8'b00000000; //  657 :   0 - 0x0
      12'h292: dout <= 8'b11111110; //  658 : 254 - 0xfe
      12'h293: dout <= 8'b11111110; //  659 : 254 - 0xfe
      12'h294: dout <= 8'b11100000; //  660 : 224 - 0xe0
      12'h295: dout <= 8'b11100000; //  661 : 224 - 0xe0
      12'h296: dout <= 8'b11111000; //  662 : 248 - 0xf8
      12'h297: dout <= 8'b11111000; //  663 : 248 - 0xf8
      12'h298: dout <= 8'b00000000; //  664 :   0 - 0x0 -- Sprite 0x53
      12'h299: dout <= 8'b00000000; //  665 :   0 - 0x0
      12'h29A: dout <= 8'b01111100; //  666 : 124 - 0x7c
      12'h29B: dout <= 8'b11111110; //  667 : 254 - 0xfe
      12'h29C: dout <= 8'b11101110; //  668 : 238 - 0xee
      12'h29D: dout <= 8'b11100000; //  669 : 224 - 0xe0
      12'h29E: dout <= 8'b11111100; //  670 : 252 - 0xfc
      12'h29F: dout <= 8'b01111110; //  671 : 126 - 0x7e
      12'h2A0: dout <= 8'b00000000; //  672 :   0 - 0x0 -- Sprite 0x54
      12'h2A1: dout <= 8'b00000000; //  673 :   0 - 0x0
      12'h2A2: dout <= 8'b11111110; //  674 : 254 - 0xfe
      12'h2A3: dout <= 8'b11111110; //  675 : 254 - 0xfe
      12'h2A4: dout <= 8'b00111000; //  676 :  56 - 0x38
      12'h2A5: dout <= 8'b00111000; //  677 :  56 - 0x38
      12'h2A6: dout <= 8'b00111000; //  678 :  56 - 0x38
      12'h2A7: dout <= 8'b00111000; //  679 :  56 - 0x38
      12'h2A8: dout <= 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      12'h2A9: dout <= 8'b00000000; //  681 :   0 - 0x0
      12'h2AA: dout <= 8'b01111100; //  682 : 124 - 0x7c
      12'h2AB: dout <= 8'b11111110; //  683 : 254 - 0xfe
      12'h2AC: dout <= 8'b11101110; //  684 : 238 - 0xee
      12'h2AD: dout <= 8'b11101110; //  685 : 238 - 0xee
      12'h2AE: dout <= 8'b11101110; //  686 : 238 - 0xee
      12'h2AF: dout <= 8'b11101110; //  687 : 238 - 0xee
      12'h2B0: dout <= 8'b00000000; //  688 :   0 - 0x0 -- Sprite 0x56
      12'h2B1: dout <= 8'b00000000; //  689 :   0 - 0x0
      12'h2B2: dout <= 8'b11100000; //  690 : 224 - 0xe0
      12'h2B3: dout <= 8'b11100000; //  691 : 224 - 0xe0
      12'h2B4: dout <= 8'b11100000; //  692 : 224 - 0xe0
      12'h2B5: dout <= 8'b11100000; //  693 : 224 - 0xe0
      12'h2B6: dout <= 8'b11100000; //  694 : 224 - 0xe0
      12'h2B7: dout <= 8'b11100000; //  695 : 224 - 0xe0
      12'h2B8: dout <= 8'b00000000; //  696 :   0 - 0x0 -- Sprite 0x57
      12'h2B9: dout <= 8'b00000000; //  697 :   0 - 0x0
      12'h2BA: dout <= 8'b11101110; //  698 : 238 - 0xee
      12'h2BB: dout <= 8'b11101110; //  699 : 238 - 0xee
      12'h2BC: dout <= 8'b11101110; //  700 : 238 - 0xee
      12'h2BD: dout <= 8'b11101110; //  701 : 238 - 0xee
      12'h2BE: dout <= 8'b11101110; //  702 : 238 - 0xee
      12'h2BF: dout <= 8'b11101110; //  703 : 238 - 0xee
      12'h2C0: dout <= 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x58
      12'h2C1: dout <= 8'b00000000; //  705 :   0 - 0x0
      12'h2C2: dout <= 8'b10001110; //  706 : 142 - 0x8e
      12'h2C3: dout <= 8'b11001110; //  707 : 206 - 0xce
      12'h2C4: dout <= 8'b11101110; //  708 : 238 - 0xee
      12'h2C5: dout <= 8'b11111110; //  709 : 254 - 0xfe
      12'h2C6: dout <= 8'b11111110; //  710 : 254 - 0xfe
      12'h2C7: dout <= 8'b11101110; //  711 : 238 - 0xee
      12'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0 -- Sprite 0x59
      12'h2C9: dout <= 8'b00000000; //  713 :   0 - 0x0
      12'h2CA: dout <= 8'b11111100; //  714 : 252 - 0xfc
      12'h2CB: dout <= 8'b11111110; //  715 : 254 - 0xfe
      12'h2CC: dout <= 8'b11101110; //  716 : 238 - 0xee
      12'h2CD: dout <= 8'b11101110; //  717 : 238 - 0xee
      12'h2CE: dout <= 8'b11101110; //  718 : 238 - 0xee
      12'h2CF: dout <= 8'b11101110; //  719 : 238 - 0xee
      12'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x5a
      12'h2D1: dout <= 8'b00000000; //  721 :   0 - 0x0
      12'h2D2: dout <= 8'b01111100; //  722 : 124 - 0x7c
      12'h2D3: dout <= 8'b11111110; //  723 : 254 - 0xfe
      12'h2D4: dout <= 8'b11101110; //  724 : 238 - 0xee
      12'h2D5: dout <= 8'b11101110; //  725 : 238 - 0xee
      12'h2D6: dout <= 8'b11101110; //  726 : 238 - 0xee
      12'h2D7: dout <= 8'b11101110; //  727 : 238 - 0xee
      12'h2D8: dout <= 8'b00000000; //  728 :   0 - 0x0 -- Sprite 0x5b
      12'h2D9: dout <= 8'b00000000; //  729 :   0 - 0x0
      12'h2DA: dout <= 8'b11111110; //  730 : 254 - 0xfe
      12'h2DB: dout <= 8'b11111110; //  731 : 254 - 0xfe
      12'h2DC: dout <= 8'b11100000; //  732 : 224 - 0xe0
      12'h2DD: dout <= 8'b11100000; //  733 : 224 - 0xe0
      12'h2DE: dout <= 8'b11111000; //  734 : 248 - 0xf8
      12'h2DF: dout <= 8'b11111000; //  735 : 248 - 0xf8
      12'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x5c
      12'h2E1: dout <= 8'b00000000; //  737 :   0 - 0x0
      12'h2E2: dout <= 8'b00000000; //  738 :   0 - 0x0
      12'h2E3: dout <= 8'b00000000; //  739 :   0 - 0x0
      12'h2E4: dout <= 8'b00000000; //  740 :   0 - 0x0
      12'h2E5: dout <= 8'b00000000; //  741 :   0 - 0x0
      12'h2E6: dout <= 8'b11001100; //  742 : 204 - 0xcc
      12'h2E7: dout <= 8'b11001100; //  743 : 204 - 0xcc
      12'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0 -- Sprite 0x5d
      12'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      12'h2EA: dout <= 8'b11111110; //  746 : 254 - 0xfe
      12'h2EB: dout <= 8'b11111110; //  747 : 254 - 0xfe
      12'h2EC: dout <= 8'b11100000; //  748 : 224 - 0xe0
      12'h2ED: dout <= 8'b11100000; //  749 : 224 - 0xe0
      12'h2EE: dout <= 8'b11111000; //  750 : 248 - 0xf8
      12'h2EF: dout <= 8'b11111000; //  751 : 248 - 0xf8
      12'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x5e
      12'h2F1: dout <= 8'b00000000; //  753 :   0 - 0x0
      12'h2F2: dout <= 8'b11101110; //  754 : 238 - 0xee
      12'h2F3: dout <= 8'b11101110; //  755 : 238 - 0xee
      12'h2F4: dout <= 8'b11101110; //  756 : 238 - 0xee
      12'h2F5: dout <= 8'b11101110; //  757 : 238 - 0xee
      12'h2F6: dout <= 8'b11101110; //  758 : 238 - 0xee
      12'h2F7: dout <= 8'b11101110; //  759 : 238 - 0xee
      12'h2F8: dout <= 8'b01111110; //  760 : 126 - 0x7e -- Sprite 0x5f
      12'h2F9: dout <= 8'b01111110; //  761 : 126 - 0x7e
      12'h2FA: dout <= 8'b01111110; //  762 : 126 - 0x7e
      12'h2FB: dout <= 8'b01111110; //  763 : 126 - 0x7e
      12'h2FC: dout <= 8'b01111110; //  764 : 126 - 0x7e
      12'h2FD: dout <= 8'b01111110; //  765 : 126 - 0x7e
      12'h2FE: dout <= 8'b01111110; //  766 : 126 - 0x7e
      12'h2FF: dout <= 8'b01111110; //  767 : 126 - 0x7e
      12'h300: dout <= 8'b11101110; //  768 : 238 - 0xee -- Sprite 0x60
      12'h301: dout <= 8'b11101110; //  769 : 238 - 0xee
      12'h302: dout <= 8'b11111110; //  770 : 254 - 0xfe
      12'h303: dout <= 8'b11111100; //  771 : 252 - 0xfc
      12'h304: dout <= 8'b11100000; //  772 : 224 - 0xe0
      12'h305: dout <= 8'b11100000; //  773 : 224 - 0xe0
      12'h306: dout <= 8'b00000000; //  774 :   0 - 0x0
      12'h307: dout <= 8'b00000000; //  775 :   0 - 0x0
      12'h308: dout <= 8'b11101110; //  776 : 238 - 0xee -- Sprite 0x61
      12'h309: dout <= 8'b11101110; //  777 : 238 - 0xee
      12'h30A: dout <= 8'b11111100; //  778 : 252 - 0xfc
      12'h30B: dout <= 8'b11111100; //  779 : 252 - 0xfc
      12'h30C: dout <= 8'b11101110; //  780 : 238 - 0xee
      12'h30D: dout <= 8'b11101110; //  781 : 238 - 0xee
      12'h30E: dout <= 8'b00000000; //  782 :   0 - 0x0
      12'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      12'h310: dout <= 8'b11100000; //  784 : 224 - 0xe0 -- Sprite 0x62
      12'h311: dout <= 8'b11100000; //  785 : 224 - 0xe0
      12'h312: dout <= 8'b11100000; //  786 : 224 - 0xe0
      12'h313: dout <= 8'b11100000; //  787 : 224 - 0xe0
      12'h314: dout <= 8'b11111110; //  788 : 254 - 0xfe
      12'h315: dout <= 8'b11111110; //  789 : 254 - 0xfe
      12'h316: dout <= 8'b00000000; //  790 :   0 - 0x0
      12'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout <= 8'b00001110; //  792 :  14 - 0xe -- Sprite 0x63
      12'h319: dout <= 8'b00001110; //  793 :  14 - 0xe
      12'h31A: dout <= 8'b00001110; //  794 :  14 - 0xe
      12'h31B: dout <= 8'b11101110; //  795 : 238 - 0xee
      12'h31C: dout <= 8'b11111110; //  796 : 254 - 0xfe
      12'h31D: dout <= 8'b01111100; //  797 : 124 - 0x7c
      12'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      12'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout <= 8'b00111000; //  800 :  56 - 0x38 -- Sprite 0x64
      12'h321: dout <= 8'b00111000; //  801 :  56 - 0x38
      12'h322: dout <= 8'b00111000; //  802 :  56 - 0x38
      12'h323: dout <= 8'b00111000; //  803 :  56 - 0x38
      12'h324: dout <= 8'b00111000; //  804 :  56 - 0x38
      12'h325: dout <= 8'b00111000; //  805 :  56 - 0x38
      12'h326: dout <= 8'b00000000; //  806 :   0 - 0x0
      12'h327: dout <= 8'b00000000; //  807 :   0 - 0x0
      12'h328: dout <= 8'b11101110; //  808 : 238 - 0xee -- Sprite 0x65
      12'h329: dout <= 8'b11101110; //  809 : 238 - 0xee
      12'h32A: dout <= 8'b11111110; //  810 : 254 - 0xfe
      12'h32B: dout <= 8'b11111110; //  811 : 254 - 0xfe
      12'h32C: dout <= 8'b11101110; //  812 : 238 - 0xee
      12'h32D: dout <= 8'b11101110; //  813 : 238 - 0xee
      12'h32E: dout <= 8'b00000000; //  814 :   0 - 0x0
      12'h32F: dout <= 8'b00000000; //  815 :   0 - 0x0
      12'h330: dout <= 8'b11100000; //  816 : 224 - 0xe0 -- Sprite 0x66
      12'h331: dout <= 8'b11100000; //  817 : 224 - 0xe0
      12'h332: dout <= 8'b11100000; //  818 : 224 - 0xe0
      12'h333: dout <= 8'b11101110; //  819 : 238 - 0xee
      12'h334: dout <= 8'b11111110; //  820 : 254 - 0xfe
      12'h335: dout <= 8'b11111110; //  821 : 254 - 0xfe
      12'h336: dout <= 8'b00000000; //  822 :   0 - 0x0
      12'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      12'h338: dout <= 8'b11101110; //  824 : 238 - 0xee -- Sprite 0x67
      12'h339: dout <= 8'b11101110; //  825 : 238 - 0xee
      12'h33A: dout <= 8'b11111110; //  826 : 254 - 0xfe
      12'h33B: dout <= 8'b11111110; //  827 : 254 - 0xfe
      12'h33C: dout <= 8'b11101110; //  828 : 238 - 0xee
      12'h33D: dout <= 8'b11000110; //  829 : 198 - 0xc6
      12'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout <= 8'b11101110; //  832 : 238 - 0xee -- Sprite 0x68
      12'h341: dout <= 8'b11101110; //  833 : 238 - 0xee
      12'h342: dout <= 8'b11101110; //  834 : 238 - 0xee
      12'h343: dout <= 8'b11101110; //  835 : 238 - 0xee
      12'h344: dout <= 8'b11101110; //  836 : 238 - 0xee
      12'h345: dout <= 8'b11101110; //  837 : 238 - 0xee
      12'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      12'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout <= 8'b11101110; //  840 : 238 - 0xee -- Sprite 0x69
      12'h349: dout <= 8'b11101110; //  841 : 238 - 0xee
      12'h34A: dout <= 8'b11101110; //  842 : 238 - 0xee
      12'h34B: dout <= 8'b11101110; //  843 : 238 - 0xee
      12'h34C: dout <= 8'b11111110; //  844 : 254 - 0xfe
      12'h34D: dout <= 8'b11111100; //  845 : 252 - 0xfc
      12'h34E: dout <= 8'b00000000; //  846 :   0 - 0x0
      12'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout <= 8'b11101110; //  848 : 238 - 0xee -- Sprite 0x6a
      12'h351: dout <= 8'b11101110; //  849 : 238 - 0xee
      12'h352: dout <= 8'b11101110; //  850 : 238 - 0xee
      12'h353: dout <= 8'b11101110; //  851 : 238 - 0xee
      12'h354: dout <= 8'b11111110; //  852 : 254 - 0xfe
      12'h355: dout <= 8'b01111100; //  853 : 124 - 0x7c
      12'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout <= 8'b11100000; //  856 : 224 - 0xe0 -- Sprite 0x6b
      12'h359: dout <= 8'b11100000; //  857 : 224 - 0xe0
      12'h35A: dout <= 8'b11100000; //  858 : 224 - 0xe0
      12'h35B: dout <= 8'b11100000; //  859 : 224 - 0xe0
      12'h35C: dout <= 8'b11111110; //  860 : 254 - 0xfe
      12'h35D: dout <= 8'b11111110; //  861 : 254 - 0xfe
      12'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout <= 8'b00011000; //  864 :  24 - 0x18 -- Sprite 0x6c
      12'h361: dout <= 8'b00011000; //  865 :  24 - 0x18
      12'h362: dout <= 8'b00110000; //  866 :  48 - 0x30
      12'h363: dout <= 8'b00110000; //  867 :  48 - 0x30
      12'h364: dout <= 8'b01100110; //  868 : 102 - 0x66
      12'h365: dout <= 8'b01100110; //  869 : 102 - 0x66
      12'h366: dout <= 8'b00000000; //  870 :   0 - 0x0
      12'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      12'h368: dout <= 8'b11100000; //  872 : 224 - 0xe0 -- Sprite 0x6d
      12'h369: dout <= 8'b11100000; //  873 : 224 - 0xe0
      12'h36A: dout <= 8'b11100000; //  874 : 224 - 0xe0
      12'h36B: dout <= 8'b11100000; //  875 : 224 - 0xe0
      12'h36C: dout <= 8'b11100000; //  876 : 224 - 0xe0
      12'h36D: dout <= 8'b11100000; //  877 : 224 - 0xe0
      12'h36E: dout <= 8'b00000000; //  878 :   0 - 0x0
      12'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout <= 8'b11101110; //  880 : 238 - 0xee -- Sprite 0x6e
      12'h371: dout <= 8'b11101110; //  881 : 238 - 0xee
      12'h372: dout <= 8'b11101110; //  882 : 238 - 0xee
      12'h373: dout <= 8'b11101110; //  883 : 238 - 0xee
      12'h374: dout <= 8'b11111110; //  884 : 254 - 0xfe
      12'h375: dout <= 8'b01111100; //  885 : 124 - 0x7c
      12'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout <= 8'b01111110; //  888 : 126 - 0x7e -- Sprite 0x6f
      12'h379: dout <= 8'b01111110; //  889 : 126 - 0x7e
      12'h37A: dout <= 8'b01111110; //  890 : 126 - 0x7e
      12'h37B: dout <= 8'b01111110; //  891 : 126 - 0x7e
      12'h37C: dout <= 8'b00111100; //  892 :  60 - 0x3c
      12'h37D: dout <= 8'b00111100; //  893 :  60 - 0x3c
      12'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b00000111; //  896 :   7 - 0x7 -- Sprite 0x70
      12'h381: dout <= 8'b00011111; //  897 :  31 - 0x1f
      12'h382: dout <= 8'b00111111; //  898 :  63 - 0x3f
      12'h383: dout <= 8'b00111111; //  899 :  63 - 0x3f
      12'h384: dout <= 8'b01111111; //  900 : 127 - 0x7f
      12'h385: dout <= 8'b01111111; //  901 : 127 - 0x7f
      12'h386: dout <= 8'b01111111; //  902 : 127 - 0x7f
      12'h387: dout <= 8'b01111110; //  903 : 126 - 0x7e
      12'h388: dout <= 8'b11100000; //  904 : 224 - 0xe0 -- Sprite 0x71
      12'h389: dout <= 8'b11111000; //  905 : 248 - 0xf8
      12'h38A: dout <= 8'b11111100; //  906 : 252 - 0xfc
      12'h38B: dout <= 8'b11111100; //  907 : 252 - 0xfc
      12'h38C: dout <= 8'b11111110; //  908 : 254 - 0xfe
      12'h38D: dout <= 8'b11111110; //  909 : 254 - 0xfe
      12'h38E: dout <= 8'b11111110; //  910 : 254 - 0xfe
      12'h38F: dout <= 8'b01111110; //  911 : 126 - 0x7e
      12'h390: dout <= 8'b01111110; //  912 : 126 - 0x7e -- Sprite 0x72
      12'h391: dout <= 8'b01111110; //  913 : 126 - 0x7e
      12'h392: dout <= 8'b01111110; //  914 : 126 - 0x7e
      12'h393: dout <= 8'b01111110; //  915 : 126 - 0x7e
      12'h394: dout <= 8'b01111110; //  916 : 126 - 0x7e
      12'h395: dout <= 8'b01111110; //  917 : 126 - 0x7e
      12'h396: dout <= 8'b01111110; //  918 : 126 - 0x7e
      12'h397: dout <= 8'b01111110; //  919 : 126 - 0x7e
      12'h398: dout <= 8'b01111110; //  920 : 126 - 0x7e -- Sprite 0x73
      12'h399: dout <= 8'b01111111; //  921 : 127 - 0x7f
      12'h39A: dout <= 8'b01111111; //  922 : 127 - 0x7f
      12'h39B: dout <= 8'b01111111; //  923 : 127 - 0x7f
      12'h39C: dout <= 8'b00111111; //  924 :  63 - 0x3f
      12'h39D: dout <= 8'b00111111; //  925 :  63 - 0x3f
      12'h39E: dout <= 8'b00011111; //  926 :  31 - 0x1f
      12'h39F: dout <= 8'b00000111; //  927 :   7 - 0x7
      12'h3A0: dout <= 8'b01111110; //  928 : 126 - 0x7e -- Sprite 0x74
      12'h3A1: dout <= 8'b11111110; //  929 : 254 - 0xfe
      12'h3A2: dout <= 8'b11111110; //  930 : 254 - 0xfe
      12'h3A3: dout <= 8'b11111110; //  931 : 254 - 0xfe
      12'h3A4: dout <= 8'b11111100; //  932 : 252 - 0xfc
      12'h3A5: dout <= 8'b11111100; //  933 : 252 - 0xfc
      12'h3A6: dout <= 8'b11111000; //  934 : 248 - 0xf8
      12'h3A7: dout <= 8'b11100000; //  935 : 224 - 0xe0
      12'h3A8: dout <= 8'b01111111; //  936 : 127 - 0x7f -- Sprite 0x75
      12'h3A9: dout <= 8'b01111111; //  937 : 127 - 0x7f
      12'h3AA: dout <= 8'b01111111; //  938 : 127 - 0x7f
      12'h3AB: dout <= 8'b01111111; //  939 : 127 - 0x7f
      12'h3AC: dout <= 8'b01111111; //  940 : 127 - 0x7f
      12'h3AD: dout <= 8'b01111111; //  941 : 127 - 0x7f
      12'h3AE: dout <= 8'b00000111; //  942 :   7 - 0x7
      12'h3AF: dout <= 8'b00000111; //  943 :   7 - 0x7
      12'h3B0: dout <= 8'b11111110; //  944 : 254 - 0xfe -- Sprite 0x76
      12'h3B1: dout <= 8'b11111110; //  945 : 254 - 0xfe
      12'h3B2: dout <= 8'b11111110; //  946 : 254 - 0xfe
      12'h3B3: dout <= 8'b11111110; //  947 : 254 - 0xfe
      12'h3B4: dout <= 8'b11111110; //  948 : 254 - 0xfe
      12'h3B5: dout <= 8'b11111110; //  949 : 254 - 0xfe
      12'h3B6: dout <= 8'b11100000; //  950 : 224 - 0xe0
      12'h3B7: dout <= 8'b11100000; //  951 : 224 - 0xe0
      12'h3B8: dout <= 8'b00000111; //  952 :   7 - 0x7 -- Sprite 0x77
      12'h3B9: dout <= 8'b00000111; //  953 :   7 - 0x7
      12'h3BA: dout <= 8'b00000111; //  954 :   7 - 0x7
      12'h3BB: dout <= 8'b00000111; //  955 :   7 - 0x7
      12'h3BC: dout <= 8'b00000111; //  956 :   7 - 0x7
      12'h3BD: dout <= 8'b00000111; //  957 :   7 - 0x7
      12'h3BE: dout <= 8'b00000111; //  958 :   7 - 0x7
      12'h3BF: dout <= 8'b00000111; //  959 :   7 - 0x7
      12'h3C0: dout <= 8'b11100000; //  960 : 224 - 0xe0 -- Sprite 0x78
      12'h3C1: dout <= 8'b11100000; //  961 : 224 - 0xe0
      12'h3C2: dout <= 8'b11100000; //  962 : 224 - 0xe0
      12'h3C3: dout <= 8'b11100000; //  963 : 224 - 0xe0
      12'h3C4: dout <= 8'b11100000; //  964 : 224 - 0xe0
      12'h3C5: dout <= 8'b11100000; //  965 : 224 - 0xe0
      12'h3C6: dout <= 8'b11100000; //  966 : 224 - 0xe0
      12'h3C7: dout <= 8'b11100000; //  967 : 224 - 0xe0
      12'h3C8: dout <= 8'b01111111; //  968 : 127 - 0x7f -- Sprite 0x79
      12'h3C9: dout <= 8'b01111111; //  969 : 127 - 0x7f
      12'h3CA: dout <= 8'b01111111; //  970 : 127 - 0x7f
      12'h3CB: dout <= 8'b01111111; //  971 : 127 - 0x7f
      12'h3CC: dout <= 8'b01111111; //  972 : 127 - 0x7f
      12'h3CD: dout <= 8'b01111111; //  973 : 127 - 0x7f
      12'h3CE: dout <= 8'b01111110; //  974 : 126 - 0x7e
      12'h3CF: dout <= 8'b01111110; //  975 : 126 - 0x7e
      12'h3D0: dout <= 8'b11111110; //  976 : 254 - 0xfe -- Sprite 0x7a
      12'h3D1: dout <= 8'b11111110; //  977 : 254 - 0xfe
      12'h3D2: dout <= 8'b11111110; //  978 : 254 - 0xfe
      12'h3D3: dout <= 8'b11111110; //  979 : 254 - 0xfe
      12'h3D4: dout <= 8'b11111110; //  980 : 254 - 0xfe
      12'h3D5: dout <= 8'b11111110; //  981 : 254 - 0xfe
      12'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout <= 8'b01111110; //  984 : 126 - 0x7e -- Sprite 0x7b
      12'h3D9: dout <= 8'b01111111; //  985 : 127 - 0x7f
      12'h3DA: dout <= 8'b01111111; //  986 : 127 - 0x7f
      12'h3DB: dout <= 8'b01111111; //  987 : 127 - 0x7f
      12'h3DC: dout <= 8'b01111111; //  988 : 127 - 0x7f
      12'h3DD: dout <= 8'b01111111; //  989 : 127 - 0x7f
      12'h3DE: dout <= 8'b01111111; //  990 : 127 - 0x7f
      12'h3DF: dout <= 8'b01111110; //  991 : 126 - 0x7e
      12'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      12'h3E1: dout <= 8'b11110000; //  993 : 240 - 0xf0
      12'h3E2: dout <= 8'b11110000; //  994 : 240 - 0xf0
      12'h3E3: dout <= 8'b11110000; //  995 : 240 - 0xf0
      12'h3E4: dout <= 8'b11110000; //  996 : 240 - 0xf0
      12'h3E5: dout <= 8'b11110000; //  997 : 240 - 0xf0
      12'h3E6: dout <= 8'b11110000; //  998 : 240 - 0xf0
      12'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      12'h3E8: dout <= 8'b01111110; // 1000 : 126 - 0x7e -- Sprite 0x7d
      12'h3E9: dout <= 8'b01111110; // 1001 : 126 - 0x7e
      12'h3EA: dout <= 8'b01111111; // 1002 : 127 - 0x7f
      12'h3EB: dout <= 8'b01111111; // 1003 : 127 - 0x7f
      12'h3EC: dout <= 8'b01111111; // 1004 : 127 - 0x7f
      12'h3ED: dout <= 8'b01111111; // 1005 : 127 - 0x7f
      12'h3EE: dout <= 8'b01111111; // 1006 : 127 - 0x7f
      12'h3EF: dout <= 8'b01111111; // 1007 : 127 - 0x7f
      12'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x7e
      12'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout <= 8'b11111110; // 1010 : 254 - 0xfe
      12'h3F3: dout <= 8'b11111110; // 1011 : 254 - 0xfe
      12'h3F4: dout <= 8'b11111110; // 1012 : 254 - 0xfe
      12'h3F5: dout <= 8'b11111110; // 1013 : 254 - 0xfe
      12'h3F6: dout <= 8'b11111110; // 1014 : 254 - 0xfe
      12'h3F7: dout <= 8'b11111110; // 1015 : 254 - 0xfe
      12'h3F8: dout <= 8'b01111110; // 1016 : 126 - 0x7e -- Sprite 0x7f
      12'h3F9: dout <= 8'b11111110; // 1017 : 254 - 0xfe
      12'h3FA: dout <= 8'b11111110; // 1018 : 254 - 0xfe
      12'h3FB: dout <= 8'b11111110; // 1019 : 254 - 0xfe
      12'h3FC: dout <= 8'b11111110; // 1020 : 254 - 0xfe
      12'h3FD: dout <= 8'b11111110; // 1021 : 254 - 0xfe
      12'h3FE: dout <= 8'b11111110; // 1022 : 254 - 0xfe
      12'h3FF: dout <= 8'b01111110; // 1023 : 126 - 0x7e
      12'h400: dout <= 8'b01000000; // 1024 :  64 - 0x40 -- Sprite 0x80
      12'h401: dout <= 8'b00001000; // 1025 :   8 - 0x8
      12'h402: dout <= 8'b00000010; // 1026 :   2 - 0x2
      12'h403: dout <= 8'b00100000; // 1027 :  32 - 0x20
      12'h404: dout <= 8'b00000100; // 1028 :   4 - 0x4
      12'h405: dout <= 8'b01000000; // 1029 :  64 - 0x40
      12'h406: dout <= 8'b00000001; // 1030 :   1 - 0x1
      12'h407: dout <= 8'b00010000; // 1031 :  16 - 0x10
      12'h408: dout <= 8'b00000000; // 1032 :   0 - 0x0 -- Sprite 0x81
      12'h409: dout <= 8'b00010001; // 1033 :  17 - 0x11
      12'h40A: dout <= 8'b00000000; // 1034 :   0 - 0x0
      12'h40B: dout <= 8'b00100000; // 1035 :  32 - 0x20
      12'h40C: dout <= 8'b10001000; // 1036 : 136 - 0x88
      12'h40D: dout <= 8'b00000010; // 1037 :   2 - 0x2
      12'h40E: dout <= 8'b00100000; // 1038 :  32 - 0x20
      12'h40F: dout <= 8'b01000000; // 1039 :  64 - 0x40
      12'h410: dout <= 8'b00000001; // 1040 :   1 - 0x1 -- Sprite 0x82
      12'h411: dout <= 8'b00010000; // 1041 :  16 - 0x10
      12'h412: dout <= 8'b01000000; // 1042 :  64 - 0x40
      12'h413: dout <= 8'b00001000; // 1043 :   8 - 0x8
      12'h414: dout <= 8'b00000010; // 1044 :   2 - 0x2
      12'h415: dout <= 8'b00100000; // 1045 :  32 - 0x20
      12'h416: dout <= 8'b00000100; // 1046 :   4 - 0x4
      12'h417: dout <= 8'b01000000; // 1047 :  64 - 0x40
      12'h418: dout <= 8'b00010000; // 1048 :  16 - 0x10 -- Sprite 0x83
      12'h419: dout <= 8'b00000000; // 1049 :   0 - 0x0
      12'h41A: dout <= 8'b01000100; // 1050 :  68 - 0x44
      12'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      12'h41C: dout <= 8'b00001000; // 1052 :   8 - 0x8
      12'h41D: dout <= 8'b00100010; // 1053 :  34 - 0x22
      12'h41E: dout <= 8'b10000000; // 1054 : 128 - 0x80
      12'h41F: dout <= 8'b00001000; // 1055 :   8 - 0x8
      12'h420: dout <= 8'b00010100; // 1056 :  20 - 0x14 -- Sprite 0x84
      12'h421: dout <= 8'b10110101; // 1057 : 181 - 0xb5
      12'h422: dout <= 8'b01000100; // 1058 :  68 - 0x44
      12'h423: dout <= 8'b01001010; // 1059 :  74 - 0x4a
      12'h424: dout <= 8'b10010010; // 1060 : 146 - 0x92
      12'h425: dout <= 8'b10010010; // 1061 : 146 - 0x92
      12'h426: dout <= 8'b01000100; // 1062 :  68 - 0x44
      12'h427: dout <= 8'b01001001; // 1063 :  73 - 0x49
      12'h428: dout <= 8'b01000010; // 1064 :  66 - 0x42 -- Sprite 0x85
      12'h429: dout <= 8'b01001010; // 1065 :  74 - 0x4a
      12'h42A: dout <= 8'b11001010; // 1066 : 202 - 0xca
      12'h42B: dout <= 8'b00101001; // 1067 :  41 - 0x29
      12'h42C: dout <= 8'b10100110; // 1068 : 166 - 0xa6
      12'h42D: dout <= 8'b10010010; // 1069 : 146 - 0x92
      12'h42E: dout <= 8'b10001001; // 1070 : 137 - 0x89
      12'h42F: dout <= 8'b00101101; // 1071 :  45 - 0x2d
      12'h430: dout <= 8'b10001000; // 1072 : 136 - 0x88 -- Sprite 0x86
      12'h431: dout <= 8'b00101001; // 1073 :  41 - 0x29
      12'h432: dout <= 8'b10000010; // 1074 : 130 - 0x82
      12'h433: dout <= 8'b10110110; // 1075 : 182 - 0xb6
      12'h434: dout <= 8'b10001000; // 1076 : 136 - 0x88
      12'h435: dout <= 8'b01001001; // 1077 :  73 - 0x49
      12'h436: dout <= 8'b01010010; // 1078 :  82 - 0x52
      12'h437: dout <= 8'b01010010; // 1079 :  82 - 0x52
      12'h438: dout <= 8'b10110010; // 1080 : 178 - 0xb2 -- Sprite 0x87
      12'h439: dout <= 8'b01001010; // 1081 :  74 - 0x4a
      12'h43A: dout <= 8'b10101001; // 1082 : 169 - 0xa9
      12'h43B: dout <= 8'b10100100; // 1083 : 164 - 0xa4
      12'h43C: dout <= 8'b01100010; // 1084 :  98 - 0x62
      12'h43D: dout <= 8'b01001011; // 1085 :  75 - 0x4b
      12'h43E: dout <= 8'b10010000; // 1086 : 144 - 0x90
      12'h43F: dout <= 8'b10010010; // 1087 : 146 - 0x92
      12'h440: dout <= 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x88
      12'h441: dout <= 8'b01100000; // 1089 :  96 - 0x60
      12'h442: dout <= 8'b11111110; // 1090 : 254 - 0xfe
      12'h443: dout <= 8'b11111111; // 1091 : 255 - 0xff
      12'h444: dout <= 8'b01111111; // 1092 : 127 - 0x7f
      12'h445: dout <= 8'b00011111; // 1093 :  31 - 0x1f
      12'h446: dout <= 8'b00001110; // 1094 :  14 - 0xe
      12'h447: dout <= 8'b00000000; // 1095 :   0 - 0x0
      12'h448: dout <= 8'b00110000; // 1096 :  48 - 0x30 -- Sprite 0x89
      12'h449: dout <= 8'b01111000; // 1097 : 120 - 0x78
      12'h44A: dout <= 8'b01111000; // 1098 : 120 - 0x78
      12'h44B: dout <= 8'b00111110; // 1099 :  62 - 0x3e
      12'h44C: dout <= 8'b00011111; // 1100 :  31 - 0x1f
      12'h44D: dout <= 8'b00011111; // 1101 :  31 - 0x1f
      12'h44E: dout <= 8'b00011111; // 1102 :  31 - 0x1f
      12'h44F: dout <= 8'b00001110; // 1103 :  14 - 0xe
      12'h450: dout <= 8'b01000000; // 1104 :  64 - 0x40 -- Sprite 0x8a
      12'h451: dout <= 8'b00001000; // 1105 :   8 - 0x8
      12'h452: dout <= 8'b00000010; // 1106 :   2 - 0x2
      12'h453: dout <= 8'b00101000; // 1107 :  40 - 0x28
      12'h454: dout <= 8'b00010100; // 1108 :  20 - 0x14
      12'h455: dout <= 8'b01010100; // 1109 :  84 - 0x54
      12'h456: dout <= 8'b00000001; // 1110 :   1 - 0x1
      12'h457: dout <= 8'b00010000; // 1111 :  16 - 0x10
      12'h458: dout <= 8'b01000000; // 1112 :  64 - 0x40 -- Sprite 0x8b
      12'h459: dout <= 8'b00000000; // 1113 :   0 - 0x0
      12'h45A: dout <= 8'b10010001; // 1114 : 145 - 0x91
      12'h45B: dout <= 8'b00010100; // 1115 :  20 - 0x14
      12'h45C: dout <= 8'b00101000; // 1116 :  40 - 0x28
      12'h45D: dout <= 8'b10001010; // 1117 : 138 - 0x8a
      12'h45E: dout <= 8'b01000000; // 1118 :  64 - 0x40
      12'h45F: dout <= 8'b00100000; // 1119 :  32 - 0x20
      12'h460: dout <= 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x8c
      12'h461: dout <= 8'b00000111; // 1121 :   7 - 0x7
      12'h462: dout <= 8'b00011111; // 1122 :  31 - 0x1f
      12'h463: dout <= 8'b00111111; // 1123 :  63 - 0x3f
      12'h464: dout <= 8'b00111111; // 1124 :  63 - 0x3f
      12'h465: dout <= 8'b01111111; // 1125 : 127 - 0x7f
      12'h466: dout <= 8'b01111111; // 1126 : 127 - 0x7f
      12'h467: dout <= 8'b01111111; // 1127 : 127 - 0x7f
      12'h468: dout <= 8'b00000000; // 1128 :   0 - 0x0 -- Sprite 0x8d
      12'h469: dout <= 8'b11100000; // 1129 : 224 - 0xe0
      12'h46A: dout <= 8'b11111000; // 1130 : 248 - 0xf8
      12'h46B: dout <= 8'b11111000; // 1131 : 248 - 0xf8
      12'h46C: dout <= 8'b11110000; // 1132 : 240 - 0xf0
      12'h46D: dout <= 8'b11111000; // 1133 : 248 - 0xf8
      12'h46E: dout <= 8'b11110100; // 1134 : 244 - 0xf4
      12'h46F: dout <= 8'b11111000; // 1135 : 248 - 0xf8
      12'h470: dout <= 8'b01111111; // 1136 : 127 - 0x7f -- Sprite 0x8e
      12'h471: dout <= 8'b00111111; // 1137 :  63 - 0x3f
      12'h472: dout <= 8'b00111111; // 1138 :  63 - 0x3f
      12'h473: dout <= 8'b00011111; // 1139 :  31 - 0x1f
      12'h474: dout <= 8'b00011111; // 1140 :  31 - 0x1f
      12'h475: dout <= 8'b00001111; // 1141 :  15 - 0xf
      12'h476: dout <= 8'b00001111; // 1142 :  15 - 0xf
      12'h477: dout <= 8'b00000111; // 1143 :   7 - 0x7
      12'h478: dout <= 8'b11111110; // 1144 : 254 - 0xfe -- Sprite 0x8f
      12'h479: dout <= 8'b11111100; // 1145 : 252 - 0xfc
      12'h47A: dout <= 8'b11111100; // 1146 : 252 - 0xfc
      12'h47B: dout <= 8'b11111000; // 1147 : 248 - 0xf8
      12'h47C: dout <= 8'b11111000; // 1148 : 248 - 0xf8
      12'h47D: dout <= 8'b11110000; // 1149 : 240 - 0xf0
      12'h47E: dout <= 8'b11110000; // 1150 : 240 - 0xf0
      12'h47F: dout <= 8'b11100000; // 1151 : 224 - 0xe0
      12'h480: dout <= 8'b01000001; // 1152 :  65 - 0x41 -- Sprite 0x90
      12'h481: dout <= 8'b00001000; // 1153 :   8 - 0x8
      12'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      12'h483: dout <= 8'b00100000; // 1155 :  32 - 0x20
      12'h484: dout <= 8'b00000100; // 1156 :   4 - 0x4
      12'h485: dout <= 8'b00000001; // 1157 :   1 - 0x1
      12'h486: dout <= 8'b01000000; // 1158 :  64 - 0x40
      12'h487: dout <= 8'b00001000; // 1159 :   8 - 0x8
      12'h488: dout <= 8'b00010001; // 1160 :  17 - 0x11 -- Sprite 0x91
      12'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      12'h48A: dout <= 8'b10000100; // 1162 : 132 - 0x84
      12'h48B: dout <= 8'b00000010; // 1163 :   2 - 0x2
      12'h48C: dout <= 8'b00010000; // 1164 :  16 - 0x10
      12'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      12'h48E: dout <= 8'b01000010; // 1166 :  66 - 0x42
      12'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout <= 8'b00000100; // 1168 :   4 - 0x4 -- Sprite 0x92
      12'h491: dout <= 8'b01000000; // 1169 :  64 - 0x40
      12'h492: dout <= 8'b00010000; // 1170 :  16 - 0x10
      12'h493: dout <= 8'b00000010; // 1171 :   2 - 0x2
      12'h494: dout <= 8'b00000000; // 1172 :   0 - 0x0
      12'h495: dout <= 8'b01000000; // 1173 :  64 - 0x40
      12'h496: dout <= 8'b00000100; // 1174 :   4 - 0x4
      12'h497: dout <= 8'b00100000; // 1175 :  32 - 0x20
      12'h498: dout <= 8'b01000010; // 1176 :  66 - 0x42 -- Sprite 0x93
      12'h499: dout <= 8'b00000000; // 1177 :   0 - 0x0
      12'h49A: dout <= 8'b10001000; // 1178 : 136 - 0x88
      12'h49B: dout <= 8'b00000001; // 1179 :   1 - 0x1
      12'h49C: dout <= 8'b00100000; // 1180 :  32 - 0x20
      12'h49D: dout <= 8'b00000100; // 1181 :   4 - 0x4
      12'h49E: dout <= 8'b00010000; // 1182 :  16 - 0x10
      12'h49F: dout <= 8'b10000000; // 1183 : 128 - 0x80
      12'h4A0: dout <= 8'b11001000; // 1184 : 200 - 0xc8 -- Sprite 0x94
      12'h4A1: dout <= 8'b00101010; // 1185 :  42 - 0x2a
      12'h4A2: dout <= 8'b10100010; // 1186 : 162 - 0xa2
      12'h4A3: dout <= 8'b10010100; // 1187 : 148 - 0x94
      12'h4A4: dout <= 8'b10010001; // 1188 : 145 - 0x91
      12'h4A5: dout <= 8'b01010101; // 1189 :  85 - 0x55
      12'h4A6: dout <= 8'b01000100; // 1190 :  68 - 0x44
      12'h4A7: dout <= 8'b00010010; // 1191 :  18 - 0x12
      12'h4A8: dout <= 8'b10101010; // 1192 : 170 - 0xaa -- Sprite 0x95
      12'h4A9: dout <= 8'b10100010; // 1193 : 162 - 0xa2
      12'h4AA: dout <= 8'b00010010; // 1194 :  18 - 0x12
      12'h4AB: dout <= 8'b01010011; // 1195 :  83 - 0x53
      12'h4AC: dout <= 8'b01001100; // 1196 :  76 - 0x4c
      12'h4AD: dout <= 8'b01010101; // 1197 :  85 - 0x55
      12'h4AE: dout <= 8'b10010001; // 1198 : 145 - 0x91
      12'h4AF: dout <= 8'b01001000; // 1199 :  72 - 0x48
      12'h4B0: dout <= 8'b01010001; // 1200 :  81 - 0x51 -- Sprite 0x96
      12'h4B1: dout <= 8'b00010101; // 1201 :  21 - 0x15
      12'h4B2: dout <= 8'b10100100; // 1202 : 164 - 0xa4
      12'h4B3: dout <= 8'b10001100; // 1203 : 140 - 0x8c
      12'h4B4: dout <= 8'b10101010; // 1204 : 170 - 0xaa
      12'h4B5: dout <= 8'b00100010; // 1205 :  34 - 0x22
      12'h4B6: dout <= 8'b10010000; // 1206 : 144 - 0x90
      12'h4B7: dout <= 8'b01000110; // 1207 :  70 - 0x46
      12'h4B8: dout <= 8'b00010011; // 1208 :  19 - 0x13 -- Sprite 0x97
      12'h4B9: dout <= 8'b01010101; // 1209 :  85 - 0x55
      12'h4BA: dout <= 8'b01100100; // 1210 : 100 - 0x64
      12'h4BB: dout <= 8'b00010010; // 1211 :  18 - 0x12
      12'h4BC: dout <= 8'b10101010; // 1212 : 170 - 0xaa
      12'h4BD: dout <= 8'b10101000; // 1213 : 168 - 0xa8
      12'h4BE: dout <= 8'b10000100; // 1214 : 132 - 0x84
      12'h4BF: dout <= 8'b11010100; // 1215 : 212 - 0xd4
      12'h4C0: dout <= 8'b00110000; // 1216 :  48 - 0x30 -- Sprite 0x98
      12'h4C1: dout <= 8'b01111000; // 1217 : 120 - 0x78
      12'h4C2: dout <= 8'b01111000; // 1218 : 120 - 0x78
      12'h4C3: dout <= 8'b00111110; // 1219 :  62 - 0x3e
      12'h4C4: dout <= 8'b00011111; // 1220 :  31 - 0x1f
      12'h4C5: dout <= 8'b00011111; // 1221 :  31 - 0x1f
      12'h4C6: dout <= 8'b00011111; // 1222 :  31 - 0x1f
      12'h4C7: dout <= 8'b00001110; // 1223 :  14 - 0xe
      12'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0 -- Sprite 0x99
      12'h4C9: dout <= 8'b01100000; // 1225 :  96 - 0x60
      12'h4CA: dout <= 8'b11111110; // 1226 : 254 - 0xfe
      12'h4CB: dout <= 8'b11111111; // 1227 : 255 - 0xff
      12'h4CC: dout <= 8'b01111111; // 1228 : 127 - 0x7f
      12'h4CD: dout <= 8'b00011111; // 1229 :  31 - 0x1f
      12'h4CE: dout <= 8'b00001110; // 1230 :  14 - 0xe
      12'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      12'h4D0: dout <= 8'b01000000; // 1232 :  64 - 0x40 -- Sprite 0x9a
      12'h4D1: dout <= 8'b00001100; // 1233 :  12 - 0xc
      12'h4D2: dout <= 8'b00000000; // 1234 :   0 - 0x0
      12'h4D3: dout <= 8'b00101000; // 1235 :  40 - 0x28
      12'h4D4: dout <= 8'b00101100; // 1236 :  44 - 0x2c
      12'h4D5: dout <= 8'b00010001; // 1237 :  17 - 0x11
      12'h4D6: dout <= 8'b01000000; // 1238 :  64 - 0x40
      12'h4D7: dout <= 8'b00001000; // 1239 :   8 - 0x8
      12'h4D8: dout <= 8'b00100000; // 1240 :  32 - 0x20 -- Sprite 0x9b
      12'h4D9: dout <= 8'b00000000; // 1241 :   0 - 0x0
      12'h4DA: dout <= 8'b10010100; // 1242 : 148 - 0x94
      12'h4DB: dout <= 8'b01001000; // 1243 :  72 - 0x48
      12'h4DC: dout <= 8'b00011000; // 1244 :  24 - 0x18
      12'h4DD: dout <= 8'b00000110; // 1245 :   6 - 0x6
      12'h4DE: dout <= 8'b01000000; // 1246 :  64 - 0x40
      12'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout <= 8'b01111111; // 1248 : 127 - 0x7f -- Sprite 0x9c
      12'h4E1: dout <= 8'b01111111; // 1249 : 127 - 0x7f
      12'h4E2: dout <= 8'b01111111; // 1250 : 127 - 0x7f
      12'h4E3: dout <= 8'b00111111; // 1251 :  63 - 0x3f
      12'h4E4: dout <= 8'b00110101; // 1252 :  53 - 0x35
      12'h4E5: dout <= 8'b00000010; // 1253 :   2 - 0x2
      12'h4E6: dout <= 8'b00000000; // 1254 :   0 - 0x0
      12'h4E7: dout <= 8'b00000000; // 1255 :   0 - 0x0
      12'h4E8: dout <= 8'b11110100; // 1256 : 244 - 0xf4 -- Sprite 0x9d
      12'h4E9: dout <= 8'b11111000; // 1257 : 248 - 0xf8
      12'h4EA: dout <= 8'b11110000; // 1258 : 240 - 0xf0
      12'h4EB: dout <= 8'b11101000; // 1259 : 232 - 0xe8
      12'h4EC: dout <= 8'b01010000; // 1260 :  80 - 0x50
      12'h4ED: dout <= 8'b10000000; // 1261 : 128 - 0x80
      12'h4EE: dout <= 8'b00000000; // 1262 :   0 - 0x0
      12'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout <= 8'b11111110; // 1264 : 254 - 0xfe -- Sprite 0x9e
      12'h4F1: dout <= 8'b11111100; // 1265 : 252 - 0xfc
      12'h4F2: dout <= 8'b11111100; // 1266 : 252 - 0xfc
      12'h4F3: dout <= 8'b11111000; // 1267 : 248 - 0xf8
      12'h4F4: dout <= 8'b11111000; // 1268 : 248 - 0xf8
      12'h4F5: dout <= 8'b11111100; // 1269 : 252 - 0xfc
      12'h4F6: dout <= 8'b11111100; // 1270 : 252 - 0xfc
      12'h4F7: dout <= 8'b11111110; // 1271 : 254 - 0xfe
      12'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0 -- Sprite 0x9f
      12'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout <= 8'b01111110; // 1274 : 126 - 0x7e
      12'h4FB: dout <= 8'b01111110; // 1275 : 126 - 0x7e
      12'h4FC: dout <= 8'b01111110; // 1276 : 126 - 0x7e
      12'h4FD: dout <= 8'b01111110; // 1277 : 126 - 0x7e
      12'h4FE: dout <= 8'b01111110; // 1278 : 126 - 0x7e
      12'h4FF: dout <= 8'b01111110; // 1279 : 126 - 0x7e
      12'h500: dout <= 8'b00010000; // 1280 :  16 - 0x10 -- Sprite 0xa0
      12'h501: dout <= 8'b00111000; // 1281 :  56 - 0x38
      12'h502: dout <= 8'b01111100; // 1282 : 124 - 0x7c
      12'h503: dout <= 8'b11111000; // 1283 : 248 - 0xf8
      12'h504: dout <= 8'b01110000; // 1284 : 112 - 0x70
      12'h505: dout <= 8'b00100010; // 1285 :  34 - 0x22
      12'h506: dout <= 8'b00000101; // 1286 :   5 - 0x5
      12'h507: dout <= 8'b00000010; // 1287 :   2 - 0x2
      12'h508: dout <= 8'b00010000; // 1288 :  16 - 0x10 -- Sprite 0xa1
      12'h509: dout <= 8'b00111000; // 1289 :  56 - 0x38
      12'h50A: dout <= 8'b01111100; // 1290 : 124 - 0x7c
      12'h50B: dout <= 8'b11100000; // 1291 : 224 - 0xe0
      12'h50C: dout <= 8'b01100000; // 1292 :  96 - 0x60
      12'h50D: dout <= 8'b00100000; // 1293 :  32 - 0x20
      12'h50E: dout <= 8'b00000000; // 1294 :   0 - 0x0
      12'h50F: dout <= 8'b00000000; // 1295 :   0 - 0x0
      12'h510: dout <= 8'b00010000; // 1296 :  16 - 0x10 -- Sprite 0xa2
      12'h511: dout <= 8'b00111000; // 1297 :  56 - 0x38
      12'h512: dout <= 8'b01111100; // 1298 : 124 - 0x7c
      12'h513: dout <= 8'b00000000; // 1299 :   0 - 0x0
      12'h514: dout <= 8'b00000000; // 1300 :   0 - 0x0
      12'h515: dout <= 8'b00000000; // 1301 :   0 - 0x0
      12'h516: dout <= 8'b00000000; // 1302 :   0 - 0x0
      12'h517: dout <= 8'b00000000; // 1303 :   0 - 0x0
      12'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0 -- Sprite 0xa3
      12'h519: dout <= 8'b00100000; // 1305 :  32 - 0x20
      12'h51A: dout <= 8'b01100000; // 1306 :  96 - 0x60
      12'h51B: dout <= 8'b11100000; // 1307 : 224 - 0xe0
      12'h51C: dout <= 8'b01100000; // 1308 :  96 - 0x60
      12'h51D: dout <= 8'b00100000; // 1309 :  32 - 0x20
      12'h51E: dout <= 8'b00000000; // 1310 :   0 - 0x0
      12'h51F: dout <= 8'b00000000; // 1311 :   0 - 0x0
      12'h520: dout <= 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0xa4
      12'h521: dout <= 8'b00100000; // 1313 :  32 - 0x20
      12'h522: dout <= 8'b01100011; // 1314 :  99 - 0x63
      12'h523: dout <= 8'b11100111; // 1315 : 231 - 0xe7
      12'h524: dout <= 8'b01100000; // 1316 :  96 - 0x60
      12'h525: dout <= 8'b00100010; // 1317 :  34 - 0x22
      12'h526: dout <= 8'b00000101; // 1318 :   5 - 0x5
      12'h527: dout <= 8'b00000010; // 1319 :   2 - 0x2
      12'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0 -- Sprite 0xa5
      12'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      12'h52A: dout <= 8'b11111111; // 1322 : 255 - 0xff
      12'h52B: dout <= 8'b11111111; // 1323 : 255 - 0xff
      12'h52C: dout <= 8'b00000000; // 1324 :   0 - 0x0
      12'h52D: dout <= 8'b00100010; // 1325 :  34 - 0x22
      12'h52E: dout <= 8'b00000101; // 1326 :   5 - 0x5
      12'h52F: dout <= 8'b00000010; // 1327 :   2 - 0x2
      12'h530: dout <= 8'b00010000; // 1328 :  16 - 0x10 -- Sprite 0xa6
      12'h531: dout <= 8'b00111000; // 1329 :  56 - 0x38
      12'h532: dout <= 8'b01111100; // 1330 : 124 - 0x7c
      12'h533: dout <= 8'b00000000; // 1331 :   0 - 0x0
      12'h534: dout <= 8'b00000000; // 1332 :   0 - 0x0
      12'h535: dout <= 8'b00010010; // 1333 :  18 - 0x12
      12'h536: dout <= 8'b00110101; // 1334 :  53 - 0x35
      12'h537: dout <= 8'b00110010; // 1335 :  50 - 0x32
      12'h538: dout <= 8'b00110000; // 1336 :  48 - 0x30 -- Sprite 0xa7
      12'h539: dout <= 8'b00110000; // 1337 :  48 - 0x30
      12'h53A: dout <= 8'b00110100; // 1338 :  52 - 0x34
      12'h53B: dout <= 8'b00110000; // 1339 :  48 - 0x30
      12'h53C: dout <= 8'b00110000; // 1340 :  48 - 0x30
      12'h53D: dout <= 8'b00110010; // 1341 :  50 - 0x32
      12'h53E: dout <= 8'b00110101; // 1342 :  53 - 0x35
      12'h53F: dout <= 8'b00110010; // 1343 :  50 - 0x32
      12'h540: dout <= 8'b00110000; // 1344 :  48 - 0x30 -- Sprite 0xa8
      12'h541: dout <= 8'b00110000; // 1345 :  48 - 0x30
      12'h542: dout <= 8'b11110100; // 1346 : 244 - 0xf4
      12'h543: dout <= 8'b11110000; // 1347 : 240 - 0xf0
      12'h544: dout <= 8'b00000000; // 1348 :   0 - 0x0
      12'h545: dout <= 8'b00100010; // 1349 :  34 - 0x22
      12'h546: dout <= 8'b00000101; // 1350 :   5 - 0x5
      12'h547: dout <= 8'b00000010; // 1351 :   2 - 0x2
      12'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0 -- Sprite 0xa9
      12'h549: dout <= 8'b00000000; // 1353 :   0 - 0x0
      12'h54A: dout <= 8'b00000000; // 1354 :   0 - 0x0
      12'h54B: dout <= 8'b00000000; // 1355 :   0 - 0x0
      12'h54C: dout <= 8'b00000000; // 1356 :   0 - 0x0
      12'h54D: dout <= 8'b00000000; // 1357 :   0 - 0x0
      12'h54E: dout <= 8'b00000000; // 1358 :   0 - 0x0
      12'h54F: dout <= 8'b00000000; // 1359 :   0 - 0x0
      12'h550: dout <= 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      12'h551: dout <= 8'b00000000; // 1361 :   0 - 0x0
      12'h552: dout <= 8'b01010000; // 1362 :  80 - 0x50
      12'h553: dout <= 8'b10101000; // 1363 : 168 - 0xa8
      12'h554: dout <= 8'b01110000; // 1364 : 112 - 0x70
      12'h555: dout <= 8'b00100010; // 1365 :  34 - 0x22
      12'h556: dout <= 8'b00000101; // 1366 :   5 - 0x5
      12'h557: dout <= 8'b00000010; // 1367 :   2 - 0x2
      12'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0 -- Sprite 0xab
      12'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      12'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      12'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      12'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      12'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      12'h560: dout <= 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      12'h561: dout <= 8'b00000000; // 1377 :   0 - 0x0
      12'h562: dout <= 8'b00000000; // 1378 :   0 - 0x0
      12'h563: dout <= 8'b00000000; // 1379 :   0 - 0x0
      12'h564: dout <= 8'b00000000; // 1380 :   0 - 0x0
      12'h565: dout <= 8'b00000000; // 1381 :   0 - 0x0
      12'h566: dout <= 8'b00000000; // 1382 :   0 - 0x0
      12'h567: dout <= 8'b00000000; // 1383 :   0 - 0x0
      12'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0 -- Sprite 0xad
      12'h569: dout <= 8'b00000000; // 1385 :   0 - 0x0
      12'h56A: dout <= 8'b11111111; // 1386 : 255 - 0xff
      12'h56B: dout <= 8'b00000000; // 1387 :   0 - 0x0
      12'h56C: dout <= 8'b00000000; // 1388 :   0 - 0x0
      12'h56D: dout <= 8'b00000000; // 1389 :   0 - 0x0
      12'h56E: dout <= 8'b00000000; // 1390 :   0 - 0x0
      12'h56F: dout <= 8'b00000000; // 1391 :   0 - 0x0
      12'h570: dout <= 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      12'h571: dout <= 8'b00000000; // 1393 :   0 - 0x0
      12'h572: dout <= 8'b00000000; // 1394 :   0 - 0x0
      12'h573: dout <= 8'b00000000; // 1395 :   0 - 0x0
      12'h574: dout <= 8'b00000000; // 1396 :   0 - 0x0
      12'h575: dout <= 8'b11111111; // 1397 : 255 - 0xff
      12'h576: dout <= 8'b00000000; // 1398 :   0 - 0x0
      12'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0 -- Sprite 0xaf
      12'h579: dout <= 8'b00000000; // 1401 :   0 - 0x0
      12'h57A: dout <= 8'b00000000; // 1402 :   0 - 0x0
      12'h57B: dout <= 8'b00000000; // 1403 :   0 - 0x0
      12'h57C: dout <= 8'b00000000; // 1404 :   0 - 0x0
      12'h57D: dout <= 8'b00000000; // 1405 :   0 - 0x0
      12'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      12'h57F: dout <= 8'b00000000; // 1407 :   0 - 0x0
      12'h580: dout <= 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      12'h581: dout <= 8'b00011111; // 1409 :  31 - 0x1f
      12'h582: dout <= 8'b00011111; // 1410 :  31 - 0x1f
      12'h583: dout <= 8'b00011111; // 1411 :  31 - 0x1f
      12'h584: dout <= 8'b00011111; // 1412 :  31 - 0x1f
      12'h585: dout <= 8'b00011111; // 1413 :  31 - 0x1f
      12'h586: dout <= 8'b00011111; // 1414 :  31 - 0x1f
      12'h587: dout <= 8'b00011111; // 1415 :  31 - 0x1f
      12'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0 -- Sprite 0xb1
      12'h589: dout <= 8'b11110000; // 1417 : 240 - 0xf0
      12'h58A: dout <= 8'b11110000; // 1418 : 240 - 0xf0
      12'h58B: dout <= 8'b11110000; // 1419 : 240 - 0xf0
      12'h58C: dout <= 8'b11110000; // 1420 : 240 - 0xf0
      12'h58D: dout <= 8'b11110000; // 1421 : 240 - 0xf0
      12'h58E: dout <= 8'b11110000; // 1422 : 240 - 0xf0
      12'h58F: dout <= 8'b11110000; // 1423 : 240 - 0xf0
      12'h590: dout <= 8'b00011111; // 1424 :  31 - 0x1f -- Sprite 0xb2
      12'h591: dout <= 8'b00011111; // 1425 :  31 - 0x1f
      12'h592: dout <= 8'b00011111; // 1426 :  31 - 0x1f
      12'h593: dout <= 8'b00011111; // 1427 :  31 - 0x1f
      12'h594: dout <= 8'b00000000; // 1428 :   0 - 0x0
      12'h595: dout <= 8'b00000000; // 1429 :   0 - 0x0
      12'h596: dout <= 8'b00000000; // 1430 :   0 - 0x0
      12'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      12'h598: dout <= 8'b11110000; // 1432 : 240 - 0xf0 -- Sprite 0xb3
      12'h599: dout <= 8'b11110000; // 1433 : 240 - 0xf0
      12'h59A: dout <= 8'b11110000; // 1434 : 240 - 0xf0
      12'h59B: dout <= 8'b11110000; // 1435 : 240 - 0xf0
      12'h59C: dout <= 8'b00000000; // 1436 :   0 - 0x0
      12'h59D: dout <= 8'b00000000; // 1437 :   0 - 0x0
      12'h59E: dout <= 8'b00000000; // 1438 :   0 - 0x0
      12'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout <= 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0xb4
      12'h5A1: dout <= 8'b00000000; // 1441 :   0 - 0x0
      12'h5A2: dout <= 8'b00111111; // 1442 :  63 - 0x3f
      12'h5A3: dout <= 8'b01111111; // 1443 : 127 - 0x7f
      12'h5A4: dout <= 8'b01111111; // 1444 : 127 - 0x7f
      12'h5A5: dout <= 8'b01111111; // 1445 : 127 - 0x7f
      12'h5A6: dout <= 8'b01111111; // 1446 : 127 - 0x7f
      12'h5A7: dout <= 8'b01111111; // 1447 : 127 - 0x7f
      12'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0 -- Sprite 0xb5
      12'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      12'h5AA: dout <= 8'b11111000; // 1450 : 248 - 0xf8
      12'h5AB: dout <= 8'b11111000; // 1451 : 248 - 0xf8
      12'h5AC: dout <= 8'b11111000; // 1452 : 248 - 0xf8
      12'h5AD: dout <= 8'b11111000; // 1453 : 248 - 0xf8
      12'h5AE: dout <= 8'b11111000; // 1454 : 248 - 0xf8
      12'h5AF: dout <= 8'b11111000; // 1455 : 248 - 0xf8
      12'h5B0: dout <= 8'b01111111; // 1456 : 127 - 0x7f -- Sprite 0xb6
      12'h5B1: dout <= 8'b01111111; // 1457 : 127 - 0x7f
      12'h5B2: dout <= 8'b01111111; // 1458 : 127 - 0x7f
      12'h5B3: dout <= 8'b01000000; // 1459 :  64 - 0x40
      12'h5B4: dout <= 8'b00000000; // 1460 :   0 - 0x0
      12'h5B5: dout <= 8'b00000000; // 1461 :   0 - 0x0
      12'h5B6: dout <= 8'b00000000; // 1462 :   0 - 0x0
      12'h5B7: dout <= 8'b00000000; // 1463 :   0 - 0x0
      12'h5B8: dout <= 8'b11111000; // 1464 : 248 - 0xf8 -- Sprite 0xb7
      12'h5B9: dout <= 8'b11111000; // 1465 : 248 - 0xf8
      12'h5BA: dout <= 8'b11111000; // 1466 : 248 - 0xf8
      12'h5BB: dout <= 8'b00000000; // 1467 :   0 - 0x0
      12'h5BC: dout <= 8'b00000000; // 1468 :   0 - 0x0
      12'h5BD: dout <= 8'b00000000; // 1469 :   0 - 0x0
      12'h5BE: dout <= 8'b00000000; // 1470 :   0 - 0x0
      12'h5BF: dout <= 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout <= 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0xb8
      12'h5C1: dout <= 8'b00000011; // 1473 :   3 - 0x3
      12'h5C2: dout <= 8'b00000111; // 1474 :   7 - 0x7
      12'h5C3: dout <= 8'b00000111; // 1475 :   7 - 0x7
      12'h5C4: dout <= 8'b00000111; // 1476 :   7 - 0x7
      12'h5C5: dout <= 8'b00000011; // 1477 :   3 - 0x3
      12'h5C6: dout <= 8'b00000000; // 1478 :   0 - 0x0
      12'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout <= 8'b00000000; // 1480 :   0 - 0x0 -- Sprite 0xb9
      12'h5C9: dout <= 8'b11000001; // 1481 : 193 - 0xc1
      12'h5CA: dout <= 8'b11100010; // 1482 : 226 - 0xe2
      12'h5CB: dout <= 8'b11001100; // 1483 : 204 - 0xcc
      12'h5CC: dout <= 8'b11000000; // 1484 : 192 - 0xc0
      12'h5CD: dout <= 8'b10000000; // 1485 : 128 - 0x80
      12'h5CE: dout <= 8'b00000001; // 1486 :   1 - 0x1
      12'h5CF: dout <= 8'b00000010; // 1487 :   2 - 0x2
      12'h5D0: dout <= 8'b11110000; // 1488 : 240 - 0xf0 -- Sprite 0xba
      12'h5D1: dout <= 8'b00000000; // 1489 :   0 - 0x0
      12'h5D2: dout <= 8'b00100000; // 1490 :  32 - 0x20
      12'h5D3: dout <= 8'b00100000; // 1491 :  32 - 0x20
      12'h5D4: dout <= 8'b00000000; // 1492 :   0 - 0x0
      12'h5D5: dout <= 8'b11110000; // 1493 : 240 - 0xf0
      12'h5D6: dout <= 8'b00000000; // 1494 :   0 - 0x0
      12'h5D7: dout <= 8'b00000000; // 1495 :   0 - 0x0
      12'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0 -- Sprite 0xbb
      12'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      12'h5DB: dout <= 8'b00000000; // 1499 :   0 - 0x0
      12'h5DC: dout <= 8'b00000000; // 1500 :   0 - 0x0
      12'h5DD: dout <= 8'b01100000; // 1501 :  96 - 0x60
      12'h5DE: dout <= 8'b01100000; // 1502 :  96 - 0x60
      12'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout <= 8'b00001100; // 1504 :  12 - 0xc -- Sprite 0xbc
      12'h5E1: dout <= 8'b00000000; // 1505 :   0 - 0x0
      12'h5E2: dout <= 8'b00000000; // 1506 :   0 - 0x0
      12'h5E3: dout <= 8'b00000000; // 1507 :   0 - 0x0
      12'h5E4: dout <= 8'b00000000; // 1508 :   0 - 0x0
      12'h5E5: dout <= 8'b00000110; // 1509 :   6 - 0x6
      12'h5E6: dout <= 8'b00000110; // 1510 :   6 - 0x6
      12'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0 -- Sprite 0xbd
      12'h5E9: dout <= 8'b10000011; // 1513 : 131 - 0x83
      12'h5EA: dout <= 8'b00000111; // 1514 :   7 - 0x7
      12'h5EB: dout <= 8'b00000111; // 1515 :   7 - 0x7
      12'h5EC: dout <= 8'b00000111; // 1516 :   7 - 0x7
      12'h5ED: dout <= 8'b00000011; // 1517 :   3 - 0x3
      12'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      12'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout <= 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      12'h5F1: dout <= 8'b11000100; // 1521 : 196 - 0xc4
      12'h5F2: dout <= 8'b11100000; // 1522 : 224 - 0xe0
      12'h5F3: dout <= 8'b11000000; // 1523 : 192 - 0xc0
      12'h5F4: dout <= 8'b11000000; // 1524 : 192 - 0xc0
      12'h5F5: dout <= 8'b10000000; // 1525 : 128 - 0x80
      12'h5F6: dout <= 8'b00000000; // 1526 :   0 - 0x0
      12'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      12'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      12'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      12'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      12'h5FC: dout <= 8'b00001000; // 1532 :   8 - 0x8
      12'h5FD: dout <= 8'b10001000; // 1533 : 136 - 0x88
      12'h5FE: dout <= 8'b00001011; // 1534 :  11 - 0xb
      12'h5FF: dout <= 8'b00001000; // 1535 :   8 - 0x8
      12'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      12'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout <= 8'b00000000; // 1538 :   0 - 0x0
      12'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      12'h604: dout <= 8'b00100000; // 1540 :  32 - 0x20
      12'h605: dout <= 8'b00100100; // 1541 :  36 - 0x24
      12'h606: dout <= 8'b10100000; // 1542 : 160 - 0xa0
      12'h607: dout <= 8'b00100000; // 1543 :  32 - 0x20
      12'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0 -- Sprite 0xc1
      12'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      12'h60A: dout <= 8'b00000000; // 1546 :   0 - 0x0
      12'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      12'h60C: dout <= 8'b00000000; // 1548 :   0 - 0x0
      12'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      12'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      12'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      12'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      12'h612: dout <= 8'b00000000; // 1554 :   0 - 0x0
      12'h613: dout <= 8'b00000000; // 1555 :   0 - 0x0
      12'h614: dout <= 8'b00000000; // 1556 :   0 - 0x0
      12'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      12'h616: dout <= 8'b00000000; // 1558 :   0 - 0x0
      12'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      12'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0 -- Sprite 0xc3
      12'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      12'h61A: dout <= 8'b00001000; // 1562 :   8 - 0x8
      12'h61B: dout <= 8'b00001011; // 1563 :  11 - 0xb
      12'h61C: dout <= 8'b00001000; // 1564 :   8 - 0x8
      12'h61D: dout <= 8'b00001000; // 1565 :   8 - 0x8
      12'h61E: dout <= 8'b00001000; // 1566 :   8 - 0x8
      12'h61F: dout <= 8'b00001000; // 1567 :   8 - 0x8
      12'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      12'h621: dout <= 8'b00000000; // 1569 :   0 - 0x0
      12'h622: dout <= 8'b00100000; // 1570 :  32 - 0x20
      12'h623: dout <= 8'b10100000; // 1571 : 160 - 0xa0
      12'h624: dout <= 8'b00100000; // 1572 :  32 - 0x20
      12'h625: dout <= 8'b00100000; // 1573 :  32 - 0x20
      12'h626: dout <= 8'b00100000; // 1574 :  32 - 0x20
      12'h627: dout <= 8'b00100000; // 1575 :  32 - 0x20
      12'h628: dout <= 8'b00001000; // 1576 :   8 - 0x8 -- Sprite 0xc5
      12'h629: dout <= 8'b11001000; // 1577 : 200 - 0xc8
      12'h62A: dout <= 8'b00000011; // 1578 :   3 - 0x3
      12'h62B: dout <= 8'b00000111; // 1579 :   7 - 0x7
      12'h62C: dout <= 8'b00000111; // 1580 :   7 - 0x7
      12'h62D: dout <= 8'b00000111; // 1581 :   7 - 0x7
      12'h62E: dout <= 8'b00000011; // 1582 :   3 - 0x3
      12'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout <= 8'b00100000; // 1584 :  32 - 0x20 -- Sprite 0xc6
      12'h631: dout <= 8'b00100110; // 1585 :  38 - 0x26
      12'h632: dout <= 8'b11000000; // 1586 : 192 - 0xc0
      12'h633: dout <= 8'b11100000; // 1587 : 224 - 0xe0
      12'h634: dout <= 8'b11000000; // 1588 : 192 - 0xc0
      12'h635: dout <= 8'b11000000; // 1589 : 192 - 0xc0
      12'h636: dout <= 8'b10000000; // 1590 : 128 - 0x80
      12'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      12'h638: dout <= 8'b00000000; // 1592 :   0 - 0x0 -- Sprite 0xc7
      12'h639: dout <= 8'b00000000; // 1593 :   0 - 0x0
      12'h63A: dout <= 8'b00000000; // 1594 :   0 - 0x0
      12'h63B: dout <= 8'b00000000; // 1595 :   0 - 0x0
      12'h63C: dout <= 8'b00000000; // 1596 :   0 - 0x0
      12'h63D: dout <= 8'b11000000; // 1597 : 192 - 0xc0
      12'h63E: dout <= 8'b00000000; // 1598 :   0 - 0x0
      12'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      12'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      12'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      12'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      12'h644: dout <= 8'b00000000; // 1604 :   0 - 0x0
      12'h645: dout <= 8'b00000110; // 1605 :   6 - 0x6
      12'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      12'h647: dout <= 8'b00000000; // 1607 :   0 - 0x0
      12'h648: dout <= 8'b00001111; // 1608 :  15 - 0xf -- Sprite 0xc9
      12'h649: dout <= 8'b00000000; // 1609 :   0 - 0x0
      12'h64A: dout <= 8'b00001000; // 1610 :   8 - 0x8
      12'h64B: dout <= 8'b00001000; // 1611 :   8 - 0x8
      12'h64C: dout <= 8'b00000000; // 1612 :   0 - 0x0
      12'h64D: dout <= 8'b00001111; // 1613 :  15 - 0xf
      12'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      12'h651: dout <= 8'b10000011; // 1617 : 131 - 0x83
      12'h652: dout <= 8'b01000111; // 1618 :  71 - 0x47
      12'h653: dout <= 8'b00110111; // 1619 :  55 - 0x37
      12'h654: dout <= 8'b00000111; // 1620 :   7 - 0x7
      12'h655: dout <= 8'b00000011; // 1621 :   3 - 0x3
      12'h656: dout <= 8'b10000000; // 1622 : 128 - 0x80
      12'h657: dout <= 8'b01000000; // 1623 :  64 - 0x40
      12'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- Sprite 0xcb
      12'h659: dout <= 8'b11000000; // 1625 : 192 - 0xc0
      12'h65A: dout <= 8'b11100000; // 1626 : 224 - 0xe0
      12'h65B: dout <= 8'b11000000; // 1627 : 192 - 0xc0
      12'h65C: dout <= 8'b11000000; // 1628 : 192 - 0xc0
      12'h65D: dout <= 8'b10000000; // 1629 : 128 - 0x80
      12'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout <= 8'b00110000; // 1632 :  48 - 0x30 -- Sprite 0xcc
      12'h661: dout <= 8'b00000000; // 1633 :   0 - 0x0
      12'h662: dout <= 8'b00000000; // 1634 :   0 - 0x0
      12'h663: dout <= 8'b00000000; // 1635 :   0 - 0x0
      12'h664: dout <= 8'b00000000; // 1636 :   0 - 0x0
      12'h665: dout <= 8'b01100000; // 1637 :  96 - 0x60
      12'h666: dout <= 8'b01100000; // 1638 :  96 - 0x60
      12'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      12'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- Sprite 0xcd
      12'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout <= 8'b00000000; // 1643 :   0 - 0x0
      12'h66C: dout <= 8'b00000000; // 1644 :   0 - 0x0
      12'h66D: dout <= 8'b00000110; // 1645 :   6 - 0x6
      12'h66E: dout <= 8'b00000110; // 1646 :   6 - 0x6
      12'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      12'h670: dout <= 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      12'h671: dout <= 8'b00000001; // 1649 :   1 - 0x1
      12'h672: dout <= 8'b00011011; // 1650 :  27 - 0x1b
      12'h673: dout <= 8'b00010011; // 1651 :  19 - 0x13
      12'h674: dout <= 8'b00011111; // 1652 :  31 - 0x1f
      12'h675: dout <= 8'b00111111; // 1653 :  63 - 0x3f
      12'h676: dout <= 8'b00111111; // 1654 :  63 - 0x3f
      12'h677: dout <= 8'b00111111; // 1655 :  63 - 0x3f
      12'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- Sprite 0xcf
      12'h679: dout <= 8'b11111000; // 1657 : 248 - 0xf8
      12'h67A: dout <= 8'b00001000; // 1658 :   8 - 0x8
      12'h67B: dout <= 8'b00001000; // 1659 :   8 - 0x8
      12'h67C: dout <= 8'b00001000; // 1660 :   8 - 0x8
      12'h67D: dout <= 8'b11111000; // 1661 : 248 - 0xf8
      12'h67E: dout <= 8'b11110000; // 1662 : 240 - 0xf0
      12'h67F: dout <= 8'b11010000; // 1663 : 208 - 0xd0
      12'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      12'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout <= 8'b01111100; // 1666 : 124 - 0x7c
      12'h683: dout <= 8'b11111110; // 1667 : 254 - 0xfe
      12'h684: dout <= 8'b11101110; // 1668 : 238 - 0xee
      12'h685: dout <= 8'b11101110; // 1669 : 238 - 0xee
      12'h686: dout <= 8'b11101110; // 1670 : 238 - 0xee
      12'h687: dout <= 8'b11101110; // 1671 : 238 - 0xee
      12'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- Sprite 0xd1
      12'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      12'h68A: dout <= 8'b00111000; // 1674 :  56 - 0x38
      12'h68B: dout <= 8'b01111000; // 1675 : 120 - 0x78
      12'h68C: dout <= 8'b01111000; // 1676 : 120 - 0x78
      12'h68D: dout <= 8'b00111000; // 1677 :  56 - 0x38
      12'h68E: dout <= 8'b00111000; // 1678 :  56 - 0x38
      12'h68F: dout <= 8'b00111000; // 1679 :  56 - 0x38
      12'h690: dout <= 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0xd2
      12'h691: dout <= 8'b00000000; // 1681 :   0 - 0x0
      12'h692: dout <= 8'b01111100; // 1682 : 124 - 0x7c
      12'h693: dout <= 8'b11111110; // 1683 : 254 - 0xfe
      12'h694: dout <= 8'b11101110; // 1684 : 238 - 0xee
      12'h695: dout <= 8'b00001110; // 1685 :  14 - 0xe
      12'h696: dout <= 8'b00001110; // 1686 :  14 - 0xe
      12'h697: dout <= 8'b01111110; // 1687 : 126 - 0x7e
      12'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0 -- Sprite 0xd3
      12'h699: dout <= 8'b00000000; // 1689 :   0 - 0x0
      12'h69A: dout <= 8'b01111100; // 1690 : 124 - 0x7c
      12'h69B: dout <= 8'b11111110; // 1691 : 254 - 0xfe
      12'h69C: dout <= 8'b11101110; // 1692 : 238 - 0xee
      12'h69D: dout <= 8'b00001110; // 1693 :  14 - 0xe
      12'h69E: dout <= 8'b00111100; // 1694 :  60 - 0x3c
      12'h69F: dout <= 8'b00111100; // 1695 :  60 - 0x3c
      12'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      12'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout <= 8'b00111110; // 1698 :  62 - 0x3e
      12'h6A3: dout <= 8'b01111110; // 1699 : 126 - 0x7e
      12'h6A4: dout <= 8'b11101110; // 1700 : 238 - 0xee
      12'h6A5: dout <= 8'b11101110; // 1701 : 238 - 0xee
      12'h6A6: dout <= 8'b11101110; // 1702 : 238 - 0xee
      12'h6A7: dout <= 8'b11101110; // 1703 : 238 - 0xee
      12'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0 -- Sprite 0xd5
      12'h6A9: dout <= 8'b00000000; // 1705 :   0 - 0x0
      12'h6AA: dout <= 8'b11111100; // 1706 : 252 - 0xfc
      12'h6AB: dout <= 8'b11111100; // 1707 : 252 - 0xfc
      12'h6AC: dout <= 8'b11100000; // 1708 : 224 - 0xe0
      12'h6AD: dout <= 8'b11100000; // 1709 : 224 - 0xe0
      12'h6AE: dout <= 8'b11111100; // 1710 : 252 - 0xfc
      12'h6AF: dout <= 8'b11111110; // 1711 : 254 - 0xfe
      12'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      12'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout <= 8'b01111100; // 1714 : 124 - 0x7c
      12'h6B3: dout <= 8'b11111100; // 1715 : 252 - 0xfc
      12'h6B4: dout <= 8'b11100000; // 1716 : 224 - 0xe0
      12'h6B5: dout <= 8'b11100000; // 1717 : 224 - 0xe0
      12'h6B6: dout <= 8'b11111100; // 1718 : 252 - 0xfc
      12'h6B7: dout <= 8'b11111110; // 1719 : 254 - 0xfe
      12'h6B8: dout <= 8'b00000000; // 1720 :   0 - 0x0 -- Sprite 0xd7
      12'h6B9: dout <= 8'b00000000; // 1721 :   0 - 0x0
      12'h6BA: dout <= 8'b11111110; // 1722 : 254 - 0xfe
      12'h6BB: dout <= 8'b11111110; // 1723 : 254 - 0xfe
      12'h6BC: dout <= 8'b11101110; // 1724 : 238 - 0xee
      12'h6BD: dout <= 8'b00001110; // 1725 :  14 - 0xe
      12'h6BE: dout <= 8'b00001110; // 1726 :  14 - 0xe
      12'h6BF: dout <= 8'b00011100; // 1727 :  28 - 0x1c
      12'h6C0: dout <= 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0xd8
      12'h6C1: dout <= 8'b00000000; // 1729 :   0 - 0x0
      12'h6C2: dout <= 8'b01111100; // 1730 : 124 - 0x7c
      12'h6C3: dout <= 8'b11111110; // 1731 : 254 - 0xfe
      12'h6C4: dout <= 8'b11101110; // 1732 : 238 - 0xee
      12'h6C5: dout <= 8'b11101110; // 1733 : 238 - 0xee
      12'h6C6: dout <= 8'b01111100; // 1734 : 124 - 0x7c
      12'h6C7: dout <= 8'b11111110; // 1735 : 254 - 0xfe
      12'h6C8: dout <= 8'b00000000; // 1736 :   0 - 0x0 -- Sprite 0xd9
      12'h6C9: dout <= 8'b00000000; // 1737 :   0 - 0x0
      12'h6CA: dout <= 8'b01111100; // 1738 : 124 - 0x7c
      12'h6CB: dout <= 8'b11111110; // 1739 : 254 - 0xfe
      12'h6CC: dout <= 8'b11101110; // 1740 : 238 - 0xee
      12'h6CD: dout <= 8'b11101110; // 1741 : 238 - 0xee
      12'h6CE: dout <= 8'b11101110; // 1742 : 238 - 0xee
      12'h6CF: dout <= 8'b11101110; // 1743 : 238 - 0xee
      12'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0xda
      12'h6D1: dout <= 8'b00100000; // 1745 :  32 - 0x20
      12'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      12'h6D3: dout <= 8'b00000010; // 1747 :   2 - 0x2
      12'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      12'h6D5: dout <= 8'b00100000; // 1749 :  32 - 0x20
      12'h6D6: dout <= 8'b00000000; // 1750 :   0 - 0x0
      12'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      12'h6D8: dout <= 8'b00100000; // 1752 :  32 - 0x20 -- Sprite 0xdb
      12'h6D9: dout <= 8'b00000000; // 1753 :   0 - 0x0
      12'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      12'h6DB: dout <= 8'b00000000; // 1755 :   0 - 0x0
      12'h6DC: dout <= 8'b10000000; // 1756 : 128 - 0x80
      12'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      12'h6DE: dout <= 8'b00000100; // 1758 :   4 - 0x4
      12'h6DF: dout <= 8'b00000000; // 1759 :   0 - 0x0
      12'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0xdc
      12'h6E1: dout <= 8'b00001000; // 1761 :   8 - 0x8
      12'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout <= 8'b00000010; // 1764 :   2 - 0x2
      12'h6E5: dout <= 8'b00000000; // 1765 :   0 - 0x0
      12'h6E6: dout <= 8'b01000000; // 1766 :  64 - 0x40
      12'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      12'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- Sprite 0xdd
      12'h6E9: dout <= 8'b01000000; // 1769 :  64 - 0x40
      12'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      12'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      12'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      12'h6ED: dout <= 8'b00000000; // 1773 :   0 - 0x0
      12'h6EE: dout <= 8'b00000010; // 1774 :   2 - 0x2
      12'h6EF: dout <= 8'b00100000; // 1775 :  32 - 0x20
      12'h6F0: dout <= 8'b00111110; // 1776 :  62 - 0x3e -- Sprite 0xde
      12'h6F1: dout <= 8'b00111111; // 1777 :  63 - 0x3f
      12'h6F2: dout <= 8'b00111110; // 1778 :  62 - 0x3e
      12'h6F3: dout <= 8'b00111100; // 1779 :  60 - 0x3c
      12'h6F4: dout <= 8'b00111111; // 1780 :  63 - 0x3f
      12'h6F5: dout <= 8'b00110000; // 1781 :  48 - 0x30
      12'h6F6: dout <= 8'b00000000; // 1782 :   0 - 0x0
      12'h6F7: dout <= 8'b00000000; // 1783 :   0 - 0x0
      12'h6F8: dout <= 8'b00010000; // 1784 :  16 - 0x10 -- Sprite 0xdf
      12'h6F9: dout <= 8'b10110000; // 1785 : 176 - 0xb0
      12'h6FA: dout <= 8'b00110000; // 1786 :  48 - 0x30
      12'h6FB: dout <= 8'b11110000; // 1787 : 240 - 0xf0
      12'h6FC: dout <= 8'b11110000; // 1788 : 240 - 0xf0
      12'h6FD: dout <= 8'b00000000; // 1789 :   0 - 0x0
      12'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      12'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout <= 8'b11101110; // 1792 : 238 - 0xee -- Sprite 0xe0
      12'h701: dout <= 8'b11101110; // 1793 : 238 - 0xee
      12'h702: dout <= 8'b11101110; // 1794 : 238 - 0xee
      12'h703: dout <= 8'b11101110; // 1795 : 238 - 0xee
      12'h704: dout <= 8'b11111110; // 1796 : 254 - 0xfe
      12'h705: dout <= 8'b01111100; // 1797 : 124 - 0x7c
      12'h706: dout <= 8'b00000000; // 1798 :   0 - 0x0
      12'h707: dout <= 8'b00000000; // 1799 :   0 - 0x0
      12'h708: dout <= 8'b00111000; // 1800 :  56 - 0x38 -- Sprite 0xe1
      12'h709: dout <= 8'b00111000; // 1801 :  56 - 0x38
      12'h70A: dout <= 8'b00111000; // 1802 :  56 - 0x38
      12'h70B: dout <= 8'b00111000; // 1803 :  56 - 0x38
      12'h70C: dout <= 8'b01111100; // 1804 : 124 - 0x7c
      12'h70D: dout <= 8'b01111100; // 1805 : 124 - 0x7c
      12'h70E: dout <= 8'b00000000; // 1806 :   0 - 0x0
      12'h70F: dout <= 8'b00000000; // 1807 :   0 - 0x0
      12'h710: dout <= 8'b11111100; // 1808 : 252 - 0xfc -- Sprite 0xe2
      12'h711: dout <= 8'b11100000; // 1809 : 224 - 0xe0
      12'h712: dout <= 8'b11100000; // 1810 : 224 - 0xe0
      12'h713: dout <= 8'b11100000; // 1811 : 224 - 0xe0
      12'h714: dout <= 8'b11111110; // 1812 : 254 - 0xfe
      12'h715: dout <= 8'b11111110; // 1813 : 254 - 0xfe
      12'h716: dout <= 8'b00000000; // 1814 :   0 - 0x0
      12'h717: dout <= 8'b00000000; // 1815 :   0 - 0x0
      12'h718: dout <= 8'b00001110; // 1816 :  14 - 0xe -- Sprite 0xe3
      12'h719: dout <= 8'b00001110; // 1817 :  14 - 0xe
      12'h71A: dout <= 8'b00001110; // 1818 :  14 - 0xe
      12'h71B: dout <= 8'b11101110; // 1819 : 238 - 0xee
      12'h71C: dout <= 8'b11111110; // 1820 : 254 - 0xfe
      12'h71D: dout <= 8'b01111100; // 1821 : 124 - 0x7c
      12'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      12'h720: dout <= 8'b11101110; // 1824 : 238 - 0xee -- Sprite 0xe4
      12'h721: dout <= 8'b11101110; // 1825 : 238 - 0xee
      12'h722: dout <= 8'b11111110; // 1826 : 254 - 0xfe
      12'h723: dout <= 8'b11111110; // 1827 : 254 - 0xfe
      12'h724: dout <= 8'b00001110; // 1828 :  14 - 0xe
      12'h725: dout <= 8'b00001110; // 1829 :  14 - 0xe
      12'h726: dout <= 8'b00000000; // 1830 :   0 - 0x0
      12'h727: dout <= 8'b00000000; // 1831 :   0 - 0x0
      12'h728: dout <= 8'b00001110; // 1832 :  14 - 0xe -- Sprite 0xe5
      12'h729: dout <= 8'b00001110; // 1833 :  14 - 0xe
      12'h72A: dout <= 8'b00001110; // 1834 :  14 - 0xe
      12'h72B: dout <= 8'b11101110; // 1835 : 238 - 0xee
      12'h72C: dout <= 8'b11111110; // 1836 : 254 - 0xfe
      12'h72D: dout <= 8'b01111100; // 1837 : 124 - 0x7c
      12'h72E: dout <= 8'b00000000; // 1838 :   0 - 0x0
      12'h72F: dout <= 8'b00000000; // 1839 :   0 - 0x0
      12'h730: dout <= 8'b11101110; // 1840 : 238 - 0xee -- Sprite 0xe6
      12'h731: dout <= 8'b11101110; // 1841 : 238 - 0xee
      12'h732: dout <= 8'b11101110; // 1842 : 238 - 0xee
      12'h733: dout <= 8'b11101110; // 1843 : 238 - 0xee
      12'h734: dout <= 8'b11111110; // 1844 : 254 - 0xfe
      12'h735: dout <= 8'b01111100; // 1845 : 124 - 0x7c
      12'h736: dout <= 8'b00000000; // 1846 :   0 - 0x0
      12'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      12'h738: dout <= 8'b00011100; // 1848 :  28 - 0x1c -- Sprite 0xe7
      12'h739: dout <= 8'b00011100; // 1849 :  28 - 0x1c
      12'h73A: dout <= 8'b00111000; // 1850 :  56 - 0x38
      12'h73B: dout <= 8'b00111000; // 1851 :  56 - 0x38
      12'h73C: dout <= 8'b00111000; // 1852 :  56 - 0x38
      12'h73D: dout <= 8'b00111000; // 1853 :  56 - 0x38
      12'h73E: dout <= 8'b00000000; // 1854 :   0 - 0x0
      12'h73F: dout <= 8'b00000000; // 1855 :   0 - 0x0
      12'h740: dout <= 8'b11101110; // 1856 : 238 - 0xee -- Sprite 0xe8
      12'h741: dout <= 8'b11101110; // 1857 : 238 - 0xee
      12'h742: dout <= 8'b11101110; // 1858 : 238 - 0xee
      12'h743: dout <= 8'b11101110; // 1859 : 238 - 0xee
      12'h744: dout <= 8'b11111110; // 1860 : 254 - 0xfe
      12'h745: dout <= 8'b01111100; // 1861 : 124 - 0x7c
      12'h746: dout <= 8'b00000000; // 1862 :   0 - 0x0
      12'h747: dout <= 8'b00000000; // 1863 :   0 - 0x0
      12'h748: dout <= 8'b11111110; // 1864 : 254 - 0xfe -- Sprite 0xe9
      12'h749: dout <= 8'b01111110; // 1865 : 126 - 0x7e
      12'h74A: dout <= 8'b00001110; // 1866 :  14 - 0xe
      12'h74B: dout <= 8'b00001110; // 1867 :  14 - 0xe
      12'h74C: dout <= 8'b01111110; // 1868 : 126 - 0x7e
      12'h74D: dout <= 8'b01111100; // 1869 : 124 - 0x7c
      12'h74E: dout <= 8'b00000000; // 1870 :   0 - 0x0
      12'h74F: dout <= 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0xea
      12'h751: dout <= 8'b01110000; // 1873 : 112 - 0x70
      12'h752: dout <= 8'b00111000; // 1874 :  56 - 0x38
      12'h753: dout <= 8'b00000000; // 1875 :   0 - 0x0
      12'h754: dout <= 8'b00000010; // 1876 :   2 - 0x2
      12'h755: dout <= 8'b00000111; // 1877 :   7 - 0x7
      12'h756: dout <= 8'b00000011; // 1878 :   3 - 0x3
      12'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout <= 8'b00000000; // 1880 :   0 - 0x0 -- Sprite 0xeb
      12'h759: dout <= 8'b00001100; // 1881 :  12 - 0xc
      12'h75A: dout <= 8'b00000110; // 1882 :   6 - 0x6
      12'h75B: dout <= 8'b00000110; // 1883 :   6 - 0x6
      12'h75C: dout <= 8'b01100000; // 1884 :  96 - 0x60
      12'h75D: dout <= 8'b01110000; // 1885 : 112 - 0x70
      12'h75E: dout <= 8'b00110000; // 1886 :  48 - 0x30
      12'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      12'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      12'h761: dout <= 8'b11000000; // 1889 : 192 - 0xc0
      12'h762: dout <= 8'b11100000; // 1890 : 224 - 0xe0
      12'h763: dout <= 8'b01100000; // 1891 :  96 - 0x60
      12'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      12'h765: dout <= 8'b00001100; // 1893 :  12 - 0xc
      12'h766: dout <= 8'b00001110; // 1894 :  14 - 0xe
      12'h767: dout <= 8'b00000110; // 1895 :   6 - 0x6
      12'h768: dout <= 8'b01100000; // 1896 :  96 - 0x60 -- Sprite 0xed
      12'h769: dout <= 8'b01110000; // 1897 : 112 - 0x70
      12'h76A: dout <= 8'b00110000; // 1898 :  48 - 0x30
      12'h76B: dout <= 8'b00000000; // 1899 :   0 - 0x0
      12'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      12'h76D: dout <= 8'b00001100; // 1901 :  12 - 0xc
      12'h76E: dout <= 8'b00001110; // 1902 :  14 - 0xe
      12'h76F: dout <= 8'b00000110; // 1903 :   6 - 0x6
      12'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0xee
      12'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout <= 8'b01000010; // 1906 :  66 - 0x42
      12'h773: dout <= 8'b00000000; // 1907 :   0 - 0x0
      12'h774: dout <= 8'b00000000; // 1908 :   0 - 0x0
      12'h775: dout <= 8'b00000100; // 1909 :   4 - 0x4
      12'h776: dout <= 8'b00000000; // 1910 :   0 - 0x0
      12'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      12'h778: dout <= 8'b00000000; // 1912 :   0 - 0x0 -- Sprite 0xef
      12'h779: dout <= 8'b00000000; // 1913 :   0 - 0x0
      12'h77A: dout <= 8'b00000100; // 1914 :   4 - 0x4
      12'h77B: dout <= 8'b00000000; // 1915 :   0 - 0x0
      12'h77C: dout <= 8'b00100000; // 1916 :  32 - 0x20
      12'h77D: dout <= 8'b00000000; // 1917 :   0 - 0x0
      12'h77E: dout <= 8'b00000000; // 1918 :   0 - 0x0
      12'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      12'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      12'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout <= 8'b10000000; // 1928 : 128 - 0x80 -- Sprite 0xf1
      12'h789: dout <= 8'b10000000; // 1929 : 128 - 0x80
      12'h78A: dout <= 8'b10000000; // 1930 : 128 - 0x80
      12'h78B: dout <= 8'b10000000; // 1931 : 128 - 0x80
      12'h78C: dout <= 8'b00000000; // 1932 :   0 - 0x0
      12'h78D: dout <= 8'b00000000; // 1933 :   0 - 0x0
      12'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      12'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout <= 8'b11000000; // 1936 : 192 - 0xc0 -- Sprite 0xf2
      12'h791: dout <= 8'b11000000; // 1937 : 192 - 0xc0
      12'h792: dout <= 8'b11000000; // 1938 : 192 - 0xc0
      12'h793: dout <= 8'b11000000; // 1939 : 192 - 0xc0
      12'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout <= 8'b11100000; // 1944 : 224 - 0xe0 -- Sprite 0xf3
      12'h799: dout <= 8'b11100000; // 1945 : 224 - 0xe0
      12'h79A: dout <= 8'b11100000; // 1946 : 224 - 0xe0
      12'h79B: dout <= 8'b11100000; // 1947 : 224 - 0xe0
      12'h79C: dout <= 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout <= 8'b00000000; // 1949 :   0 - 0x0
      12'h79E: dout <= 8'b00000000; // 1950 :   0 - 0x0
      12'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      12'h7A0: dout <= 8'b11110000; // 1952 : 240 - 0xf0 -- Sprite 0xf4
      12'h7A1: dout <= 8'b11110000; // 1953 : 240 - 0xf0
      12'h7A2: dout <= 8'b11110000; // 1954 : 240 - 0xf0
      12'h7A3: dout <= 8'b11110000; // 1955 : 240 - 0xf0
      12'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      12'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      12'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout <= 8'b11111000; // 1960 : 248 - 0xf8 -- Sprite 0xf5
      12'h7A9: dout <= 8'b11111000; // 1961 : 248 - 0xf8
      12'h7AA: dout <= 8'b11111000; // 1962 : 248 - 0xf8
      12'h7AB: dout <= 8'b11111000; // 1963 : 248 - 0xf8
      12'h7AC: dout <= 8'b00000000; // 1964 :   0 - 0x0
      12'h7AD: dout <= 8'b00000000; // 1965 :   0 - 0x0
      12'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      12'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout <= 8'b11111100; // 1968 : 252 - 0xfc -- Sprite 0xf6
      12'h7B1: dout <= 8'b11111100; // 1969 : 252 - 0xfc
      12'h7B2: dout <= 8'b11111100; // 1970 : 252 - 0xfc
      12'h7B3: dout <= 8'b11111100; // 1971 : 252 - 0xfc
      12'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      12'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      12'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout <= 8'b11111110; // 1976 : 254 - 0xfe -- Sprite 0xf7
      12'h7B9: dout <= 8'b11111110; // 1977 : 254 - 0xfe
      12'h7BA: dout <= 8'b11111110; // 1978 : 254 - 0xfe
      12'h7BB: dout <= 8'b11111110; // 1979 : 254 - 0xfe
      12'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout <= 8'b00000000; // 1982 :   0 - 0x0
      12'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout <= 8'b11111111; // 1984 : 255 - 0xff -- Sprite 0xf8
      12'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      12'h7C2: dout <= 8'b11111111; // 1986 : 255 - 0xff
      12'h7C3: dout <= 8'b11111111; // 1987 : 255 - 0xff
      12'h7C4: dout <= 8'b00000000; // 1988 :   0 - 0x0
      12'h7C5: dout <= 8'b00000000; // 1989 :   0 - 0x0
      12'h7C6: dout <= 8'b00000000; // 1990 :   0 - 0x0
      12'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      12'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0 -- Sprite 0xf9
      12'h7C9: dout <= 8'b00000000; // 1993 :   0 - 0x0
      12'h7CA: dout <= 8'b00000000; // 1994 :   0 - 0x0
      12'h7CB: dout <= 8'b00000000; // 1995 :   0 - 0x0
      12'h7CC: dout <= 8'b01111111; // 1996 : 127 - 0x7f
      12'h7CD: dout <= 8'b01000000; // 1997 :  64 - 0x40
      12'h7CE: dout <= 8'b01000000; // 1998 :  64 - 0x40
      12'h7CF: dout <= 8'b01000000; // 1999 :  64 - 0x40
      12'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0xfa
      12'h7D1: dout <= 8'b00000000; // 2001 :   0 - 0x0
      12'h7D2: dout <= 8'b00000000; // 2002 :   0 - 0x0
      12'h7D3: dout <= 8'b00000000; // 2003 :   0 - 0x0
      12'h7D4: dout <= 8'b11111111; // 2004 : 255 - 0xff
      12'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      12'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      12'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      12'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0 -- Sprite 0xfb
      12'h7D9: dout <= 8'b00000000; // 2009 :   0 - 0x0
      12'h7DA: dout <= 8'b00000000; // 2010 :   0 - 0x0
      12'h7DB: dout <= 8'b00000000; // 2011 :   0 - 0x0
      12'h7DC: dout <= 8'b11111110; // 2012 : 254 - 0xfe
      12'h7DD: dout <= 8'b00000010; // 2013 :   2 - 0x2
      12'h7DE: dout <= 8'b00000010; // 2014 :   2 - 0x2
      12'h7DF: dout <= 8'b00000010; // 2015 :   2 - 0x2
      12'h7E0: dout <= 8'b01000000; // 2016 :  64 - 0x40 -- Sprite 0xfc
      12'h7E1: dout <= 8'b01000000; // 2017 :  64 - 0x40
      12'h7E2: dout <= 8'b01000000; // 2018 :  64 - 0x40
      12'h7E3: dout <= 8'b01111111; // 2019 : 127 - 0x7f
      12'h7E4: dout <= 8'b00000000; // 2020 :   0 - 0x0
      12'h7E5: dout <= 8'b00000000; // 2021 :   0 - 0x0
      12'h7E6: dout <= 8'b00000000; // 2022 :   0 - 0x0
      12'h7E7: dout <= 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0 -- Sprite 0xfd
      12'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout <= 8'b00000000; // 2026 :   0 - 0x0
      12'h7EB: dout <= 8'b11111111; // 2027 : 255 - 0xff
      12'h7EC: dout <= 8'b00000000; // 2028 :   0 - 0x0
      12'h7ED: dout <= 8'b00000000; // 2029 :   0 - 0x0
      12'h7EE: dout <= 8'b00000000; // 2030 :   0 - 0x0
      12'h7EF: dout <= 8'b00000000; // 2031 :   0 - 0x0
      12'h7F0: dout <= 8'b00000010; // 2032 :   2 - 0x2 -- Sprite 0xfe
      12'h7F1: dout <= 8'b00000010; // 2033 :   2 - 0x2
      12'h7F2: dout <= 8'b00000010; // 2034 :   2 - 0x2
      12'h7F3: dout <= 8'b11111110; // 2035 : 254 - 0xfe
      12'h7F4: dout <= 8'b00000000; // 2036 :   0 - 0x0
      12'h7F5: dout <= 8'b00000000; // 2037 :   0 - 0x0
      12'h7F6: dout <= 8'b00000000; // 2038 :   0 - 0x0
      12'h7F7: dout <= 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      12'h7F9: dout <= 8'b00000000; // 2041 :   0 - 0x0
      12'h7FA: dout <= 8'b00000000; // 2042 :   0 - 0x0
      12'h7FB: dout <= 8'b00000000; // 2043 :   0 - 0x0
      12'h7FC: dout <= 8'b00000000; // 2044 :   0 - 0x0
      12'h7FD: dout <= 8'b00000000; // 2045 :   0 - 0x0
      12'h7FE: dout <= 8'b00000000; // 2046 :   0 - 0x0
      12'h7FF: dout <= 8'b00000000; // 2047 :   0 - 0x0
          // Background pattern Table
      12'h800: dout <= 8'b00000101; // 2048 :   5 - 0x5 -- Background 0x0
      12'h801: dout <= 8'b01010101; // 2049 :  85 - 0x55
      12'h802: dout <= 8'b01010101; // 2050 :  85 - 0x55
      12'h803: dout <= 8'b01010000; // 2051 :  80 - 0x50
      12'h804: dout <= 8'b00000000; // 2052 :   0 - 0x0
      12'h805: dout <= 8'b00000000; // 2053 :   0 - 0x0
      12'h806: dout <= 8'b00000000; // 2054 :   0 - 0x0
      12'h807: dout <= 8'b00000000; // 2055 :   0 - 0x0
      12'h808: dout <= 8'b00000101; // 2056 :   5 - 0x5 -- Background 0x1
      12'h809: dout <= 8'b01010101; // 2057 :  85 - 0x55
      12'h80A: dout <= 8'b01010101; // 2058 :  85 - 0x55
      12'h80B: dout <= 8'b01010000; // 2059 :  80 - 0x50
      12'h80C: dout <= 8'b00000000; // 2060 :   0 - 0x0
      12'h80D: dout <= 8'b00000000; // 2061 :   0 - 0x0
      12'h80E: dout <= 8'b00000000; // 2062 :   0 - 0x0
      12'h80F: dout <= 8'b00000000; // 2063 :   0 - 0x0
      12'h810: dout <= 8'b00000101; // 2064 :   5 - 0x5 -- Background 0x2
      12'h811: dout <= 8'b01010000; // 2065 :  80 - 0x50
      12'h812: dout <= 8'b00000101; // 2066 :   5 - 0x5
      12'h813: dout <= 8'b01010000; // 2067 :  80 - 0x50
      12'h814: dout <= 8'b00000000; // 2068 :   0 - 0x0
      12'h815: dout <= 8'b00000000; // 2069 :   0 - 0x0
      12'h816: dout <= 8'b00000000; // 2070 :   0 - 0x0
      12'h817: dout <= 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout <= 8'b00000101; // 2072 :   5 - 0x5 -- Background 0x3
      12'h819: dout <= 8'b01010101; // 2073 :  85 - 0x55
      12'h81A: dout <= 8'b01010101; // 2074 :  85 - 0x55
      12'h81B: dout <= 8'b01010000; // 2075 :  80 - 0x50
      12'h81C: dout <= 8'b00000000; // 2076 :   0 - 0x0
      12'h81D: dout <= 8'b00000000; // 2077 :   0 - 0x0
      12'h81E: dout <= 8'b00000000; // 2078 :   0 - 0x0
      12'h81F: dout <= 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout <= 8'b00000101; // 2080 :   5 - 0x5 -- Background 0x4
      12'h821: dout <= 8'b01010101; // 2081 :  85 - 0x55
      12'h822: dout <= 8'b01010101; // 2082 :  85 - 0x55
      12'h823: dout <= 8'b01010000; // 2083 :  80 - 0x50
      12'h824: dout <= 8'b00000000; // 2084 :   0 - 0x0
      12'h825: dout <= 8'b00000000; // 2085 :   0 - 0x0
      12'h826: dout <= 8'b00000000; // 2086 :   0 - 0x0
      12'h827: dout <= 8'b00000000; // 2087 :   0 - 0x0
      12'h828: dout <= 8'b00001110; // 2088 :  14 - 0xe -- Background 0x5
      12'h829: dout <= 8'b00000111; // 2089 :   7 - 0x7
      12'h82A: dout <= 8'b00001000; // 2090 :   8 - 0x8
      12'h82B: dout <= 8'b01100000; // 2091 :  96 - 0x60
      12'h82C: dout <= 8'b00000000; // 2092 :   0 - 0x0
      12'h82D: dout <= 8'b00001010; // 2093 :  10 - 0xa
      12'h82E: dout <= 8'b00000001; // 2094 :   1 - 0x1
      12'h82F: dout <= 8'b00010101; // 2095 :  21 - 0x15
      12'h830: dout <= 8'b01010101; // 2096 :  85 - 0x55 -- Background 0x6
      12'h831: dout <= 8'b01010101; // 2097 :  85 - 0x55
      12'h832: dout <= 8'b01010100; // 2098 :  84 - 0x54
      12'h833: dout <= 8'b00000000; // 2099 :   0 - 0x0
      12'h834: dout <= 8'b00000000; // 2100 :   0 - 0x0
      12'h835: dout <= 8'b00000000; // 2101 :   0 - 0x0
      12'h836: dout <= 8'b00000000; // 2102 :   0 - 0x0
      12'h837: dout <= 8'b00010110; // 2103 :  22 - 0x16
      12'h838: dout <= 8'b01010101; // 2104 :  85 - 0x55 -- Background 0x7
      12'h839: dout <= 8'b01010101; // 2105 :  85 - 0x55
      12'h83A: dout <= 8'b10010100; // 2106 : 148 - 0x94
      12'h83B: dout <= 8'b00000000; // 2107 :   0 - 0x0
      12'h83C: dout <= 8'b00000000; // 2108 :   0 - 0x0
      12'h83D: dout <= 8'b00000000; // 2109 :   0 - 0x0
      12'h83E: dout <= 8'b00000000; // 2110 :   0 - 0x0
      12'h83F: dout <= 8'b00010110; // 2111 :  22 - 0x16
      12'h840: dout <= 8'b01010000; // 2112 :  80 - 0x50 -- Background 0x8
      12'h841: dout <= 8'b00000101; // 2113 :   5 - 0x5
      12'h842: dout <= 8'b01010100; // 2114 :  84 - 0x54
      12'h843: dout <= 8'b00000000; // 2115 :   0 - 0x0
      12'h844: dout <= 8'b00000000; // 2116 :   0 - 0x0
      12'h845: dout <= 8'b00000000; // 2117 :   0 - 0x0
      12'h846: dout <= 8'b00000000; // 2118 :   0 - 0x0
      12'h847: dout <= 8'b00010110; // 2119 :  22 - 0x16
      12'h848: dout <= 8'b01010101; // 2120 :  85 - 0x55 -- Background 0x9
      12'h849: dout <= 8'b01010101; // 2121 :  85 - 0x55
      12'h84A: dout <= 8'b10010100; // 2122 : 148 - 0x94
      12'h84B: dout <= 8'b00000000; // 2123 :   0 - 0x0
      12'h84C: dout <= 8'b00000000; // 2124 :   0 - 0x0
      12'h84D: dout <= 8'b00000000; // 2125 :   0 - 0x0
      12'h84E: dout <= 8'b00000000; // 2126 :   0 - 0x0
      12'h84F: dout <= 8'b00010110; // 2127 :  22 - 0x16
      12'h850: dout <= 8'b01010101; // 2128 :  85 - 0x55 -- Background 0xa
      12'h851: dout <= 8'b01010101; // 2129 :  85 - 0x55
      12'h852: dout <= 8'b01010100; // 2130 :  84 - 0x54
      12'h853: dout <= 8'b00000000; // 2131 :   0 - 0x0
      12'h854: dout <= 8'b00000000; // 2132 :   0 - 0x0
      12'h855: dout <= 8'b00000000; // 2133 :   0 - 0x0
      12'h856: dout <= 8'b00000000; // 2134 :   0 - 0x0
      12'h857: dout <= 8'b00010101; // 2135 :  21 - 0x15
      12'h858: dout <= 8'b00000111; // 2136 :   7 - 0x7 -- Background 0xb
      12'h859: dout <= 8'b00001000; // 2137 :   8 - 0x8
      12'h85A: dout <= 8'b01110100; // 2138 : 116 - 0x74
      12'h85B: dout <= 8'b00000000; // 2139 :   0 - 0x0
      12'h85C: dout <= 8'b11011100; // 2140 : 220 - 0xdc
      12'h85D: dout <= 8'b00000000; // 2141 :   0 - 0x0
      12'h85E: dout <= 8'b00010101; // 2142 :  21 - 0x15
      12'h85F: dout <= 8'b01010101; // 2143 :  85 - 0x55
      12'h860: dout <= 8'b01110110; // 2144 : 118 - 0x76 -- Background 0xc
      12'h861: dout <= 8'b10100100; // 2145 : 164 - 0xa4
      12'h862: dout <= 8'b00000000; // 2146 :   0 - 0x0
      12'h863: dout <= 8'b00000000; // 2147 :   0 - 0x0
      12'h864: dout <= 8'b00000000; // 2148 :   0 - 0x0
      12'h865: dout <= 8'b00000000; // 2149 :   0 - 0x0
      12'h866: dout <= 8'b00010101; // 2150 :  21 - 0x15
      12'h867: dout <= 8'b01010101; // 2151 :  85 - 0x55
      12'h868: dout <= 8'b01010101; // 2152 :  85 - 0x55 -- Background 0xd
      12'h869: dout <= 8'b11010100; // 2153 : 212 - 0xd4
      12'h86A: dout <= 8'b00000000; // 2154 :   0 - 0x0
      12'h86B: dout <= 8'b00000000; // 2155 :   0 - 0x0
      12'h86C: dout <= 8'b00000000; // 2156 :   0 - 0x0
      12'h86D: dout <= 8'b00000000; // 2157 :   0 - 0x0
      12'h86E: dout <= 8'b00010101; // 2158 :  21 - 0x15
      12'h86F: dout <= 8'b01010000; // 2159 :  80 - 0x50
      12'h870: dout <= 8'b00000101; // 2160 :   5 - 0x5 -- Background 0xe
      12'h871: dout <= 8'b01010100; // 2161 :  84 - 0x54
      12'h872: dout <= 8'b00000000; // 2162 :   0 - 0x0
      12'h873: dout <= 8'b00000000; // 2163 :   0 - 0x0
      12'h874: dout <= 8'b00000000; // 2164 :   0 - 0x0
      12'h875: dout <= 8'b00000000; // 2165 :   0 - 0x0
      12'h876: dout <= 8'b00010101; // 2166 :  21 - 0x15
      12'h877: dout <= 8'b01010000; // 2167 :  80 - 0x50
      12'h878: dout <= 8'b01010101; // 2168 :  85 - 0x55 -- Background 0xf
      12'h879: dout <= 8'b11010100; // 2169 : 212 - 0xd4
      12'h87A: dout <= 8'b00000000; // 2170 :   0 - 0x0
      12'h87B: dout <= 8'b00000000; // 2171 :   0 - 0x0
      12'h87C: dout <= 8'b00000000; // 2172 :   0 - 0x0
      12'h87D: dout <= 8'b00000000; // 2173 :   0 - 0x0
      12'h87E: dout <= 8'b00010101; // 2174 :  21 - 0x15
      12'h87F: dout <= 8'b01010101; // 2175 :  85 - 0x55
      12'h880: dout <= 8'b01110110; // 2176 : 118 - 0x76 -- Background 0x10
      12'h881: dout <= 8'b10100100; // 2177 : 164 - 0xa4
      12'h882: dout <= 8'b00000000; // 2178 :   0 - 0x0
      12'h883: dout <= 8'b00000000; // 2179 :   0 - 0x0
      12'h884: dout <= 8'b00000000; // 2180 :   0 - 0x0
      12'h885: dout <= 8'b00000000; // 2181 :   0 - 0x0
      12'h886: dout <= 8'b00010101; // 2182 :  21 - 0x15
      12'h887: dout <= 8'b01010101; // 2183 :  85 - 0x55
      12'h888: dout <= 8'b00001000; // 2184 :   8 - 0x8 -- Background 0x11
      12'h889: dout <= 8'b01111010; // 2185 : 122 - 0x7a
      12'h88A: dout <= 8'b00000000; // 2186 :   0 - 0x0
      12'h88B: dout <= 8'b11010001; // 2187 : 209 - 0xd1
      12'h88C: dout <= 8'b00000000; // 2188 :   0 - 0x0
      12'h88D: dout <= 8'b00010101; // 2189 :  21 - 0x15
      12'h88E: dout <= 8'b01010101; // 2190 :  85 - 0x55
      12'h88F: dout <= 8'b01010101; // 2191 :  85 - 0x55
      12'h890: dout <= 8'b01010101; // 2192 :  85 - 0x55 -- Background 0x12
      12'h891: dout <= 8'b01010101; // 2193 :  85 - 0x55
      12'h892: dout <= 8'b01000000; // 2194 :  64 - 0x40
      12'h893: dout <= 8'b00000000; // 2195 :   0 - 0x0
      12'h894: dout <= 8'b00000000; // 2196 :   0 - 0x0
      12'h895: dout <= 8'b00010110; // 2197 :  22 - 0x16
      12'h896: dout <= 8'b10100101; // 2198 : 165 - 0xa5
      12'h897: dout <= 8'b01010101; // 2199 :  85 - 0x55
      12'h898: dout <= 8'b10010101; // 2200 : 149 - 0x95 -- Background 0x13
      12'h899: dout <= 8'b01011001; // 2201 :  89 - 0x59
      12'h89A: dout <= 8'b01000000; // 2202 :  64 - 0x40
      12'h89B: dout <= 8'b00000000; // 2203 :   0 - 0x0
      12'h89C: dout <= 8'b00000000; // 2204 :   0 - 0x0
      12'h89D: dout <= 8'b00010110; // 2205 :  22 - 0x16
      12'h89E: dout <= 8'b01000000; // 2206 :  64 - 0x40
      12'h89F: dout <= 8'b01010101; // 2207 :  85 - 0x55
      12'h8A0: dout <= 8'b01010101; // 2208 :  85 - 0x55 -- Background 0x14
      12'h8A1: dout <= 8'b01010101; // 2209 :  85 - 0x55
      12'h8A2: dout <= 8'b01000000; // 2210 :  64 - 0x40
      12'h8A3: dout <= 8'b00000000; // 2211 :   0 - 0x0
      12'h8A4: dout <= 8'b00000000; // 2212 :   0 - 0x0
      12'h8A5: dout <= 8'b00010110; // 2213 :  22 - 0x16
      12'h8A6: dout <= 8'b01000000; // 2214 :  64 - 0x40
      12'h8A7: dout <= 8'b01010101; // 2215 :  85 - 0x55
      12'h8A8: dout <= 8'b10010101; // 2216 : 149 - 0x95 -- Background 0x15
      12'h8A9: dout <= 8'b01011001; // 2217 :  89 - 0x59
      12'h8AA: dout <= 8'b01000000; // 2218 :  64 - 0x40
      12'h8AB: dout <= 8'b00000000; // 2219 :   0 - 0x0
      12'h8AC: dout <= 8'b00000000; // 2220 :   0 - 0x0
      12'h8AD: dout <= 8'b00010110; // 2221 :  22 - 0x16
      12'h8AE: dout <= 8'b10100101; // 2222 : 165 - 0xa5
      12'h8AF: dout <= 8'b01010101; // 2223 :  85 - 0x55
      12'h8B0: dout <= 8'b01010101; // 2224 :  85 - 0x55 -- Background 0x16
      12'h8B1: dout <= 8'b01010101; // 2225 :  85 - 0x55
      12'h8B2: dout <= 8'b01000000; // 2226 :  64 - 0x40
      12'h8B3: dout <= 8'b00000000; // 2227 :   0 - 0x0
      12'h8B4: dout <= 8'b00000000; // 2228 :   0 - 0x0
      12'h8B5: dout <= 8'b00010101; // 2229 :  21 - 0x15
      12'h8B6: dout <= 8'b01010101; // 2230 :  85 - 0x55
      12'h8B7: dout <= 8'b01010101; // 2231 :  85 - 0x55
      12'h8B8: dout <= 8'b10110111; // 2232 : 183 - 0xb7 -- Background 0x17
      12'h8B9: dout <= 8'b00000000; // 2233 :   0 - 0x0
      12'h8BA: dout <= 8'b10001011; // 2234 : 139 - 0x8b
      12'h8BB: dout <= 8'b00000000; // 2235 :   0 - 0x0
      12'h8BC: dout <= 8'b00010101; // 2236 :  21 - 0x15
      12'h8BD: dout <= 8'b01010101; // 2237 :  85 - 0x55
      12'h8BE: dout <= 8'b01010101; // 2238 :  85 - 0x55
      12'h8BF: dout <= 8'b01010101; // 2239 :  85 - 0x55
      12'h8C0: dout <= 8'b01011010; // 2240 :  90 - 0x5a -- Background 0x18
      12'h8C1: dout <= 8'b01000000; // 2241 :  64 - 0x40
      12'h8C2: dout <= 8'b00000000; // 2242 :   0 - 0x0
      12'h8C3: dout <= 8'b00000000; // 2243 :   0 - 0x0
      12'h8C4: dout <= 8'b00011010; // 2244 :  26 - 0x1a
      12'h8C5: dout <= 8'b01010111; // 2245 :  87 - 0x57
      12'h8C6: dout <= 8'b01010101; // 2246 :  85 - 0x55
      12'h8C7: dout <= 8'b01011101; // 2247 :  93 - 0x5d
      12'h8C8: dout <= 8'b01010101; // 2248 :  85 - 0x55 -- Background 0x19
      12'h8C9: dout <= 8'b01000000; // 2249 :  64 - 0x40
      12'h8CA: dout <= 8'b00000000; // 2250 :   0 - 0x0
      12'h8CB: dout <= 8'b00000000; // 2251 :   0 - 0x0
      12'h8CC: dout <= 8'b00010000; // 2252 :  16 - 0x10
      12'h8CD: dout <= 8'b00010101; // 2253 :  21 - 0x15
      12'h8CE: dout <= 8'b01011010; // 2254 :  90 - 0x5a
      12'h8CF: dout <= 8'b01010101; // 2255 :  85 - 0x55
      12'h8D0: dout <= 8'b01010101; // 2256 :  85 - 0x55 -- Background 0x1a
      12'h8D1: dout <= 8'b01000000; // 2257 :  64 - 0x40
      12'h8D2: dout <= 8'b00000000; // 2258 :   0 - 0x0
      12'h8D3: dout <= 8'b00000000; // 2259 :   0 - 0x0
      12'h8D4: dout <= 8'b00010000; // 2260 :  16 - 0x10
      12'h8D5: dout <= 8'b00010101; // 2261 :  21 - 0x15
      12'h8D6: dout <= 8'b01011010; // 2262 :  90 - 0x5a
      12'h8D7: dout <= 8'b01010101; // 2263 :  85 - 0x55
      12'h8D8: dout <= 8'b01010101; // 2264 :  85 - 0x55 -- Background 0x1b
      12'h8D9: dout <= 8'b01000000; // 2265 :  64 - 0x40
      12'h8DA: dout <= 8'b00000000; // 2266 :   0 - 0x0
      12'h8DB: dout <= 8'b00000000; // 2267 :   0 - 0x0
      12'h8DC: dout <= 8'b00011010; // 2268 :  26 - 0x1a
      12'h8DD: dout <= 8'b01010111; // 2269 :  87 - 0x57
      12'h8DE: dout <= 8'b01010101; // 2270 :  85 - 0x55
      12'h8DF: dout <= 8'b01011101; // 2271 :  93 - 0x5d
      12'h8E0: dout <= 8'b01011010; // 2272 :  90 - 0x5a -- Background 0x1c
      12'h8E1: dout <= 8'b01000000; // 2273 :  64 - 0x40
      12'h8E2: dout <= 8'b00000000; // 2274 :   0 - 0x0
      12'h8E3: dout <= 8'b00000000; // 2275 :   0 - 0x0
      12'h8E4: dout <= 8'b00010101; // 2276 :  21 - 0x15
      12'h8E5: dout <= 8'b01010101; // 2277 :  85 - 0x55
      12'h8E6: dout <= 8'b01010101; // 2278 :  85 - 0x55
      12'h8E7: dout <= 8'b01010101; // 2279 :  85 - 0x55
      12'h8E8: dout <= 8'b00000000; // 2280 :   0 - 0x0 -- Background 0x1d
      12'h8E9: dout <= 8'b10010011; // 2281 : 147 - 0x93
      12'h8EA: dout <= 8'b00000000; // 2282 :   0 - 0x0
      12'h8EB: dout <= 8'b00010101; // 2283 :  21 - 0x15
      12'h8EC: dout <= 8'b01010101; // 2284 :  85 - 0x55
      12'h8ED: dout <= 8'b01010101; // 2285 :  85 - 0x55
      12'h8EE: dout <= 8'b01010101; // 2286 :  85 - 0x55
      12'h8EF: dout <= 8'b01010101; // 2287 :  85 - 0x55
      12'h8F0: dout <= 8'b01010111; // 2288 :  87 - 0x57 -- Background 0x1e
      12'h8F1: dout <= 8'b01010000; // 2289 :  80 - 0x50
      12'h8F2: dout <= 8'b00000000; // 2290 :   0 - 0x0
      12'h8F3: dout <= 8'b00011101; // 2291 :  29 - 0x1d
      12'h8F4: dout <= 8'b01010101; // 2292 :  85 - 0x55
      12'h8F5: dout <= 8'b01110101; // 2293 : 117 - 0x75
      12'h8F6: dout <= 8'b01010101; // 2294 :  85 - 0x55
      12'h8F7: dout <= 8'b01011101; // 2295 :  93 - 0x5d
      12'h8F8: dout <= 8'b01110101; // 2296 : 117 - 0x75 -- Background 0x1f
      12'h8F9: dout <= 8'b01010000; // 2297 :  80 - 0x50
      12'h8FA: dout <= 8'b00000000; // 2298 :   0 - 0x0
      12'h8FB: dout <= 8'b00010101; // 2299 :  21 - 0x15
      12'h8FC: dout <= 8'b01010101; // 2300 :  85 - 0x55
      12'h8FD: dout <= 8'b01010101; // 2301 :  85 - 0x55
      12'h8FE: dout <= 8'b00000001; // 2302 :   1 - 0x1
      12'h8FF: dout <= 8'b01010101; // 2303 :  85 - 0x55
      12'h900: dout <= 8'b01010101; // 2304 :  85 - 0x55 -- Background 0x20
      12'h901: dout <= 8'b01010000; // 2305 :  80 - 0x50
      12'h902: dout <= 8'b00000000; // 2306 :   0 - 0x0
      12'h903: dout <= 8'b00010101; // 2307 :  21 - 0x15
      12'h904: dout <= 8'b01011101; // 2308 :  93 - 0x5d
      12'h905: dout <= 8'b01010101; // 2309 :  85 - 0x55
      12'h906: dout <= 8'b00000001; // 2310 :   1 - 0x1
      12'h907: dout <= 8'b01010101; // 2311 :  85 - 0x55
      12'h908: dout <= 8'b01110101; // 2312 : 117 - 0x75 -- Background 0x21
      12'h909: dout <= 8'b01010000; // 2313 :  80 - 0x50
      12'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout <= 8'b00011101; // 2315 :  29 - 0x1d
      12'h90C: dout <= 8'b01010101; // 2316 :  85 - 0x55
      12'h90D: dout <= 8'b01010101; // 2317 :  85 - 0x55
      12'h90E: dout <= 8'b01010101; // 2318 :  85 - 0x55
      12'h90F: dout <= 8'b01110101; // 2319 : 117 - 0x75
      12'h910: dout <= 8'b01010111; // 2320 :  87 - 0x57 -- Background 0x22
      12'h911: dout <= 8'b01010000; // 2321 :  80 - 0x50
      12'h912: dout <= 8'b00000000; // 2322 :   0 - 0x0
      12'h913: dout <= 8'b00010101; // 2323 :  21 - 0x15
      12'h914: dout <= 8'b01010101; // 2324 :  85 - 0x55
      12'h915: dout <= 8'b01010101; // 2325 :  85 - 0x55
      12'h916: dout <= 8'b01010101; // 2326 :  85 - 0x55
      12'h917: dout <= 8'b01010101; // 2327 :  85 - 0x55
      12'h918: dout <= 8'b01100111; // 2328 : 103 - 0x67 -- Background 0x23
      12'h919: dout <= 8'b00000000; // 2329 :   0 - 0x0
      12'h91A: dout <= 8'b00010101; // 2330 :  21 - 0x15
      12'h91B: dout <= 8'b01010101; // 2331 :  85 - 0x55
      12'h91C: dout <= 8'b01010101; // 2332 :  85 - 0x55
      12'h91D: dout <= 8'b01010101; // 2333 :  85 - 0x55
      12'h91E: dout <= 8'b01010101; // 2334 :  85 - 0x55
      12'h91F: dout <= 8'b01010101; // 2335 :  85 - 0x55
      12'h920: dout <= 8'b10010000; // 2336 : 144 - 0x90 -- Background 0x24
      12'h921: dout <= 8'b00000000; // 2337 :   0 - 0x0
      12'h922: dout <= 8'b00011001; // 2338 :  25 - 0x19
      12'h923: dout <= 8'b01011001; // 2339 :  89 - 0x59
      12'h924: dout <= 8'b10010101; // 2340 : 149 - 0x95
      12'h925: dout <= 8'b10011001; // 2341 : 153 - 0x99
      12'h926: dout <= 8'b01011001; // 2342 :  89 - 0x59
      12'h927: dout <= 8'b10010101; // 2343 : 149 - 0x95
      12'h928: dout <= 8'b01010000; // 2344 :  80 - 0x50 -- Background 0x25
      12'h929: dout <= 8'b00000000; // 2345 :   0 - 0x0
      12'h92A: dout <= 8'b00010000; // 2346 :  16 - 0x10
      12'h92B: dout <= 8'b00010101; // 2347 :  21 - 0x15
      12'h92C: dout <= 8'b10010101; // 2348 : 149 - 0x95
      12'h92D: dout <= 8'b10011010; // 2349 : 154 - 0x9a
      12'h92E: dout <= 8'b10101001; // 2350 : 169 - 0xa9
      12'h92F: dout <= 8'b01010101; // 2351 :  85 - 0x55
      12'h930: dout <= 8'b01010000; // 2352 :  80 - 0x50 -- Background 0x26
      12'h931: dout <= 8'b00000000; // 2353 :   0 - 0x0
      12'h932: dout <= 8'b00010000; // 2354 :  16 - 0x10
      12'h933: dout <= 8'b00010101; // 2355 :  21 - 0x15
      12'h934: dout <= 8'b10101010; // 2356 : 170 - 0xaa
      12'h935: dout <= 8'b10011001; // 2357 : 153 - 0x99
      12'h936: dout <= 8'b01011001; // 2358 :  89 - 0x59
      12'h937: dout <= 8'b01010101; // 2359 :  85 - 0x55
      12'h938: dout <= 8'b01010000; // 2360 :  80 - 0x50 -- Background 0x27
      12'h939: dout <= 8'b00000000; // 2361 :   0 - 0x0
      12'h93A: dout <= 8'b00011001; // 2362 :  25 - 0x19
      12'h93B: dout <= 8'b01011001; // 2363 :  89 - 0x59
      12'h93C: dout <= 8'b10010101; // 2364 : 149 - 0x95
      12'h93D: dout <= 8'b10011001; // 2365 : 153 - 0x99
      12'h93E: dout <= 8'b01011001; // 2366 :  89 - 0x59
      12'h93F: dout <= 8'b10010101; // 2367 : 149 - 0x95
      12'h940: dout <= 8'b10010000; // 2368 : 144 - 0x90 -- Background 0x28
      12'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout <= 8'b00010101; // 2370 :  21 - 0x15
      12'h943: dout <= 8'b01010101; // 2371 :  85 - 0x55
      12'h944: dout <= 8'b01010101; // 2372 :  85 - 0x55
      12'h945: dout <= 8'b01010101; // 2373 :  85 - 0x55
      12'h946: dout <= 8'b01010101; // 2374 :  85 - 0x55
      12'h947: dout <= 8'b01010101; // 2375 :  85 - 0x55
      12'h948: dout <= 8'b00000000; // 2376 :   0 - 0x0 -- Background 0x29
      12'h949: dout <= 8'b00010101; // 2377 :  21 - 0x15
      12'h94A: dout <= 8'b01010111; // 2378 :  87 - 0x57
      12'h94B: dout <= 8'b01010101; // 2379 :  85 - 0x55
      12'h94C: dout <= 8'b01010101; // 2380 :  85 - 0x55
      12'h94D: dout <= 8'b01010111; // 2381 :  87 - 0x57
      12'h94E: dout <= 8'b01010101; // 2382 :  85 - 0x55
      12'h94F: dout <= 8'b01010000; // 2383 :  80 - 0x50
      12'h950: dout <= 8'b00000000; // 2384 :   0 - 0x0 -- Background 0x2a
      12'h951: dout <= 8'b00010101; // 2385 :  21 - 0x15
      12'h952: dout <= 8'b01010111; // 2386 :  87 - 0x57
      12'h953: dout <= 8'b01101010; // 2387 : 106 - 0x6a
      12'h954: dout <= 8'b01010110; // 2388 :  86 - 0x56
      12'h955: dout <= 8'b10100111; // 2389 : 167 - 0xa7
      12'h956: dout <= 8'b01010101; // 2390 :  85 - 0x55
      12'h957: dout <= 8'b01010000; // 2391 :  80 - 0x50
      12'h958: dout <= 8'b00000000; // 2392 :   0 - 0x0 -- Background 0x2b
      12'h959: dout <= 8'b00010000; // 2393 :  16 - 0x10
      12'h95A: dout <= 8'b00010101; // 2394 :  21 - 0x15
      12'h95B: dout <= 8'b01010101; // 2395 :  85 - 0x55
      12'h95C: dout <= 8'b01110101; // 2396 : 117 - 0x75
      12'h95D: dout <= 8'b01010101; // 2397 :  85 - 0x55
      12'h95E: dout <= 8'b01010101; // 2398 :  85 - 0x55
      12'h95F: dout <= 8'b01010000; // 2399 :  80 - 0x50
      12'h960: dout <= 8'b00000000; // 2400 :   0 - 0x0 -- Background 0x2c
      12'h961: dout <= 8'b00010000; // 2401 :  16 - 0x10
      12'h962: dout <= 8'b00010101; // 2402 :  21 - 0x15
      12'h963: dout <= 8'b01010101; // 2403 :  85 - 0x55
      12'h964: dout <= 8'b01110101; // 2404 : 117 - 0x75
      12'h965: dout <= 8'b01010101; // 2405 :  85 - 0x55
      12'h966: dout <= 8'b01010101; // 2406 :  85 - 0x55
      12'h967: dout <= 8'b01010000; // 2407 :  80 - 0x50
      12'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0 -- Background 0x2d
      12'h969: dout <= 8'b00010101; // 2409 :  21 - 0x15
      12'h96A: dout <= 8'b01010111; // 2410 :  87 - 0x57
      12'h96B: dout <= 8'b01101010; // 2411 : 106 - 0x6a
      12'h96C: dout <= 8'b01010110; // 2412 :  86 - 0x56
      12'h96D: dout <= 8'b10100111; // 2413 : 167 - 0xa7
      12'h96E: dout <= 8'b01010101; // 2414 :  85 - 0x55
      12'h96F: dout <= 8'b01010000; // 2415 :  80 - 0x50
      12'h970: dout <= 8'b00000000; // 2416 :   0 - 0x0 -- Background 0x2e
      12'h971: dout <= 8'b00010101; // 2417 :  21 - 0x15
      12'h972: dout <= 8'b01010111; // 2418 :  87 - 0x57
      12'h973: dout <= 8'b01010101; // 2419 :  85 - 0x55
      12'h974: dout <= 8'b01010101; // 2420 :  85 - 0x55
      12'h975: dout <= 8'b01010111; // 2421 :  87 - 0x57
      12'h976: dout <= 8'b01010101; // 2422 :  85 - 0x55
      12'h977: dout <= 8'b01010000; // 2423 :  80 - 0x50
      12'h978: dout <= 8'b00010101; // 2424 :  21 - 0x15 -- Background 0x2f
      12'h979: dout <= 8'b01010101; // 2425 :  85 - 0x55
      12'h97A: dout <= 8'b01010101; // 2426 :  85 - 0x55
      12'h97B: dout <= 8'b01010101; // 2427 :  85 - 0x55
      12'h97C: dout <= 8'b01010101; // 2428 :  85 - 0x55
      12'h97D: dout <= 8'b01010101; // 2429 :  85 - 0x55
      12'h97E: dout <= 8'b01010101; // 2430 :  85 - 0x55
      12'h97F: dout <= 8'b01010100; // 2431 :  84 - 0x54
      12'h980: dout <= 8'b00011001; // 2432 :  25 - 0x19 -- Background 0x30
      12'h981: dout <= 8'b01100101; // 2433 : 101 - 0x65
      12'h982: dout <= 8'b10010101; // 2434 : 149 - 0x95
      12'h983: dout <= 8'b01010101; // 2435 :  85 - 0x55
      12'h984: dout <= 8'b01010101; // 2436 :  85 - 0x55
      12'h985: dout <= 8'b01010110; // 2437 :  86 - 0x56
      12'h986: dout <= 8'b01011001; // 2438 :  89 - 0x59
      12'h987: dout <= 8'b01100100; // 2439 : 100 - 0x64
      12'h988: dout <= 8'b00010101; // 2440 :  21 - 0x15 -- Background 0x31
      12'h989: dout <= 8'b01010101; // 2441 :  85 - 0x55
      12'h98A: dout <= 8'b01010101; // 2442 :  85 - 0x55
      12'h98B: dout <= 8'b01010000; // 2443 :  80 - 0x50
      12'h98C: dout <= 8'b00000101; // 2444 :   5 - 0x5
      12'h98D: dout <= 8'b01010101; // 2445 :  85 - 0x55
      12'h98E: dout <= 8'b01010101; // 2446 :  85 - 0x55
      12'h98F: dout <= 8'b01010100; // 2447 :  84 - 0x54
      12'h990: dout <= 8'b00010101; // 2448 :  21 - 0x15 -- Background 0x32
      12'h991: dout <= 8'b01010101; // 2449 :  85 - 0x55
      12'h992: dout <= 8'b01010101; // 2450 :  85 - 0x55
      12'h993: dout <= 8'b01010000; // 2451 :  80 - 0x50
      12'h994: dout <= 8'b00000101; // 2452 :   5 - 0x5
      12'h995: dout <= 8'b01010101; // 2453 :  85 - 0x55
      12'h996: dout <= 8'b01010101; // 2454 :  85 - 0x55
      12'h997: dout <= 8'b01010100; // 2455 :  84 - 0x54
      12'h998: dout <= 8'b00011001; // 2456 :  25 - 0x19 -- Background 0x33
      12'h999: dout <= 8'b01100101; // 2457 : 101 - 0x65
      12'h99A: dout <= 8'b10010101; // 2458 : 149 - 0x95
      12'h99B: dout <= 8'b01010101; // 2459 :  85 - 0x55
      12'h99C: dout <= 8'b01010101; // 2460 :  85 - 0x55
      12'h99D: dout <= 8'b01010110; // 2461 :  86 - 0x56
      12'h99E: dout <= 8'b01011001; // 2462 :  89 - 0x59
      12'h99F: dout <= 8'b01100100; // 2463 : 100 - 0x64
      12'h9A0: dout <= 8'b00010101; // 2464 :  21 - 0x15 -- Background 0x34
      12'h9A1: dout <= 8'b01010101; // 2465 :  85 - 0x55
      12'h9A2: dout <= 8'b01010101; // 2466 :  85 - 0x55
      12'h9A3: dout <= 8'b01010101; // 2467 :  85 - 0x55
      12'h9A4: dout <= 8'b01010101; // 2468 :  85 - 0x55
      12'h9A5: dout <= 8'b01010101; // 2469 :  85 - 0x55
      12'h9A6: dout <= 8'b01010101; // 2470 :  85 - 0x55
      12'h9A7: dout <= 8'b01010100; // 2471 :  84 - 0x54
      12'h9A8: dout <= 8'b01010101; // 2472 :  85 - 0x55 -- Background 0x35
      12'h9A9: dout <= 8'b01010101; // 2473 :  85 - 0x55
      12'h9AA: dout <= 8'b01010101; // 2474 :  85 - 0x55
      12'h9AB: dout <= 8'b01010101; // 2475 :  85 - 0x55
      12'h9AC: dout <= 8'b01010101; // 2476 :  85 - 0x55
      12'h9AD: dout <= 8'b01010101; // 2477 :  85 - 0x55
      12'h9AE: dout <= 8'b01010100; // 2478 :  84 - 0x54
      12'h9AF: dout <= 8'b00010111; // 2479 :  23 - 0x17
      12'h9B0: dout <= 8'b01010101; // 2480 :  85 - 0x55 -- Background 0x36
      12'h9B1: dout <= 8'b01110110; // 2481 : 118 - 0x76
      12'h9B2: dout <= 8'b10100101; // 2482 : 165 - 0xa5
      12'h9B3: dout <= 8'b01011010; // 2483 :  90 - 0x5a
      12'h9B4: dout <= 8'b10011101; // 2484 : 157 - 0x9d
      12'h9B5: dout <= 8'b01010101; // 2485 :  85 - 0x55
      12'h9B6: dout <= 8'b01010100; // 2486 :  84 - 0x54
      12'h9B7: dout <= 8'b00010111; // 2487 :  23 - 0x17
      12'h9B8: dout <= 8'b01101010; // 2488 : 106 - 0x6a -- Background 0x37
      12'h9B9: dout <= 8'b01110101; // 2489 : 117 - 0x75
      12'h9BA: dout <= 8'b01010000; // 2490 :  80 - 0x50
      12'h9BB: dout <= 8'b00000101; // 2491 :   5 - 0x5
      12'h9BC: dout <= 8'b01011101; // 2492 :  93 - 0x5d
      12'h9BD: dout <= 8'b10101001; // 2493 : 169 - 0xa9
      12'h9BE: dout <= 8'b01010100; // 2494 :  84 - 0x54
      12'h9BF: dout <= 8'b00010101; // 2495 :  21 - 0x15
      12'h9C0: dout <= 8'b01101010; // 2496 : 106 - 0x6a -- Background 0x38
      12'h9C1: dout <= 8'b01110101; // 2497 : 117 - 0x75
      12'h9C2: dout <= 8'b01010000; // 2498 :  80 - 0x50
      12'h9C3: dout <= 8'b00000101; // 2499 :   5 - 0x5
      12'h9C4: dout <= 8'b01011101; // 2500 :  93 - 0x5d
      12'h9C5: dout <= 8'b10101001; // 2501 : 169 - 0xa9
      12'h9C6: dout <= 8'b01010100; // 2502 :  84 - 0x54
      12'h9C7: dout <= 8'b00010111; // 2503 :  23 - 0x17
      12'h9C8: dout <= 8'b01010101; // 2504 :  85 - 0x55 -- Background 0x39
      12'h9C9: dout <= 8'b01110101; // 2505 : 117 - 0x75
      12'h9CA: dout <= 8'b10101010; // 2506 : 170 - 0xaa
      12'h9CB: dout <= 8'b10101010; // 2507 : 170 - 0xaa
      12'h9CC: dout <= 8'b01011101; // 2508 :  93 - 0x5d
      12'h9CD: dout <= 8'b01010101; // 2509 :  85 - 0x55
      12'h9CE: dout <= 8'b01010100; // 2510 :  84 - 0x54
      12'h9CF: dout <= 8'b00010111; // 2511 :  23 - 0x17
      12'h9D0: dout <= 8'b01010101; // 2512 :  85 - 0x55 -- Background 0x3a
      12'h9D1: dout <= 8'b01010101; // 2513 :  85 - 0x55
      12'h9D2: dout <= 8'b01010101; // 2514 :  85 - 0x55
      12'h9D3: dout <= 8'b01010101; // 2515 :  85 - 0x55
      12'h9D4: dout <= 8'b01010101; // 2516 :  85 - 0x55
      12'h9D5: dout <= 8'b01010101; // 2517 :  85 - 0x55
      12'h9D6: dout <= 8'b01010100; // 2518 :  84 - 0x54
      12'h9D7: dout <= 8'b00011110; // 2519 :  30 - 0x1e
      12'h9D8: dout <= 8'b00000000; // 2520 :   0 - 0x0 -- Background 0x3b
      12'h9D9: dout <= 8'b00000000; // 2521 :   0 - 0x0
      12'h9DA: dout <= 8'b00000000; // 2522 :   0 - 0x0
      12'h9DB: dout <= 8'b00000000; // 2523 :   0 - 0x0
      12'h9DC: dout <= 8'b00000000; // 2524 :   0 - 0x0
      12'h9DD: dout <= 8'b00000000; // 2525 :   0 - 0x0
      12'h9DE: dout <= 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout <= 8'b00000000; // 2528 :   0 - 0x0 -- Background 0x3c
      12'h9E1: dout <= 8'b00000000; // 2529 :   0 - 0x0
      12'h9E2: dout <= 8'b00000000; // 2530 :   0 - 0x0
      12'h9E3: dout <= 8'b00000000; // 2531 :   0 - 0x0
      12'h9E4: dout <= 8'b00000000; // 2532 :   0 - 0x0
      12'h9E5: dout <= 8'b00000000; // 2533 :   0 - 0x0
      12'h9E6: dout <= 8'b00000000; // 2534 :   0 - 0x0
      12'h9E7: dout <= 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0 -- Background 0x3d
      12'h9E9: dout <= 8'b00000000; // 2537 :   0 - 0x0
      12'h9EA: dout <= 8'b00000000; // 2538 :   0 - 0x0
      12'h9EB: dout <= 8'b00000000; // 2539 :   0 - 0x0
      12'h9EC: dout <= 8'b00000000; // 2540 :   0 - 0x0
      12'h9ED: dout <= 8'b00000000; // 2541 :   0 - 0x0
      12'h9EE: dout <= 8'b00000000; // 2542 :   0 - 0x0
      12'h9EF: dout <= 8'b00000000; // 2543 :   0 - 0x0
      12'h9F0: dout <= 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x3e
      12'h9F1: dout <= 8'b00000000; // 2545 :   0 - 0x0
      12'h9F2: dout <= 8'b00000000; // 2546 :   0 - 0x0
      12'h9F3: dout <= 8'b00000000; // 2547 :   0 - 0x0
      12'h9F4: dout <= 8'b00000000; // 2548 :   0 - 0x0
      12'h9F5: dout <= 8'b00000000; // 2549 :   0 - 0x0
      12'h9F6: dout <= 8'b00000000; // 2550 :   0 - 0x0
      12'h9F7: dout <= 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- Background 0x3f
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout <= 8'b00000000; // 2560 :   0 - 0x0 -- Background 0x40
      12'hA01: dout <= 8'b00000000; // 2561 :   0 - 0x0
      12'hA02: dout <= 8'b00000000; // 2562 :   0 - 0x0
      12'hA03: dout <= 8'b00000000; // 2563 :   0 - 0x0
      12'hA04: dout <= 8'b00000000; // 2564 :   0 - 0x0
      12'hA05: dout <= 8'b00000000; // 2565 :   0 - 0x0
      12'hA06: dout <= 8'b00000000; // 2566 :   0 - 0x0
      12'hA07: dout <= 8'b00000000; // 2567 :   0 - 0x0
      12'hA08: dout <= 8'b00000000; // 2568 :   0 - 0x0 -- Background 0x41
      12'hA09: dout <= 8'b00000000; // 2569 :   0 - 0x0
      12'hA0A: dout <= 8'b00000000; // 2570 :   0 - 0x0
      12'hA0B: dout <= 8'b00000000; // 2571 :   0 - 0x0
      12'hA0C: dout <= 8'b00000000; // 2572 :   0 - 0x0
      12'hA0D: dout <= 8'b00000000; // 2573 :   0 - 0x0
      12'hA0E: dout <= 8'b00000000; // 2574 :   0 - 0x0
      12'hA0F: dout <= 8'b00000000; // 2575 :   0 - 0x0
      12'hA10: dout <= 8'b00000000; // 2576 :   0 - 0x0 -- Background 0x42
      12'hA11: dout <= 8'b00000000; // 2577 :   0 - 0x0
      12'hA12: dout <= 8'b00000000; // 2578 :   0 - 0x0
      12'hA13: dout <= 8'b00000000; // 2579 :   0 - 0x0
      12'hA14: dout <= 8'b00000000; // 2580 :   0 - 0x0
      12'hA15: dout <= 8'b00000000; // 2581 :   0 - 0x0
      12'hA16: dout <= 8'b00000000; // 2582 :   0 - 0x0
      12'hA17: dout <= 8'b00000000; // 2583 :   0 - 0x0
      12'hA18: dout <= 8'b00000000; // 2584 :   0 - 0x0 -- Background 0x43
      12'hA19: dout <= 8'b00000000; // 2585 :   0 - 0x0
      12'hA1A: dout <= 8'b00000000; // 2586 :   0 - 0x0
      12'hA1B: dout <= 8'b00000000; // 2587 :   0 - 0x0
      12'hA1C: dout <= 8'b00000000; // 2588 :   0 - 0x0
      12'hA1D: dout <= 8'b00000000; // 2589 :   0 - 0x0
      12'hA1E: dout <= 8'b00000000; // 2590 :   0 - 0x0
      12'hA1F: dout <= 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout <= 8'b00000000; // 2592 :   0 - 0x0 -- Background 0x44
      12'hA21: dout <= 8'b00000000; // 2593 :   0 - 0x0
      12'hA22: dout <= 8'b00000000; // 2594 :   0 - 0x0
      12'hA23: dout <= 8'b00000000; // 2595 :   0 - 0x0
      12'hA24: dout <= 8'b00000000; // 2596 :   0 - 0x0
      12'hA25: dout <= 8'b00000000; // 2597 :   0 - 0x0
      12'hA26: dout <= 8'b00000000; // 2598 :   0 - 0x0
      12'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0 -- Background 0x45
      12'hA29: dout <= 8'b00000000; // 2601 :   0 - 0x0
      12'hA2A: dout <= 8'b00000000; // 2602 :   0 - 0x0
      12'hA2B: dout <= 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout <= 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout <= 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout <= 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout <= 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout <= 8'b00000000; // 2608 :   0 - 0x0 -- Background 0x46
      12'hA31: dout <= 8'b00000000; // 2609 :   0 - 0x0
      12'hA32: dout <= 8'b00000000; // 2610 :   0 - 0x0
      12'hA33: dout <= 8'b00000000; // 2611 :   0 - 0x0
      12'hA34: dout <= 8'b00000000; // 2612 :   0 - 0x0
      12'hA35: dout <= 8'b00000000; // 2613 :   0 - 0x0
      12'hA36: dout <= 8'b00000000; // 2614 :   0 - 0x0
      12'hA37: dout <= 8'b00000000; // 2615 :   0 - 0x0
      12'hA38: dout <= 8'b00000000; // 2616 :   0 - 0x0 -- Background 0x47
      12'hA39: dout <= 8'b00000000; // 2617 :   0 - 0x0
      12'hA3A: dout <= 8'b00000000; // 2618 :   0 - 0x0
      12'hA3B: dout <= 8'b00000000; // 2619 :   0 - 0x0
      12'hA3C: dout <= 8'b00000000; // 2620 :   0 - 0x0
      12'hA3D: dout <= 8'b00000000; // 2621 :   0 - 0x0
      12'hA3E: dout <= 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout <= 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout <= 8'b00000000; // 2624 :   0 - 0x0 -- Background 0x48
      12'hA41: dout <= 8'b00000000; // 2625 :   0 - 0x0
      12'hA42: dout <= 8'b00000000; // 2626 :   0 - 0x0
      12'hA43: dout <= 8'b00000000; // 2627 :   0 - 0x0
      12'hA44: dout <= 8'b00000000; // 2628 :   0 - 0x0
      12'hA45: dout <= 8'b00000000; // 2629 :   0 - 0x0
      12'hA46: dout <= 8'b00000000; // 2630 :   0 - 0x0
      12'hA47: dout <= 8'b00000000; // 2631 :   0 - 0x0
      12'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0 -- Background 0x49
      12'hA49: dout <= 8'b00000000; // 2633 :   0 - 0x0
      12'hA4A: dout <= 8'b00000000; // 2634 :   0 - 0x0
      12'hA4B: dout <= 8'b00000000; // 2635 :   0 - 0x0
      12'hA4C: dout <= 8'b00000000; // 2636 :   0 - 0x0
      12'hA4D: dout <= 8'b00000000; // 2637 :   0 - 0x0
      12'hA4E: dout <= 8'b00000000; // 2638 :   0 - 0x0
      12'hA4F: dout <= 8'b00000000; // 2639 :   0 - 0x0
      12'hA50: dout <= 8'b00000000; // 2640 :   0 - 0x0 -- Background 0x4a
      12'hA51: dout <= 8'b00000000; // 2641 :   0 - 0x0
      12'hA52: dout <= 8'b00000000; // 2642 :   0 - 0x0
      12'hA53: dout <= 8'b00000000; // 2643 :   0 - 0x0
      12'hA54: dout <= 8'b00000000; // 2644 :   0 - 0x0
      12'hA55: dout <= 8'b00000000; // 2645 :   0 - 0x0
      12'hA56: dout <= 8'b00000000; // 2646 :   0 - 0x0
      12'hA57: dout <= 8'b00000000; // 2647 :   0 - 0x0
      12'hA58: dout <= 8'b00000000; // 2648 :   0 - 0x0 -- Background 0x4b
      12'hA59: dout <= 8'b00000000; // 2649 :   0 - 0x0
      12'hA5A: dout <= 8'b00000000; // 2650 :   0 - 0x0
      12'hA5B: dout <= 8'b00000000; // 2651 :   0 - 0x0
      12'hA5C: dout <= 8'b00000000; // 2652 :   0 - 0x0
      12'hA5D: dout <= 8'b00000000; // 2653 :   0 - 0x0
      12'hA5E: dout <= 8'b00000000; // 2654 :   0 - 0x0
      12'hA5F: dout <= 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout <= 8'b00000000; // 2656 :   0 - 0x0 -- Background 0x4c
      12'hA61: dout <= 8'b00000000; // 2657 :   0 - 0x0
      12'hA62: dout <= 8'b00000000; // 2658 :   0 - 0x0
      12'hA63: dout <= 8'b00000000; // 2659 :   0 - 0x0
      12'hA64: dout <= 8'b00000000; // 2660 :   0 - 0x0
      12'hA65: dout <= 8'b00000000; // 2661 :   0 - 0x0
      12'hA66: dout <= 8'b00000000; // 2662 :   0 - 0x0
      12'hA67: dout <= 8'b00000000; // 2663 :   0 - 0x0
      12'hA68: dout <= 8'b00000000; // 2664 :   0 - 0x0 -- Background 0x4d
      12'hA69: dout <= 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout <= 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout <= 8'b00000000; // 2667 :   0 - 0x0
      12'hA6C: dout <= 8'b00000000; // 2668 :   0 - 0x0
      12'hA6D: dout <= 8'b00000000; // 2669 :   0 - 0x0
      12'hA6E: dout <= 8'b00000000; // 2670 :   0 - 0x0
      12'hA6F: dout <= 8'b00000000; // 2671 :   0 - 0x0
      12'hA70: dout <= 8'b00000000; // 2672 :   0 - 0x0 -- Background 0x4e
      12'hA71: dout <= 8'b00000000; // 2673 :   0 - 0x0
      12'hA72: dout <= 8'b00000000; // 2674 :   0 - 0x0
      12'hA73: dout <= 8'b00000000; // 2675 :   0 - 0x0
      12'hA74: dout <= 8'b00000000; // 2676 :   0 - 0x0
      12'hA75: dout <= 8'b00000000; // 2677 :   0 - 0x0
      12'hA76: dout <= 8'b00000000; // 2678 :   0 - 0x0
      12'hA77: dout <= 8'b00000000; // 2679 :   0 - 0x0
      12'hA78: dout <= 8'b00000000; // 2680 :   0 - 0x0 -- Background 0x4f
      12'hA79: dout <= 8'b00000000; // 2681 :   0 - 0x0
      12'hA7A: dout <= 8'b00000000; // 2682 :   0 - 0x0
      12'hA7B: dout <= 8'b00000000; // 2683 :   0 - 0x0
      12'hA7C: dout <= 8'b00000000; // 2684 :   0 - 0x0
      12'hA7D: dout <= 8'b00000000; // 2685 :   0 - 0x0
      12'hA7E: dout <= 8'b00000000; // 2686 :   0 - 0x0
      12'hA7F: dout <= 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout <= 8'b00000000; // 2688 :   0 - 0x0 -- Background 0x50
      12'hA81: dout <= 8'b00000000; // 2689 :   0 - 0x0
      12'hA82: dout <= 8'b00000000; // 2690 :   0 - 0x0
      12'hA83: dout <= 8'b00000000; // 2691 :   0 - 0x0
      12'hA84: dout <= 8'b00000000; // 2692 :   0 - 0x0
      12'hA85: dout <= 8'b00000000; // 2693 :   0 - 0x0
      12'hA86: dout <= 8'b00000000; // 2694 :   0 - 0x0
      12'hA87: dout <= 8'b00000000; // 2695 :   0 - 0x0
      12'hA88: dout <= 8'b00000000; // 2696 :   0 - 0x0 -- Background 0x51
      12'hA89: dout <= 8'b00000000; // 2697 :   0 - 0x0
      12'hA8A: dout <= 8'b00000000; // 2698 :   0 - 0x0
      12'hA8B: dout <= 8'b00000000; // 2699 :   0 - 0x0
      12'hA8C: dout <= 8'b00000000; // 2700 :   0 - 0x0
      12'hA8D: dout <= 8'b00000000; // 2701 :   0 - 0x0
      12'hA8E: dout <= 8'b00000000; // 2702 :   0 - 0x0
      12'hA8F: dout <= 8'b00000000; // 2703 :   0 - 0x0
      12'hA90: dout <= 8'b00000000; // 2704 :   0 - 0x0 -- Background 0x52
      12'hA91: dout <= 8'b00000000; // 2705 :   0 - 0x0
      12'hA92: dout <= 8'b00000000; // 2706 :   0 - 0x0
      12'hA93: dout <= 8'b00000000; // 2707 :   0 - 0x0
      12'hA94: dout <= 8'b00000000; // 2708 :   0 - 0x0
      12'hA95: dout <= 8'b00000000; // 2709 :   0 - 0x0
      12'hA96: dout <= 8'b00000000; // 2710 :   0 - 0x0
      12'hA97: dout <= 8'b00000000; // 2711 :   0 - 0x0
      12'hA98: dout <= 8'b00000000; // 2712 :   0 - 0x0 -- Background 0x53
      12'hA99: dout <= 8'b00000000; // 2713 :   0 - 0x0
      12'hA9A: dout <= 8'b00000000; // 2714 :   0 - 0x0
      12'hA9B: dout <= 8'b00000000; // 2715 :   0 - 0x0
      12'hA9C: dout <= 8'b00000000; // 2716 :   0 - 0x0
      12'hA9D: dout <= 8'b00000000; // 2717 :   0 - 0x0
      12'hA9E: dout <= 8'b00000000; // 2718 :   0 - 0x0
      12'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout <= 8'b00000000; // 2720 :   0 - 0x0 -- Background 0x54
      12'hAA1: dout <= 8'b00000000; // 2721 :   0 - 0x0
      12'hAA2: dout <= 8'b00000000; // 2722 :   0 - 0x0
      12'hAA3: dout <= 8'b00000000; // 2723 :   0 - 0x0
      12'hAA4: dout <= 8'b00000000; // 2724 :   0 - 0x0
      12'hAA5: dout <= 8'b00000000; // 2725 :   0 - 0x0
      12'hAA6: dout <= 8'b00000000; // 2726 :   0 - 0x0
      12'hAA7: dout <= 8'b00000000; // 2727 :   0 - 0x0
      12'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0 -- Background 0x55
      12'hAA9: dout <= 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout <= 8'b00000000; // 2730 :   0 - 0x0
      12'hAAB: dout <= 8'b00000000; // 2731 :   0 - 0x0
      12'hAAC: dout <= 8'b00000000; // 2732 :   0 - 0x0
      12'hAAD: dout <= 8'b00000000; // 2733 :   0 - 0x0
      12'hAAE: dout <= 8'b00000000; // 2734 :   0 - 0x0
      12'hAAF: dout <= 8'b00000000; // 2735 :   0 - 0x0
      12'hAB0: dout <= 8'b00000000; // 2736 :   0 - 0x0 -- Background 0x56
      12'hAB1: dout <= 8'b00000000; // 2737 :   0 - 0x0
      12'hAB2: dout <= 8'b00000000; // 2738 :   0 - 0x0
      12'hAB3: dout <= 8'b00000000; // 2739 :   0 - 0x0
      12'hAB4: dout <= 8'b00000000; // 2740 :   0 - 0x0
      12'hAB5: dout <= 8'b00000000; // 2741 :   0 - 0x0
      12'hAB6: dout <= 8'b00000000; // 2742 :   0 - 0x0
      12'hAB7: dout <= 8'b00000000; // 2743 :   0 - 0x0
      12'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0 -- Background 0x57
      12'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout <= 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout <= 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout <= 8'b00000000; // 2752 :   0 - 0x0 -- Background 0x58
      12'hAC1: dout <= 8'b00000000; // 2753 :   0 - 0x0
      12'hAC2: dout <= 8'b00000000; // 2754 :   0 - 0x0
      12'hAC3: dout <= 8'b00000000; // 2755 :   0 - 0x0
      12'hAC4: dout <= 8'b00000000; // 2756 :   0 - 0x0
      12'hAC5: dout <= 8'b00000000; // 2757 :   0 - 0x0
      12'hAC6: dout <= 8'b00000000; // 2758 :   0 - 0x0
      12'hAC7: dout <= 8'b00000000; // 2759 :   0 - 0x0
      12'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0 -- Background 0x59
      12'hAC9: dout <= 8'b00000000; // 2761 :   0 - 0x0
      12'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout <= 8'b00000000; // 2763 :   0 - 0x0
      12'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      12'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout <= 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout <= 8'b00000000; // 2768 :   0 - 0x0 -- Background 0x5a
      12'hAD1: dout <= 8'b00000000; // 2769 :   0 - 0x0
      12'hAD2: dout <= 8'b00000000; // 2770 :   0 - 0x0
      12'hAD3: dout <= 8'b00000000; // 2771 :   0 - 0x0
      12'hAD4: dout <= 8'b00000000; // 2772 :   0 - 0x0
      12'hAD5: dout <= 8'b00000000; // 2773 :   0 - 0x0
      12'hAD6: dout <= 8'b00000000; // 2774 :   0 - 0x0
      12'hAD7: dout <= 8'b00000000; // 2775 :   0 - 0x0
      12'hAD8: dout <= 8'b00000000; // 2776 :   0 - 0x0 -- Background 0x5b
      12'hAD9: dout <= 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout <= 8'b00000000; // 2778 :   0 - 0x0
      12'hADB: dout <= 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout <= 8'b00000000; // 2780 :   0 - 0x0
      12'hADD: dout <= 8'b00000000; // 2781 :   0 - 0x0
      12'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      12'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout <= 8'b00000000; // 2784 :   0 - 0x0 -- Background 0x5c
      12'hAE1: dout <= 8'b00000000; // 2785 :   0 - 0x0
      12'hAE2: dout <= 8'b00000000; // 2786 :   0 - 0x0
      12'hAE3: dout <= 8'b00000000; // 2787 :   0 - 0x0
      12'hAE4: dout <= 8'b00000000; // 2788 :   0 - 0x0
      12'hAE5: dout <= 8'b00000000; // 2789 :   0 - 0x0
      12'hAE6: dout <= 8'b00000000; // 2790 :   0 - 0x0
      12'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0 -- Background 0x5d
      12'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout <= 8'b00000000; // 2794 :   0 - 0x0
      12'hAEB: dout <= 8'b00000000; // 2795 :   0 - 0x0
      12'hAEC: dout <= 8'b00000000; // 2796 :   0 - 0x0
      12'hAED: dout <= 8'b00000000; // 2797 :   0 - 0x0
      12'hAEE: dout <= 8'b00000000; // 2798 :   0 - 0x0
      12'hAEF: dout <= 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout <= 8'b00000000; // 2800 :   0 - 0x0 -- Background 0x5e
      12'hAF1: dout <= 8'b00000000; // 2801 :   0 - 0x0
      12'hAF2: dout <= 8'b00000000; // 2802 :   0 - 0x0
      12'hAF3: dout <= 8'b00000000; // 2803 :   0 - 0x0
      12'hAF4: dout <= 8'b00000000; // 2804 :   0 - 0x0
      12'hAF5: dout <= 8'b00000000; // 2805 :   0 - 0x0
      12'hAF6: dout <= 8'b00000000; // 2806 :   0 - 0x0
      12'hAF7: dout <= 8'b00000000; // 2807 :   0 - 0x0
      12'hAF8: dout <= 8'b00000000; // 2808 :   0 - 0x0 -- Background 0x5f
      12'hAF9: dout <= 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout <= 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout <= 8'b00000000; // 2811 :   0 - 0x0
      12'hAFC: dout <= 8'b00000000; // 2812 :   0 - 0x0
      12'hAFD: dout <= 8'b00000000; // 2813 :   0 - 0x0
      12'hAFE: dout <= 8'b00000000; // 2814 :   0 - 0x0
      12'hAFF: dout <= 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout <= 8'b00000000; // 2816 :   0 - 0x0 -- Background 0x60
      12'hB01: dout <= 8'b00000000; // 2817 :   0 - 0x0
      12'hB02: dout <= 8'b00000000; // 2818 :   0 - 0x0
      12'hB03: dout <= 8'b00000000; // 2819 :   0 - 0x0
      12'hB04: dout <= 8'b00000000; // 2820 :   0 - 0x0
      12'hB05: dout <= 8'b00000000; // 2821 :   0 - 0x0
      12'hB06: dout <= 8'b00000000; // 2822 :   0 - 0x0
      12'hB07: dout <= 8'b00000000; // 2823 :   0 - 0x0
      12'hB08: dout <= 8'b00000000; // 2824 :   0 - 0x0 -- Background 0x61
      12'hB09: dout <= 8'b00000000; // 2825 :   0 - 0x0
      12'hB0A: dout <= 8'b00000000; // 2826 :   0 - 0x0
      12'hB0B: dout <= 8'b00000000; // 2827 :   0 - 0x0
      12'hB0C: dout <= 8'b00000000; // 2828 :   0 - 0x0
      12'hB0D: dout <= 8'b00000000; // 2829 :   0 - 0x0
      12'hB0E: dout <= 8'b00000000; // 2830 :   0 - 0x0
      12'hB0F: dout <= 8'b00000000; // 2831 :   0 - 0x0
      12'hB10: dout <= 8'b00000000; // 2832 :   0 - 0x0 -- Background 0x62
      12'hB11: dout <= 8'b00000000; // 2833 :   0 - 0x0
      12'hB12: dout <= 8'b00000000; // 2834 :   0 - 0x0
      12'hB13: dout <= 8'b00000000; // 2835 :   0 - 0x0
      12'hB14: dout <= 8'b00000000; // 2836 :   0 - 0x0
      12'hB15: dout <= 8'b00000000; // 2837 :   0 - 0x0
      12'hB16: dout <= 8'b00000000; // 2838 :   0 - 0x0
      12'hB17: dout <= 8'b00000000; // 2839 :   0 - 0x0
      12'hB18: dout <= 8'b00000000; // 2840 :   0 - 0x0 -- Background 0x63
      12'hB19: dout <= 8'b00000000; // 2841 :   0 - 0x0
      12'hB1A: dout <= 8'b00000000; // 2842 :   0 - 0x0
      12'hB1B: dout <= 8'b00000000; // 2843 :   0 - 0x0
      12'hB1C: dout <= 8'b00000000; // 2844 :   0 - 0x0
      12'hB1D: dout <= 8'b00000000; // 2845 :   0 - 0x0
      12'hB1E: dout <= 8'b00000000; // 2846 :   0 - 0x0
      12'hB1F: dout <= 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout <= 8'b00000000; // 2848 :   0 - 0x0 -- Background 0x64
      12'hB21: dout <= 8'b00000000; // 2849 :   0 - 0x0
      12'hB22: dout <= 8'b00000000; // 2850 :   0 - 0x0
      12'hB23: dout <= 8'b00000000; // 2851 :   0 - 0x0
      12'hB24: dout <= 8'b00000000; // 2852 :   0 - 0x0
      12'hB25: dout <= 8'b00000000; // 2853 :   0 - 0x0
      12'hB26: dout <= 8'b00000000; // 2854 :   0 - 0x0
      12'hB27: dout <= 8'b00000000; // 2855 :   0 - 0x0
      12'hB28: dout <= 8'b00000000; // 2856 :   0 - 0x0 -- Background 0x65
      12'hB29: dout <= 8'b00000000; // 2857 :   0 - 0x0
      12'hB2A: dout <= 8'b00000000; // 2858 :   0 - 0x0
      12'hB2B: dout <= 8'b00000000; // 2859 :   0 - 0x0
      12'hB2C: dout <= 8'b00000000; // 2860 :   0 - 0x0
      12'hB2D: dout <= 8'b00000000; // 2861 :   0 - 0x0
      12'hB2E: dout <= 8'b00000000; // 2862 :   0 - 0x0
      12'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout <= 8'b00000000; // 2864 :   0 - 0x0 -- Background 0x66
      12'hB31: dout <= 8'b00000000; // 2865 :   0 - 0x0
      12'hB32: dout <= 8'b00000000; // 2866 :   0 - 0x0
      12'hB33: dout <= 8'b00000000; // 2867 :   0 - 0x0
      12'hB34: dout <= 8'b00000000; // 2868 :   0 - 0x0
      12'hB35: dout <= 8'b00000000; // 2869 :   0 - 0x0
      12'hB36: dout <= 8'b00000000; // 2870 :   0 - 0x0
      12'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      12'hB38: dout <= 8'b00000000; // 2872 :   0 - 0x0 -- Background 0x67
      12'hB39: dout <= 8'b00000000; // 2873 :   0 - 0x0
      12'hB3A: dout <= 8'b00000000; // 2874 :   0 - 0x0
      12'hB3B: dout <= 8'b00000000; // 2875 :   0 - 0x0
      12'hB3C: dout <= 8'b00000000; // 2876 :   0 - 0x0
      12'hB3D: dout <= 8'b00000000; // 2877 :   0 - 0x0
      12'hB3E: dout <= 8'b00000000; // 2878 :   0 - 0x0
      12'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout <= 8'b00000000; // 2880 :   0 - 0x0 -- Background 0x68
      12'hB41: dout <= 8'b00000000; // 2881 :   0 - 0x0
      12'hB42: dout <= 8'b00000000; // 2882 :   0 - 0x0
      12'hB43: dout <= 8'b00000000; // 2883 :   0 - 0x0
      12'hB44: dout <= 8'b00000000; // 2884 :   0 - 0x0
      12'hB45: dout <= 8'b00000000; // 2885 :   0 - 0x0
      12'hB46: dout <= 8'b00000000; // 2886 :   0 - 0x0
      12'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout <= 8'b00000000; // 2888 :   0 - 0x0 -- Background 0x69
      12'hB49: dout <= 8'b00000000; // 2889 :   0 - 0x0
      12'hB4A: dout <= 8'b00000000; // 2890 :   0 - 0x0
      12'hB4B: dout <= 8'b00000000; // 2891 :   0 - 0x0
      12'hB4C: dout <= 8'b00000000; // 2892 :   0 - 0x0
      12'hB4D: dout <= 8'b00000000; // 2893 :   0 - 0x0
      12'hB4E: dout <= 8'b00000000; // 2894 :   0 - 0x0
      12'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout <= 8'b00000000; // 2896 :   0 - 0x0 -- Background 0x6a
      12'hB51: dout <= 8'b00000000; // 2897 :   0 - 0x0
      12'hB52: dout <= 8'b00000000; // 2898 :   0 - 0x0
      12'hB53: dout <= 8'b00000000; // 2899 :   0 - 0x0
      12'hB54: dout <= 8'b00000000; // 2900 :   0 - 0x0
      12'hB55: dout <= 8'b00000000; // 2901 :   0 - 0x0
      12'hB56: dout <= 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout <= 8'b00000000; // 2904 :   0 - 0x0 -- Background 0x6b
      12'hB59: dout <= 8'b00000000; // 2905 :   0 - 0x0
      12'hB5A: dout <= 8'b00000000; // 2906 :   0 - 0x0
      12'hB5B: dout <= 8'b00000000; // 2907 :   0 - 0x0
      12'hB5C: dout <= 8'b00000000; // 2908 :   0 - 0x0
      12'hB5D: dout <= 8'b00000000; // 2909 :   0 - 0x0
      12'hB5E: dout <= 8'b00000000; // 2910 :   0 - 0x0
      12'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout <= 8'b00000000; // 2912 :   0 - 0x0 -- Background 0x6c
      12'hB61: dout <= 8'b00000000; // 2913 :   0 - 0x0
      12'hB62: dout <= 8'b00000000; // 2914 :   0 - 0x0
      12'hB63: dout <= 8'b00000000; // 2915 :   0 - 0x0
      12'hB64: dout <= 8'b00000000; // 2916 :   0 - 0x0
      12'hB65: dout <= 8'b00000000; // 2917 :   0 - 0x0
      12'hB66: dout <= 8'b00000000; // 2918 :   0 - 0x0
      12'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout <= 8'b00000000; // 2920 :   0 - 0x0 -- Background 0x6d
      12'hB69: dout <= 8'b00000000; // 2921 :   0 - 0x0
      12'hB6A: dout <= 8'b00000000; // 2922 :   0 - 0x0
      12'hB6B: dout <= 8'b00000000; // 2923 :   0 - 0x0
      12'hB6C: dout <= 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout <= 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout <= 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout <= 8'b00000000; // 2928 :   0 - 0x0 -- Background 0x6e
      12'hB71: dout <= 8'b00000000; // 2929 :   0 - 0x0
      12'hB72: dout <= 8'b00000000; // 2930 :   0 - 0x0
      12'hB73: dout <= 8'b00000000; // 2931 :   0 - 0x0
      12'hB74: dout <= 8'b00000000; // 2932 :   0 - 0x0
      12'hB75: dout <= 8'b00000000; // 2933 :   0 - 0x0
      12'hB76: dout <= 8'b00000000; // 2934 :   0 - 0x0
      12'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout <= 8'b00000000; // 2936 :   0 - 0x0 -- Background 0x6f
      12'hB79: dout <= 8'b00000000; // 2937 :   0 - 0x0
      12'hB7A: dout <= 8'b00000000; // 2938 :   0 - 0x0
      12'hB7B: dout <= 8'b00000000; // 2939 :   0 - 0x0
      12'hB7C: dout <= 8'b00000000; // 2940 :   0 - 0x0
      12'hB7D: dout <= 8'b00000000; // 2941 :   0 - 0x0
      12'hB7E: dout <= 8'b00000000; // 2942 :   0 - 0x0
      12'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout <= 8'b00000000; // 2944 :   0 - 0x0 -- Background 0x70
      12'hB81: dout <= 8'b00000000; // 2945 :   0 - 0x0
      12'hB82: dout <= 8'b00000000; // 2946 :   0 - 0x0
      12'hB83: dout <= 8'b00000000; // 2947 :   0 - 0x0
      12'hB84: dout <= 8'b00000000; // 2948 :   0 - 0x0
      12'hB85: dout <= 8'b00000000; // 2949 :   0 - 0x0
      12'hB86: dout <= 8'b00000000; // 2950 :   0 - 0x0
      12'hB87: dout <= 8'b00000000; // 2951 :   0 - 0x0
      12'hB88: dout <= 8'b00000000; // 2952 :   0 - 0x0 -- Background 0x71
      12'hB89: dout <= 8'b00000000; // 2953 :   0 - 0x0
      12'hB8A: dout <= 8'b00000000; // 2954 :   0 - 0x0
      12'hB8B: dout <= 8'b00000000; // 2955 :   0 - 0x0
      12'hB8C: dout <= 8'b00000000; // 2956 :   0 - 0x0
      12'hB8D: dout <= 8'b00000000; // 2957 :   0 - 0x0
      12'hB8E: dout <= 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b00000000; // 2960 :   0 - 0x0 -- Background 0x72
      12'hB91: dout <= 8'b00000000; // 2961 :   0 - 0x0
      12'hB92: dout <= 8'b00000000; // 2962 :   0 - 0x0
      12'hB93: dout <= 8'b00000000; // 2963 :   0 - 0x0
      12'hB94: dout <= 8'b00000000; // 2964 :   0 - 0x0
      12'hB95: dout <= 8'b00000000; // 2965 :   0 - 0x0
      12'hB96: dout <= 8'b00000000; // 2966 :   0 - 0x0
      12'hB97: dout <= 8'b00000000; // 2967 :   0 - 0x0
      12'hB98: dout <= 8'b00000000; // 2968 :   0 - 0x0 -- Background 0x73
      12'hB99: dout <= 8'b00000000; // 2969 :   0 - 0x0
      12'hB9A: dout <= 8'b00000000; // 2970 :   0 - 0x0
      12'hB9B: dout <= 8'b00000000; // 2971 :   0 - 0x0
      12'hB9C: dout <= 8'b00000000; // 2972 :   0 - 0x0
      12'hB9D: dout <= 8'b00000000; // 2973 :   0 - 0x0
      12'hB9E: dout <= 8'b00000000; // 2974 :   0 - 0x0
      12'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout <= 8'b00000000; // 2976 :   0 - 0x0 -- Background 0x74
      12'hBA1: dout <= 8'b00000000; // 2977 :   0 - 0x0
      12'hBA2: dout <= 8'b00000000; // 2978 :   0 - 0x0
      12'hBA3: dout <= 8'b00000000; // 2979 :   0 - 0x0
      12'hBA4: dout <= 8'b00000000; // 2980 :   0 - 0x0
      12'hBA5: dout <= 8'b00000000; // 2981 :   0 - 0x0
      12'hBA6: dout <= 8'b00000000; // 2982 :   0 - 0x0
      12'hBA7: dout <= 8'b00000000; // 2983 :   0 - 0x0
      12'hBA8: dout <= 8'b00000000; // 2984 :   0 - 0x0 -- Background 0x75
      12'hBA9: dout <= 8'b00000000; // 2985 :   0 - 0x0
      12'hBAA: dout <= 8'b00000000; // 2986 :   0 - 0x0
      12'hBAB: dout <= 8'b00000000; // 2987 :   0 - 0x0
      12'hBAC: dout <= 8'b00000000; // 2988 :   0 - 0x0
      12'hBAD: dout <= 8'b00000000; // 2989 :   0 - 0x0
      12'hBAE: dout <= 8'b00000000; // 2990 :   0 - 0x0
      12'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout <= 8'b00000000; // 2992 :   0 - 0x0 -- Background 0x76
      12'hBB1: dout <= 8'b00000000; // 2993 :   0 - 0x0
      12'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      12'hBB3: dout <= 8'b00000000; // 2995 :   0 - 0x0
      12'hBB4: dout <= 8'b00000000; // 2996 :   0 - 0x0
      12'hBB5: dout <= 8'b00000000; // 2997 :   0 - 0x0
      12'hBB6: dout <= 8'b00000000; // 2998 :   0 - 0x0
      12'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0 -- Background 0x77
      12'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      12'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      12'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      12'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      12'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b00000000; // 3008 :   0 - 0x0 -- Background 0x78
      12'hBC1: dout <= 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout <= 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout <= 8'b00000000; // 3011 :   0 - 0x0
      12'hBC4: dout <= 8'b00000000; // 3012 :   0 - 0x0
      12'hBC5: dout <= 8'b00000000; // 3013 :   0 - 0x0
      12'hBC6: dout <= 8'b00000000; // 3014 :   0 - 0x0
      12'hBC7: dout <= 8'b00000000; // 3015 :   0 - 0x0
      12'hBC8: dout <= 8'b00000000; // 3016 :   0 - 0x0 -- Background 0x79
      12'hBC9: dout <= 8'b00000000; // 3017 :   0 - 0x0
      12'hBCA: dout <= 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout <= 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout <= 8'b00000000; // 3021 :   0 - 0x0
      12'hBCE: dout <= 8'b00000000; // 3022 :   0 - 0x0
      12'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout <= 8'b00000000; // 3024 :   0 - 0x0 -- Background 0x7a
      12'hBD1: dout <= 8'b00000000; // 3025 :   0 - 0x0
      12'hBD2: dout <= 8'b00000000; // 3026 :   0 - 0x0
      12'hBD3: dout <= 8'b00000000; // 3027 :   0 - 0x0
      12'hBD4: dout <= 8'b00000000; // 3028 :   0 - 0x0
      12'hBD5: dout <= 8'b00000000; // 3029 :   0 - 0x0
      12'hBD6: dout <= 8'b00000000; // 3030 :   0 - 0x0
      12'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0 -- Background 0x7b
      12'hBD9: dout <= 8'b00000000; // 3033 :   0 - 0x0
      12'hBDA: dout <= 8'b00000000; // 3034 :   0 - 0x0
      12'hBDB: dout <= 8'b00000000; // 3035 :   0 - 0x0
      12'hBDC: dout <= 8'b00000000; // 3036 :   0 - 0x0
      12'hBDD: dout <= 8'b00000000; // 3037 :   0 - 0x0
      12'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout <= 8'b00000000; // 3040 :   0 - 0x0 -- Background 0x7c
      12'hBE1: dout <= 8'b00000000; // 3041 :   0 - 0x0
      12'hBE2: dout <= 8'b00000000; // 3042 :   0 - 0x0
      12'hBE3: dout <= 8'b00000000; // 3043 :   0 - 0x0
      12'hBE4: dout <= 8'b00000000; // 3044 :   0 - 0x0
      12'hBE5: dout <= 8'b00000000; // 3045 :   0 - 0x0
      12'hBE6: dout <= 8'b00000000; // 3046 :   0 - 0x0
      12'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      12'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0 -- Background 0x7d
      12'hBE9: dout <= 8'b00000000; // 3049 :   0 - 0x0
      12'hBEA: dout <= 8'b00000000; // 3050 :   0 - 0x0
      12'hBEB: dout <= 8'b00000000; // 3051 :   0 - 0x0
      12'hBEC: dout <= 8'b00000000; // 3052 :   0 - 0x0
      12'hBED: dout <= 8'b00000000; // 3053 :   0 - 0x0
      12'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      12'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Background 0x7e
      12'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      12'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      12'hBF4: dout <= 8'b00000000; // 3060 :   0 - 0x0
      12'hBF5: dout <= 8'b00000000; // 3061 :   0 - 0x0
      12'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      12'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0 -- Background 0x7f
      12'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      12'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      12'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      12'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout <= 8'b01000000; // 3072 :  64 - 0x40 -- Background 0x80
      12'hC01: dout <= 8'b00001000; // 3073 :   8 - 0x8
      12'hC02: dout <= 8'b00000010; // 3074 :   2 - 0x2
      12'hC03: dout <= 8'b00100000; // 3075 :  32 - 0x20
      12'hC04: dout <= 8'b00000100; // 3076 :   4 - 0x4
      12'hC05: dout <= 8'b01000000; // 3077 :  64 - 0x40
      12'hC06: dout <= 8'b00000001; // 3078 :   1 - 0x1
      12'hC07: dout <= 8'b00010000; // 3079 :  16 - 0x10
      12'hC08: dout <= 8'b00000000; // 3080 :   0 - 0x0 -- Background 0x81
      12'hC09: dout <= 8'b00010001; // 3081 :  17 - 0x11
      12'hC0A: dout <= 8'b00000000; // 3082 :   0 - 0x0
      12'hC0B: dout <= 8'b00100000; // 3083 :  32 - 0x20
      12'hC0C: dout <= 8'b10001000; // 3084 : 136 - 0x88
      12'hC0D: dout <= 8'b00000010; // 3085 :   2 - 0x2
      12'hC0E: dout <= 8'b00100000; // 3086 :  32 - 0x20
      12'hC0F: dout <= 8'b01000000; // 3087 :  64 - 0x40
      12'hC10: dout <= 8'b00000001; // 3088 :   1 - 0x1 -- Background 0x82
      12'hC11: dout <= 8'b00010000; // 3089 :  16 - 0x10
      12'hC12: dout <= 8'b01000000; // 3090 :  64 - 0x40
      12'hC13: dout <= 8'b00001000; // 3091 :   8 - 0x8
      12'hC14: dout <= 8'b00000010; // 3092 :   2 - 0x2
      12'hC15: dout <= 8'b00100000; // 3093 :  32 - 0x20
      12'hC16: dout <= 8'b00000100; // 3094 :   4 - 0x4
      12'hC17: dout <= 8'b01000000; // 3095 :  64 - 0x40
      12'hC18: dout <= 8'b00010000; // 3096 :  16 - 0x10 -- Background 0x83
      12'hC19: dout <= 8'b00000000; // 3097 :   0 - 0x0
      12'hC1A: dout <= 8'b01000100; // 3098 :  68 - 0x44
      12'hC1B: dout <= 8'b00000000; // 3099 :   0 - 0x0
      12'hC1C: dout <= 8'b00001000; // 3100 :   8 - 0x8
      12'hC1D: dout <= 8'b00100010; // 3101 :  34 - 0x22
      12'hC1E: dout <= 8'b10000000; // 3102 : 128 - 0x80
      12'hC1F: dout <= 8'b00001000; // 3103 :   8 - 0x8
      12'hC20: dout <= 8'b00010100; // 3104 :  20 - 0x14 -- Background 0x84
      12'hC21: dout <= 8'b10110101; // 3105 : 181 - 0xb5
      12'hC22: dout <= 8'b01000100; // 3106 :  68 - 0x44
      12'hC23: dout <= 8'b01001010; // 3107 :  74 - 0x4a
      12'hC24: dout <= 8'b10010010; // 3108 : 146 - 0x92
      12'hC25: dout <= 8'b10010010; // 3109 : 146 - 0x92
      12'hC26: dout <= 8'b01000100; // 3110 :  68 - 0x44
      12'hC27: dout <= 8'b01001001; // 3111 :  73 - 0x49
      12'hC28: dout <= 8'b01000010; // 3112 :  66 - 0x42 -- Background 0x85
      12'hC29: dout <= 8'b01001010; // 3113 :  74 - 0x4a
      12'hC2A: dout <= 8'b11001010; // 3114 : 202 - 0xca
      12'hC2B: dout <= 8'b00101001; // 3115 :  41 - 0x29
      12'hC2C: dout <= 8'b10100110; // 3116 : 166 - 0xa6
      12'hC2D: dout <= 8'b10010010; // 3117 : 146 - 0x92
      12'hC2E: dout <= 8'b10001001; // 3118 : 137 - 0x89
      12'hC2F: dout <= 8'b00101101; // 3119 :  45 - 0x2d
      12'hC30: dout <= 8'b10001000; // 3120 : 136 - 0x88 -- Background 0x86
      12'hC31: dout <= 8'b00101001; // 3121 :  41 - 0x29
      12'hC32: dout <= 8'b10000010; // 3122 : 130 - 0x82
      12'hC33: dout <= 8'b10110110; // 3123 : 182 - 0xb6
      12'hC34: dout <= 8'b10001000; // 3124 : 136 - 0x88
      12'hC35: dout <= 8'b01001001; // 3125 :  73 - 0x49
      12'hC36: dout <= 8'b01010010; // 3126 :  82 - 0x52
      12'hC37: dout <= 8'b01010010; // 3127 :  82 - 0x52
      12'hC38: dout <= 8'b10110010; // 3128 : 178 - 0xb2 -- Background 0x87
      12'hC39: dout <= 8'b01001010; // 3129 :  74 - 0x4a
      12'hC3A: dout <= 8'b10101001; // 3130 : 169 - 0xa9
      12'hC3B: dout <= 8'b10100100; // 3131 : 164 - 0xa4
      12'hC3C: dout <= 8'b01100010; // 3132 :  98 - 0x62
      12'hC3D: dout <= 8'b01001011; // 3133 :  75 - 0x4b
      12'hC3E: dout <= 8'b10010000; // 3134 : 144 - 0x90
      12'hC3F: dout <= 8'b10010010; // 3135 : 146 - 0x92
      12'hC40: dout <= 8'b01100000; // 3136 :  96 - 0x60 -- Background 0x88
      12'hC41: dout <= 8'b11110000; // 3137 : 240 - 0xf0
      12'hC42: dout <= 8'b11110000; // 3138 : 240 - 0xf0
      12'hC43: dout <= 8'b01101110; // 3139 : 110 - 0x6e
      12'hC44: dout <= 8'b00011111; // 3140 :  31 - 0x1f
      12'hC45: dout <= 8'b00011111; // 3141 :  31 - 0x1f
      12'hC46: dout <= 8'b00011111; // 3142 :  31 - 0x1f
      12'hC47: dout <= 8'b00001110; // 3143 :  14 - 0xe
      12'hC48: dout <= 8'b01100000; // 3144 :  96 - 0x60 -- Background 0x89
      12'hC49: dout <= 8'b11110000; // 3145 : 240 - 0xf0
      12'hC4A: dout <= 8'b11111110; // 3146 : 254 - 0xfe
      12'hC4B: dout <= 8'b01111111; // 3147 : 127 - 0x7f
      12'hC4C: dout <= 8'b00011111; // 3148 :  31 - 0x1f
      12'hC4D: dout <= 8'b00011111; // 3149 :  31 - 0x1f
      12'hC4E: dout <= 8'b00001110; // 3150 :  14 - 0xe
      12'hC4F: dout <= 8'b00000000; // 3151 :   0 - 0x0
      12'hC50: dout <= 8'b01000000; // 3152 :  64 - 0x40 -- Background 0x8a
      12'hC51: dout <= 8'b00001000; // 3153 :   8 - 0x8
      12'hC52: dout <= 8'b00000010; // 3154 :   2 - 0x2
      12'hC53: dout <= 8'b00101000; // 3155 :  40 - 0x28
      12'hC54: dout <= 8'b00010100; // 3156 :  20 - 0x14
      12'hC55: dout <= 8'b01010100; // 3157 :  84 - 0x54
      12'hC56: dout <= 8'b00000001; // 3158 :   1 - 0x1
      12'hC57: dout <= 8'b00010000; // 3159 :  16 - 0x10
      12'hC58: dout <= 8'b01000000; // 3160 :  64 - 0x40 -- Background 0x8b
      12'hC59: dout <= 8'b00000000; // 3161 :   0 - 0x0
      12'hC5A: dout <= 8'b10010001; // 3162 : 145 - 0x91
      12'hC5B: dout <= 8'b00010100; // 3163 :  20 - 0x14
      12'hC5C: dout <= 8'b00101000; // 3164 :  40 - 0x28
      12'hC5D: dout <= 8'b10001010; // 3165 : 138 - 0x8a
      12'hC5E: dout <= 8'b01000000; // 3166 :  64 - 0x40
      12'hC5F: dout <= 8'b00100000; // 3167 :  32 - 0x20
      12'hC60: dout <= 8'b00000000; // 3168 :   0 - 0x0 -- Background 0x8c
      12'hC61: dout <= 8'b00000111; // 3169 :   7 - 0x7
      12'hC62: dout <= 8'b00011111; // 3170 :  31 - 0x1f
      12'hC63: dout <= 8'b00111111; // 3171 :  63 - 0x3f
      12'hC64: dout <= 8'b00111111; // 3172 :  63 - 0x3f
      12'hC65: dout <= 8'b01111111; // 3173 : 127 - 0x7f
      12'hC66: dout <= 8'b01111111; // 3174 : 127 - 0x7f
      12'hC67: dout <= 8'b01111111; // 3175 : 127 - 0x7f
      12'hC68: dout <= 8'b00000000; // 3176 :   0 - 0x0 -- Background 0x8d
      12'hC69: dout <= 8'b11100000; // 3177 : 224 - 0xe0
      12'hC6A: dout <= 8'b11111000; // 3178 : 248 - 0xf8
      12'hC6B: dout <= 8'b11111000; // 3179 : 248 - 0xf8
      12'hC6C: dout <= 8'b11110000; // 3180 : 240 - 0xf0
      12'hC6D: dout <= 8'b11111000; // 3181 : 248 - 0xf8
      12'hC6E: dout <= 8'b11110100; // 3182 : 244 - 0xf4
      12'hC6F: dout <= 8'b11111000; // 3183 : 248 - 0xf8
      12'hC70: dout <= 8'b01111111; // 3184 : 127 - 0x7f -- Background 0x8e
      12'hC71: dout <= 8'b00111111; // 3185 :  63 - 0x3f
      12'hC72: dout <= 8'b00111111; // 3186 :  63 - 0x3f
      12'hC73: dout <= 8'b00011111; // 3187 :  31 - 0x1f
      12'hC74: dout <= 8'b00011111; // 3188 :  31 - 0x1f
      12'hC75: dout <= 8'b00001111; // 3189 :  15 - 0xf
      12'hC76: dout <= 8'b00001111; // 3190 :  15 - 0xf
      12'hC77: dout <= 8'b00000111; // 3191 :   7 - 0x7
      12'hC78: dout <= 8'b11111110; // 3192 : 254 - 0xfe -- Background 0x8f
      12'hC79: dout <= 8'b11111100; // 3193 : 252 - 0xfc
      12'hC7A: dout <= 8'b11111100; // 3194 : 252 - 0xfc
      12'hC7B: dout <= 8'b11111000; // 3195 : 248 - 0xf8
      12'hC7C: dout <= 8'b11111000; // 3196 : 248 - 0xf8
      12'hC7D: dout <= 8'b11110000; // 3197 : 240 - 0xf0
      12'hC7E: dout <= 8'b11110000; // 3198 : 240 - 0xf0
      12'hC7F: dout <= 8'b11100000; // 3199 : 224 - 0xe0
      12'hC80: dout <= 8'b01000001; // 3200 :  65 - 0x41 -- Background 0x90
      12'hC81: dout <= 8'b00001000; // 3201 :   8 - 0x8
      12'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      12'hC83: dout <= 8'b00100000; // 3203 :  32 - 0x20
      12'hC84: dout <= 8'b00000100; // 3204 :   4 - 0x4
      12'hC85: dout <= 8'b00000001; // 3205 :   1 - 0x1
      12'hC86: dout <= 8'b01000000; // 3206 :  64 - 0x40
      12'hC87: dout <= 8'b00001000; // 3207 :   8 - 0x8
      12'hC88: dout <= 8'b00010001; // 3208 :  17 - 0x11 -- Background 0x91
      12'hC89: dout <= 8'b00000000; // 3209 :   0 - 0x0
      12'hC8A: dout <= 8'b10000100; // 3210 : 132 - 0x84
      12'hC8B: dout <= 8'b00000010; // 3211 :   2 - 0x2
      12'hC8C: dout <= 8'b00010000; // 3212 :  16 - 0x10
      12'hC8D: dout <= 8'b00000000; // 3213 :   0 - 0x0
      12'hC8E: dout <= 8'b01000010; // 3214 :  66 - 0x42
      12'hC8F: dout <= 8'b00000000; // 3215 :   0 - 0x0
      12'hC90: dout <= 8'b00000100; // 3216 :   4 - 0x4 -- Background 0x92
      12'hC91: dout <= 8'b01000000; // 3217 :  64 - 0x40
      12'hC92: dout <= 8'b00010000; // 3218 :  16 - 0x10
      12'hC93: dout <= 8'b00000010; // 3219 :   2 - 0x2
      12'hC94: dout <= 8'b00000000; // 3220 :   0 - 0x0
      12'hC95: dout <= 8'b01000000; // 3221 :  64 - 0x40
      12'hC96: dout <= 8'b00000100; // 3222 :   4 - 0x4
      12'hC97: dout <= 8'b00100000; // 3223 :  32 - 0x20
      12'hC98: dout <= 8'b01000010; // 3224 :  66 - 0x42 -- Background 0x93
      12'hC99: dout <= 8'b00000000; // 3225 :   0 - 0x0
      12'hC9A: dout <= 8'b10001000; // 3226 : 136 - 0x88
      12'hC9B: dout <= 8'b00000001; // 3227 :   1 - 0x1
      12'hC9C: dout <= 8'b00100000; // 3228 :  32 - 0x20
      12'hC9D: dout <= 8'b00000100; // 3229 :   4 - 0x4
      12'hC9E: dout <= 8'b00010000; // 3230 :  16 - 0x10
      12'hC9F: dout <= 8'b10000000; // 3231 : 128 - 0x80
      12'hCA0: dout <= 8'b11001000; // 3232 : 200 - 0xc8 -- Background 0x94
      12'hCA1: dout <= 8'b00101010; // 3233 :  42 - 0x2a
      12'hCA2: dout <= 8'b10100010; // 3234 : 162 - 0xa2
      12'hCA3: dout <= 8'b10010100; // 3235 : 148 - 0x94
      12'hCA4: dout <= 8'b10010001; // 3236 : 145 - 0x91
      12'hCA5: dout <= 8'b01010101; // 3237 :  85 - 0x55
      12'hCA6: dout <= 8'b01000100; // 3238 :  68 - 0x44
      12'hCA7: dout <= 8'b00010010; // 3239 :  18 - 0x12
      12'hCA8: dout <= 8'b10101010; // 3240 : 170 - 0xaa -- Background 0x95
      12'hCA9: dout <= 8'b10100010; // 3241 : 162 - 0xa2
      12'hCAA: dout <= 8'b00010010; // 3242 :  18 - 0x12
      12'hCAB: dout <= 8'b01010011; // 3243 :  83 - 0x53
      12'hCAC: dout <= 8'b01001100; // 3244 :  76 - 0x4c
      12'hCAD: dout <= 8'b01010101; // 3245 :  85 - 0x55
      12'hCAE: dout <= 8'b10010001; // 3246 : 145 - 0x91
      12'hCAF: dout <= 8'b01001000; // 3247 :  72 - 0x48
      12'hCB0: dout <= 8'b01010001; // 3248 :  81 - 0x51 -- Background 0x96
      12'hCB1: dout <= 8'b00010101; // 3249 :  21 - 0x15
      12'hCB2: dout <= 8'b10100100; // 3250 : 164 - 0xa4
      12'hCB3: dout <= 8'b10001100; // 3251 : 140 - 0x8c
      12'hCB4: dout <= 8'b10101010; // 3252 : 170 - 0xaa
      12'hCB5: dout <= 8'b00100010; // 3253 :  34 - 0x22
      12'hCB6: dout <= 8'b10010000; // 3254 : 144 - 0x90
      12'hCB7: dout <= 8'b01000110; // 3255 :  70 - 0x46
      12'hCB8: dout <= 8'b00010011; // 3256 :  19 - 0x13 -- Background 0x97
      12'hCB9: dout <= 8'b01010101; // 3257 :  85 - 0x55
      12'hCBA: dout <= 8'b01100100; // 3258 : 100 - 0x64
      12'hCBB: dout <= 8'b00010010; // 3259 :  18 - 0x12
      12'hCBC: dout <= 8'b10101010; // 3260 : 170 - 0xaa
      12'hCBD: dout <= 8'b10101000; // 3261 : 168 - 0xa8
      12'hCBE: dout <= 8'b10000100; // 3262 : 132 - 0x84
      12'hCBF: dout <= 8'b11010100; // 3263 : 212 - 0xd4
      12'hCC0: dout <= 8'b01100000; // 3264 :  96 - 0x60 -- Background 0x98
      12'hCC1: dout <= 8'b11110000; // 3265 : 240 - 0xf0
      12'hCC2: dout <= 8'b11111110; // 3266 : 254 - 0xfe
      12'hCC3: dout <= 8'b01111111; // 3267 : 127 - 0x7f
      12'hCC4: dout <= 8'b00011111; // 3268 :  31 - 0x1f
      12'hCC5: dout <= 8'b00011111; // 3269 :  31 - 0x1f
      12'hCC6: dout <= 8'b00001110; // 3270 :  14 - 0xe
      12'hCC7: dout <= 8'b00000000; // 3271 :   0 - 0x0
      12'hCC8: dout <= 8'b01100000; // 3272 :  96 - 0x60 -- Background 0x99
      12'hCC9: dout <= 8'b11110000; // 3273 : 240 - 0xf0
      12'hCCA: dout <= 8'b11110000; // 3274 : 240 - 0xf0
      12'hCCB: dout <= 8'b01101110; // 3275 : 110 - 0x6e
      12'hCCC: dout <= 8'b00011111; // 3276 :  31 - 0x1f
      12'hCCD: dout <= 8'b00011111; // 3277 :  31 - 0x1f
      12'hCCE: dout <= 8'b00011111; // 3278 :  31 - 0x1f
      12'hCCF: dout <= 8'b00001110; // 3279 :  14 - 0xe
      12'hCD0: dout <= 8'b01000000; // 3280 :  64 - 0x40 -- Background 0x9a
      12'hCD1: dout <= 8'b00001100; // 3281 :  12 - 0xc
      12'hCD2: dout <= 8'b00000000; // 3282 :   0 - 0x0
      12'hCD3: dout <= 8'b00101000; // 3283 :  40 - 0x28
      12'hCD4: dout <= 8'b00101100; // 3284 :  44 - 0x2c
      12'hCD5: dout <= 8'b00010001; // 3285 :  17 - 0x11
      12'hCD6: dout <= 8'b01000000; // 3286 :  64 - 0x40
      12'hCD7: dout <= 8'b00001000; // 3287 :   8 - 0x8
      12'hCD8: dout <= 8'b00100000; // 3288 :  32 - 0x20 -- Background 0x9b
      12'hCD9: dout <= 8'b00000000; // 3289 :   0 - 0x0
      12'hCDA: dout <= 8'b10010100; // 3290 : 148 - 0x94
      12'hCDB: dout <= 8'b01001000; // 3291 :  72 - 0x48
      12'hCDC: dout <= 8'b00011000; // 3292 :  24 - 0x18
      12'hCDD: dout <= 8'b00000110; // 3293 :   6 - 0x6
      12'hCDE: dout <= 8'b01000000; // 3294 :  64 - 0x40
      12'hCDF: dout <= 8'b00000000; // 3295 :   0 - 0x0
      12'hCE0: dout <= 8'b01111111; // 3296 : 127 - 0x7f -- Background 0x9c
      12'hCE1: dout <= 8'b01111111; // 3297 : 127 - 0x7f
      12'hCE2: dout <= 8'b01111111; // 3298 : 127 - 0x7f
      12'hCE3: dout <= 8'b00111111; // 3299 :  63 - 0x3f
      12'hCE4: dout <= 8'b00110101; // 3300 :  53 - 0x35
      12'hCE5: dout <= 8'b00000010; // 3301 :   2 - 0x2
      12'hCE6: dout <= 8'b00000000; // 3302 :   0 - 0x0
      12'hCE7: dout <= 8'b00000000; // 3303 :   0 - 0x0
      12'hCE8: dout <= 8'b11110100; // 3304 : 244 - 0xf4 -- Background 0x9d
      12'hCE9: dout <= 8'b11111000; // 3305 : 248 - 0xf8
      12'hCEA: dout <= 8'b11110000; // 3306 : 240 - 0xf0
      12'hCEB: dout <= 8'b11101000; // 3307 : 232 - 0xe8
      12'hCEC: dout <= 8'b01010000; // 3308 :  80 - 0x50
      12'hCED: dout <= 8'b10000000; // 3309 : 128 - 0x80
      12'hCEE: dout <= 8'b00000000; // 3310 :   0 - 0x0
      12'hCEF: dout <= 8'b00000000; // 3311 :   0 - 0x0
      12'hCF0: dout <= 8'b11111110; // 3312 : 254 - 0xfe -- Background 0x9e
      12'hCF1: dout <= 8'b11111100; // 3313 : 252 - 0xfc
      12'hCF2: dout <= 8'b11111100; // 3314 : 252 - 0xfc
      12'hCF3: dout <= 8'b11111000; // 3315 : 248 - 0xf8
      12'hCF4: dout <= 8'b11111000; // 3316 : 248 - 0xf8
      12'hCF5: dout <= 8'b11111100; // 3317 : 252 - 0xfc
      12'hCF6: dout <= 8'b11111100; // 3318 : 252 - 0xfc
      12'hCF7: dout <= 8'b11111110; // 3319 : 254 - 0xfe
      12'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0 -- Background 0x9f
      12'hCF9: dout <= 8'b00000000; // 3321 :   0 - 0x0
      12'hCFA: dout <= 8'b01111110; // 3322 : 126 - 0x7e
      12'hCFB: dout <= 8'b01111110; // 3323 : 126 - 0x7e
      12'hCFC: dout <= 8'b01111110; // 3324 : 126 - 0x7e
      12'hCFD: dout <= 8'b01111110; // 3325 : 126 - 0x7e
      12'hCFE: dout <= 8'b01111110; // 3326 : 126 - 0x7e
      12'hCFF: dout <= 8'b01111110; // 3327 : 126 - 0x7e
      12'hD00: dout <= 8'b00010000; // 3328 :  16 - 0x10 -- Background 0xa0
      12'hD01: dout <= 8'b00111000; // 3329 :  56 - 0x38
      12'hD02: dout <= 8'b01111100; // 3330 : 124 - 0x7c
      12'hD03: dout <= 8'b11111000; // 3331 : 248 - 0xf8
      12'hD04: dout <= 8'b01110000; // 3332 : 112 - 0x70
      12'hD05: dout <= 8'b00100010; // 3333 :  34 - 0x22
      12'hD06: dout <= 8'b00000101; // 3334 :   5 - 0x5
      12'hD07: dout <= 8'b00000010; // 3335 :   2 - 0x2
      12'hD08: dout <= 8'b00010000; // 3336 :  16 - 0x10 -- Background 0xa1
      12'hD09: dout <= 8'b00111000; // 3337 :  56 - 0x38
      12'hD0A: dout <= 8'b01111100; // 3338 : 124 - 0x7c
      12'hD0B: dout <= 8'b11100000; // 3339 : 224 - 0xe0
      12'hD0C: dout <= 8'b01100000; // 3340 :  96 - 0x60
      12'hD0D: dout <= 8'b00100000; // 3341 :  32 - 0x20
      12'hD0E: dout <= 8'b00000000; // 3342 :   0 - 0x0
      12'hD0F: dout <= 8'b00000000; // 3343 :   0 - 0x0
      12'hD10: dout <= 8'b00010000; // 3344 :  16 - 0x10 -- Background 0xa2
      12'hD11: dout <= 8'b00111000; // 3345 :  56 - 0x38
      12'hD12: dout <= 8'b01111100; // 3346 : 124 - 0x7c
      12'hD13: dout <= 8'b00000000; // 3347 :   0 - 0x0
      12'hD14: dout <= 8'b00000000; // 3348 :   0 - 0x0
      12'hD15: dout <= 8'b00000000; // 3349 :   0 - 0x0
      12'hD16: dout <= 8'b00000000; // 3350 :   0 - 0x0
      12'hD17: dout <= 8'b00000000; // 3351 :   0 - 0x0
      12'hD18: dout <= 8'b00000000; // 3352 :   0 - 0x0 -- Background 0xa3
      12'hD19: dout <= 8'b00100000; // 3353 :  32 - 0x20
      12'hD1A: dout <= 8'b01100000; // 3354 :  96 - 0x60
      12'hD1B: dout <= 8'b11100000; // 3355 : 224 - 0xe0
      12'hD1C: dout <= 8'b01100000; // 3356 :  96 - 0x60
      12'hD1D: dout <= 8'b00100000; // 3357 :  32 - 0x20
      12'hD1E: dout <= 8'b00000000; // 3358 :   0 - 0x0
      12'hD1F: dout <= 8'b00000000; // 3359 :   0 - 0x0
      12'hD20: dout <= 8'b00000000; // 3360 :   0 - 0x0 -- Background 0xa4
      12'hD21: dout <= 8'b00100000; // 3361 :  32 - 0x20
      12'hD22: dout <= 8'b01100011; // 3362 :  99 - 0x63
      12'hD23: dout <= 8'b11100111; // 3363 : 231 - 0xe7
      12'hD24: dout <= 8'b01100000; // 3364 :  96 - 0x60
      12'hD25: dout <= 8'b00100010; // 3365 :  34 - 0x22
      12'hD26: dout <= 8'b00000101; // 3366 :   5 - 0x5
      12'hD27: dout <= 8'b00000010; // 3367 :   2 - 0x2
      12'hD28: dout <= 8'b00000000; // 3368 :   0 - 0x0 -- Background 0xa5
      12'hD29: dout <= 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout <= 8'b11111111; // 3370 : 255 - 0xff
      12'hD2B: dout <= 8'b11111111; // 3371 : 255 - 0xff
      12'hD2C: dout <= 8'b00000000; // 3372 :   0 - 0x0
      12'hD2D: dout <= 8'b00100010; // 3373 :  34 - 0x22
      12'hD2E: dout <= 8'b00000101; // 3374 :   5 - 0x5
      12'hD2F: dout <= 8'b00000010; // 3375 :   2 - 0x2
      12'hD30: dout <= 8'b00010000; // 3376 :  16 - 0x10 -- Background 0xa6
      12'hD31: dout <= 8'b00111000; // 3377 :  56 - 0x38
      12'hD32: dout <= 8'b01111100; // 3378 : 124 - 0x7c
      12'hD33: dout <= 8'b00000000; // 3379 :   0 - 0x0
      12'hD34: dout <= 8'b00000000; // 3380 :   0 - 0x0
      12'hD35: dout <= 8'b00010010; // 3381 :  18 - 0x12
      12'hD36: dout <= 8'b00110101; // 3382 :  53 - 0x35
      12'hD37: dout <= 8'b00110010; // 3383 :  50 - 0x32
      12'hD38: dout <= 8'b00110000; // 3384 :  48 - 0x30 -- Background 0xa7
      12'hD39: dout <= 8'b00110000; // 3385 :  48 - 0x30
      12'hD3A: dout <= 8'b00110100; // 3386 :  52 - 0x34
      12'hD3B: dout <= 8'b00110000; // 3387 :  48 - 0x30
      12'hD3C: dout <= 8'b00110000; // 3388 :  48 - 0x30
      12'hD3D: dout <= 8'b00110010; // 3389 :  50 - 0x32
      12'hD3E: dout <= 8'b00110101; // 3390 :  53 - 0x35
      12'hD3F: dout <= 8'b00110010; // 3391 :  50 - 0x32
      12'hD40: dout <= 8'b00110000; // 3392 :  48 - 0x30 -- Background 0xa8
      12'hD41: dout <= 8'b00110000; // 3393 :  48 - 0x30
      12'hD42: dout <= 8'b11110100; // 3394 : 244 - 0xf4
      12'hD43: dout <= 8'b11110000; // 3395 : 240 - 0xf0
      12'hD44: dout <= 8'b00000000; // 3396 :   0 - 0x0
      12'hD45: dout <= 8'b00100010; // 3397 :  34 - 0x22
      12'hD46: dout <= 8'b00000101; // 3398 :   5 - 0x5
      12'hD47: dout <= 8'b00000010; // 3399 :   2 - 0x2
      12'hD48: dout <= 8'b00000000; // 3400 :   0 - 0x0 -- Background 0xa9
      12'hD49: dout <= 8'b00000000; // 3401 :   0 - 0x0
      12'hD4A: dout <= 8'b00000000; // 3402 :   0 - 0x0
      12'hD4B: dout <= 8'b00000000; // 3403 :   0 - 0x0
      12'hD4C: dout <= 8'b00000000; // 3404 :   0 - 0x0
      12'hD4D: dout <= 8'b00000000; // 3405 :   0 - 0x0
      12'hD4E: dout <= 8'b00000000; // 3406 :   0 - 0x0
      12'hD4F: dout <= 8'b00000000; // 3407 :   0 - 0x0
      12'hD50: dout <= 8'b00000000; // 3408 :   0 - 0x0 -- Background 0xaa
      12'hD51: dout <= 8'b00000000; // 3409 :   0 - 0x0
      12'hD52: dout <= 8'b01010000; // 3410 :  80 - 0x50
      12'hD53: dout <= 8'b10101000; // 3411 : 168 - 0xa8
      12'hD54: dout <= 8'b01110000; // 3412 : 112 - 0x70
      12'hD55: dout <= 8'b00100010; // 3413 :  34 - 0x22
      12'hD56: dout <= 8'b00000101; // 3414 :   5 - 0x5
      12'hD57: dout <= 8'b00000010; // 3415 :   2 - 0x2
      12'hD58: dout <= 8'b00000000; // 3416 :   0 - 0x0 -- Background 0xab
      12'hD59: dout <= 8'b00000000; // 3417 :   0 - 0x0
      12'hD5A: dout <= 8'b00000000; // 3418 :   0 - 0x0
      12'hD5B: dout <= 8'b00000000; // 3419 :   0 - 0x0
      12'hD5C: dout <= 8'b00000000; // 3420 :   0 - 0x0
      12'hD5D: dout <= 8'b00000000; // 3421 :   0 - 0x0
      12'hD5E: dout <= 8'b00000000; // 3422 :   0 - 0x0
      12'hD5F: dout <= 8'b00000000; // 3423 :   0 - 0x0
      12'hD60: dout <= 8'b00000000; // 3424 :   0 - 0x0 -- Background 0xac
      12'hD61: dout <= 8'b00000000; // 3425 :   0 - 0x0
      12'hD62: dout <= 8'b00000000; // 3426 :   0 - 0x0
      12'hD63: dout <= 8'b00000000; // 3427 :   0 - 0x0
      12'hD64: dout <= 8'b00000000; // 3428 :   0 - 0x0
      12'hD65: dout <= 8'b00000000; // 3429 :   0 - 0x0
      12'hD66: dout <= 8'b00000000; // 3430 :   0 - 0x0
      12'hD67: dout <= 8'b00000000; // 3431 :   0 - 0x0
      12'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0 -- Background 0xad
      12'hD69: dout <= 8'b00000000; // 3433 :   0 - 0x0
      12'hD6A: dout <= 8'b11111111; // 3434 : 255 - 0xff
      12'hD6B: dout <= 8'b00000000; // 3435 :   0 - 0x0
      12'hD6C: dout <= 8'b00000000; // 3436 :   0 - 0x0
      12'hD6D: dout <= 8'b00000000; // 3437 :   0 - 0x0
      12'hD6E: dout <= 8'b00000000; // 3438 :   0 - 0x0
      12'hD6F: dout <= 8'b00000000; // 3439 :   0 - 0x0
      12'hD70: dout <= 8'b00000000; // 3440 :   0 - 0x0 -- Background 0xae
      12'hD71: dout <= 8'b00000000; // 3441 :   0 - 0x0
      12'hD72: dout <= 8'b00000000; // 3442 :   0 - 0x0
      12'hD73: dout <= 8'b00000000; // 3443 :   0 - 0x0
      12'hD74: dout <= 8'b00000000; // 3444 :   0 - 0x0
      12'hD75: dout <= 8'b11111111; // 3445 : 255 - 0xff
      12'hD76: dout <= 8'b00000000; // 3446 :   0 - 0x0
      12'hD77: dout <= 8'b00000000; // 3447 :   0 - 0x0
      12'hD78: dout <= 8'b00000000; // 3448 :   0 - 0x0 -- Background 0xaf
      12'hD79: dout <= 8'b00000000; // 3449 :   0 - 0x0
      12'hD7A: dout <= 8'b00000000; // 3450 :   0 - 0x0
      12'hD7B: dout <= 8'b00000000; // 3451 :   0 - 0x0
      12'hD7C: dout <= 8'b00000000; // 3452 :   0 - 0x0
      12'hD7D: dout <= 8'b00000000; // 3453 :   0 - 0x0
      12'hD7E: dout <= 8'b00000000; // 3454 :   0 - 0x0
      12'hD7F: dout <= 8'b00000000; // 3455 :   0 - 0x0
      12'hD80: dout <= 8'b00000000; // 3456 :   0 - 0x0 -- Background 0xb0
      12'hD81: dout <= 8'b00000000; // 3457 :   0 - 0x0
      12'hD82: dout <= 8'b00011111; // 3458 :  31 - 0x1f
      12'hD83: dout <= 8'b00011111; // 3459 :  31 - 0x1f
      12'hD84: dout <= 8'b00011111; // 3460 :  31 - 0x1f
      12'hD85: dout <= 8'b00011111; // 3461 :  31 - 0x1f
      12'hD86: dout <= 8'b00011111; // 3462 :  31 - 0x1f
      12'hD87: dout <= 8'b00011111; // 3463 :  31 - 0x1f
      12'hD88: dout <= 8'b00000000; // 3464 :   0 - 0x0 -- Background 0xb1
      12'hD89: dout <= 8'b00000000; // 3465 :   0 - 0x0
      12'hD8A: dout <= 8'b11110000; // 3466 : 240 - 0xf0
      12'hD8B: dout <= 8'b11110000; // 3467 : 240 - 0xf0
      12'hD8C: dout <= 8'b11110000; // 3468 : 240 - 0xf0
      12'hD8D: dout <= 8'b11110000; // 3469 : 240 - 0xf0
      12'hD8E: dout <= 8'b11110000; // 3470 : 240 - 0xf0
      12'hD8F: dout <= 8'b11110000; // 3471 : 240 - 0xf0
      12'hD90: dout <= 8'b00011111; // 3472 :  31 - 0x1f -- Background 0xb2
      12'hD91: dout <= 8'b00011111; // 3473 :  31 - 0x1f
      12'hD92: dout <= 8'b00011111; // 3474 :  31 - 0x1f
      12'hD93: dout <= 8'b00011111; // 3475 :  31 - 0x1f
      12'hD94: dout <= 8'b00011111; // 3476 :  31 - 0x1f
      12'hD95: dout <= 8'b00000000; // 3477 :   0 - 0x0
      12'hD96: dout <= 8'b00000000; // 3478 :   0 - 0x0
      12'hD97: dout <= 8'b00000000; // 3479 :   0 - 0x0
      12'hD98: dout <= 8'b11110000; // 3480 : 240 - 0xf0 -- Background 0xb3
      12'hD99: dout <= 8'b11110000; // 3481 : 240 - 0xf0
      12'hD9A: dout <= 8'b11110000; // 3482 : 240 - 0xf0
      12'hD9B: dout <= 8'b11110000; // 3483 : 240 - 0xf0
      12'hD9C: dout <= 8'b11110000; // 3484 : 240 - 0xf0
      12'hD9D: dout <= 8'b00000000; // 3485 :   0 - 0x0
      12'hD9E: dout <= 8'b00000000; // 3486 :   0 - 0x0
      12'hD9F: dout <= 8'b00000000; // 3487 :   0 - 0x0
      12'hDA0: dout <= 8'b00000000; // 3488 :   0 - 0x0 -- Background 0xb4
      12'hDA1: dout <= 8'b00000000; // 3489 :   0 - 0x0
      12'hDA2: dout <= 8'b00000000; // 3490 :   0 - 0x0
      12'hDA3: dout <= 8'b00111111; // 3491 :  63 - 0x3f
      12'hDA4: dout <= 8'b01111111; // 3492 : 127 - 0x7f
      12'hDA5: dout <= 8'b01111111; // 3493 : 127 - 0x7f
      12'hDA6: dout <= 8'b01111111; // 3494 : 127 - 0x7f
      12'hDA7: dout <= 8'b01111111; // 3495 : 127 - 0x7f
      12'hDA8: dout <= 8'b00000000; // 3496 :   0 - 0x0 -- Background 0xb5
      12'hDA9: dout <= 8'b00000000; // 3497 :   0 - 0x0
      12'hDAA: dout <= 8'b00000000; // 3498 :   0 - 0x0
      12'hDAB: dout <= 8'b11111000; // 3499 : 248 - 0xf8
      12'hDAC: dout <= 8'b11111000; // 3500 : 248 - 0xf8
      12'hDAD: dout <= 8'b11111000; // 3501 : 248 - 0xf8
      12'hDAE: dout <= 8'b11111000; // 3502 : 248 - 0xf8
      12'hDAF: dout <= 8'b11111000; // 3503 : 248 - 0xf8
      12'hDB0: dout <= 8'b01111111; // 3504 : 127 - 0x7f -- Background 0xb6
      12'hDB1: dout <= 8'b01111111; // 3505 : 127 - 0x7f
      12'hDB2: dout <= 8'b01111111; // 3506 : 127 - 0x7f
      12'hDB3: dout <= 8'b01111111; // 3507 : 127 - 0x7f
      12'hDB4: dout <= 8'b01000000; // 3508 :  64 - 0x40
      12'hDB5: dout <= 8'b00000000; // 3509 :   0 - 0x0
      12'hDB6: dout <= 8'b00000000; // 3510 :   0 - 0x0
      12'hDB7: dout <= 8'b00000000; // 3511 :   0 - 0x0
      12'hDB8: dout <= 8'b11111000; // 3512 : 248 - 0xf8 -- Background 0xb7
      12'hDB9: dout <= 8'b11111000; // 3513 : 248 - 0xf8
      12'hDBA: dout <= 8'b11111000; // 3514 : 248 - 0xf8
      12'hDBB: dout <= 8'b11111000; // 3515 : 248 - 0xf8
      12'hDBC: dout <= 8'b00000000; // 3516 :   0 - 0x0
      12'hDBD: dout <= 8'b00000000; // 3517 :   0 - 0x0
      12'hDBE: dout <= 8'b00000000; // 3518 :   0 - 0x0
      12'hDBF: dout <= 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout <= 8'b00000000; // 3520 :   0 - 0x0 -- Background 0xb8
      12'hDC1: dout <= 8'b00000000; // 3521 :   0 - 0x0
      12'hDC2: dout <= 8'b00000011; // 3522 :   3 - 0x3
      12'hDC3: dout <= 8'b00000111; // 3523 :   7 - 0x7
      12'hDC4: dout <= 8'b00000111; // 3524 :   7 - 0x7
      12'hDC5: dout <= 8'b00000111; // 3525 :   7 - 0x7
      12'hDC6: dout <= 8'b00000011; // 3526 :   3 - 0x3
      12'hDC7: dout <= 8'b00000000; // 3527 :   0 - 0x0
      12'hDC8: dout <= 8'b00000000; // 3528 :   0 - 0x0 -- Background 0xb9
      12'hDC9: dout <= 8'b00000000; // 3529 :   0 - 0x0
      12'hDCA: dout <= 8'b11000001; // 3530 : 193 - 0xc1
      12'hDCB: dout <= 8'b11100010; // 3531 : 226 - 0xe2
      12'hDCC: dout <= 8'b11001100; // 3532 : 204 - 0xcc
      12'hDCD: dout <= 8'b11000000; // 3533 : 192 - 0xc0
      12'hDCE: dout <= 8'b10000000; // 3534 : 128 - 0x80
      12'hDCF: dout <= 8'b00000001; // 3535 :   1 - 0x1
      12'hDD0: dout <= 8'b00000000; // 3536 :   0 - 0x0 -- Background 0xba
      12'hDD1: dout <= 8'b11110000; // 3537 : 240 - 0xf0
      12'hDD2: dout <= 8'b00000000; // 3538 :   0 - 0x0
      12'hDD3: dout <= 8'b00100000; // 3539 :  32 - 0x20
      12'hDD4: dout <= 8'b00100000; // 3540 :  32 - 0x20
      12'hDD5: dout <= 8'b00000000; // 3541 :   0 - 0x0
      12'hDD6: dout <= 8'b11110000; // 3542 : 240 - 0xf0
      12'hDD7: dout <= 8'b00000000; // 3543 :   0 - 0x0
      12'hDD8: dout <= 8'b00000000; // 3544 :   0 - 0x0 -- Background 0xbb
      12'hDD9: dout <= 8'b00000000; // 3545 :   0 - 0x0
      12'hDDA: dout <= 8'b00000000; // 3546 :   0 - 0x0
      12'hDDB: dout <= 8'b00000000; // 3547 :   0 - 0x0
      12'hDDC: dout <= 8'b00000000; // 3548 :   0 - 0x0
      12'hDDD: dout <= 8'b01100000; // 3549 :  96 - 0x60
      12'hDDE: dout <= 8'b01100000; // 3550 :  96 - 0x60
      12'hDDF: dout <= 8'b00000000; // 3551 :   0 - 0x0
      12'hDE0: dout <= 8'b00000010; // 3552 :   2 - 0x2 -- Background 0xbc
      12'hDE1: dout <= 8'b00001100; // 3553 :  12 - 0xc
      12'hDE2: dout <= 8'b00000000; // 3554 :   0 - 0x0
      12'hDE3: dout <= 8'b00000000; // 3555 :   0 - 0x0
      12'hDE4: dout <= 8'b00000000; // 3556 :   0 - 0x0
      12'hDE5: dout <= 8'b00000110; // 3557 :   6 - 0x6
      12'hDE6: dout <= 8'b00000110; // 3558 :   6 - 0x6
      12'hDE7: dout <= 8'b00000000; // 3559 :   0 - 0x0
      12'hDE8: dout <= 8'b00000000; // 3560 :   0 - 0x0 -- Background 0xbd
      12'hDE9: dout <= 8'b10000000; // 3561 : 128 - 0x80
      12'hDEA: dout <= 8'b00000011; // 3562 :   3 - 0x3
      12'hDEB: dout <= 8'b00000111; // 3563 :   7 - 0x7
      12'hDEC: dout <= 8'b00000111; // 3564 :   7 - 0x7
      12'hDED: dout <= 8'b00000111; // 3565 :   7 - 0x7
      12'hDEE: dout <= 8'b00000011; // 3566 :   3 - 0x3
      12'hDEF: dout <= 8'b00000000; // 3567 :   0 - 0x0
      12'hDF0: dout <= 8'b00000000; // 3568 :   0 - 0x0 -- Background 0xbe
      12'hDF1: dout <= 8'b00000100; // 3569 :   4 - 0x4
      12'hDF2: dout <= 8'b11000000; // 3570 : 192 - 0xc0
      12'hDF3: dout <= 8'b11100000; // 3571 : 224 - 0xe0
      12'hDF4: dout <= 8'b11000000; // 3572 : 192 - 0xc0
      12'hDF5: dout <= 8'b11000000; // 3573 : 192 - 0xc0
      12'hDF6: dout <= 8'b10000000; // 3574 : 128 - 0x80
      12'hDF7: dout <= 8'b00000000; // 3575 :   0 - 0x0
      12'hDF8: dout <= 8'b00000000; // 3576 :   0 - 0x0 -- Background 0xbf
      12'hDF9: dout <= 8'b00000000; // 3577 :   0 - 0x0
      12'hDFA: dout <= 8'b00000000; // 3578 :   0 - 0x0
      12'hDFB: dout <= 8'b00000000; // 3579 :   0 - 0x0
      12'hDFC: dout <= 8'b00000000; // 3580 :   0 - 0x0
      12'hDFD: dout <= 8'b10001000; // 3581 : 136 - 0x88
      12'hDFE: dout <= 8'b00001000; // 3582 :   8 - 0x8
      12'hDFF: dout <= 8'b00001011; // 3583 :  11 - 0xb
      12'hE00: dout <= 8'b00000000; // 3584 :   0 - 0x0 -- Background 0xc0
      12'hE01: dout <= 8'b00000000; // 3585 :   0 - 0x0
      12'hE02: dout <= 8'b00000000; // 3586 :   0 - 0x0
      12'hE03: dout <= 8'b00000000; // 3587 :   0 - 0x0
      12'hE04: dout <= 8'b00000000; // 3588 :   0 - 0x0
      12'hE05: dout <= 8'b00100100; // 3589 :  36 - 0x24
      12'hE06: dout <= 8'b00100000; // 3590 :  32 - 0x20
      12'hE07: dout <= 8'b10100000; // 3591 : 160 - 0xa0
      12'hE08: dout <= 8'b00000000; // 3592 :   0 - 0x0 -- Background 0xc1
      12'hE09: dout <= 8'b00000000; // 3593 :   0 - 0x0
      12'hE0A: dout <= 8'b00000000; // 3594 :   0 - 0x0
      12'hE0B: dout <= 8'b00000000; // 3595 :   0 - 0x0
      12'hE0C: dout <= 8'b00000000; // 3596 :   0 - 0x0
      12'hE0D: dout <= 8'b00000000; // 3597 :   0 - 0x0
      12'hE0E: dout <= 8'b00000000; // 3598 :   0 - 0x0
      12'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout <= 8'b00000000; // 3600 :   0 - 0x0 -- Background 0xc2
      12'hE11: dout <= 8'b00000000; // 3601 :   0 - 0x0
      12'hE12: dout <= 8'b00000000; // 3602 :   0 - 0x0
      12'hE13: dout <= 8'b00000000; // 3603 :   0 - 0x0
      12'hE14: dout <= 8'b00000000; // 3604 :   0 - 0x0
      12'hE15: dout <= 8'b00000000; // 3605 :   0 - 0x0
      12'hE16: dout <= 8'b00000000; // 3606 :   0 - 0x0
      12'hE17: dout <= 8'b00000000; // 3607 :   0 - 0x0
      12'hE18: dout <= 8'b00000000; // 3608 :   0 - 0x0 -- Background 0xc3
      12'hE19: dout <= 8'b00000000; // 3609 :   0 - 0x0
      12'hE1A: dout <= 8'b00000000; // 3610 :   0 - 0x0
      12'hE1B: dout <= 8'b00001000; // 3611 :   8 - 0x8
      12'hE1C: dout <= 8'b00001011; // 3612 :  11 - 0xb
      12'hE1D: dout <= 8'b00001000; // 3613 :   8 - 0x8
      12'hE1E: dout <= 8'b00001000; // 3614 :   8 - 0x8
      12'hE1F: dout <= 8'b00001000; // 3615 :   8 - 0x8
      12'hE20: dout <= 8'b00000000; // 3616 :   0 - 0x0 -- Background 0xc4
      12'hE21: dout <= 8'b00000000; // 3617 :   0 - 0x0
      12'hE22: dout <= 8'b00000000; // 3618 :   0 - 0x0
      12'hE23: dout <= 8'b00100000; // 3619 :  32 - 0x20
      12'hE24: dout <= 8'b10100000; // 3620 : 160 - 0xa0
      12'hE25: dout <= 8'b00100000; // 3621 :  32 - 0x20
      12'hE26: dout <= 8'b00100000; // 3622 :  32 - 0x20
      12'hE27: dout <= 8'b00100000; // 3623 :  32 - 0x20
      12'hE28: dout <= 8'b00001000; // 3624 :   8 - 0x8 -- Background 0xc5
      12'hE29: dout <= 8'b11001000; // 3625 : 200 - 0xc8
      12'hE2A: dout <= 8'b00001000; // 3626 :   8 - 0x8
      12'hE2B: dout <= 8'b00000011; // 3627 :   3 - 0x3
      12'hE2C: dout <= 8'b00000111; // 3628 :   7 - 0x7
      12'hE2D: dout <= 8'b00000111; // 3629 :   7 - 0x7
      12'hE2E: dout <= 8'b00000111; // 3630 :   7 - 0x7
      12'hE2F: dout <= 8'b00000011; // 3631 :   3 - 0x3
      12'hE30: dout <= 8'b00100000; // 3632 :  32 - 0x20 -- Background 0xc6
      12'hE31: dout <= 8'b00100110; // 3633 :  38 - 0x26
      12'hE32: dout <= 8'b00100000; // 3634 :  32 - 0x20
      12'hE33: dout <= 8'b11000000; // 3635 : 192 - 0xc0
      12'hE34: dout <= 8'b11100000; // 3636 : 224 - 0xe0
      12'hE35: dout <= 8'b11000000; // 3637 : 192 - 0xc0
      12'hE36: dout <= 8'b11000000; // 3638 : 192 - 0xc0
      12'hE37: dout <= 8'b10000000; // 3639 : 128 - 0x80
      12'hE38: dout <= 8'b00000000; // 3640 :   0 - 0x0 -- Background 0xc7
      12'hE39: dout <= 8'b00000000; // 3641 :   0 - 0x0
      12'hE3A: dout <= 8'b00000000; // 3642 :   0 - 0x0
      12'hE3B: dout <= 8'b00000000; // 3643 :   0 - 0x0
      12'hE3C: dout <= 8'b00000000; // 3644 :   0 - 0x0
      12'hE3D: dout <= 8'b11000000; // 3645 : 192 - 0xc0
      12'hE3E: dout <= 8'b00000000; // 3646 :   0 - 0x0
      12'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout <= 8'b00000000; // 3648 :   0 - 0x0 -- Background 0xc8
      12'hE41: dout <= 8'b00000000; // 3649 :   0 - 0x0
      12'hE42: dout <= 8'b00000000; // 3650 :   0 - 0x0
      12'hE43: dout <= 8'b00000000; // 3651 :   0 - 0x0
      12'hE44: dout <= 8'b00000000; // 3652 :   0 - 0x0
      12'hE45: dout <= 8'b00000110; // 3653 :   6 - 0x6
      12'hE46: dout <= 8'b00000000; // 3654 :   0 - 0x0
      12'hE47: dout <= 8'b00000000; // 3655 :   0 - 0x0
      12'hE48: dout <= 8'b00000000; // 3656 :   0 - 0x0 -- Background 0xc9
      12'hE49: dout <= 8'b00001111; // 3657 :  15 - 0xf
      12'hE4A: dout <= 8'b00000000; // 3658 :   0 - 0x0
      12'hE4B: dout <= 8'b00001000; // 3659 :   8 - 0x8
      12'hE4C: dout <= 8'b00001000; // 3660 :   8 - 0x8
      12'hE4D: dout <= 8'b00000000; // 3661 :   0 - 0x0
      12'hE4E: dout <= 8'b00001111; // 3662 :  15 - 0xf
      12'hE4F: dout <= 8'b00000000; // 3663 :   0 - 0x0
      12'hE50: dout <= 8'b00000000; // 3664 :   0 - 0x0 -- Background 0xca
      12'hE51: dout <= 8'b00000000; // 3665 :   0 - 0x0
      12'hE52: dout <= 8'b10000011; // 3666 : 131 - 0x83
      12'hE53: dout <= 8'b01000111; // 3667 :  71 - 0x47
      12'hE54: dout <= 8'b00110111; // 3668 :  55 - 0x37
      12'hE55: dout <= 8'b00000111; // 3669 :   7 - 0x7
      12'hE56: dout <= 8'b00000011; // 3670 :   3 - 0x3
      12'hE57: dout <= 8'b10000000; // 3671 : 128 - 0x80
      12'hE58: dout <= 8'b00000000; // 3672 :   0 - 0x0 -- Background 0xcb
      12'hE59: dout <= 8'b00000000; // 3673 :   0 - 0x0
      12'hE5A: dout <= 8'b11000000; // 3674 : 192 - 0xc0
      12'hE5B: dout <= 8'b11100000; // 3675 : 224 - 0xe0
      12'hE5C: dout <= 8'b11000000; // 3676 : 192 - 0xc0
      12'hE5D: dout <= 8'b11000000; // 3677 : 192 - 0xc0
      12'hE5E: dout <= 8'b10000000; // 3678 : 128 - 0x80
      12'hE5F: dout <= 8'b00000000; // 3679 :   0 - 0x0
      12'hE60: dout <= 8'b01000000; // 3680 :  64 - 0x40 -- Background 0xcc
      12'hE61: dout <= 8'b00110000; // 3681 :  48 - 0x30
      12'hE62: dout <= 8'b00000000; // 3682 :   0 - 0x0
      12'hE63: dout <= 8'b00000000; // 3683 :   0 - 0x0
      12'hE64: dout <= 8'b00000000; // 3684 :   0 - 0x0
      12'hE65: dout <= 8'b01100000; // 3685 :  96 - 0x60
      12'hE66: dout <= 8'b01100000; // 3686 :  96 - 0x60
      12'hE67: dout <= 8'b00000000; // 3687 :   0 - 0x0
      12'hE68: dout <= 8'b00000000; // 3688 :   0 - 0x0 -- Background 0xcd
      12'hE69: dout <= 8'b00000000; // 3689 :   0 - 0x0
      12'hE6A: dout <= 8'b00000000; // 3690 :   0 - 0x0
      12'hE6B: dout <= 8'b00000000; // 3691 :   0 - 0x0
      12'hE6C: dout <= 8'b00000000; // 3692 :   0 - 0x0
      12'hE6D: dout <= 8'b00000110; // 3693 :   6 - 0x6
      12'hE6E: dout <= 8'b00000110; // 3694 :   6 - 0x6
      12'hE6F: dout <= 8'b00000000; // 3695 :   0 - 0x0
      12'hE70: dout <= 8'b00000000; // 3696 :   0 - 0x0 -- Background 0xce
      12'hE71: dout <= 8'b00000001; // 3697 :   1 - 0x1
      12'hE72: dout <= 8'b00011011; // 3698 :  27 - 0x1b
      12'hE73: dout <= 8'b00010011; // 3699 :  19 - 0x13
      12'hE74: dout <= 8'b00011111; // 3700 :  31 - 0x1f
      12'hE75: dout <= 8'b00111111; // 3701 :  63 - 0x3f
      12'hE76: dout <= 8'b00111111; // 3702 :  63 - 0x3f
      12'hE77: dout <= 8'b00111111; // 3703 :  63 - 0x3f
      12'hE78: dout <= 8'b00000000; // 3704 :   0 - 0x0 -- Background 0xcf
      12'hE79: dout <= 8'b11111000; // 3705 : 248 - 0xf8
      12'hE7A: dout <= 8'b00001000; // 3706 :   8 - 0x8
      12'hE7B: dout <= 8'b00001000; // 3707 :   8 - 0x8
      12'hE7C: dout <= 8'b00001000; // 3708 :   8 - 0x8
      12'hE7D: dout <= 8'b11111000; // 3709 : 248 - 0xf8
      12'hE7E: dout <= 8'b11110000; // 3710 : 240 - 0xf0
      12'hE7F: dout <= 8'b11010000; // 3711 : 208 - 0xd0
      12'hE80: dout <= 8'b00000000; // 3712 :   0 - 0x0 -- Background 0xd0
      12'hE81: dout <= 8'b00000000; // 3713 :   0 - 0x0
      12'hE82: dout <= 8'b01111100; // 3714 : 124 - 0x7c
      12'hE83: dout <= 8'b11111110; // 3715 : 254 - 0xfe
      12'hE84: dout <= 8'b11101110; // 3716 : 238 - 0xee
      12'hE85: dout <= 8'b11101110; // 3717 : 238 - 0xee
      12'hE86: dout <= 8'b11101110; // 3718 : 238 - 0xee
      12'hE87: dout <= 8'b11101110; // 3719 : 238 - 0xee
      12'hE88: dout <= 8'b00000000; // 3720 :   0 - 0x0 -- Background 0xd1
      12'hE89: dout <= 8'b00000000; // 3721 :   0 - 0x0
      12'hE8A: dout <= 8'b00111000; // 3722 :  56 - 0x38
      12'hE8B: dout <= 8'b01111000; // 3723 : 120 - 0x78
      12'hE8C: dout <= 8'b01111000; // 3724 : 120 - 0x78
      12'hE8D: dout <= 8'b00111000; // 3725 :  56 - 0x38
      12'hE8E: dout <= 8'b00111000; // 3726 :  56 - 0x38
      12'hE8F: dout <= 8'b00111000; // 3727 :  56 - 0x38
      12'hE90: dout <= 8'b00000000; // 3728 :   0 - 0x0 -- Background 0xd2
      12'hE91: dout <= 8'b00000000; // 3729 :   0 - 0x0
      12'hE92: dout <= 8'b01111100; // 3730 : 124 - 0x7c
      12'hE93: dout <= 8'b11111110; // 3731 : 254 - 0xfe
      12'hE94: dout <= 8'b11101110; // 3732 : 238 - 0xee
      12'hE95: dout <= 8'b00001110; // 3733 :  14 - 0xe
      12'hE96: dout <= 8'b00001110; // 3734 :  14 - 0xe
      12'hE97: dout <= 8'b01111110; // 3735 : 126 - 0x7e
      12'hE98: dout <= 8'b00000000; // 3736 :   0 - 0x0 -- Background 0xd3
      12'hE99: dout <= 8'b00000000; // 3737 :   0 - 0x0
      12'hE9A: dout <= 8'b01111100; // 3738 : 124 - 0x7c
      12'hE9B: dout <= 8'b11111110; // 3739 : 254 - 0xfe
      12'hE9C: dout <= 8'b11101110; // 3740 : 238 - 0xee
      12'hE9D: dout <= 8'b00001110; // 3741 :  14 - 0xe
      12'hE9E: dout <= 8'b00111100; // 3742 :  60 - 0x3c
      12'hE9F: dout <= 8'b00111100; // 3743 :  60 - 0x3c
      12'hEA0: dout <= 8'b00000000; // 3744 :   0 - 0x0 -- Background 0xd4
      12'hEA1: dout <= 8'b00000000; // 3745 :   0 - 0x0
      12'hEA2: dout <= 8'b00111110; // 3746 :  62 - 0x3e
      12'hEA3: dout <= 8'b01111110; // 3747 : 126 - 0x7e
      12'hEA4: dout <= 8'b11101110; // 3748 : 238 - 0xee
      12'hEA5: dout <= 8'b11101110; // 3749 : 238 - 0xee
      12'hEA6: dout <= 8'b11101110; // 3750 : 238 - 0xee
      12'hEA7: dout <= 8'b11101110; // 3751 : 238 - 0xee
      12'hEA8: dout <= 8'b00000000; // 3752 :   0 - 0x0 -- Background 0xd5
      12'hEA9: dout <= 8'b00000000; // 3753 :   0 - 0x0
      12'hEAA: dout <= 8'b11111100; // 3754 : 252 - 0xfc
      12'hEAB: dout <= 8'b11111100; // 3755 : 252 - 0xfc
      12'hEAC: dout <= 8'b11100000; // 3756 : 224 - 0xe0
      12'hEAD: dout <= 8'b11100000; // 3757 : 224 - 0xe0
      12'hEAE: dout <= 8'b11111100; // 3758 : 252 - 0xfc
      12'hEAF: dout <= 8'b11111110; // 3759 : 254 - 0xfe
      12'hEB0: dout <= 8'b00000000; // 3760 :   0 - 0x0 -- Background 0xd6
      12'hEB1: dout <= 8'b00000000; // 3761 :   0 - 0x0
      12'hEB2: dout <= 8'b01111100; // 3762 : 124 - 0x7c
      12'hEB3: dout <= 8'b11111100; // 3763 : 252 - 0xfc
      12'hEB4: dout <= 8'b11100000; // 3764 : 224 - 0xe0
      12'hEB5: dout <= 8'b11100000; // 3765 : 224 - 0xe0
      12'hEB6: dout <= 8'b11111100; // 3766 : 252 - 0xfc
      12'hEB7: dout <= 8'b11111110; // 3767 : 254 - 0xfe
      12'hEB8: dout <= 8'b00000000; // 3768 :   0 - 0x0 -- Background 0xd7
      12'hEB9: dout <= 8'b00000000; // 3769 :   0 - 0x0
      12'hEBA: dout <= 8'b11111110; // 3770 : 254 - 0xfe
      12'hEBB: dout <= 8'b11111110; // 3771 : 254 - 0xfe
      12'hEBC: dout <= 8'b11101110; // 3772 : 238 - 0xee
      12'hEBD: dout <= 8'b00001110; // 3773 :  14 - 0xe
      12'hEBE: dout <= 8'b00001110; // 3774 :  14 - 0xe
      12'hEBF: dout <= 8'b00011100; // 3775 :  28 - 0x1c
      12'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Background 0xd8
      12'hEC1: dout <= 8'b00000000; // 3777 :   0 - 0x0
      12'hEC2: dout <= 8'b01111100; // 3778 : 124 - 0x7c
      12'hEC3: dout <= 8'b11111110; // 3779 : 254 - 0xfe
      12'hEC4: dout <= 8'b11101110; // 3780 : 238 - 0xee
      12'hEC5: dout <= 8'b11101110; // 3781 : 238 - 0xee
      12'hEC6: dout <= 8'b01111100; // 3782 : 124 - 0x7c
      12'hEC7: dout <= 8'b11111110; // 3783 : 254 - 0xfe
      12'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0 -- Background 0xd9
      12'hEC9: dout <= 8'b00000000; // 3785 :   0 - 0x0
      12'hECA: dout <= 8'b01111100; // 3786 : 124 - 0x7c
      12'hECB: dout <= 8'b11111110; // 3787 : 254 - 0xfe
      12'hECC: dout <= 8'b11101110; // 3788 : 238 - 0xee
      12'hECD: dout <= 8'b11101110; // 3789 : 238 - 0xee
      12'hECE: dout <= 8'b11101110; // 3790 : 238 - 0xee
      12'hECF: dout <= 8'b11101110; // 3791 : 238 - 0xee
      12'hED0: dout <= 8'b00000000; // 3792 :   0 - 0x0 -- Background 0xda
      12'hED1: dout <= 8'b00100000; // 3793 :  32 - 0x20
      12'hED2: dout <= 8'b00000000; // 3794 :   0 - 0x0
      12'hED3: dout <= 8'b00000010; // 3795 :   2 - 0x2
      12'hED4: dout <= 8'b00000000; // 3796 :   0 - 0x0
      12'hED5: dout <= 8'b00100000; // 3797 :  32 - 0x20
      12'hED6: dout <= 8'b00000000; // 3798 :   0 - 0x0
      12'hED7: dout <= 8'b00000000; // 3799 :   0 - 0x0
      12'hED8: dout <= 8'b00100000; // 3800 :  32 - 0x20 -- Background 0xdb
      12'hED9: dout <= 8'b00000000; // 3801 :   0 - 0x0
      12'hEDA: dout <= 8'b00000000; // 3802 :   0 - 0x0
      12'hEDB: dout <= 8'b00000000; // 3803 :   0 - 0x0
      12'hEDC: dout <= 8'b10000000; // 3804 : 128 - 0x80
      12'hEDD: dout <= 8'b00000000; // 3805 :   0 - 0x0
      12'hEDE: dout <= 8'b00000100; // 3806 :   4 - 0x4
      12'hEDF: dout <= 8'b00000000; // 3807 :   0 - 0x0
      12'hEE0: dout <= 8'b00000000; // 3808 :   0 - 0x0 -- Background 0xdc
      12'hEE1: dout <= 8'b00001000; // 3809 :   8 - 0x8
      12'hEE2: dout <= 8'b00000000; // 3810 :   0 - 0x0
      12'hEE3: dout <= 8'b00000000; // 3811 :   0 - 0x0
      12'hEE4: dout <= 8'b00000010; // 3812 :   2 - 0x2
      12'hEE5: dout <= 8'b00000000; // 3813 :   0 - 0x0
      12'hEE6: dout <= 8'b01000000; // 3814 :  64 - 0x40
      12'hEE7: dout <= 8'b00000000; // 3815 :   0 - 0x0
      12'hEE8: dout <= 8'b00000000; // 3816 :   0 - 0x0 -- Background 0xdd
      12'hEE9: dout <= 8'b01000000; // 3817 :  64 - 0x40
      12'hEEA: dout <= 8'b00000000; // 3818 :   0 - 0x0
      12'hEEB: dout <= 8'b00000000; // 3819 :   0 - 0x0
      12'hEEC: dout <= 8'b00000000; // 3820 :   0 - 0x0
      12'hEED: dout <= 8'b00000000; // 3821 :   0 - 0x0
      12'hEEE: dout <= 8'b00000010; // 3822 :   2 - 0x2
      12'hEEF: dout <= 8'b00100000; // 3823 :  32 - 0x20
      12'hEF0: dout <= 8'b00111110; // 3824 :  62 - 0x3e -- Background 0xde
      12'hEF1: dout <= 8'b00111111; // 3825 :  63 - 0x3f
      12'hEF2: dout <= 8'b00111110; // 3826 :  62 - 0x3e
      12'hEF3: dout <= 8'b00111100; // 3827 :  60 - 0x3c
      12'hEF4: dout <= 8'b00111111; // 3828 :  63 - 0x3f
      12'hEF5: dout <= 8'b00110000; // 3829 :  48 - 0x30
      12'hEF6: dout <= 8'b00000000; // 3830 :   0 - 0x0
      12'hEF7: dout <= 8'b00000000; // 3831 :   0 - 0x0
      12'hEF8: dout <= 8'b00010000; // 3832 :  16 - 0x10 -- Background 0xdf
      12'hEF9: dout <= 8'b10110000; // 3833 : 176 - 0xb0
      12'hEFA: dout <= 8'b00110000; // 3834 :  48 - 0x30
      12'hEFB: dout <= 8'b11110000; // 3835 : 240 - 0xf0
      12'hEFC: dout <= 8'b11110000; // 3836 : 240 - 0xf0
      12'hEFD: dout <= 8'b00000000; // 3837 :   0 - 0x0
      12'hEFE: dout <= 8'b00000000; // 3838 :   0 - 0x0
      12'hEFF: dout <= 8'b00000000; // 3839 :   0 - 0x0
      12'hF00: dout <= 8'b11101110; // 3840 : 238 - 0xee -- Background 0xe0
      12'hF01: dout <= 8'b11101110; // 3841 : 238 - 0xee
      12'hF02: dout <= 8'b11101110; // 3842 : 238 - 0xee
      12'hF03: dout <= 8'b11101110; // 3843 : 238 - 0xee
      12'hF04: dout <= 8'b11111110; // 3844 : 254 - 0xfe
      12'hF05: dout <= 8'b01111100; // 3845 : 124 - 0x7c
      12'hF06: dout <= 8'b00000000; // 3846 :   0 - 0x0
      12'hF07: dout <= 8'b00000000; // 3847 :   0 - 0x0
      12'hF08: dout <= 8'b00111000; // 3848 :  56 - 0x38 -- Background 0xe1
      12'hF09: dout <= 8'b00111000; // 3849 :  56 - 0x38
      12'hF0A: dout <= 8'b00111000; // 3850 :  56 - 0x38
      12'hF0B: dout <= 8'b00111000; // 3851 :  56 - 0x38
      12'hF0C: dout <= 8'b01111100; // 3852 : 124 - 0x7c
      12'hF0D: dout <= 8'b01111100; // 3853 : 124 - 0x7c
      12'hF0E: dout <= 8'b00000000; // 3854 :   0 - 0x0
      12'hF0F: dout <= 8'b00000000; // 3855 :   0 - 0x0
      12'hF10: dout <= 8'b11111100; // 3856 : 252 - 0xfc -- Background 0xe2
      12'hF11: dout <= 8'b11100000; // 3857 : 224 - 0xe0
      12'hF12: dout <= 8'b11100000; // 3858 : 224 - 0xe0
      12'hF13: dout <= 8'b11100000; // 3859 : 224 - 0xe0
      12'hF14: dout <= 8'b11111110; // 3860 : 254 - 0xfe
      12'hF15: dout <= 8'b11111110; // 3861 : 254 - 0xfe
      12'hF16: dout <= 8'b00000000; // 3862 :   0 - 0x0
      12'hF17: dout <= 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout <= 8'b00001110; // 3864 :  14 - 0xe -- Background 0xe3
      12'hF19: dout <= 8'b00001110; // 3865 :  14 - 0xe
      12'hF1A: dout <= 8'b00001110; // 3866 :  14 - 0xe
      12'hF1B: dout <= 8'b11101110; // 3867 : 238 - 0xee
      12'hF1C: dout <= 8'b11111110; // 3868 : 254 - 0xfe
      12'hF1D: dout <= 8'b01111100; // 3869 : 124 - 0x7c
      12'hF1E: dout <= 8'b00000000; // 3870 :   0 - 0x0
      12'hF1F: dout <= 8'b00000000; // 3871 :   0 - 0x0
      12'hF20: dout <= 8'b11101110; // 3872 : 238 - 0xee -- Background 0xe4
      12'hF21: dout <= 8'b11101110; // 3873 : 238 - 0xee
      12'hF22: dout <= 8'b11111110; // 3874 : 254 - 0xfe
      12'hF23: dout <= 8'b11111110; // 3875 : 254 - 0xfe
      12'hF24: dout <= 8'b00001110; // 3876 :  14 - 0xe
      12'hF25: dout <= 8'b00001110; // 3877 :  14 - 0xe
      12'hF26: dout <= 8'b00000000; // 3878 :   0 - 0x0
      12'hF27: dout <= 8'b00000000; // 3879 :   0 - 0x0
      12'hF28: dout <= 8'b00001110; // 3880 :  14 - 0xe -- Background 0xe5
      12'hF29: dout <= 8'b00001110; // 3881 :  14 - 0xe
      12'hF2A: dout <= 8'b00001110; // 3882 :  14 - 0xe
      12'hF2B: dout <= 8'b11101110; // 3883 : 238 - 0xee
      12'hF2C: dout <= 8'b11111110; // 3884 : 254 - 0xfe
      12'hF2D: dout <= 8'b01111100; // 3885 : 124 - 0x7c
      12'hF2E: dout <= 8'b00000000; // 3886 :   0 - 0x0
      12'hF2F: dout <= 8'b00000000; // 3887 :   0 - 0x0
      12'hF30: dout <= 8'b11101110; // 3888 : 238 - 0xee -- Background 0xe6
      12'hF31: dout <= 8'b11101110; // 3889 : 238 - 0xee
      12'hF32: dout <= 8'b11101110; // 3890 : 238 - 0xee
      12'hF33: dout <= 8'b11101110; // 3891 : 238 - 0xee
      12'hF34: dout <= 8'b11111110; // 3892 : 254 - 0xfe
      12'hF35: dout <= 8'b01111100; // 3893 : 124 - 0x7c
      12'hF36: dout <= 8'b00000000; // 3894 :   0 - 0x0
      12'hF37: dout <= 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout <= 8'b00011100; // 3896 :  28 - 0x1c -- Background 0xe7
      12'hF39: dout <= 8'b00011100; // 3897 :  28 - 0x1c
      12'hF3A: dout <= 8'b00111000; // 3898 :  56 - 0x38
      12'hF3B: dout <= 8'b00111000; // 3899 :  56 - 0x38
      12'hF3C: dout <= 8'b00111000; // 3900 :  56 - 0x38
      12'hF3D: dout <= 8'b00111000; // 3901 :  56 - 0x38
      12'hF3E: dout <= 8'b00000000; // 3902 :   0 - 0x0
      12'hF3F: dout <= 8'b00000000; // 3903 :   0 - 0x0
      12'hF40: dout <= 8'b11101110; // 3904 : 238 - 0xee -- Background 0xe8
      12'hF41: dout <= 8'b11101110; // 3905 : 238 - 0xee
      12'hF42: dout <= 8'b11101110; // 3906 : 238 - 0xee
      12'hF43: dout <= 8'b11101110; // 3907 : 238 - 0xee
      12'hF44: dout <= 8'b11111110; // 3908 : 254 - 0xfe
      12'hF45: dout <= 8'b01111100; // 3909 : 124 - 0x7c
      12'hF46: dout <= 8'b00000000; // 3910 :   0 - 0x0
      12'hF47: dout <= 8'b00000000; // 3911 :   0 - 0x0
      12'hF48: dout <= 8'b11111110; // 3912 : 254 - 0xfe -- Background 0xe9
      12'hF49: dout <= 8'b01111110; // 3913 : 126 - 0x7e
      12'hF4A: dout <= 8'b00001110; // 3914 :  14 - 0xe
      12'hF4B: dout <= 8'b00001110; // 3915 :  14 - 0xe
      12'hF4C: dout <= 8'b01111110; // 3916 : 126 - 0x7e
      12'hF4D: dout <= 8'b01111100; // 3917 : 124 - 0x7c
      12'hF4E: dout <= 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout <= 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout <= 8'b00000000; // 3920 :   0 - 0x0 -- Background 0xea
      12'hF51: dout <= 8'b01110000; // 3921 : 112 - 0x70
      12'hF52: dout <= 8'b00111000; // 3922 :  56 - 0x38
      12'hF53: dout <= 8'b00000000; // 3923 :   0 - 0x0
      12'hF54: dout <= 8'b00000010; // 3924 :   2 - 0x2
      12'hF55: dout <= 8'b00000111; // 3925 :   7 - 0x7
      12'hF56: dout <= 8'b00000011; // 3926 :   3 - 0x3
      12'hF57: dout <= 8'b00000000; // 3927 :   0 - 0x0
      12'hF58: dout <= 8'b00000000; // 3928 :   0 - 0x0 -- Background 0xeb
      12'hF59: dout <= 8'b00001100; // 3929 :  12 - 0xc
      12'hF5A: dout <= 8'b00000110; // 3930 :   6 - 0x6
      12'hF5B: dout <= 8'b00000110; // 3931 :   6 - 0x6
      12'hF5C: dout <= 8'b01100000; // 3932 :  96 - 0x60
      12'hF5D: dout <= 8'b01110000; // 3933 : 112 - 0x70
      12'hF5E: dout <= 8'b00110000; // 3934 :  48 - 0x30
      12'hF5F: dout <= 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Background 0xec
      12'hF61: dout <= 8'b11000000; // 3937 : 192 - 0xc0
      12'hF62: dout <= 8'b11100000; // 3938 : 224 - 0xe0
      12'hF63: dout <= 8'b01100000; // 3939 :  96 - 0x60
      12'hF64: dout <= 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout <= 8'b00001100; // 3941 :  12 - 0xc
      12'hF66: dout <= 8'b00001110; // 3942 :  14 - 0xe
      12'hF67: dout <= 8'b00000110; // 3943 :   6 - 0x6
      12'hF68: dout <= 8'b01100000; // 3944 :  96 - 0x60 -- Background 0xed
      12'hF69: dout <= 8'b01110000; // 3945 : 112 - 0x70
      12'hF6A: dout <= 8'b00110000; // 3946 :  48 - 0x30
      12'hF6B: dout <= 8'b00000000; // 3947 :   0 - 0x0
      12'hF6C: dout <= 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout <= 8'b00001100; // 3949 :  12 - 0xc
      12'hF6E: dout <= 8'b00001110; // 3950 :  14 - 0xe
      12'hF6F: dout <= 8'b00000110; // 3951 :   6 - 0x6
      12'hF70: dout <= 8'b00000000; // 3952 :   0 - 0x0 -- Background 0xee
      12'hF71: dout <= 8'b00000000; // 3953 :   0 - 0x0
      12'hF72: dout <= 8'b01000010; // 3954 :  66 - 0x42
      12'hF73: dout <= 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout <= 8'b00000000; // 3956 :   0 - 0x0
      12'hF75: dout <= 8'b00000100; // 3957 :   4 - 0x4
      12'hF76: dout <= 8'b00000000; // 3958 :   0 - 0x0
      12'hF77: dout <= 8'b00000000; // 3959 :   0 - 0x0
      12'hF78: dout <= 8'b00000000; // 3960 :   0 - 0x0 -- Background 0xef
      12'hF79: dout <= 8'b00000000; // 3961 :   0 - 0x0
      12'hF7A: dout <= 8'b00000100; // 3962 :   4 - 0x4
      12'hF7B: dout <= 8'b00000000; // 3963 :   0 - 0x0
      12'hF7C: dout <= 8'b00100000; // 3964 :  32 - 0x20
      12'hF7D: dout <= 8'b00000000; // 3965 :   0 - 0x0
      12'hF7E: dout <= 8'b00000000; // 3966 :   0 - 0x0
      12'hF7F: dout <= 8'b00000000; // 3967 :   0 - 0x0
      12'hF80: dout <= 8'b00000000; // 3968 :   0 - 0x0 -- Background 0xf0
      12'hF81: dout <= 8'b00000000; // 3969 :   0 - 0x0
      12'hF82: dout <= 8'b00000000; // 3970 :   0 - 0x0
      12'hF83: dout <= 8'b00000000; // 3971 :   0 - 0x0
      12'hF84: dout <= 8'b00000000; // 3972 :   0 - 0x0
      12'hF85: dout <= 8'b00000000; // 3973 :   0 - 0x0
      12'hF86: dout <= 8'b00000000; // 3974 :   0 - 0x0
      12'hF87: dout <= 8'b00000000; // 3975 :   0 - 0x0
      12'hF88: dout <= 8'b10000000; // 3976 : 128 - 0x80 -- Background 0xf1
      12'hF89: dout <= 8'b10000000; // 3977 : 128 - 0x80
      12'hF8A: dout <= 8'b10000000; // 3978 : 128 - 0x80
      12'hF8B: dout <= 8'b10000000; // 3979 : 128 - 0x80
      12'hF8C: dout <= 8'b00000000; // 3980 :   0 - 0x0
      12'hF8D: dout <= 8'b00000000; // 3981 :   0 - 0x0
      12'hF8E: dout <= 8'b00000000; // 3982 :   0 - 0x0
      12'hF8F: dout <= 8'b00000000; // 3983 :   0 - 0x0
      12'hF90: dout <= 8'b11000000; // 3984 : 192 - 0xc0 -- Background 0xf2
      12'hF91: dout <= 8'b11000000; // 3985 : 192 - 0xc0
      12'hF92: dout <= 8'b11000000; // 3986 : 192 - 0xc0
      12'hF93: dout <= 8'b11000000; // 3987 : 192 - 0xc0
      12'hF94: dout <= 8'b00000000; // 3988 :   0 - 0x0
      12'hF95: dout <= 8'b00000000; // 3989 :   0 - 0x0
      12'hF96: dout <= 8'b00000000; // 3990 :   0 - 0x0
      12'hF97: dout <= 8'b00000000; // 3991 :   0 - 0x0
      12'hF98: dout <= 8'b11100000; // 3992 : 224 - 0xe0 -- Background 0xf3
      12'hF99: dout <= 8'b11100000; // 3993 : 224 - 0xe0
      12'hF9A: dout <= 8'b11100000; // 3994 : 224 - 0xe0
      12'hF9B: dout <= 8'b11100000; // 3995 : 224 - 0xe0
      12'hF9C: dout <= 8'b00000000; // 3996 :   0 - 0x0
      12'hF9D: dout <= 8'b00000000; // 3997 :   0 - 0x0
      12'hF9E: dout <= 8'b00000000; // 3998 :   0 - 0x0
      12'hF9F: dout <= 8'b00000000; // 3999 :   0 - 0x0
      12'hFA0: dout <= 8'b11110000; // 4000 : 240 - 0xf0 -- Background 0xf4
      12'hFA1: dout <= 8'b11110000; // 4001 : 240 - 0xf0
      12'hFA2: dout <= 8'b11110000; // 4002 : 240 - 0xf0
      12'hFA3: dout <= 8'b11110000; // 4003 : 240 - 0xf0
      12'hFA4: dout <= 8'b00000000; // 4004 :   0 - 0x0
      12'hFA5: dout <= 8'b00000000; // 4005 :   0 - 0x0
      12'hFA6: dout <= 8'b00000000; // 4006 :   0 - 0x0
      12'hFA7: dout <= 8'b00000000; // 4007 :   0 - 0x0
      12'hFA8: dout <= 8'b11111000; // 4008 : 248 - 0xf8 -- Background 0xf5
      12'hFA9: dout <= 8'b11111000; // 4009 : 248 - 0xf8
      12'hFAA: dout <= 8'b11111000; // 4010 : 248 - 0xf8
      12'hFAB: dout <= 8'b11111000; // 4011 : 248 - 0xf8
      12'hFAC: dout <= 8'b00000000; // 4012 :   0 - 0x0
      12'hFAD: dout <= 8'b00000000; // 4013 :   0 - 0x0
      12'hFAE: dout <= 8'b00000000; // 4014 :   0 - 0x0
      12'hFAF: dout <= 8'b00000000; // 4015 :   0 - 0x0
      12'hFB0: dout <= 8'b11111100; // 4016 : 252 - 0xfc -- Background 0xf6
      12'hFB1: dout <= 8'b11111100; // 4017 : 252 - 0xfc
      12'hFB2: dout <= 8'b11111100; // 4018 : 252 - 0xfc
      12'hFB3: dout <= 8'b11111100; // 4019 : 252 - 0xfc
      12'hFB4: dout <= 8'b00000000; // 4020 :   0 - 0x0
      12'hFB5: dout <= 8'b00000000; // 4021 :   0 - 0x0
      12'hFB6: dout <= 8'b00000000; // 4022 :   0 - 0x0
      12'hFB7: dout <= 8'b00000000; // 4023 :   0 - 0x0
      12'hFB8: dout <= 8'b11111110; // 4024 : 254 - 0xfe -- Background 0xf7
      12'hFB9: dout <= 8'b11111110; // 4025 : 254 - 0xfe
      12'hFBA: dout <= 8'b11111110; // 4026 : 254 - 0xfe
      12'hFBB: dout <= 8'b11111110; // 4027 : 254 - 0xfe
      12'hFBC: dout <= 8'b00000000; // 4028 :   0 - 0x0
      12'hFBD: dout <= 8'b00000000; // 4029 :   0 - 0x0
      12'hFBE: dout <= 8'b00000000; // 4030 :   0 - 0x0
      12'hFBF: dout <= 8'b00000000; // 4031 :   0 - 0x0
      12'hFC0: dout <= 8'b11111111; // 4032 : 255 - 0xff -- Background 0xf8
      12'hFC1: dout <= 8'b11111111; // 4033 : 255 - 0xff
      12'hFC2: dout <= 8'b11111111; // 4034 : 255 - 0xff
      12'hFC3: dout <= 8'b11111111; // 4035 : 255 - 0xff
      12'hFC4: dout <= 8'b00000000; // 4036 :   0 - 0x0
      12'hFC5: dout <= 8'b00000000; // 4037 :   0 - 0x0
      12'hFC6: dout <= 8'b00000000; // 4038 :   0 - 0x0
      12'hFC7: dout <= 8'b00000000; // 4039 :   0 - 0x0
      12'hFC8: dout <= 8'b00000000; // 4040 :   0 - 0x0 -- Background 0xf9
      12'hFC9: dout <= 8'b00000000; // 4041 :   0 - 0x0
      12'hFCA: dout <= 8'b00000000; // 4042 :   0 - 0x0
      12'hFCB: dout <= 8'b00000000; // 4043 :   0 - 0x0
      12'hFCC: dout <= 8'b01111111; // 4044 : 127 - 0x7f
      12'hFCD: dout <= 8'b01000000; // 4045 :  64 - 0x40
      12'hFCE: dout <= 8'b01000000; // 4046 :  64 - 0x40
      12'hFCF: dout <= 8'b01000000; // 4047 :  64 - 0x40
      12'hFD0: dout <= 8'b00000000; // 4048 :   0 - 0x0 -- Background 0xfa
      12'hFD1: dout <= 8'b00000000; // 4049 :   0 - 0x0
      12'hFD2: dout <= 8'b00000000; // 4050 :   0 - 0x0
      12'hFD3: dout <= 8'b00000000; // 4051 :   0 - 0x0
      12'hFD4: dout <= 8'b11111111; // 4052 : 255 - 0xff
      12'hFD5: dout <= 8'b00000000; // 4053 :   0 - 0x0
      12'hFD6: dout <= 8'b00000000; // 4054 :   0 - 0x0
      12'hFD7: dout <= 8'b00000000; // 4055 :   0 - 0x0
      12'hFD8: dout <= 8'b00000000; // 4056 :   0 - 0x0 -- Background 0xfb
      12'hFD9: dout <= 8'b00000000; // 4057 :   0 - 0x0
      12'hFDA: dout <= 8'b00000000; // 4058 :   0 - 0x0
      12'hFDB: dout <= 8'b00000000; // 4059 :   0 - 0x0
      12'hFDC: dout <= 8'b11111110; // 4060 : 254 - 0xfe
      12'hFDD: dout <= 8'b00000010; // 4061 :   2 - 0x2
      12'hFDE: dout <= 8'b00000010; // 4062 :   2 - 0x2
      12'hFDF: dout <= 8'b00000010; // 4063 :   2 - 0x2
      12'hFE0: dout <= 8'b01000000; // 4064 :  64 - 0x40 -- Background 0xfc
      12'hFE1: dout <= 8'b01000000; // 4065 :  64 - 0x40
      12'hFE2: dout <= 8'b01000000; // 4066 :  64 - 0x40
      12'hFE3: dout <= 8'b01111111; // 4067 : 127 - 0x7f
      12'hFE4: dout <= 8'b00000000; // 4068 :   0 - 0x0
      12'hFE5: dout <= 8'b00000000; // 4069 :   0 - 0x0
      12'hFE6: dout <= 8'b00000000; // 4070 :   0 - 0x0
      12'hFE7: dout <= 8'b00000000; // 4071 :   0 - 0x0
      12'hFE8: dout <= 8'b00000000; // 4072 :   0 - 0x0 -- Background 0xfd
      12'hFE9: dout <= 8'b00000000; // 4073 :   0 - 0x0
      12'hFEA: dout <= 8'b00000000; // 4074 :   0 - 0x0
      12'hFEB: dout <= 8'b11111111; // 4075 : 255 - 0xff
      12'hFEC: dout <= 8'b00000000; // 4076 :   0 - 0x0
      12'hFED: dout <= 8'b00000000; // 4077 :   0 - 0x0
      12'hFEE: dout <= 8'b00000000; // 4078 :   0 - 0x0
      12'hFEF: dout <= 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout <= 8'b00000010; // 4080 :   2 - 0x2 -- Background 0xfe
      12'hFF1: dout <= 8'b00000010; // 4081 :   2 - 0x2
      12'hFF2: dout <= 8'b00000010; // 4082 :   2 - 0x2
      12'hFF3: dout <= 8'b11111110; // 4083 : 254 - 0xfe
      12'hFF4: dout <= 8'b00000000; // 4084 :   0 - 0x0
      12'hFF5: dout <= 8'b00000000; // 4085 :   0 - 0x0
      12'hFF6: dout <= 8'b00000000; // 4086 :   0 - 0x0
      12'hFF7: dout <= 8'b00000000; // 4087 :   0 - 0x0
      12'hFF8: dout <= 8'b00000000; // 4088 :   0 - 0x0 -- Background 0xff
      12'hFF9: dout <= 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout <= 8'b00000000; // 4090 :   0 - 0x0
      12'hFFB: dout <= 8'b00000000; // 4091 :   0 - 0x0
      12'hFFC: dout <= 8'b00000000; // 4092 :   0 - 0x0
      12'hFFD: dout <= 8'b00000000; // 4093 :   0 - 0x0
      12'hFFE: dout <= 8'b00000000; // 4094 :   0 - 0x0
      12'hFFF: dout <= 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
