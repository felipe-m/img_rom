---   Background Pattern table BOTH COLOR PLANES
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: nova_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_NOVA_BG is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_NOVA_BG;

architecture BEHAVIORAL of ROM_PTABLE_NOVA_BG is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table both color planes
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Background 0x0
    "00001111", --    1 -  0x1  :   15 - 0xf
    "00000100", --    2 -  0x2  :    4 - 0x4
    "00000011", --    3 -  0x3  :    3 - 0x3
    "00000011", --    4 -  0x4  :    3 - 0x3
    "00000011", --    5 -  0x5  :    3 - 0x3
    "00000100", --    6 -  0x6  :    4 - 0x4
    "00111010", --    7 -  0x7  :   58 - 0x3a
    "00000000", --    8 -  0x8  :    0 - 0x0 -- plane 1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000011", --   10 -  0xa  :    3 - 0x3
    "00000001", --   11 -  0xb  :    1 - 0x1
    "00000001", --   12 -  0xc  :    1 - 0x1
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000011", --   14 -  0xe  :    3 - 0x3
    "00000001", --   15 -  0xf  :    1 - 0x1
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Background 0x1
    "00111000", --   17 - 0x11  :   56 - 0x38
    "11000110", --   18 - 0x12  :  198 - 0xc6
    "11001011", --   19 - 0x13  :  203 - 0xcb
    "11011100", --   20 - 0x14  :  220 - 0xdc
    "00111010", --   21 - 0x15  :   58 - 0x3a
    "10011010", --   22 - 0x16  :  154 - 0x9a
    "10000001", --   23 - 0x17  :  129 - 0x81
    "00000000", --   24 - 0x18  :    0 - 0x0 -- plane 1
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00111000", --   26 - 0x1a  :   56 - 0x38
    "10110100", --   27 - 0x1b  :  180 - 0xb4
    "10101000", --   28 - 0x1c  :  168 - 0xa8
    "11010100", --   29 - 0x1d  :  212 - 0xd4
    "01110100", --   30 - 0x1e  :  116 - 0x74
    "01111110", --   31 - 0x1f  :  126 - 0x7e
    "01000101", --   32 - 0x20  :   69 - 0x45 -- Background 0x2
    "10000111", --   33 - 0x21  :  135 - 0x87
    "10000011", --   34 - 0x22  :  131 - 0x83
    "10000001", --   35 - 0x23  :  129 - 0x81
    "10000001", --   36 - 0x24  :  129 - 0x81
    "10000001", --   37 - 0x25  :  129 - 0x81
    "01000001", --   38 - 0x26  :   65 - 0x41
    "00100001", --   39 - 0x27  :   33 - 0x21
    "00111000", --   40 - 0x28  :   56 - 0x38 -- plane 1
    "01111000", --   41 - 0x29  :  120 - 0x78
    "01111100", --   42 - 0x2a  :  124 - 0x7c
    "01111110", --   43 - 0x2b  :  126 - 0x7e
    "01111110", --   44 - 0x2c  :  126 - 0x7e
    "01111110", --   45 - 0x2d  :  126 - 0x7e
    "00111110", --   46 - 0x2e  :   62 - 0x3e
    "00011110", --   47 - 0x2f  :   30 - 0x1e
    "01111111", --   48 - 0x30  :  127 - 0x7f -- Background 0x3
    "01111110", --   49 - 0x31  :  126 - 0x7e
    "11111100", --   50 - 0x32  :  252 - 0xfc
    "00111000", --   51 - 0x33  :   56 - 0x38
    "00011000", --   52 - 0x34  :   24 - 0x18
    "10001100", --   53 - 0x35  :  140 - 0x8c
    "11000100", --   54 - 0x36  :  196 - 0xc4
    "11111100", --   55 - 0x37  :  252 - 0xfc
    "11110110", --   56 - 0x38  :  246 - 0xf6 -- plane 1
    "11110000", --   57 - 0x39  :  240 - 0xf0
    "00111000", --   58 - 0x3a  :   56 - 0x38
    "11010000", --   59 - 0x3b  :  208 - 0xd0
    "11100000", --   60 - 0x3c  :  224 - 0xe0
    "01110000", --   61 - 0x3d  :  112 - 0x70
    "10111000", --   62 - 0x3e  :  184 - 0xb8
    "01000000", --   63 - 0x3f  :   64 - 0x40
    "00100011", --   64 - 0x40  :   35 - 0x23 -- Background 0x4
    "00100011", --   65 - 0x41  :   35 - 0x23
    "00100001", --   66 - 0x42  :   33 - 0x21
    "00100000", --   67 - 0x43  :   32 - 0x20
    "00010011", --   68 - 0x44  :   19 - 0x13
    "00001100", --   69 - 0x45  :   12 - 0xc
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00011100", --   72 - 0x48  :   28 - 0x1c -- plane 1
    "00011100", --   73 - 0x49  :   28 - 0x1c
    "00011110", --   74 - 0x4a  :   30 - 0x1e
    "00011111", --   75 - 0x4b  :   31 - 0x1f
    "00001100", --   76 - 0x4c  :   12 - 0xc
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "11111100", --   80 - 0x50  :  252 - 0xfc -- Background 0x5
    "11111100", --   81 - 0x51  :  252 - 0xfc
    "11111100", --   82 - 0x52  :  252 - 0xfc
    "11111100", --   83 - 0x53  :  252 - 0xfc
    "10010000", --   84 - 0x54  :  144 - 0x90
    "10010000", --   85 - 0x55  :  144 - 0x90
    "10001000", --   86 - 0x56  :  136 - 0x88
    "11111000", --   87 - 0x57  :  248 - 0xf8
    "10101000", --   88 - 0x58  :  168 - 0xa8 -- plane 1
    "01010000", --   89 - 0x59  :   80 - 0x50
    "10101000", --   90 - 0x5a  :  168 - 0xa8
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "01100000", --   92 - 0x5c  :   96 - 0x60
    "01100000", --   93 - 0x5d  :   96 - 0x60
    "01110000", --   94 - 0x5e  :  112 - 0x70
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00100011", --   96 - 0x60  :   35 - 0x23 -- Background 0x6
    "00100011", --   97 - 0x61  :   35 - 0x23
    "00100001", --   98 - 0x62  :   33 - 0x21
    "00100000", --   99 - 0x63  :   32 - 0x20
    "00010011", --  100 - 0x64  :   19 - 0x13
    "00001101", --  101 - 0x65  :   13 - 0xd
    "00000010", --  102 - 0x66  :    2 - 0x2
    "00000001", --  103 - 0x67  :    1 - 0x1
    "00011100", --  104 - 0x68  :   28 - 0x1c -- plane 1
    "00011100", --  105 - 0x69  :   28 - 0x1c
    "00011110", --  106 - 0x6a  :   30 - 0x1e
    "00011111", --  107 - 0x6b  :   31 - 0x1f
    "00001100", --  108 - 0x6c  :   12 - 0xc
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000001", --  110 - 0x6e  :    1 - 0x1
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "11111100", --  112 - 0x70  :  252 - 0xfc -- Background 0x7
    "11111100", --  113 - 0x71  :  252 - 0xfc
    "11111100", --  114 - 0x72  :  252 - 0xfc
    "11111100", --  115 - 0x73  :  252 - 0xfc
    "10100100", --  116 - 0x74  :  164 - 0xa4
    "00100100", --  117 - 0x75  :   36 - 0x24
    "01010010", --  118 - 0x76  :   82 - 0x52
    "11101110", --  119 - 0x77  :  238 - 0xee
    "10101000", --  120 - 0x78  :  168 - 0xa8 -- plane 1
    "01010000", --  121 - 0x79  :   80 - 0x50
    "10101000", --  122 - 0x7a  :  168 - 0xa8
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "01011000", --  124 - 0x7c  :   88 - 0x58
    "11011000", --  125 - 0x7d  :  216 - 0xd8
    "10001100", --  126 - 0x7e  :  140 - 0x8c
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00100011", --  128 - 0x80  :   35 - 0x23 -- Background 0x8
    "00100011", --  129 - 0x81  :   35 - 0x23
    "00100001", --  130 - 0x82  :   33 - 0x21
    "00100000", --  131 - 0x83  :   32 - 0x20
    "00010011", --  132 - 0x84  :   19 - 0x13
    "00001101", --  133 - 0x85  :   13 - 0xd
    "00000001", --  134 - 0x86  :    1 - 0x1
    "00000001", --  135 - 0x87  :    1 - 0x1
    "00011100", --  136 - 0x88  :   28 - 0x1c -- plane 1
    "00011100", --  137 - 0x89  :   28 - 0x1c
    "00011110", --  138 - 0x8a  :   30 - 0x1e
    "00011111", --  139 - 0x8b  :   31 - 0x1f
    "00001100", --  140 - 0x8c  :   12 - 0xc
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "11111110", --  144 - 0x90  :  254 - 0xfe -- Background 0x9
    "11111110", --  145 - 0x91  :  254 - 0xfe
    "11111110", --  146 - 0x92  :  254 - 0xfe
    "11111111", --  147 - 0x93  :  255 - 0xff
    "10010001", --  148 - 0x94  :  145 - 0x91
    "00101111", --  149 - 0x95  :   47 - 0x2f
    "01000000", --  150 - 0x96  :   64 - 0x40
    "11100000", --  151 - 0x97  :  224 - 0xe0
    "10101000", --  152 - 0x98  :  168 - 0xa8 -- plane 1
    "01010100", --  153 - 0x99  :   84 - 0x54
    "10101000", --  154 - 0x9a  :  168 - 0xa8
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "01101110", --  156 - 0x9c  :  110 - 0x6e
    "11000000", --  157 - 0x9d  :  192 - 0xc0
    "10000000", --  158 - 0x9e  :  128 - 0x80
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00100011", --  160 - 0xa0  :   35 - 0x23 -- Background 0xa
    "00100011", --  161 - 0xa1  :   35 - 0x23
    "00100001", --  162 - 0xa2  :   33 - 0x21
    "00100000", --  163 - 0xa3  :   32 - 0x20
    "00010011", --  164 - 0xa4  :   19 - 0x13
    "00001110", --  165 - 0xa5  :   14 - 0xe
    "00000001", --  166 - 0xa6  :    1 - 0x1
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00011100", --  168 - 0xa8  :   28 - 0x1c -- plane 1
    "00011100", --  169 - 0xa9  :   28 - 0x1c
    "00011110", --  170 - 0xaa  :   30 - 0x1e
    "00011111", --  171 - 0xab  :   31 - 0x1f
    "00001100", --  172 - 0xac  :   12 - 0xc
    "00000001", --  173 - 0xad  :    1 - 0x1
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "11111110", --  176 - 0xb0  :  254 - 0xfe -- Background 0xb
    "11111110", --  177 - 0xb1  :  254 - 0xfe
    "11111110", --  178 - 0xb2  :  254 - 0xfe
    "11111100", --  179 - 0xb3  :  252 - 0xfc
    "00100100", --  180 - 0xb4  :   36 - 0x24
    "00100010", --  181 - 0xb5  :   34 - 0x22
    "11010010", --  182 - 0xb6  :  210 - 0xd2
    "00001111", --  183 - 0xb7  :   15 - 0xf
    "10101000", --  184 - 0xb8  :  168 - 0xa8 -- plane 1
    "01010100", --  185 - 0xb9  :   84 - 0x54
    "10101000", --  186 - 0xba  :  168 - 0xa8
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "11011000", --  188 - 0xbc  :  216 - 0xd8
    "11011100", --  189 - 0xbd  :  220 - 0xdc
    "00001100", --  190 - 0xbe  :   12 - 0xc
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "01111111", --  192 - 0xc0  :  127 - 0x7f -- Background 0xc
    "01111110", --  193 - 0xc1  :  126 - 0x7e
    "11111100", --  194 - 0xc2  :  252 - 0xfc
    "00000010", --  195 - 0xc3  :    2 - 0x2
    "00000100", --  196 - 0xc4  :    4 - 0x4
    "11111100", --  197 - 0xc5  :  252 - 0xfc
    "11111100", --  198 - 0xc6  :  252 - 0xfc
    "11111110", --  199 - 0xc7  :  254 - 0xfe
    "11110110", --  200 - 0xc8  :  246 - 0xf6 -- plane 1
    "11110000", --  201 - 0xc9  :  240 - 0xf0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "11111100", --  203 - 0xcb  :  252 - 0xfc
    "11111000", --  204 - 0xcc  :  248 - 0xf8
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "10101000", --  206 - 0xce  :  168 - 0xa8
    "01010100", --  207 - 0xcf  :   84 - 0x54
    "01000101", --  208 - 0xd0  :   69 - 0x45 -- Background 0xd
    "10000111", --  209 - 0xd1  :  135 - 0x87
    "10000011", --  210 - 0xd2  :  131 - 0x83
    "10000010", --  211 - 0xd3  :  130 - 0x82
    "10000010", --  212 - 0xd4  :  130 - 0x82
    "10000100", --  213 - 0xd5  :  132 - 0x84
    "01000100", --  214 - 0xd6  :   68 - 0x44
    "00100100", --  215 - 0xd7  :   36 - 0x24
    "00111000", --  216 - 0xd8  :   56 - 0x38 -- plane 1
    "01111000", --  217 - 0xd9  :  120 - 0x78
    "01111100", --  218 - 0xda  :  124 - 0x7c
    "01111101", --  219 - 0xdb  :  125 - 0x7d
    "01111101", --  220 - 0xdc  :  125 - 0x7d
    "01111011", --  221 - 0xdd  :  123 - 0x7b
    "00111011", --  222 - 0xde  :   59 - 0x3b
    "00011011", --  223 - 0xdf  :   27 - 0x1b
    "01111111", --  224 - 0xe0  :  127 - 0x7f -- Background 0xe
    "01111110", --  225 - 0xe1  :  126 - 0x7e
    "11111100", --  226 - 0xe2  :  252 - 0xfc
    "11111000", --  227 - 0xe3  :  248 - 0xf8
    "01111000", --  228 - 0xe4  :  120 - 0x78
    "01111100", --  229 - 0xe5  :  124 - 0x7c
    "11111100", --  230 - 0xe6  :  252 - 0xfc
    "11111110", --  231 - 0xe7  :  254 - 0xfe
    "11110110", --  232 - 0xe8  :  246 - 0xf6 -- plane 1
    "11110000", --  233 - 0xe9  :  240 - 0xf0
    "01111000", --  234 - 0xea  :  120 - 0x78
    "01110000", --  235 - 0xeb  :  112 - 0x70
    "10100000", --  236 - 0xec  :  160 - 0xa0
    "10010000", --  237 - 0xed  :  144 - 0x90
    "00101000", --  238 - 0xee  :   40 - 0x28
    "01010100", --  239 - 0xef  :   84 - 0x54
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Background 0xf
    "00001111", --  241 - 0xf1  :   15 - 0xf
    "00000100", --  242 - 0xf2  :    4 - 0x4
    "00000011", --  243 - 0xf3  :    3 - 0x3
    "00000011", --  244 - 0xf4  :    3 - 0x3
    "00000011", --  245 - 0xf5  :    3 - 0x3
    "00000100", --  246 - 0xf6  :    4 - 0x4
    "00000010", --  247 - 0xf7  :    2 - 0x2
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- plane 1
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000011", --  250 - 0xfa  :    3 - 0x3
    "00000001", --  251 - 0xfb  :    1 - 0x1
    "00000001", --  252 - 0xfc  :    1 - 0x1
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000011", --  254 - 0xfe  :    3 - 0x3
    "00000001", --  255 - 0xff  :    1 - 0x1
    "00000111", --  256 - 0x100  :    7 - 0x7 -- Background 0x10
    "00001100", --  257 - 0x101  :   12 - 0xc
    "00010000", --  258 - 0x102  :   16 - 0x10
    "00010000", --  259 - 0x103  :   16 - 0x10
    "00010000", --  260 - 0x104  :   16 - 0x10
    "00100000", --  261 - 0x105  :   32 - 0x20
    "00100000", --  262 - 0x106  :   32 - 0x20
    "00100001", --  263 - 0x107  :   33 - 0x21
    "00000000", --  264 - 0x108  :    0 - 0x0 -- plane 1
    "00000011", --  265 - 0x109  :    3 - 0x3
    "00001111", --  266 - 0x10a  :   15 - 0xf
    "00001111", --  267 - 0x10b  :   15 - 0xf
    "00001111", --  268 - 0x10c  :   15 - 0xf
    "00011111", --  269 - 0x10d  :   31 - 0x1f
    "00011111", --  270 - 0x10e  :   31 - 0x1f
    "00011110", --  271 - 0x10f  :   30 - 0x1e
    "11111111", --  272 - 0x110  :  255 - 0xff -- Background 0x11
    "01111110", --  273 - 0x111  :  126 - 0x7e
    "01111100", --  274 - 0x112  :  124 - 0x7c
    "01111000", --  275 - 0x113  :  120 - 0x78
    "01011000", --  276 - 0x114  :   88 - 0x58
    "10001100", --  277 - 0x115  :  140 - 0x8c
    "11000100", --  278 - 0x116  :  196 - 0xc4
    "11111100", --  279 - 0x117  :  252 - 0xfc
    "00110110", --  280 - 0x118  :   54 - 0x36 -- plane 1
    "10110000", --  281 - 0x119  :  176 - 0xb0
    "10111000", --  282 - 0x11a  :  184 - 0xb8
    "10010000", --  283 - 0x11b  :  144 - 0x90
    "10100000", --  284 - 0x11c  :  160 - 0xa0
    "01110000", --  285 - 0x11d  :  112 - 0x70
    "00111000", --  286 - 0x11e  :   56 - 0x38
    "01000000", --  287 - 0x11f  :   64 - 0x40
    "00100011", --  288 - 0x120  :   35 - 0x23 -- Background 0x12
    "00100011", --  289 - 0x121  :   35 - 0x23
    "00100001", --  290 - 0x122  :   33 - 0x21
    "00100000", --  291 - 0x123  :   32 - 0x20
    "00010011", --  292 - 0x124  :   19 - 0x13
    "00001100", --  293 - 0x125  :   12 - 0xc
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00011100", --  296 - 0x128  :   28 - 0x1c -- plane 1
    "00011100", --  297 - 0x129  :   28 - 0x1c
    "00011110", --  298 - 0x12a  :   30 - 0x1e
    "00011111", --  299 - 0x12b  :   31 - 0x1f
    "00001100", --  300 - 0x12c  :   12 - 0xc
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000001", --  304 - 0x130  :    1 - 0x1 -- Background 0x13
    "00000001", --  305 - 0x131  :    1 - 0x1
    "00000011", --  306 - 0x132  :    3 - 0x3
    "00000100", --  307 - 0x133  :    4 - 0x4
    "00001000", --  308 - 0x134  :    8 - 0x8
    "00010000", --  309 - 0x135  :   16 - 0x10
    "00010000", --  310 - 0x136  :   16 - 0x10
    "00100000", --  311 - 0x137  :   32 - 0x20
    "00000000", --  312 - 0x138  :    0 - 0x0 -- plane 1
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000011", --  315 - 0x13b  :    3 - 0x3
    "00000111", --  316 - 0x13c  :    7 - 0x7
    "00001111", --  317 - 0x13d  :   15 - 0xf
    "00001111", --  318 - 0x13e  :   15 - 0xf
    "00011111", --  319 - 0x13f  :   31 - 0x1f
    "01111111", --  320 - 0x140  :  127 - 0x7f -- Background 0x14
    "11111110", --  321 - 0x141  :  254 - 0xfe
    "00000110", --  322 - 0x142  :    6 - 0x6
    "00000001", --  323 - 0x143  :    1 - 0x1
    "00000001", --  324 - 0x144  :    1 - 0x1
    "00000001", --  325 - 0x145  :    1 - 0x1
    "00000111", --  326 - 0x146  :    7 - 0x7
    "11111110", --  327 - 0x147  :  254 - 0xfe
    "11110110", --  328 - 0x148  :  246 - 0xf6 -- plane 1
    "00000000", --  329 - 0x149  :    0 - 0x0
    "11111000", --  330 - 0x14a  :  248 - 0xf8
    "11111110", --  331 - 0x14b  :  254 - 0xfe
    "11111110", --  332 - 0x14c  :  254 - 0xfe
    "11111110", --  333 - 0x14d  :  254 - 0xfe
    "11111000", --  334 - 0x14e  :  248 - 0xf8
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00000101", --  336 - 0x150  :    5 - 0x5 -- Background 0x15
    "00000101", --  337 - 0x151  :    5 - 0x5
    "00000111", --  338 - 0x152  :    7 - 0x7
    "00000100", --  339 - 0x153  :    4 - 0x4
    "00000100", --  340 - 0x154  :    4 - 0x4
    "00001111", --  341 - 0x155  :   15 - 0xf
    "00110000", --  342 - 0x156  :   48 - 0x30
    "01000000", --  343 - 0x157  :   64 - 0x40
    "00000011", --  344 - 0x158  :    3 - 0x3 -- plane 1
    "00000011", --  345 - 0x159  :    3 - 0x3
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000011", --  347 - 0x15b  :    3 - 0x3
    "00000011", --  348 - 0x15c  :    3 - 0x3
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00001111", --  350 - 0x15e  :   15 - 0xf
    "00111111", --  351 - 0x15f  :   63 - 0x3f
    "11111100", --  352 - 0x160  :  252 - 0xfc -- Background 0x16
    "11111000", --  353 - 0x161  :  248 - 0xf8
    "11110000", --  354 - 0x162  :  240 - 0xf0
    "11100000", --  355 - 0x163  :  224 - 0xe0
    "01100000", --  356 - 0x164  :   96 - 0x60
    "11110000", --  357 - 0x165  :  240 - 0xf0
    "00011100", --  358 - 0x166  :   28 - 0x1c
    "00000010", --  359 - 0x167  :    2 - 0x2
    "11011000", --  360 - 0x168  :  216 - 0xd8 -- plane 1
    "11000000", --  361 - 0x169  :  192 - 0xc0
    "11100000", --  362 - 0x16a  :  224 - 0xe0
    "01000000", --  363 - 0x16b  :   64 - 0x40
    "10000000", --  364 - 0x16c  :  128 - 0x80
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "11100000", --  366 - 0x16e  :  224 - 0xe0
    "11111100", --  367 - 0x16f  :  252 - 0xfc
    "10000000", --  368 - 0x170  :  128 - 0x80 -- Background 0x17
    "10000000", --  369 - 0x171  :  128 - 0x80
    "10000000", --  370 - 0x172  :  128 - 0x80
    "10000011", --  371 - 0x173  :  131 - 0x83
    "01001111", --  372 - 0x174  :   79 - 0x4f
    "00110010", --  373 - 0x175  :   50 - 0x32
    "00000010", --  374 - 0x176  :    2 - 0x2
    "00000011", --  375 - 0x177  :    3 - 0x3
    "01111111", --  376 - 0x178  :  127 - 0x7f -- plane 1
    "01111111", --  377 - 0x179  :  127 - 0x7f
    "01111111", --  378 - 0x17a  :  127 - 0x7f
    "01111100", --  379 - 0x17b  :  124 - 0x7c
    "00110000", --  380 - 0x17c  :   48 - 0x30
    "00000001", --  381 - 0x17d  :    1 - 0x1
    "00000001", --  382 - 0x17e  :    1 - 0x1
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000010", --  384 - 0x180  :    2 - 0x2 -- Background 0x18
    "00000001", --  385 - 0x181  :    1 - 0x1
    "00000010", --  386 - 0x182  :    2 - 0x2
    "11111100", --  387 - 0x183  :  252 - 0xfc
    "11000000", --  388 - 0x184  :  192 - 0xc0
    "01000000", --  389 - 0x185  :   64 - 0x40
    "00100000", --  390 - 0x186  :   32 - 0x20
    "11100000", --  391 - 0x187  :  224 - 0xe0
    "11111100", --  392 - 0x188  :  252 - 0xfc -- plane 1
    "11111110", --  393 - 0x189  :  254 - 0xfe
    "11111100", --  394 - 0x18a  :  252 - 0xfc
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "10000000", --  397 - 0x18d  :  128 - 0x80
    "11000000", --  398 - 0x18e  :  192 - 0xc0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00001011", --  400 - 0x190  :   11 - 0xb -- Background 0x19
    "00001011", --  401 - 0x191  :   11 - 0xb
    "00001111", --  402 - 0x192  :   15 - 0xf
    "00001001", --  403 - 0x193  :    9 - 0x9
    "00001000", --  404 - 0x194  :    8 - 0x8
    "00001001", --  405 - 0x195  :    9 - 0x9
    "00001111", --  406 - 0x196  :   15 - 0xf
    "00110000", --  407 - 0x197  :   48 - 0x30
    "00000111", --  408 - 0x198  :    7 - 0x7 -- plane 1
    "00000111", --  409 - 0x199  :    7 - 0x7
    "00000001", --  410 - 0x19a  :    1 - 0x1
    "00000110", --  411 - 0x19b  :    6 - 0x6
    "00000111", --  412 - 0x19c  :    7 - 0x7
    "00000110", --  413 - 0x19d  :    6 - 0x6
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00001111", --  415 - 0x19f  :   15 - 0xf
    "11111000", --  416 - 0x1a0  :  248 - 0xf8 -- Background 0x1a
    "11110000", --  417 - 0x1a1  :  240 - 0xf0
    "11100000", --  418 - 0x1a2  :  224 - 0xe0
    "11000000", --  419 - 0x1a3  :  192 - 0xc0
    "11000000", --  420 - 0x1a4  :  192 - 0xc0
    "11000000", --  421 - 0x1a5  :  192 - 0xc0
    "11111000", --  422 - 0x1a6  :  248 - 0xf8
    "00011111", --  423 - 0x1a7  :   31 - 0x1f
    "10110000", --  424 - 0x1a8  :  176 - 0xb0 -- plane 1
    "10000000", --  425 - 0x1a9  :  128 - 0x80
    "11000000", --  426 - 0x1aa  :  192 - 0xc0
    "10000000", --  427 - 0x1ab  :  128 - 0x80
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "11100000", --  431 - 0x1af  :  224 - 0xe0
    "01000000", --  432 - 0x1b0  :   64 - 0x40 -- Background 0x1b
    "01000000", --  433 - 0x1b1  :   64 - 0x40
    "10000000", --  434 - 0x1b2  :  128 - 0x80
    "10000000", --  435 - 0x1b3  :  128 - 0x80
    "01000000", --  436 - 0x1b4  :   64 - 0x40
    "00111111", --  437 - 0x1b5  :   63 - 0x3f
    "00000100", --  438 - 0x1b6  :    4 - 0x4
    "00000111", --  439 - 0x1b7  :    7 - 0x7
    "00111111", --  440 - 0x1b8  :   63 - 0x3f -- plane 1
    "00111111", --  441 - 0x1b9  :   63 - 0x3f
    "01111111", --  442 - 0x1ba  :  127 - 0x7f
    "01111111", --  443 - 0x1bb  :  127 - 0x7f
    "00111111", --  444 - 0x1bc  :   63 - 0x3f
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000011", --  446 - 0x1be  :    3 - 0x3
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Background 0x1c
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "11111111", --  453 - 0x1c5  :  255 - 0xff
    "01000000", --  454 - 0x1c6  :   64 - 0x40
    "11000000", --  455 - 0x1c7  :  192 - 0xc0
    "11111111", --  456 - 0x1c8  :  255 - 0xff -- plane 1
    "11111111", --  457 - 0x1c9  :  255 - 0xff
    "11111111", --  458 - 0x1ca  :  255 - 0xff
    "11111111", --  459 - 0x1cb  :  255 - 0xff
    "11111111", --  460 - 0x1cc  :  255 - 0xff
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "10000000", --  462 - 0x1ce  :  128 - 0x80
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "11000000", --  464 - 0x1d0  :  192 - 0xc0 -- Background 0x1d
    "00100000", --  465 - 0x1d1  :   32 - 0x20
    "00100000", --  466 - 0x1d2  :   32 - 0x20
    "00100000", --  467 - 0x1d3  :   32 - 0x20
    "01000000", --  468 - 0x1d4  :   64 - 0x40
    "10000000", --  469 - 0x1d5  :  128 - 0x80
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- plane 1
    "11000000", --  473 - 0x1d9  :  192 - 0xc0
    "11000000", --  474 - 0x1da  :  192 - 0xc0
    "11000000", --  475 - 0x1db  :  192 - 0xc0
    "10000000", --  476 - 0x1dc  :  128 - 0x80
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "01111111", --  480 - 0x1e0  :  127 - 0x7f -- Background 0x1e
    "01100010", --  481 - 0x1e1  :   98 - 0x62
    "11000100", --  482 - 0x1e2  :  196 - 0xc4
    "00011000", --  483 - 0x1e3  :   24 - 0x18
    "00111100", --  484 - 0x1e4  :   60 - 0x3c
    "11111110", --  485 - 0x1e5  :  254 - 0xfe
    "11111110", --  486 - 0x1e6  :  254 - 0xfe
    "11111110", --  487 - 0x1e7  :  254 - 0xfe
    "11100000", --  488 - 0x1e8  :  224 - 0xe0 -- plane 1
    "10011100", --  489 - 0x1e9  :  156 - 0x9c
    "00111000", --  490 - 0x1ea  :   56 - 0x38
    "11100000", --  491 - 0x1eb  :  224 - 0xe0
    "11001000", --  492 - 0x1ec  :  200 - 0xc8
    "00010100", --  493 - 0x1ed  :   20 - 0x14
    "10101000", --  494 - 0x1ee  :  168 - 0xa8
    "01010100", --  495 - 0x1ef  :   84 - 0x54
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Background 0x1f
    "00111000", --  497 - 0x1f1  :   56 - 0x38
    "11000110", --  498 - 0x1f2  :  198 - 0xc6
    "11001011", --  499 - 0x1f3  :  203 - 0xcb
    "11011100", --  500 - 0x1f4  :  220 - 0xdc
    "00111010", --  501 - 0x1f5  :   58 - 0x3a
    "10011010", --  502 - 0x1f6  :  154 - 0x9a
    "11100001", --  503 - 0x1f7  :  225 - 0xe1
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- plane 1
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00111000", --  506 - 0x1fa  :   56 - 0x38
    "10110100", --  507 - 0x1fb  :  180 - 0xb4
    "10101000", --  508 - 0x1fc  :  168 - 0xa8
    "11010100", --  509 - 0x1fd  :  212 - 0xd4
    "01110100", --  510 - 0x1fe  :  116 - 0x74
    "00011110", --  511 - 0x1ff  :   30 - 0x1e
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Background 0x20
    "00011100", --  513 - 0x201  :   28 - 0x1c
    "00010011", --  514 - 0x202  :   19 - 0x13
    "00001000", --  515 - 0x203  :    8 - 0x8
    "00010000", --  516 - 0x204  :   16 - 0x10
    "00001000", --  517 - 0x205  :    8 - 0x8
    "00010000", --  518 - 0x206  :   16 - 0x10
    "00010000", --  519 - 0x207  :   16 - 0x10
    "00000000", --  520 - 0x208  :    0 - 0x0 -- plane 1
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00001100", --  522 - 0x20a  :   12 - 0xc
    "00000111", --  523 - 0x20b  :    7 - 0x7
    "00001111", --  524 - 0x20c  :   15 - 0xf
    "00000111", --  525 - 0x20d  :    7 - 0x7
    "00001111", --  526 - 0x20e  :   15 - 0xf
    "00001111", --  527 - 0x20f  :   15 - 0xf
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Background 0x21
    "00111000", --  529 - 0x211  :   56 - 0x38
    "11001000", --  530 - 0x212  :  200 - 0xc8
    "00010000", --  531 - 0x213  :   16 - 0x10
    "00001000", --  532 - 0x214  :    8 - 0x8
    "00010000", --  533 - 0x215  :   16 - 0x10
    "00001000", --  534 - 0x216  :    8 - 0x8
    "00001000", --  535 - 0x217  :    8 - 0x8
    "00000000", --  536 - 0x218  :    0 - 0x0 -- plane 1
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00110000", --  538 - 0x21a  :   48 - 0x30
    "11100000", --  539 - 0x21b  :  224 - 0xe0
    "11110000", --  540 - 0x21c  :  240 - 0xf0
    "11100000", --  541 - 0x21d  :  224 - 0xe0
    "11110000", --  542 - 0x21e  :  240 - 0xf0
    "11110000", --  543 - 0x21f  :  240 - 0xf0
    "00001000", --  544 - 0x220  :    8 - 0x8 -- Background 0x22
    "00011100", --  545 - 0x221  :   28 - 0x1c
    "00100111", --  546 - 0x222  :   39 - 0x27
    "00101111", --  547 - 0x223  :   47 - 0x2f
    "00011111", --  548 - 0x224  :   31 - 0x1f
    "00001111", --  549 - 0x225  :   15 - 0xf
    "00001111", --  550 - 0x226  :   15 - 0xf
    "00001111", --  551 - 0x227  :   15 - 0xf
    "00000111", --  552 - 0x228  :    7 - 0x7 -- plane 1
    "00000011", --  553 - 0x229  :    3 - 0x3
    "00011000", --  554 - 0x22a  :   24 - 0x18
    "00010101", --  555 - 0x22b  :   21 - 0x15
    "00000010", --  556 - 0x22c  :    2 - 0x2
    "00000101", --  557 - 0x22d  :    5 - 0x5
    "00000010", --  558 - 0x22e  :    2 - 0x2
    "00000100", --  559 - 0x22f  :    4 - 0x4
    "00010000", --  560 - 0x230  :   16 - 0x10 -- Background 0x23
    "00111100", --  561 - 0x231  :   60 - 0x3c
    "11000010", --  562 - 0x232  :  194 - 0xc2
    "10000010", --  563 - 0x233  :  130 - 0x82
    "10000010", --  564 - 0x234  :  130 - 0x82
    "10000010", --  565 - 0x235  :  130 - 0x82
    "00010010", --  566 - 0x236  :   18 - 0x12
    "00011100", --  567 - 0x237  :   28 - 0x1c
    "11100000", --  568 - 0x238  :  224 - 0xe0 -- plane 1
    "11000000", --  569 - 0x239  :  192 - 0xc0
    "00111100", --  570 - 0x23a  :   60 - 0x3c
    "01111100", --  571 - 0x23b  :  124 - 0x7c
    "01111100", --  572 - 0x23c  :  124 - 0x7c
    "01111100", --  573 - 0x23d  :  124 - 0x7c
    "11101100", --  574 - 0x23e  :  236 - 0xec
    "11100000", --  575 - 0x23f  :  224 - 0xe0
    "00001111", --  576 - 0x240  :   15 - 0xf -- Background 0x24
    "00001110", --  577 - 0x241  :   14 - 0xe
    "00010100", --  578 - 0x242  :   20 - 0x14
    "00010100", --  579 - 0x243  :   20 - 0x14
    "00010010", --  580 - 0x244  :   18 - 0x12
    "00100101", --  581 - 0x245  :   37 - 0x25
    "01000100", --  582 - 0x246  :   68 - 0x44
    "00111000", --  583 - 0x247  :   56 - 0x38
    "00000010", --  584 - 0x248  :    2 - 0x2 -- plane 1
    "00000101", --  585 - 0x249  :    5 - 0x5
    "00001011", --  586 - 0x24a  :   11 - 0xb
    "00001011", --  587 - 0x24b  :   11 - 0xb
    "00001101", --  588 - 0x24c  :   13 - 0xd
    "00011000", --  589 - 0x24d  :   24 - 0x18
    "00111000", --  590 - 0x24e  :   56 - 0x38
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00010000", --  592 - 0x250  :   16 - 0x10 -- Background 0x25
    "00010000", --  593 - 0x251  :   16 - 0x10
    "00010000", --  594 - 0x252  :   16 - 0x10
    "00101100", --  595 - 0x253  :   44 - 0x2c
    "01000100", --  596 - 0x254  :   68 - 0x44
    "11000100", --  597 - 0x255  :  196 - 0xc4
    "00111000", --  598 - 0x256  :   56 - 0x38
    "00000000", --  599 - 0x257  :    0 - 0x0
    "11100000", --  600 - 0x258  :  224 - 0xe0 -- plane 1
    "11100000", --  601 - 0x259  :  224 - 0xe0
    "11100000", --  602 - 0x25a  :  224 - 0xe0
    "11010000", --  603 - 0x25b  :  208 - 0xd0
    "10111000", --  604 - 0x25c  :  184 - 0xb8
    "00111000", --  605 - 0x25d  :   56 - 0x38
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Background 0x26
    "00000000", --  609 - 0x261  :    0 - 0x0
    "00000000", --  610 - 0x262  :    0 - 0x0
    "00000000", --  611 - 0x263  :    0 - 0x0
    "00000000", --  612 - 0x264  :    0 - 0x0
    "00000000", --  613 - 0x265  :    0 - 0x0
    "00000000", --  614 - 0x266  :    0 - 0x0
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0 -- plane 1
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Background 0x27
    "00000000", --  625 - 0x271  :    0 - 0x0
    "00000000", --  626 - 0x272  :    0 - 0x0
    "00000000", --  627 - 0x273  :    0 - 0x0
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000000", --  629 - 0x275  :    0 - 0x0
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0 -- plane 1
    "00000000", --  633 - 0x279  :    0 - 0x0
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "00000000", --  635 - 0x27b  :    0 - 0x0
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Background 0x28
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- plane 1
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00100000", --  656 - 0x290  :   32 - 0x20 -- Background 0x29
    "00100000", --  657 - 0x291  :   32 - 0x20
    "00100000", --  658 - 0x292  :   32 - 0x20
    "00100000", --  659 - 0x293  :   32 - 0x20
    "00010011", --  660 - 0x294  :   19 - 0x13
    "00001101", --  661 - 0x295  :   13 - 0xd
    "00000010", --  662 - 0x296  :    2 - 0x2
    "00000001", --  663 - 0x297  :    1 - 0x1
    "00011111", --  664 - 0x298  :   31 - 0x1f -- plane 1
    "00011111", --  665 - 0x299  :   31 - 0x1f
    "00011111", --  666 - 0x29a  :   31 - 0x1f
    "00011111", --  667 - 0x29b  :   31 - 0x1f
    "00001100", --  668 - 0x29c  :   12 - 0xc
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000001", --  670 - 0x29e  :    1 - 0x1
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00100000", --  672 - 0x2a0  :   32 - 0x20 -- Background 0x2a
    "00100000", --  673 - 0x2a1  :   32 - 0x20
    "00100000", --  674 - 0x2a2  :   32 - 0x20
    "00100000", --  675 - 0x2a3  :   32 - 0x20
    "00010011", --  676 - 0x2a4  :   19 - 0x13
    "00001101", --  677 - 0x2a5  :   13 - 0xd
    "00000001", --  678 - 0x2a6  :    1 - 0x1
    "00000001", --  679 - 0x2a7  :    1 - 0x1
    "00011111", --  680 - 0x2a8  :   31 - 0x1f -- plane 1
    "00011111", --  681 - 0x2a9  :   31 - 0x1f
    "00011111", --  682 - 0x2aa  :   31 - 0x1f
    "00011111", --  683 - 0x2ab  :   31 - 0x1f
    "00001100", --  684 - 0x2ac  :   12 - 0xc
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "00000000", --  686 - 0x2ae  :    0 - 0x0
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "00000000", --  688 - 0x2b0  :    0 - 0x0 -- Background 0x2b
    "00000000", --  689 - 0x2b1  :    0 - 0x0
    "00000000", --  690 - 0x2b2  :    0 - 0x0
    "00000000", --  691 - 0x2b3  :    0 - 0x0
    "00000000", --  692 - 0x2b4  :    0 - 0x0
    "00000000", --  693 - 0x2b5  :    0 - 0x0
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "00000000", --  696 - 0x2b8  :    0 - 0x0 -- plane 1
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Background 0x2c
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "00000000", --  707 - 0x2c3  :    0 - 0x0
    "00000000", --  708 - 0x2c4  :    0 - 0x0
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0 -- plane 1
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00111100", --  720 - 0x2d0  :   60 - 0x3c -- Background 0x2d
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "10000001", --  722 - 0x2d2  :  129 - 0x81
    "10011001", --  723 - 0x2d3  :  153 - 0x99
    "10011001", --  724 - 0x2d4  :  153 - 0x99
    "10000001", --  725 - 0x2d5  :  129 - 0x81
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00111100", --  727 - 0x2d7  :   60 - 0x3c
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- plane 1
    "01111110", --  729 - 0x2d9  :  126 - 0x7e
    "01000010", --  730 - 0x2da  :   66 - 0x42
    "01000010", --  731 - 0x2db  :   66 - 0x42
    "01000010", --  732 - 0x2dc  :   66 - 0x42
    "01000010", --  733 - 0x2dd  :   66 - 0x42
    "01111110", --  734 - 0x2de  :  126 - 0x7e
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Background 0x2e
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- plane 1
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "10011111", --  752 - 0x2f0  :  159 - 0x9f -- Background 0x2f
    "10011110", --  753 - 0x2f1  :  158 - 0x9e
    "10011100", --  754 - 0x2f2  :  156 - 0x9c
    "00011000", --  755 - 0x2f3  :   24 - 0x18
    "00111000", --  756 - 0x2f4  :   56 - 0x38
    "11111100", --  757 - 0x2f5  :  252 - 0xfc
    "11111100", --  758 - 0x2f6  :  252 - 0xfc
    "11111100", --  759 - 0x2f7  :  252 - 0xfc
    "01100110", --  760 - 0x2f8  :  102 - 0x66 -- plane 1
    "01100000", --  761 - 0x2f9  :   96 - 0x60
    "01101000", --  762 - 0x2fa  :  104 - 0x68
    "11100000", --  763 - 0x2fb  :  224 - 0xe0
    "11000000", --  764 - 0x2fc  :  192 - 0xc0
    "00010000", --  765 - 0x2fd  :   16 - 0x10
    "00101000", --  766 - 0x2fe  :   40 - 0x28
    "01010000", --  767 - 0x2ff  :   80 - 0x50
    "01111111", --  768 - 0x300  :  127 - 0x7f -- Background 0x30
    "01111110", --  769 - 0x301  :  126 - 0x7e
    "11111100", --  770 - 0x302  :  252 - 0xfc
    "00111000", --  771 - 0x303  :   56 - 0x38
    "00111000", --  772 - 0x304  :   56 - 0x38
    "00000100", --  773 - 0x305  :    4 - 0x4
    "10000100", --  774 - 0x306  :  132 - 0x84
    "11111100", --  775 - 0x307  :  252 - 0xfc
    "11110110", --  776 - 0x308  :  246 - 0xf6 -- plane 1
    "11110000", --  777 - 0x309  :  240 - 0xf0
    "00111000", --  778 - 0x30a  :   56 - 0x38
    "11010000", --  779 - 0x30b  :  208 - 0xd0
    "11000000", --  780 - 0x30c  :  192 - 0xc0
    "11111000", --  781 - 0x30d  :  248 - 0xf8
    "01111000", --  782 - 0x30e  :  120 - 0x78
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "01111111", --  784 - 0x310  :  127 - 0x7f -- Background 0x31
    "01111110", --  785 - 0x311  :  126 - 0x7e
    "11111100", --  786 - 0x312  :  252 - 0xfc
    "00111000", --  787 - 0x313  :   56 - 0x38
    "00111000", --  788 - 0x314  :   56 - 0x38
    "00011100", --  789 - 0x315  :   28 - 0x1c
    "10000100", --  790 - 0x316  :  132 - 0x84
    "11000100", --  791 - 0x317  :  196 - 0xc4
    "11110110", --  792 - 0x318  :  246 - 0xf6 -- plane 1
    "11110000", --  793 - 0x319  :  240 - 0xf0
    "00111000", --  794 - 0x31a  :   56 - 0x38
    "11010000", --  795 - 0x31b  :  208 - 0xd0
    "11000000", --  796 - 0x31c  :  192 - 0xc0
    "11100000", --  797 - 0x31d  :  224 - 0xe0
    "01111000", --  798 - 0x31e  :  120 - 0x78
    "00111000", --  799 - 0x31f  :   56 - 0x38
    "01111111", --  800 - 0x320  :  127 - 0x7f -- Background 0x32
    "01111110", --  801 - 0x321  :  126 - 0x7e
    "11111100", --  802 - 0x322  :  252 - 0xfc
    "00111000", --  803 - 0x323  :   56 - 0x38
    "00100100", --  804 - 0x324  :   36 - 0x24
    "00000100", --  805 - 0x325  :    4 - 0x4
    "10011100", --  806 - 0x326  :  156 - 0x9c
    "11111100", --  807 - 0x327  :  252 - 0xfc
    "11110110", --  808 - 0x328  :  246 - 0xf6 -- plane 1
    "11110000", --  809 - 0x329  :  240 - 0xf0
    "00111000", --  810 - 0x32a  :   56 - 0x38
    "11000000", --  811 - 0x32b  :  192 - 0xc0
    "11011000", --  812 - 0x32c  :  216 - 0xd8
    "11111000", --  813 - 0x32d  :  248 - 0xf8
    "01100000", --  814 - 0x32e  :   96 - 0x60
    "00010000", --  815 - 0x32f  :   16 - 0x10
    "00100011", --  816 - 0x330  :   35 - 0x23 -- Background 0x33
    "00100011", --  817 - 0x331  :   35 - 0x23
    "00100001", --  818 - 0x332  :   33 - 0x21
    "00100000", --  819 - 0x333  :   32 - 0x20
    "00010011", --  820 - 0x334  :   19 - 0x13
    "00001101", --  821 - 0x335  :   13 - 0xd
    "00000001", --  822 - 0x336  :    1 - 0x1
    "00000001", --  823 - 0x337  :    1 - 0x1
    "00011100", --  824 - 0x338  :   28 - 0x1c -- plane 1
    "00011100", --  825 - 0x339  :   28 - 0x1c
    "00011110", --  826 - 0x33a  :   30 - 0x1e
    "00011111", --  827 - 0x33b  :   31 - 0x1f
    "00001100", --  828 - 0x33c  :   12 - 0xc
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "11111100", --  832 - 0x340  :  252 - 0xfc -- Background 0x34
    "11111100", --  833 - 0x341  :  252 - 0xfc
    "11111100", --  834 - 0x342  :  252 - 0xfc
    "11111100", --  835 - 0x343  :  252 - 0xfc
    "10100100", --  836 - 0x344  :  164 - 0xa4
    "00100100", --  837 - 0x345  :   36 - 0x24
    "00010010", --  838 - 0x346  :   18 - 0x12
    "11101110", --  839 - 0x347  :  238 - 0xee
    "10000000", --  840 - 0x348  :  128 - 0x80 -- plane 1
    "01010000", --  841 - 0x349  :   80 - 0x50
    "10101000", --  842 - 0x34a  :  168 - 0xa8
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "01011000", --  844 - 0x34c  :   88 - 0x58
    "11011000", --  845 - 0x34d  :  216 - 0xd8
    "11101100", --  846 - 0x34e  :  236 - 0xec
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00100011", --  848 - 0x350  :   35 - 0x23 -- Background 0x35
    "00100011", --  849 - 0x351  :   35 - 0x23
    "00100001", --  850 - 0x352  :   33 - 0x21
    "00100000", --  851 - 0x353  :   32 - 0x20
    "00010011", --  852 - 0x354  :   19 - 0x13
    "00001110", --  853 - 0x355  :   14 - 0xe
    "00000010", --  854 - 0x356  :    2 - 0x2
    "00000001", --  855 - 0x357  :    1 - 0x1
    "00011100", --  856 - 0x358  :   28 - 0x1c -- plane 1
    "00011100", --  857 - 0x359  :   28 - 0x1c
    "00011110", --  858 - 0x35a  :   30 - 0x1e
    "00011111", --  859 - 0x35b  :   31 - 0x1f
    "00001100", --  860 - 0x35c  :   12 - 0xc
    "00000001", --  861 - 0x35d  :    1 - 0x1
    "00000001", --  862 - 0x35e  :    1 - 0x1
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "11111100", --  864 - 0x360  :  252 - 0xfc -- Background 0x36
    "11111100", --  865 - 0x361  :  252 - 0xfc
    "11111100", --  866 - 0x362  :  252 - 0xfc
    "11111100", --  867 - 0x363  :  252 - 0xfc
    "10100110", --  868 - 0x364  :  166 - 0xa6
    "00110001", --  869 - 0x365  :   49 - 0x31
    "01001001", --  870 - 0x366  :   73 - 0x49
    "11000110", --  871 - 0x367  :  198 - 0xc6
    "10101000", --  872 - 0x368  :  168 - 0xa8 -- plane 1
    "01010000", --  873 - 0x369  :   80 - 0x50
    "10101000", --  874 - 0x36a  :  168 - 0xa8
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "01011000", --  876 - 0x36c  :   88 - 0x58
    "11001110", --  877 - 0x36d  :  206 - 0xce
    "10000110", --  878 - 0x36e  :  134 - 0x86
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "11111100", --  880 - 0x370  :  252 - 0xfc -- Background 0x37
    "11111100", --  881 - 0x371  :  252 - 0xfc
    "11111100", --  882 - 0x372  :  252 - 0xfc
    "11111100", --  883 - 0x373  :  252 - 0xfc
    "10100100", --  884 - 0x374  :  164 - 0xa4
    "00100100", --  885 - 0x375  :   36 - 0x24
    "00010010", --  886 - 0x376  :   18 - 0x12
    "11101110", --  887 - 0x377  :  238 - 0xee
    "10101000", --  888 - 0x378  :  168 - 0xa8 -- plane 1
    "01010000", --  889 - 0x379  :   80 - 0x50
    "10101000", --  890 - 0x37a  :  168 - 0xa8
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "01011000", --  892 - 0x37c  :   88 - 0x58
    "11011000", --  893 - 0x37d  :  216 - 0xd8
    "11101100", --  894 - 0x37e  :  236 - 0xec
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Background 0x38
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0 -- plane 1
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Background 0x39
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0 -- plane 1
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Background 0x3a
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- plane 1
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Background 0x3b
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- plane 1
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Background 0x3c
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- plane 1
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Background 0x3d
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- plane 1
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Background 0x3e
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- plane 1
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Background 0x40
    "00111110", -- 1025 - 0x401  :   62 - 0x3e
    "01111111", -- 1026 - 0x402  :  127 - 0x7f
    "01111111", -- 1027 - 0x403  :  127 - 0x7f
    "01111111", -- 1028 - 0x404  :  127 - 0x7f
    "01111111", -- 1029 - 0x405  :  127 - 0x7f
    "01111111", -- 1030 - 0x406  :  127 - 0x7f
    "00111110", -- 1031 - 0x407  :   62 - 0x3e
    "00111100", -- 1032 - 0x408  :   60 - 0x3c -- plane 1
    "01111100", -- 1033 - 0x409  :  124 - 0x7c
    "11100110", -- 1034 - 0x40a  :  230 - 0xe6
    "11101110", -- 1035 - 0x40b  :  238 - 0xee
    "11110110", -- 1036 - 0x40c  :  246 - 0xf6
    "11100110", -- 1037 - 0x40d  :  230 - 0xe6
    "00111100", -- 1038 - 0x40e  :   60 - 0x3c
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Background 0x41
    "00111100", -- 1041 - 0x411  :   60 - 0x3c
    "00011100", -- 1042 - 0x412  :   28 - 0x1c
    "00011100", -- 1043 - 0x413  :   28 - 0x1c
    "00011100", -- 1044 - 0x414  :   28 - 0x1c
    "00011100", -- 1045 - 0x415  :   28 - 0x1c
    "00011100", -- 1046 - 0x416  :   28 - 0x1c
    "00011100", -- 1047 - 0x417  :   28 - 0x1c
    "00111000", -- 1048 - 0x418  :   56 - 0x38 -- plane 1
    "01111000", -- 1049 - 0x419  :  120 - 0x78
    "00111000", -- 1050 - 0x41a  :   56 - 0x38
    "00111000", -- 1051 - 0x41b  :   56 - 0x38
    "00111000", -- 1052 - 0x41c  :   56 - 0x38
    "00111000", -- 1053 - 0x41d  :   56 - 0x38
    "00111000", -- 1054 - 0x41e  :   56 - 0x38
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- Background 0x42
    "01111100", -- 1057 - 0x421  :  124 - 0x7c
    "01111111", -- 1058 - 0x422  :  127 - 0x7f
    "01100111", -- 1059 - 0x423  :  103 - 0x67
    "00111111", -- 1060 - 0x424  :   63 - 0x3f
    "01111110", -- 1061 - 0x425  :  126 - 0x7e
    "01111111", -- 1062 - 0x426  :  127 - 0x7f
    "01111111", -- 1063 - 0x427  :  127 - 0x7f
    "01111100", -- 1064 - 0x428  :  124 - 0x7c -- plane 1
    "11111110", -- 1065 - 0x429  :  254 - 0xfe
    "11100110", -- 1066 - 0x42a  :  230 - 0xe6
    "00011110", -- 1067 - 0x42b  :   30 - 0x1e
    "01111100", -- 1068 - 0x42c  :  124 - 0x7c
    "11100000", -- 1069 - 0x42d  :  224 - 0xe0
    "11111110", -- 1070 - 0x42e  :  254 - 0xfe
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Background 0x43
    "01111110", -- 1073 - 0x431  :  126 - 0x7e
    "01111111", -- 1074 - 0x432  :  127 - 0x7f
    "01111111", -- 1075 - 0x433  :  127 - 0x7f
    "00011111", -- 1076 - 0x434  :   31 - 0x1f
    "01110111", -- 1077 - 0x435  :  119 - 0x77
    "01111111", -- 1078 - 0x436  :  127 - 0x7f
    "01111110", -- 1079 - 0x437  :  126 - 0x7e
    "01111100", -- 1080 - 0x438  :  124 - 0x7c -- plane 1
    "11111100", -- 1081 - 0x439  :  252 - 0xfc
    "11100110", -- 1082 - 0x43a  :  230 - 0xe6
    "00011100", -- 1083 - 0x43b  :   28 - 0x1c
    "01100110", -- 1084 - 0x43c  :  102 - 0x66
    "11101110", -- 1085 - 0x43d  :  238 - 0xee
    "11111100", -- 1086 - 0x43e  :  252 - 0xfc
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Background 0x44
    "00001110", -- 1089 - 0x441  :   14 - 0xe
    "00011110", -- 1090 - 0x442  :   30 - 0x1e
    "00111110", -- 1091 - 0x443  :   62 - 0x3e
    "01111110", -- 1092 - 0x444  :  126 - 0x7e
    "01111111", -- 1093 - 0x445  :  127 - 0x7f
    "01111110", -- 1094 - 0x446  :  126 - 0x7e
    "00001100", -- 1095 - 0x447  :   12 - 0xc
    "00001100", -- 1096 - 0x448  :   12 - 0xc -- plane 1
    "00011100", -- 1097 - 0x449  :   28 - 0x1c
    "00111100", -- 1098 - 0x44a  :   60 - 0x3c
    "01111100", -- 1099 - 0x44b  :  124 - 0x7c
    "11101100", -- 1100 - 0x44c  :  236 - 0xec
    "11111110", -- 1101 - 0x44d  :  254 - 0xfe
    "00001100", -- 1102 - 0x44e  :   12 - 0xc
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Background 0x45
    "01111111", -- 1105 - 0x451  :  127 - 0x7f
    "01111111", -- 1106 - 0x452  :  127 - 0x7f
    "01111111", -- 1107 - 0x453  :  127 - 0x7f
    "01111111", -- 1108 - 0x454  :  127 - 0x7f
    "01110111", -- 1109 - 0x455  :  119 - 0x77
    "01111111", -- 1110 - 0x456  :  127 - 0x7f
    "01111110", -- 1111 - 0x457  :  126 - 0x7e
    "11111110", -- 1112 - 0x458  :  254 - 0xfe -- plane 1
    "11111110", -- 1113 - 0x459  :  254 - 0xfe
    "11100000", -- 1114 - 0x45a  :  224 - 0xe0
    "11111110", -- 1115 - 0x45b  :  254 - 0xfe
    "00000110", -- 1116 - 0x45c  :    6 - 0x6
    "11101110", -- 1117 - 0x45d  :  238 - 0xee
    "11111100", -- 1118 - 0x45e  :  252 - 0xfc
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Background 0x46
    "00111110", -- 1121 - 0x461  :   62 - 0x3e
    "01111110", -- 1122 - 0x462  :  126 - 0x7e
    "01111111", -- 1123 - 0x463  :  127 - 0x7f
    "01111111", -- 1124 - 0x464  :  127 - 0x7f
    "01110111", -- 1125 - 0x465  :  119 - 0x77
    "01111111", -- 1126 - 0x466  :  127 - 0x7f
    "00111110", -- 1127 - 0x467  :   62 - 0x3e
    "00111100", -- 1128 - 0x468  :   60 - 0x3c -- plane 1
    "01111100", -- 1129 - 0x469  :  124 - 0x7c
    "11100000", -- 1130 - 0x46a  :  224 - 0xe0
    "11111110", -- 1131 - 0x46b  :  254 - 0xfe
    "11100110", -- 1132 - 0x46c  :  230 - 0xe6
    "11101110", -- 1133 - 0x46d  :  238 - 0xee
    "00111100", -- 1134 - 0x46e  :   60 - 0x3c
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0 -- Background 0x47
    "01111110", -- 1137 - 0x471  :  126 - 0x7e
    "01111110", -- 1138 - 0x472  :  126 - 0x7e
    "00011110", -- 1139 - 0x473  :   30 - 0x1e
    "00011100", -- 1140 - 0x474  :   28 - 0x1c
    "00111100", -- 1141 - 0x475  :   60 - 0x3c
    "00111000", -- 1142 - 0x476  :   56 - 0x38
    "00111000", -- 1143 - 0x477  :   56 - 0x38
    "11111110", -- 1144 - 0x478  :  254 - 0xfe -- plane 1
    "11111100", -- 1145 - 0x479  :  252 - 0xfc
    "00001100", -- 1146 - 0x47a  :   12 - 0xc
    "00111000", -- 1147 - 0x47b  :   56 - 0x38
    "00111000", -- 1148 - 0x47c  :   56 - 0x38
    "01110000", -- 1149 - 0x47d  :  112 - 0x70
    "01110000", -- 1150 - 0x47e  :  112 - 0x70
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Background 0x48
    "00111110", -- 1153 - 0x481  :   62 - 0x3e
    "01111111", -- 1154 - 0x482  :  127 - 0x7f
    "01111111", -- 1155 - 0x483  :  127 - 0x7f
    "01111111", -- 1156 - 0x484  :  127 - 0x7f
    "01111111", -- 1157 - 0x485  :  127 - 0x7f
    "01111111", -- 1158 - 0x486  :  127 - 0x7f
    "00111110", -- 1159 - 0x487  :   62 - 0x3e
    "00111110", -- 1160 - 0x488  :   62 - 0x3e -- plane 1
    "01111100", -- 1161 - 0x489  :  124 - 0x7c
    "11100110", -- 1162 - 0x48a  :  230 - 0xe6
    "10111100", -- 1163 - 0x48b  :  188 - 0xbc
    "11100110", -- 1164 - 0x48c  :  230 - 0xe6
    "11101110", -- 1165 - 0x48d  :  238 - 0xee
    "00111100", -- 1166 - 0x48e  :   60 - 0x3c
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0 -- Background 0x49
    "00111110", -- 1169 - 0x491  :   62 - 0x3e
    "01111111", -- 1170 - 0x492  :  127 - 0x7f
    "01110111", -- 1171 - 0x493  :  119 - 0x77
    "01111111", -- 1172 - 0x494  :  127 - 0x7f
    "01111111", -- 1173 - 0x495  :  127 - 0x7f
    "00111111", -- 1174 - 0x496  :   63 - 0x3f
    "00111110", -- 1175 - 0x497  :   62 - 0x3e
    "00111100", -- 1176 - 0x498  :   60 - 0x3c -- plane 1
    "01111100", -- 1177 - 0x499  :  124 - 0x7c
    "11100110", -- 1178 - 0x49a  :  230 - 0xe6
    "11101110", -- 1179 - 0x49b  :  238 - 0xee
    "11111110", -- 1180 - 0x49c  :  254 - 0xfe
    "10000110", -- 1181 - 0x49d  :  134 - 0x86
    "01111100", -- 1182 - 0x49e  :  124 - 0x7c
    "01000000", -- 1183 - 0x49f  :   64 - 0x40
    "11111111", -- 1184 - 0x4a0  :  255 - 0xff -- Background 0x4a
    "10011001", -- 1185 - 0x4a1  :  153 - 0x99
    "10011001", -- 1186 - 0x4a2  :  153 - 0x99
    "10011001", -- 1187 - 0x4a3  :  153 - 0x99
    "10011001", -- 1188 - 0x4a4  :  153 - 0x99
    "10011001", -- 1189 - 0x4a5  :  153 - 0x99
    "10011001", -- 1190 - 0x4a6  :  153 - 0x99
    "11111111", -- 1191 - 0x4a7  :  255 - 0xff
    "11101110", -- 1192 - 0x4a8  :  238 - 0xee -- plane 1
    "11101110", -- 1193 - 0x4a9  :  238 - 0xee
    "11101110", -- 1194 - 0x4aa  :  238 - 0xee
    "11101110", -- 1195 - 0x4ab  :  238 - 0xee
    "11101110", -- 1196 - 0x4ac  :  238 - 0xee
    "11101110", -- 1197 - 0x4ad  :  238 - 0xee
    "11101110", -- 1198 - 0x4ae  :  238 - 0xee
    "10001000", -- 1199 - 0x4af  :  136 - 0x88
    "11110000", -- 1200 - 0x4b0  :  240 - 0xf0 -- Background 0x4b
    "10010000", -- 1201 - 0x4b1  :  144 - 0x90
    "10010000", -- 1202 - 0x4b2  :  144 - 0x90
    "10010000", -- 1203 - 0x4b3  :  144 - 0x90
    "10010000", -- 1204 - 0x4b4  :  144 - 0x90
    "10010000", -- 1205 - 0x4b5  :  144 - 0x90
    "10010000", -- 1206 - 0x4b6  :  144 - 0x90
    "11110000", -- 1207 - 0x4b7  :  240 - 0xf0
    "11100000", -- 1208 - 0x4b8  :  224 - 0xe0 -- plane 1
    "11100000", -- 1209 - 0x4b9  :  224 - 0xe0
    "11100000", -- 1210 - 0x4ba  :  224 - 0xe0
    "11100000", -- 1211 - 0x4bb  :  224 - 0xe0
    "11100000", -- 1212 - 0x4bc  :  224 - 0xe0
    "11100000", -- 1213 - 0x4bd  :  224 - 0xe0
    "11100000", -- 1214 - 0x4be  :  224 - 0xe0
    "10000000", -- 1215 - 0x4bf  :  128 - 0x80
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Background 0x4c
    "11111111", -- 1217 - 0x4c1  :  255 - 0xff
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111111", -- 1219 - 0x4c3  :  255 - 0xff
    "11111111", -- 1220 - 0x4c4  :  255 - 0xff
    "11111111", -- 1221 - 0x4c5  :  255 - 0xff
    "11111111", -- 1222 - 0x4c6  :  255 - 0xff
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0 -- plane 1
    "01111111", -- 1225 - 0x4c9  :  127 - 0x7f
    "01111111", -- 1226 - 0x4ca  :  127 - 0x7f
    "01111111", -- 1227 - 0x4cb  :  127 - 0x7f
    "01111111", -- 1228 - 0x4cc  :  127 - 0x7f
    "01111111", -- 1229 - 0x4cd  :  127 - 0x7f
    "01111111", -- 1230 - 0x4ce  :  127 - 0x7f
    "01111111", -- 1231 - 0x4cf  :  127 - 0x7f
    "11111111", -- 1232 - 0x4d0  :  255 - 0xff -- Background 0x4d
    "11111111", -- 1233 - 0x4d1  :  255 - 0xff
    "11111111", -- 1234 - 0x4d2  :  255 - 0xff
    "11111111", -- 1235 - 0x4d3  :  255 - 0xff
    "11111111", -- 1236 - 0x4d4  :  255 - 0xff
    "11111111", -- 1237 - 0x4d5  :  255 - 0xff
    "11111111", -- 1238 - 0x4d6  :  255 - 0xff
    "11111111", -- 1239 - 0x4d7  :  255 - 0xff
    "01111111", -- 1240 - 0x4d8  :  127 - 0x7f -- plane 1
    "01111111", -- 1241 - 0x4d9  :  127 - 0x7f
    "01111111", -- 1242 - 0x4da  :  127 - 0x7f
    "01111111", -- 1243 - 0x4db  :  127 - 0x7f
    "01111111", -- 1244 - 0x4dc  :  127 - 0x7f
    "01111111", -- 1245 - 0x4dd  :  127 - 0x7f
    "01111111", -- 1246 - 0x4de  :  127 - 0x7f
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "11111111", -- 1248 - 0x4e0  :  255 - 0xff -- Background 0x4e
    "11111111", -- 1249 - 0x4e1  :  255 - 0xff
    "11111111", -- 1250 - 0x4e2  :  255 - 0xff
    "11111111", -- 1251 - 0x4e3  :  255 - 0xff
    "11111111", -- 1252 - 0x4e4  :  255 - 0xff
    "11111111", -- 1253 - 0x4e5  :  255 - 0xff
    "11111111", -- 1254 - 0x4e6  :  255 - 0xff
    "11111111", -- 1255 - 0x4e7  :  255 - 0xff
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0 -- plane 1
    "11111110", -- 1257 - 0x4e9  :  254 - 0xfe
    "11111110", -- 1258 - 0x4ea  :  254 - 0xfe
    "11111110", -- 1259 - 0x4eb  :  254 - 0xfe
    "11111110", -- 1260 - 0x4ec  :  254 - 0xfe
    "11111110", -- 1261 - 0x4ed  :  254 - 0xfe
    "11111110", -- 1262 - 0x4ee  :  254 - 0xfe
    "11111110", -- 1263 - 0x4ef  :  254 - 0xfe
    "11111111", -- 1264 - 0x4f0  :  255 - 0xff -- Background 0x4f
    "11111111", -- 1265 - 0x4f1  :  255 - 0xff
    "11111111", -- 1266 - 0x4f2  :  255 - 0xff
    "11111111", -- 1267 - 0x4f3  :  255 - 0xff
    "11111111", -- 1268 - 0x4f4  :  255 - 0xff
    "11111111", -- 1269 - 0x4f5  :  255 - 0xff
    "11111111", -- 1270 - 0x4f6  :  255 - 0xff
    "11111111", -- 1271 - 0x4f7  :  255 - 0xff
    "11111110", -- 1272 - 0x4f8  :  254 - 0xfe -- plane 1
    "11111110", -- 1273 - 0x4f9  :  254 - 0xfe
    "11111110", -- 1274 - 0x4fa  :  254 - 0xfe
    "11111110", -- 1275 - 0x4fb  :  254 - 0xfe
    "11111110", -- 1276 - 0x4fc  :  254 - 0xfe
    "11111110", -- 1277 - 0x4fd  :  254 - 0xfe
    "11111110", -- 1278 - 0x4fe  :  254 - 0xfe
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00010000", -- 1280 - 0x500  :   16 - 0x10 -- Background 0x50
    "00101000", -- 1281 - 0x501  :   40 - 0x28
    "11101110", -- 1282 - 0x502  :  238 - 0xee
    "10000010", -- 1283 - 0x503  :  130 - 0x82
    "01000100", -- 1284 - 0x504  :   68 - 0x44
    "01000100", -- 1285 - 0x505  :   68 - 0x44
    "10010010", -- 1286 - 0x506  :  146 - 0x92
    "11101110", -- 1287 - 0x507  :  238 - 0xee
    "00000000", -- 1288 - 0x508  :    0 - 0x0 -- plane 1
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00000000", -- 1290 - 0x50a  :    0 - 0x0
    "00000000", -- 1291 - 0x50b  :    0 - 0x0
    "00000000", -- 1292 - 0x50c  :    0 - 0x0
    "00000000", -- 1293 - 0x50d  :    0 - 0x0
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00010000", -- 1296 - 0x510  :   16 - 0x10 -- Background 0x51
    "00101000", -- 1297 - 0x511  :   40 - 0x28
    "11101110", -- 1298 - 0x512  :  238 - 0xee
    "10000010", -- 1299 - 0x513  :  130 - 0x82
    "01000100", -- 1300 - 0x514  :   68 - 0x44
    "01000100", -- 1301 - 0x515  :   68 - 0x44
    "10010010", -- 1302 - 0x516  :  146 - 0x92
    "11101110", -- 1303 - 0x517  :  238 - 0xee
    "00000000", -- 1304 - 0x518  :    0 - 0x0 -- plane 1
    "00010000", -- 1305 - 0x519  :   16 - 0x10
    "00010000", -- 1306 - 0x51a  :   16 - 0x10
    "01111100", -- 1307 - 0x51b  :  124 - 0x7c
    "00111000", -- 1308 - 0x51c  :   56 - 0x38
    "00111000", -- 1309 - 0x51d  :   56 - 0x38
    "01101100", -- 1310 - 0x51e  :  108 - 0x6c
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00010000", -- 1312 - 0x520  :   16 - 0x10 -- Background 0x52
    "00111000", -- 1313 - 0x521  :   56 - 0x38
    "11111110", -- 1314 - 0x522  :  254 - 0xfe
    "11111110", -- 1315 - 0x523  :  254 - 0xfe
    "01111100", -- 1316 - 0x524  :  124 - 0x7c
    "01111100", -- 1317 - 0x525  :  124 - 0x7c
    "11111110", -- 1318 - 0x526  :  254 - 0xfe
    "11101110", -- 1319 - 0x527  :  238 - 0xee
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- plane 1
    "00010000", -- 1321 - 0x529  :   16 - 0x10
    "00010000", -- 1322 - 0x52a  :   16 - 0x10
    "01111100", -- 1323 - 0x52b  :  124 - 0x7c
    "00111000", -- 1324 - 0x52c  :   56 - 0x38
    "00111000", -- 1325 - 0x52d  :   56 - 0x38
    "01101100", -- 1326 - 0x52e  :  108 - 0x6c
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "11111111", -- 1328 - 0x530  :  255 - 0xff -- Background 0x53
    "11111111", -- 1329 - 0x531  :  255 - 0xff
    "11111111", -- 1330 - 0x532  :  255 - 0xff
    "11111111", -- 1331 - 0x533  :  255 - 0xff
    "11111111", -- 1332 - 0x534  :  255 - 0xff
    "11111111", -- 1333 - 0x535  :  255 - 0xff
    "11111111", -- 1334 - 0x536  :  255 - 0xff
    "11111111", -- 1335 - 0x537  :  255 - 0xff
    "00000000", -- 1336 - 0x538  :    0 - 0x0 -- plane 1
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "00000000", -- 1338 - 0x53a  :    0 - 0x0
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Background 0x54
    "00000000", -- 1345 - 0x541  :    0 - 0x0
    "00000000", -- 1346 - 0x542  :    0 - 0x0
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00000000", -- 1349 - 0x545  :    0 - 0x0
    "00000000", -- 1350 - 0x546  :    0 - 0x0
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "11111111", -- 1352 - 0x548  :  255 - 0xff -- plane 1
    "11111111", -- 1353 - 0x549  :  255 - 0xff
    "11111111", -- 1354 - 0x54a  :  255 - 0xff
    "11111111", -- 1355 - 0x54b  :  255 - 0xff
    "11111111", -- 1356 - 0x54c  :  255 - 0xff
    "11111111", -- 1357 - 0x54d  :  255 - 0xff
    "11111111", -- 1358 - 0x54e  :  255 - 0xff
    "11111111", -- 1359 - 0x54f  :  255 - 0xff
    "11111111", -- 1360 - 0x550  :  255 - 0xff -- Background 0x55
    "11111111", -- 1361 - 0x551  :  255 - 0xff
    "11111111", -- 1362 - 0x552  :  255 - 0xff
    "11111111", -- 1363 - 0x553  :  255 - 0xff
    "11111111", -- 1364 - 0x554  :  255 - 0xff
    "11111111", -- 1365 - 0x555  :  255 - 0xff
    "11111111", -- 1366 - 0x556  :  255 - 0xff
    "11111111", -- 1367 - 0x557  :  255 - 0xff
    "11111111", -- 1368 - 0x558  :  255 - 0xff -- plane 1
    "11111111", -- 1369 - 0x559  :  255 - 0xff
    "11111111", -- 1370 - 0x55a  :  255 - 0xff
    "11111111", -- 1371 - 0x55b  :  255 - 0xff
    "11111111", -- 1372 - 0x55c  :  255 - 0xff
    "11111111", -- 1373 - 0x55d  :  255 - 0xff
    "11111111", -- 1374 - 0x55e  :  255 - 0xff
    "11111111", -- 1375 - 0x55f  :  255 - 0xff
    "00101010", -- 1376 - 0x560  :   42 - 0x2a -- Background 0x56
    "01000101", -- 1377 - 0x561  :   69 - 0x45
    "00001000", -- 1378 - 0x562  :    8 - 0x8
    "00010101", -- 1379 - 0x563  :   21 - 0x15
    "00100000", -- 1380 - 0x564  :   32 - 0x20
    "01000101", -- 1381 - 0x565  :   69 - 0x45
    "10101000", -- 1382 - 0x566  :  168 - 0xa8
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000010", -- 1384 - 0x568  :    2 - 0x2 -- plane 1
    "00000101", -- 1385 - 0x569  :    5 - 0x5
    "10101010", -- 1386 - 0x56a  :  170 - 0xaa
    "01010001", -- 1387 - 0x56b  :   81 - 0x51
    "10101010", -- 1388 - 0x56c  :  170 - 0xaa
    "01010001", -- 1389 - 0x56d  :   81 - 0x51
    "10100010", -- 1390 - 0x56e  :  162 - 0xa2
    "00000100", -- 1391 - 0x56f  :    4 - 0x4
    "00001000", -- 1392 - 0x570  :    8 - 0x8 -- Background 0x57
    "01010101", -- 1393 - 0x571  :   85 - 0x55
    "10100000", -- 1394 - 0x572  :  160 - 0xa0
    "00010000", -- 1395 - 0x573  :   16 - 0x10
    "10000000", -- 1396 - 0x574  :  128 - 0x80
    "00010100", -- 1397 - 0x575  :   20 - 0x14
    "00100010", -- 1398 - 0x576  :   34 - 0x22
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00001000", -- 1400 - 0x578  :    8 - 0x8 -- plane 1
    "01010101", -- 1401 - 0x579  :   85 - 0x55
    "00101010", -- 1402 - 0x57a  :   42 - 0x2a
    "01010101", -- 1403 - 0x57b  :   85 - 0x55
    "00101010", -- 1404 - 0x57c  :   42 - 0x2a
    "01000101", -- 1405 - 0x57d  :   69 - 0x45
    "00001010", -- 1406 - 0x57e  :   10 - 0xa
    "00010000", -- 1407 - 0x57f  :   16 - 0x10
    "11111111", -- 1408 - 0x580  :  255 - 0xff -- Background 0x58
    "11010101", -- 1409 - 0x581  :  213 - 0xd5
    "10100000", -- 1410 - 0x582  :  160 - 0xa0
    "11010000", -- 1411 - 0x583  :  208 - 0xd0
    "10001111", -- 1412 - 0x584  :  143 - 0x8f
    "11001000", -- 1413 - 0x585  :  200 - 0xc8
    "10001000", -- 1414 - 0x586  :  136 - 0x88
    "11001000", -- 1415 - 0x587  :  200 - 0xc8
    "00000000", -- 1416 - 0x588  :    0 - 0x0 -- plane 1
    "00111111", -- 1417 - 0x589  :   63 - 0x3f
    "01011111", -- 1418 - 0x58a  :   95 - 0x5f
    "01101111", -- 1419 - 0x58b  :  111 - 0x6f
    "01110000", -- 1420 - 0x58c  :  112 - 0x70
    "01110111", -- 1421 - 0x58d  :  119 - 0x77
    "01110111", -- 1422 - 0x58e  :  119 - 0x77
    "01110111", -- 1423 - 0x58f  :  119 - 0x77
    "10001000", -- 1424 - 0x590  :  136 - 0x88 -- Background 0x59
    "11001000", -- 1425 - 0x591  :  200 - 0xc8
    "10001000", -- 1426 - 0x592  :  136 - 0x88
    "11001111", -- 1427 - 0x593  :  207 - 0xcf
    "10010000", -- 1428 - 0x594  :  144 - 0x90
    "11100000", -- 1429 - 0x595  :  224 - 0xe0
    "11101010", -- 1430 - 0x596  :  234 - 0xea
    "11111111", -- 1431 - 0x597  :  255 - 0xff
    "01110111", -- 1432 - 0x598  :  119 - 0x77 -- plane 1
    "01110111", -- 1433 - 0x599  :  119 - 0x77
    "01110111", -- 1434 - 0x59a  :  119 - 0x77
    "01110000", -- 1435 - 0x59b  :  112 - 0x70
    "01101111", -- 1436 - 0x59c  :  111 - 0x6f
    "01011111", -- 1437 - 0x59d  :   95 - 0x5f
    "00010101", -- 1438 - 0x59e  :   21 - 0x15
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "11111111", -- 1440 - 0x5a0  :  255 - 0xff -- Background 0x5a
    "01011011", -- 1441 - 0x5a1  :   91 - 0x5b
    "00000111", -- 1442 - 0x5a2  :    7 - 0x7
    "00001001", -- 1443 - 0x5a3  :    9 - 0x9
    "11110011", -- 1444 - 0x5a4  :  243 - 0xf3
    "00010001", -- 1445 - 0x5a5  :   17 - 0x11
    "00010011", -- 1446 - 0x5a6  :   19 - 0x13
    "00010001", -- 1447 - 0x5a7  :   17 - 0x11
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0 -- plane 1
    "11111100", -- 1449 - 0x5a9  :  252 - 0xfc
    "11111000", -- 1450 - 0x5aa  :  248 - 0xf8
    "11110110", -- 1451 - 0x5ab  :  246 - 0xf6
    "00001100", -- 1452 - 0x5ac  :   12 - 0xc
    "11101110", -- 1453 - 0x5ad  :  238 - 0xee
    "11101100", -- 1454 - 0x5ae  :  236 - 0xec
    "11101110", -- 1455 - 0x5af  :  238 - 0xee
    "00010011", -- 1456 - 0x5b0  :   19 - 0x13 -- Background 0x5b
    "00010001", -- 1457 - 0x5b1  :   17 - 0x11
    "00010011", -- 1458 - 0x5b2  :   19 - 0x13
    "11110001", -- 1459 - 0x5b3  :  241 - 0xf1
    "00001011", -- 1460 - 0x5b4  :   11 - 0xb
    "00000101", -- 1461 - 0x5b5  :    5 - 0x5
    "10101011", -- 1462 - 0x5b6  :  171 - 0xab
    "11111111", -- 1463 - 0x5b7  :  255 - 0xff
    "11101100", -- 1464 - 0x5b8  :  236 - 0xec -- plane 1
    "11101110", -- 1465 - 0x5b9  :  238 - 0xee
    "11101100", -- 1466 - 0x5ba  :  236 - 0xec
    "00001110", -- 1467 - 0x5bb  :   14 - 0xe
    "11110100", -- 1468 - 0x5bc  :  244 - 0xf4
    "11111010", -- 1469 - 0x5bd  :  250 - 0xfa
    "01010100", -- 1470 - 0x5be  :   84 - 0x54
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00011100", -- 1472 - 0x5c0  :   28 - 0x1c -- Background 0x5c
    "00100010", -- 1473 - 0x5c1  :   34 - 0x22
    "01000001", -- 1474 - 0x5c2  :   65 - 0x41
    "01000001", -- 1475 - 0x5c3  :   65 - 0x41
    "01000001", -- 1476 - 0x5c4  :   65 - 0x41
    "00100010", -- 1477 - 0x5c5  :   34 - 0x22
    "00100010", -- 1478 - 0x5c6  :   34 - 0x22
    "00011100", -- 1479 - 0x5c7  :   28 - 0x1c
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0 -- plane 1
    "00011100", -- 1481 - 0x5c9  :   28 - 0x1c
    "00111110", -- 1482 - 0x5ca  :   62 - 0x3e
    "00111110", -- 1483 - 0x5cb  :   62 - 0x3e
    "00111110", -- 1484 - 0x5cc  :   62 - 0x3e
    "00011100", -- 1485 - 0x5cd  :   28 - 0x1c
    "00011100", -- 1486 - 0x5ce  :   28 - 0x1c
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00001000", -- 1488 - 0x5d0  :    8 - 0x8 -- Background 0x5d
    "00010000", -- 1489 - 0x5d1  :   16 - 0x10
    "00010000", -- 1490 - 0x5d2  :   16 - 0x10
    "00001000", -- 1491 - 0x5d3  :    8 - 0x8
    "00000100", -- 1492 - 0x5d4  :    4 - 0x4
    "00000100", -- 1493 - 0x5d5  :    4 - 0x4
    "00001000", -- 1494 - 0x5d6  :    8 - 0x8
    "00010000", -- 1495 - 0x5d7  :   16 - 0x10
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0 -- plane 1
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00110110", -- 1504 - 0x5e0  :   54 - 0x36 -- Background 0x5e
    "01101011", -- 1505 - 0x5e1  :  107 - 0x6b
    "01001001", -- 1506 - 0x5e2  :   73 - 0x49
    "01000001", -- 1507 - 0x5e3  :   65 - 0x41
    "01000001", -- 1508 - 0x5e4  :   65 - 0x41
    "00100010", -- 1509 - 0x5e5  :   34 - 0x22
    "00010100", -- 1510 - 0x5e6  :   20 - 0x14
    "00001000", -- 1511 - 0x5e7  :    8 - 0x8
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- plane 1
    "00010100", -- 1513 - 0x5e9  :   20 - 0x14
    "00110110", -- 1514 - 0x5ea  :   54 - 0x36
    "00111110", -- 1515 - 0x5eb  :   62 - 0x3e
    "00111110", -- 1516 - 0x5ec  :   62 - 0x3e
    "00011100", -- 1517 - 0x5ed  :   28 - 0x1c
    "00001000", -- 1518 - 0x5ee  :    8 - 0x8
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00111110", -- 1520 - 0x5f0  :   62 - 0x3e -- Background 0x5f
    "01101011", -- 1521 - 0x5f1  :  107 - 0x6b
    "00100010", -- 1522 - 0x5f2  :   34 - 0x22
    "01100011", -- 1523 - 0x5f3  :   99 - 0x63
    "00100010", -- 1524 - 0x5f4  :   34 - 0x22
    "01100011", -- 1525 - 0x5f5  :   99 - 0x63
    "00100010", -- 1526 - 0x5f6  :   34 - 0x22
    "01111111", -- 1527 - 0x5f7  :  127 - 0x7f
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- plane 1
    "00010100", -- 1529 - 0x5f9  :   20 - 0x14
    "00011100", -- 1530 - 0x5fa  :   28 - 0x1c
    "00011100", -- 1531 - 0x5fb  :   28 - 0x1c
    "00011100", -- 1532 - 0x5fc  :   28 - 0x1c
    "00011100", -- 1533 - 0x5fd  :   28 - 0x1c
    "00011100", -- 1534 - 0x5fe  :   28 - 0x1c
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "11111111", -- 1536 - 0x600  :  255 - 0xff -- Background 0x60
    "11111111", -- 1537 - 0x601  :  255 - 0xff
    "11111111", -- 1538 - 0x602  :  255 - 0xff
    "11111111", -- 1539 - 0x603  :  255 - 0xff
    "11010101", -- 1540 - 0x604  :  213 - 0xd5
    "10101010", -- 1541 - 0x605  :  170 - 0xaa
    "11010101", -- 1542 - 0x606  :  213 - 0xd5
    "11111111", -- 1543 - 0x607  :  255 - 0xff
    "00000000", -- 1544 - 0x608  :    0 - 0x0 -- plane 1
    "01111111", -- 1545 - 0x609  :  127 - 0x7f
    "01111111", -- 1546 - 0x60a  :  127 - 0x7f
    "01111111", -- 1547 - 0x60b  :  127 - 0x7f
    "01111111", -- 1548 - 0x60c  :  127 - 0x7f
    "01111111", -- 1549 - 0x60d  :  127 - 0x7f
    "00101010", -- 1550 - 0x60e  :   42 - 0x2a
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "11111111", -- 1552 - 0x610  :  255 - 0xff -- Background 0x61
    "11111111", -- 1553 - 0x611  :  255 - 0xff
    "11111111", -- 1554 - 0x612  :  255 - 0xff
    "11111111", -- 1555 - 0x613  :  255 - 0xff
    "01010101", -- 1556 - 0x614  :   85 - 0x55
    "10101010", -- 1557 - 0x615  :  170 - 0xaa
    "01010101", -- 1558 - 0x616  :   85 - 0x55
    "11111111", -- 1559 - 0x617  :  255 - 0xff
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- plane 1
    "11111111", -- 1561 - 0x619  :  255 - 0xff
    "11111111", -- 1562 - 0x61a  :  255 - 0xff
    "11111111", -- 1563 - 0x61b  :  255 - 0xff
    "11111111", -- 1564 - 0x61c  :  255 - 0xff
    "11111111", -- 1565 - 0x61d  :  255 - 0xff
    "10101010", -- 1566 - 0x61e  :  170 - 0xaa
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "11111111", -- 1568 - 0x620  :  255 - 0xff -- Background 0x62
    "11111111", -- 1569 - 0x621  :  255 - 0xff
    "11111111", -- 1570 - 0x622  :  255 - 0xff
    "11111111", -- 1571 - 0x623  :  255 - 0xff
    "01010101", -- 1572 - 0x624  :   85 - 0x55
    "10101011", -- 1573 - 0x625  :  171 - 0xab
    "01010101", -- 1574 - 0x626  :   85 - 0x55
    "11111111", -- 1575 - 0x627  :  255 - 0xff
    "00000000", -- 1576 - 0x628  :    0 - 0x0 -- plane 1
    "11111110", -- 1577 - 0x629  :  254 - 0xfe
    "11111110", -- 1578 - 0x62a  :  254 - 0xfe
    "11111110", -- 1579 - 0x62b  :  254 - 0xfe
    "11111110", -- 1580 - 0x62c  :  254 - 0xfe
    "11111110", -- 1581 - 0x62d  :  254 - 0xfe
    "10101010", -- 1582 - 0x62e  :  170 - 0xaa
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "00000000", -- 1584 - 0x630  :    0 - 0x0 -- Background 0x63
    "00000000", -- 1585 - 0x631  :    0 - 0x0
    "00000000", -- 1586 - 0x632  :    0 - 0x0
    "00000000", -- 1587 - 0x633  :    0 - 0x0
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "00000000", -- 1589 - 0x635  :    0 - 0x0
    "00000000", -- 1590 - 0x636  :    0 - 0x0
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00000000", -- 1592 - 0x638  :    0 - 0x0 -- plane 1
    "00000000", -- 1593 - 0x639  :    0 - 0x0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "00000000", -- 1596 - 0x63c  :    0 - 0x0
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000001", -- 1600 - 0x640  :    1 - 0x1 -- Background 0x64
    "00000001", -- 1601 - 0x641  :    1 - 0x1
    "00000011", -- 1602 - 0x642  :    3 - 0x3
    "00000011", -- 1603 - 0x643  :    3 - 0x3
    "00000110", -- 1604 - 0x644  :    6 - 0x6
    "00000110", -- 1605 - 0x645  :    6 - 0x6
    "00001100", -- 1606 - 0x646  :   12 - 0xc
    "00001100", -- 1607 - 0x647  :   12 - 0xc
    "00000000", -- 1608 - 0x648  :    0 - 0x0 -- plane 1
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000001", -- 1610 - 0x64a  :    1 - 0x1
    "00000001", -- 1611 - 0x64b  :    1 - 0x1
    "00000011", -- 1612 - 0x64c  :    3 - 0x3
    "00000011", -- 1613 - 0x64d  :    3 - 0x3
    "00000111", -- 1614 - 0x64e  :    7 - 0x7
    "00000111", -- 1615 - 0x64f  :    7 - 0x7
    "00011000", -- 1616 - 0x650  :   24 - 0x18 -- Background 0x65
    "00011000", -- 1617 - 0x651  :   24 - 0x18
    "00110000", -- 1618 - 0x652  :   48 - 0x30
    "00110000", -- 1619 - 0x653  :   48 - 0x30
    "01100000", -- 1620 - 0x654  :   96 - 0x60
    "01100000", -- 1621 - 0x655  :   96 - 0x60
    "11101010", -- 1622 - 0x656  :  234 - 0xea
    "11111111", -- 1623 - 0x657  :  255 - 0xff
    "00001111", -- 1624 - 0x658  :   15 - 0xf -- plane 1
    "00001111", -- 1625 - 0x659  :   15 - 0xf
    "00011111", -- 1626 - 0x65a  :   31 - 0x1f
    "00011111", -- 1627 - 0x65b  :   31 - 0x1f
    "00111111", -- 1628 - 0x65c  :   63 - 0x3f
    "00111111", -- 1629 - 0x65d  :   63 - 0x3f
    "01010101", -- 1630 - 0x65e  :   85 - 0x55
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "10000000", -- 1632 - 0x660  :  128 - 0x80 -- Background 0x66
    "10000000", -- 1633 - 0x661  :  128 - 0x80
    "11000000", -- 1634 - 0x662  :  192 - 0xc0
    "01000000", -- 1635 - 0x663  :   64 - 0x40
    "10100000", -- 1636 - 0x664  :  160 - 0xa0
    "01100000", -- 1637 - 0x665  :   96 - 0x60
    "00110000", -- 1638 - 0x666  :   48 - 0x30
    "00010000", -- 1639 - 0x667  :   16 - 0x10
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- plane 1
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "10000000", -- 1643 - 0x66b  :  128 - 0x80
    "01000000", -- 1644 - 0x66c  :   64 - 0x40
    "10000000", -- 1645 - 0x66d  :  128 - 0x80
    "11000000", -- 1646 - 0x66e  :  192 - 0xc0
    "11100000", -- 1647 - 0x66f  :  224 - 0xe0
    "00101000", -- 1648 - 0x670  :   40 - 0x28 -- Background 0x67
    "00011000", -- 1649 - 0x671  :   24 - 0x18
    "00001100", -- 1650 - 0x672  :   12 - 0xc
    "00010100", -- 1651 - 0x673  :   20 - 0x14
    "00001010", -- 1652 - 0x674  :   10 - 0xa
    "00000110", -- 1653 - 0x675  :    6 - 0x6
    "10101011", -- 1654 - 0x676  :  171 - 0xab
    "11111111", -- 1655 - 0x677  :  255 - 0xff
    "11010000", -- 1656 - 0x678  :  208 - 0xd0 -- plane 1
    "11100000", -- 1657 - 0x679  :  224 - 0xe0
    "11110000", -- 1658 - 0x67a  :  240 - 0xf0
    "11101000", -- 1659 - 0x67b  :  232 - 0xe8
    "11110100", -- 1660 - 0x67c  :  244 - 0xf4
    "11111000", -- 1661 - 0x67d  :  248 - 0xf8
    "01010100", -- 1662 - 0x67e  :   84 - 0x54
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Background 0x68
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- plane 1
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00000000", -- 1680 - 0x690  :    0 - 0x0 -- Background 0x69
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00000000", -- 1685 - 0x695  :    0 - 0x0
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00000000", -- 1688 - 0x698  :    0 - 0x0 -- plane 1
    "00000000", -- 1689 - 0x699  :    0 - 0x0
    "00000000", -- 1690 - 0x69a  :    0 - 0x0
    "00000000", -- 1691 - 0x69b  :    0 - 0x0
    "00000000", -- 1692 - 0x69c  :    0 - 0x0
    "00000000", -- 1693 - 0x69d  :    0 - 0x0
    "00000000", -- 1694 - 0x69e  :    0 - 0x0
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Background 0x6a
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1705 - 0x6a9  :    0 - 0x0
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Background 0x6b
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "00000000", -- 1715 - 0x6b3  :    0 - 0x0
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "00000000", -- 1720 - 0x6b8  :    0 - 0x0 -- plane 1
    "00000000", -- 1721 - 0x6b9  :    0 - 0x0
    "00000000", -- 1722 - 0x6ba  :    0 - 0x0
    "00000000", -- 1723 - 0x6bb  :    0 - 0x0
    "00000000", -- 1724 - 0x6bc  :    0 - 0x0
    "00000000", -- 1725 - 0x6bd  :    0 - 0x0
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Background 0x6c
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000000", -- 1734 - 0x6c6  :    0 - 0x0
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0 -- plane 1
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "00000000", -- 1738 - 0x6ca  :    0 - 0x0
    "00000000", -- 1739 - 0x6cb  :    0 - 0x0
    "00000000", -- 1740 - 0x6cc  :    0 - 0x0
    "00000000", -- 1741 - 0x6cd  :    0 - 0x0
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Background 0x6d
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0 -- plane 1
    "00000000", -- 1753 - 0x6d9  :    0 - 0x0
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "00000000", -- 1755 - 0x6db  :    0 - 0x0
    "00000000", -- 1756 - 0x6dc  :    0 - 0x0
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00000000", -- 1773 - 0x6ed  :    0 - 0x0
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0 -- Background 0x6f
    "00000000", -- 1777 - 0x6f1  :    0 - 0x0
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00000000", -- 1779 - 0x6f3  :    0 - 0x0
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "00000000", -- 1781 - 0x6f5  :    0 - 0x0
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "00000000", -- 1784 - 0x6f8  :    0 - 0x0 -- plane 1
    "00000000", -- 1785 - 0x6f9  :    0 - 0x0
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "00000000", -- 1787 - 0x6fb  :    0 - 0x0
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "00000000", -- 1789 - 0x6fd  :    0 - 0x0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Background 0x70
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0 -- plane 1
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0 -- Background 0x71
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000000", -- 1816 - 0x718  :    0 - 0x0 -- plane 1
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Background 0x72
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000000", -- 1828 - 0x724  :    0 - 0x0
    "00000000", -- 1829 - 0x725  :    0 - 0x0
    "00000000", -- 1830 - 0x726  :    0 - 0x0
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- plane 1
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "00000000", -- 1840 - 0x730  :    0 - 0x0 -- Background 0x73
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "00000000", -- 1845 - 0x735  :    0 - 0x0
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0 -- plane 1
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Background 0x74
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0 -- plane 1
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Background 0x75
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- plane 1
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Background 0x76
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0 -- plane 1
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Background 0x77
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- plane 1
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Background 0x78
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- plane 1
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Background 0x79
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- plane 1
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Background 0x7a
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Background 0x7b
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- plane 1
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Background 0x7c
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- plane 1
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Background 0x7d
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- plane 1
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- plane 1
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Background 0x7f
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- plane 1
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000", -- 2047 - 0x7ff  :    0 - 0x0
    "00000011", -- 2048 - 0x800  :    3 - 0x3 -- Background 0x80
    "00001111", -- 2049 - 0x801  :   15 - 0xf
    "00011100", -- 2050 - 0x802  :   28 - 0x1c
    "00110000", -- 2051 - 0x803  :   48 - 0x30
    "00100000", -- 2052 - 0x804  :   32 - 0x20
    "01000000", -- 2053 - 0x805  :   64 - 0x40
    "01000000", -- 2054 - 0x806  :   64 - 0x40
    "01111111", -- 2055 - 0x807  :  127 - 0x7f
    "00000000", -- 2056 - 0x808  :    0 - 0x0 -- plane 1
    "00000011", -- 2057 - 0x809  :    3 - 0x3
    "00001111", -- 2058 - 0x80a  :   15 - 0xf
    "00011111", -- 2059 - 0x80b  :   31 - 0x1f
    "00011111", -- 2060 - 0x80c  :   31 - 0x1f
    "00111111", -- 2061 - 0x80d  :   63 - 0x3f
    "00111111", -- 2062 - 0x80e  :   63 - 0x3f
    "00000000", -- 2063 - 0x80f  :    0 - 0x0
    "00000001", -- 2064 - 0x810  :    1 - 0x1 -- Background 0x81
    "00000001", -- 2065 - 0x811  :    1 - 0x1
    "00000001", -- 2066 - 0x812  :    1 - 0x1
    "00000001", -- 2067 - 0x813  :    1 - 0x1
    "00000001", -- 2068 - 0x814  :    1 - 0x1
    "00000001", -- 2069 - 0x815  :    1 - 0x1
    "00000011", -- 2070 - 0x816  :    3 - 0x3
    "00000011", -- 2071 - 0x817  :    3 - 0x3
    "00000000", -- 2072 - 0x818  :    0 - 0x0 -- plane 1
    "00000000", -- 2073 - 0x819  :    0 - 0x0
    "00000000", -- 2074 - 0x81a  :    0 - 0x0
    "00000000", -- 2075 - 0x81b  :    0 - 0x0
    "00000000", -- 2076 - 0x81c  :    0 - 0x0
    "00000000", -- 2077 - 0x81d  :    0 - 0x0
    "00000000", -- 2078 - 0x81e  :    0 - 0x0
    "00000000", -- 2079 - 0x81f  :    0 - 0x0
    "11000000", -- 2080 - 0x820  :  192 - 0xc0 -- Background 0x82
    "11110000", -- 2081 - 0x821  :  240 - 0xf0
    "00111000", -- 2082 - 0x822  :   56 - 0x38
    "00001110", -- 2083 - 0x823  :   14 - 0xe
    "00011110", -- 2084 - 0x824  :   30 - 0x1e
    "00011110", -- 2085 - 0x825  :   30 - 0x1e
    "00000010", -- 2086 - 0x826  :    2 - 0x2
    "11111110", -- 2087 - 0x827  :  254 - 0xfe
    "00000000", -- 2088 - 0x828  :    0 - 0x0 -- plane 1
    "11000000", -- 2089 - 0x829  :  192 - 0xc0
    "11110000", -- 2090 - 0x82a  :  240 - 0xf0
    "11110000", -- 2091 - 0x82b  :  240 - 0xf0
    "11101100", -- 2092 - 0x82c  :  236 - 0xec
    "11100000", -- 2093 - 0x82d  :  224 - 0xe0
    "11111100", -- 2094 - 0x82e  :  252 - 0xfc
    "00000000", -- 2095 - 0x82f  :    0 - 0x0
    "10000000", -- 2096 - 0x830  :  128 - 0x80 -- Background 0x83
    "10000000", -- 2097 - 0x831  :  128 - 0x80
    "10000000", -- 2098 - 0x832  :  128 - 0x80
    "10000000", -- 2099 - 0x833  :  128 - 0x80
    "10000000", -- 2100 - 0x834  :  128 - 0x80
    "11100000", -- 2101 - 0x835  :  224 - 0xe0
    "00010000", -- 2102 - 0x836  :   16 - 0x10
    "11110000", -- 2103 - 0x837  :  240 - 0xf0
    "00000000", -- 2104 - 0x838  :    0 - 0x0 -- plane 1
    "00000000", -- 2105 - 0x839  :    0 - 0x0
    "00000000", -- 2106 - 0x83a  :    0 - 0x0
    "00000000", -- 2107 - 0x83b  :    0 - 0x0
    "00000000", -- 2108 - 0x83c  :    0 - 0x0
    "00000000", -- 2109 - 0x83d  :    0 - 0x0
    "11100000", -- 2110 - 0x83e  :  224 - 0xe0
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "00000011", -- 2112 - 0x840  :    3 - 0x3 -- Background 0x84
    "00001111", -- 2113 - 0x841  :   15 - 0xf
    "00011100", -- 2114 - 0x842  :   28 - 0x1c
    "00110000", -- 2115 - 0x843  :   48 - 0x30
    "00100000", -- 2116 - 0x844  :   32 - 0x20
    "01000000", -- 2117 - 0x845  :   64 - 0x40
    "01000000", -- 2118 - 0x846  :   64 - 0x40
    "01111111", -- 2119 - 0x847  :  127 - 0x7f
    "00000000", -- 2120 - 0x848  :    0 - 0x0 -- plane 1
    "00000011", -- 2121 - 0x849  :    3 - 0x3
    "00001111", -- 2122 - 0x84a  :   15 - 0xf
    "00011111", -- 2123 - 0x84b  :   31 - 0x1f
    "00011111", -- 2124 - 0x84c  :   31 - 0x1f
    "00111111", -- 2125 - 0x84d  :   63 - 0x3f
    "00111111", -- 2126 - 0x84e  :   63 - 0x3f
    "00000000", -- 2127 - 0x84f  :    0 - 0x0
    "00000011", -- 2128 - 0x850  :    3 - 0x3 -- Background 0x85
    "00000110", -- 2129 - 0x851  :    6 - 0x6
    "00000110", -- 2130 - 0x852  :    6 - 0x6
    "00011100", -- 2131 - 0x853  :   28 - 0x1c
    "00011000", -- 2132 - 0x854  :   24 - 0x18
    "00110110", -- 2133 - 0x855  :   54 - 0x36
    "00110001", -- 2134 - 0x856  :   49 - 0x31
    "00001111", -- 2135 - 0x857  :   15 - 0xf
    "00000000", -- 2136 - 0x858  :    0 - 0x0 -- plane 1
    "00000000", -- 2137 - 0x859  :    0 - 0x0
    "00000000", -- 2138 - 0x85a  :    0 - 0x0
    "00000000", -- 2139 - 0x85b  :    0 - 0x0
    "00000000", -- 2140 - 0x85c  :    0 - 0x0
    "00001000", -- 2141 - 0x85d  :    8 - 0x8
    "00001110", -- 2142 - 0x85e  :   14 - 0xe
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "11000000", -- 2144 - 0x860  :  192 - 0xc0 -- Background 0x86
    "11110000", -- 2145 - 0x861  :  240 - 0xf0
    "00111000", -- 2146 - 0x862  :   56 - 0x38
    "00001110", -- 2147 - 0x863  :   14 - 0xe
    "00011110", -- 2148 - 0x864  :   30 - 0x1e
    "00011110", -- 2149 - 0x865  :   30 - 0x1e
    "00000010", -- 2150 - 0x866  :    2 - 0x2
    "11111110", -- 2151 - 0x867  :  254 - 0xfe
    "00000000", -- 2152 - 0x868  :    0 - 0x0 -- plane 1
    "11000000", -- 2153 - 0x869  :  192 - 0xc0
    "11110000", -- 2154 - 0x86a  :  240 - 0xf0
    "11110000", -- 2155 - 0x86b  :  240 - 0xf0
    "11101100", -- 2156 - 0x86c  :  236 - 0xec
    "11100000", -- 2157 - 0x86d  :  224 - 0xe0
    "11111100", -- 2158 - 0x86e  :  252 - 0xfc
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "11000000", -- 2160 - 0x870  :  192 - 0xc0 -- Background 0x87
    "01100000", -- 2161 - 0x871  :   96 - 0x60
    "01100000", -- 2162 - 0x872  :   96 - 0x60
    "00110000", -- 2163 - 0x873  :   48 - 0x30
    "00111110", -- 2164 - 0x874  :   62 - 0x3e
    "00011001", -- 2165 - 0x875  :   25 - 0x19
    "00110011", -- 2166 - 0x876  :   51 - 0x33
    "00111100", -- 2167 - 0x877  :   60 - 0x3c
    "00000000", -- 2168 - 0x878  :    0 - 0x0 -- plane 1
    "00000000", -- 2169 - 0x879  :    0 - 0x0
    "00000000", -- 2170 - 0x87a  :    0 - 0x0
    "00000000", -- 2171 - 0x87b  :    0 - 0x0
    "00000000", -- 2172 - 0x87c  :    0 - 0x0
    "00000110", -- 2173 - 0x87d  :    6 - 0x6
    "00001100", -- 2174 - 0x87e  :   12 - 0xc
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "00000011", -- 2176 - 0x880  :    3 - 0x3 -- Background 0x88
    "00000111", -- 2177 - 0x881  :    7 - 0x7
    "00000111", -- 2178 - 0x882  :    7 - 0x7
    "00001011", -- 2179 - 0x883  :   11 - 0xb
    "00010000", -- 2180 - 0x884  :   16 - 0x10
    "01100000", -- 2181 - 0x885  :   96 - 0x60
    "11110000", -- 2182 - 0x886  :  240 - 0xf0
    "11110000", -- 2183 - 0x887  :  240 - 0xf0
    "00000000", -- 2184 - 0x888  :    0 - 0x0 -- plane 1
    "00000011", -- 2185 - 0x889  :    3 - 0x3
    "00000011", -- 2186 - 0x88a  :    3 - 0x3
    "00000100", -- 2187 - 0x88b  :    4 - 0x4
    "00001111", -- 2188 - 0x88c  :   15 - 0xf
    "00011111", -- 2189 - 0x88d  :   31 - 0x1f
    "01101111", -- 2190 - 0x88e  :  111 - 0x6f
    "01101111", -- 2191 - 0x88f  :  111 - 0x6f
    "11110000", -- 2192 - 0x890  :  240 - 0xf0 -- Background 0x89
    "11110000", -- 2193 - 0x891  :  240 - 0xf0
    "01100000", -- 2194 - 0x892  :   96 - 0x60
    "00010000", -- 2195 - 0x893  :   16 - 0x10
    "00001011", -- 2196 - 0x894  :   11 - 0xb
    "00000111", -- 2197 - 0x895  :    7 - 0x7
    "00000111", -- 2198 - 0x896  :    7 - 0x7
    "00000011", -- 2199 - 0x897  :    3 - 0x3
    "01101111", -- 2200 - 0x898  :  111 - 0x6f -- plane 1
    "01101111", -- 2201 - 0x899  :  111 - 0x6f
    "00011111", -- 2202 - 0x89a  :   31 - 0x1f
    "00001111", -- 2203 - 0x89b  :   15 - 0xf
    "00000100", -- 2204 - 0x89c  :    4 - 0x4
    "00000011", -- 2205 - 0x89d  :    3 - 0x3
    "00000011", -- 2206 - 0x89e  :    3 - 0x3
    "00000000", -- 2207 - 0x89f  :    0 - 0x0
    "00000000", -- 2208 - 0x8a0  :    0 - 0x0 -- Background 0x8a
    "00011100", -- 2209 - 0x8a1  :   28 - 0x1c
    "00111111", -- 2210 - 0x8a2  :   63 - 0x3f
    "01111000", -- 2211 - 0x8a3  :  120 - 0x78
    "01110000", -- 2212 - 0x8a4  :  112 - 0x70
    "01100000", -- 2213 - 0x8a5  :   96 - 0x60
    "00100000", -- 2214 - 0x8a6  :   32 - 0x20
    "00100000", -- 2215 - 0x8a7  :   32 - 0x20
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0 -- plane 1
    "00000000", -- 2217 - 0x8a9  :    0 - 0x0
    "00011000", -- 2218 - 0x8aa  :   24 - 0x18
    "00110111", -- 2219 - 0x8ab  :   55 - 0x37
    "00101111", -- 2220 - 0x8ac  :   47 - 0x2f
    "00011111", -- 2221 - 0x8ad  :   31 - 0x1f
    "00011111", -- 2222 - 0x8ae  :   31 - 0x1f
    "00011111", -- 2223 - 0x8af  :   31 - 0x1f
    "00100000", -- 2224 - 0x8b0  :   32 - 0x20 -- Background 0x8b
    "00100000", -- 2225 - 0x8b1  :   32 - 0x20
    "01100000", -- 2226 - 0x8b2  :   96 - 0x60
    "01110000", -- 2227 - 0x8b3  :  112 - 0x70
    "01111000", -- 2228 - 0x8b4  :  120 - 0x78
    "00111111", -- 2229 - 0x8b5  :   63 - 0x3f
    "00011100", -- 2230 - 0x8b6  :   28 - 0x1c
    "00000000", -- 2231 - 0x8b7  :    0 - 0x0
    "00011111", -- 2232 - 0x8b8  :   31 - 0x1f -- plane 1
    "00011111", -- 2233 - 0x8b9  :   31 - 0x1f
    "00011111", -- 2234 - 0x8ba  :   31 - 0x1f
    "00101111", -- 2235 - 0x8bb  :   47 - 0x2f
    "00110111", -- 2236 - 0x8bc  :   55 - 0x37
    "00011000", -- 2237 - 0x8bd  :   24 - 0x18
    "00000000", -- 2238 - 0x8be  :    0 - 0x0
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "00000011", -- 2240 - 0x8c0  :    3 - 0x3 -- Background 0x8c
    "00001100", -- 2241 - 0x8c1  :   12 - 0xc
    "00011110", -- 2242 - 0x8c2  :   30 - 0x1e
    "00100110", -- 2243 - 0x8c3  :   38 - 0x26
    "01000110", -- 2244 - 0x8c4  :   70 - 0x46
    "01100100", -- 2245 - 0x8c5  :  100 - 0x64
    "01110000", -- 2246 - 0x8c6  :  112 - 0x70
    "11110000", -- 2247 - 0x8c7  :  240 - 0xf0
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0 -- plane 1
    "00000011", -- 2249 - 0x8c9  :    3 - 0x3
    "00000001", -- 2250 - 0x8ca  :    1 - 0x1
    "00011001", -- 2251 - 0x8cb  :   25 - 0x19
    "00111001", -- 2252 - 0x8cc  :   57 - 0x39
    "00011011", -- 2253 - 0x8cd  :   27 - 0x1b
    "00001111", -- 2254 - 0x8ce  :   15 - 0xf
    "00001111", -- 2255 - 0x8cf  :   15 - 0xf
    "10101010", -- 2256 - 0x8d0  :  170 - 0xaa -- Background 0x8d
    "11111111", -- 2257 - 0x8d1  :  255 - 0xff
    "01111111", -- 2258 - 0x8d2  :  127 - 0x7f
    "00111001", -- 2259 - 0x8d3  :   57 - 0x39
    "00011001", -- 2260 - 0x8d4  :   25 - 0x19
    "00001011", -- 2261 - 0x8d5  :   11 - 0xb
    "00001000", -- 2262 - 0x8d6  :    8 - 0x8
    "00000111", -- 2263 - 0x8d7  :    7 - 0x7
    "01111111", -- 2264 - 0x8d8  :  127 - 0x7f -- plane 1
    "01111111", -- 2265 - 0x8d9  :  127 - 0x7f
    "00111111", -- 2266 - 0x8da  :   63 - 0x3f
    "00010111", -- 2267 - 0x8db  :   23 - 0x17
    "00000110", -- 2268 - 0x8dc  :    6 - 0x6
    "00000100", -- 2269 - 0x8dd  :    4 - 0x4
    "00000111", -- 2270 - 0x8de  :    7 - 0x7
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "11000000", -- 2272 - 0x8e0  :  192 - 0xc0 -- Background 0x8e
    "00110000", -- 2273 - 0x8e1  :   48 - 0x30
    "00001000", -- 2274 - 0x8e2  :    8 - 0x8
    "01000100", -- 2275 - 0x8e3  :   68 - 0x44
    "01100010", -- 2276 - 0x8e4  :   98 - 0x62
    "01100010", -- 2277 - 0x8e5  :   98 - 0x62
    "00000001", -- 2278 - 0x8e6  :    1 - 0x1
    "00111111", -- 2279 - 0x8e7  :   63 - 0x3f
    "00000000", -- 2280 - 0x8e8  :    0 - 0x0 -- plane 1
    "11000000", -- 2281 - 0x8e9  :  192 - 0xc0
    "11110000", -- 2282 - 0x8ea  :  240 - 0xf0
    "10111000", -- 2283 - 0x8eb  :  184 - 0xb8
    "10011100", -- 2284 - 0x8ec  :  156 - 0x9c
    "11111100", -- 2285 - 0x8ed  :  252 - 0xfc
    "11111110", -- 2286 - 0x8ee  :  254 - 0xfe
    "11000000", -- 2287 - 0x8ef  :  192 - 0xc0
    "10001011", -- 2288 - 0x8f0  :  139 - 0x8b -- Background 0x8f
    "11000001", -- 2289 - 0x8f1  :  193 - 0xc1
    "11111110", -- 2290 - 0x8f2  :  254 - 0xfe
    "11111100", -- 2291 - 0x8f3  :  252 - 0xfc
    "11110000", -- 2292 - 0x8f4  :  240 - 0xf0
    "11110000", -- 2293 - 0x8f5  :  240 - 0xf0
    "11111000", -- 2294 - 0x8f6  :  248 - 0xf8
    "11110000", -- 2295 - 0x8f7  :  240 - 0xf0
    "11111110", -- 2296 - 0x8f8  :  254 - 0xfe -- plane 1
    "11111110", -- 2297 - 0x8f9  :  254 - 0xfe
    "11111000", -- 2298 - 0x8fa  :  248 - 0xf8
    "11110000", -- 2299 - 0x8fb  :  240 - 0xf0
    "11000000", -- 2300 - 0x8fc  :  192 - 0xc0
    "00000000", -- 2301 - 0x8fd  :    0 - 0x0
    "00000000", -- 2302 - 0x8fe  :    0 - 0x0
    "10000000", -- 2303 - 0x8ff  :  128 - 0x80
    "00000011", -- 2304 - 0x900  :    3 - 0x3 -- Background 0x90
    "00001110", -- 2305 - 0x901  :   14 - 0xe
    "00010110", -- 2306 - 0x902  :   22 - 0x16
    "00100110", -- 2307 - 0x903  :   38 - 0x26
    "01100011", -- 2308 - 0x904  :   99 - 0x63
    "01110010", -- 2309 - 0x905  :  114 - 0x72
    "01110000", -- 2310 - 0x906  :  112 - 0x70
    "11010000", -- 2311 - 0x907  :  208 - 0xd0
    "00000000", -- 2312 - 0x908  :    0 - 0x0 -- plane 1
    "00000001", -- 2313 - 0x909  :    1 - 0x1
    "00001001", -- 2314 - 0x90a  :    9 - 0x9
    "00011001", -- 2315 - 0x90b  :   25 - 0x19
    "00011100", -- 2316 - 0x90c  :   28 - 0x1c
    "00001101", -- 2317 - 0x90d  :   13 - 0xd
    "00001111", -- 2318 - 0x90e  :   15 - 0xf
    "00101111", -- 2319 - 0x90f  :   47 - 0x2f
    "10101010", -- 2320 - 0x910  :  170 - 0xaa -- Background 0x91
    "11111111", -- 2321 - 0x911  :  255 - 0xff
    "01111111", -- 2322 - 0x912  :  127 - 0x7f
    "00111100", -- 2323 - 0x913  :   60 - 0x3c
    "00011100", -- 2324 - 0x914  :   28 - 0x1c
    "00000100", -- 2325 - 0x915  :    4 - 0x4
    "00000010", -- 2326 - 0x916  :    2 - 0x2
    "00000001", -- 2327 - 0x917  :    1 - 0x1
    "01111111", -- 2328 - 0x918  :  127 - 0x7f -- plane 1
    "01111111", -- 2329 - 0x919  :  127 - 0x7f
    "00111111", -- 2330 - 0x91a  :   63 - 0x3f
    "00011011", -- 2331 - 0x91b  :   27 - 0x1b
    "00000011", -- 2332 - 0x91c  :    3 - 0x3
    "00000011", -- 2333 - 0x91d  :    3 - 0x3
    "00000001", -- 2334 - 0x91e  :    1 - 0x1
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "11000000", -- 2336 - 0x920  :  192 - 0xc0 -- Background 0x92
    "00110000", -- 2337 - 0x921  :   48 - 0x30
    "00001000", -- 2338 - 0x922  :    8 - 0x8
    "00100100", -- 2339 - 0x923  :   36 - 0x24
    "00110010", -- 2340 - 0x924  :   50 - 0x32
    "00110010", -- 2341 - 0x925  :   50 - 0x32
    "00000001", -- 2342 - 0x926  :    1 - 0x1
    "00011111", -- 2343 - 0x927  :   31 - 0x1f
    "00000000", -- 2344 - 0x928  :    0 - 0x0 -- plane 1
    "11000000", -- 2345 - 0x929  :  192 - 0xc0
    "11110000", -- 2346 - 0x92a  :  240 - 0xf0
    "11011000", -- 2347 - 0x92b  :  216 - 0xd8
    "11001100", -- 2348 - 0x92c  :  204 - 0xcc
    "11111100", -- 2349 - 0x92d  :  252 - 0xfc
    "11111110", -- 2350 - 0x92e  :  254 - 0xfe
    "11100000", -- 2351 - 0x92f  :  224 - 0xe0
    "10001011", -- 2352 - 0x930  :  139 - 0x8b -- Background 0x93
    "11000001", -- 2353 - 0x931  :  193 - 0xc1
    "11111110", -- 2354 - 0x932  :  254 - 0xfe
    "11111100", -- 2355 - 0x933  :  252 - 0xfc
    "11110000", -- 2356 - 0x934  :  240 - 0xf0
    "11000000", -- 2357 - 0x935  :  192 - 0xc0
    "00100000", -- 2358 - 0x936  :   32 - 0x20
    "11100000", -- 2359 - 0x937  :  224 - 0xe0
    "11111110", -- 2360 - 0x938  :  254 - 0xfe -- plane 1
    "11111110", -- 2361 - 0x939  :  254 - 0xfe
    "11111000", -- 2362 - 0x93a  :  248 - 0xf8
    "01110000", -- 2363 - 0x93b  :  112 - 0x70
    "01000000", -- 2364 - 0x93c  :   64 - 0x40
    "00000000", -- 2365 - 0x93d  :    0 - 0x0
    "11000000", -- 2366 - 0x93e  :  192 - 0xc0
    "00100000", -- 2367 - 0x93f  :   32 - 0x20
    "00000011", -- 2368 - 0x940  :    3 - 0x3 -- Background 0x94
    "00001111", -- 2369 - 0x941  :   15 - 0xf
    "00010011", -- 2370 - 0x942  :   19 - 0x13
    "00110001", -- 2371 - 0x943  :   49 - 0x31
    "01111001", -- 2372 - 0x944  :  121 - 0x79
    "01011001", -- 2373 - 0x945  :   89 - 0x59
    "01001000", -- 2374 - 0x946  :   72 - 0x48
    "11001100", -- 2375 - 0x947  :  204 - 0xcc
    "00000000", -- 2376 - 0x948  :    0 - 0x0 -- plane 1
    "00000000", -- 2377 - 0x949  :    0 - 0x0
    "00001100", -- 2378 - 0x94a  :   12 - 0xc
    "00001110", -- 2379 - 0x94b  :   14 - 0xe
    "00000110", -- 2380 - 0x94c  :    6 - 0x6
    "00100110", -- 2381 - 0x94d  :   38 - 0x26
    "00110111", -- 2382 - 0x94e  :   55 - 0x37
    "00110011", -- 2383 - 0x94f  :   51 - 0x33
    "10010101", -- 2384 - 0x950  :  149 - 0x95 -- Background 0x95
    "11111111", -- 2385 - 0x951  :  255 - 0xff
    "01111111", -- 2386 - 0x952  :  127 - 0x7f
    "00111110", -- 2387 - 0x953  :   62 - 0x3e
    "00011111", -- 2388 - 0x954  :   31 - 0x1f
    "00001111", -- 2389 - 0x955  :   15 - 0xf
    "00001111", -- 2390 - 0x956  :   15 - 0xf
    "00000111", -- 2391 - 0x957  :    7 - 0x7
    "01111111", -- 2392 - 0x958  :  127 - 0x7f -- plane 1
    "01111111", -- 2393 - 0x959  :  127 - 0x7f
    "00111111", -- 2394 - 0x95a  :   63 - 0x3f
    "00011111", -- 2395 - 0x95b  :   31 - 0x1f
    "00001110", -- 2396 - 0x95c  :   14 - 0xe
    "00000000", -- 2397 - 0x95d  :    0 - 0x0
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "11000000", -- 2400 - 0x960  :  192 - 0xc0 -- Background 0x96
    "00110000", -- 2401 - 0x961  :   48 - 0x30
    "00001000", -- 2402 - 0x962  :    8 - 0x8
    "10010100", -- 2403 - 0x963  :  148 - 0x94
    "10011010", -- 2404 - 0x964  :  154 - 0x9a
    "00011010", -- 2405 - 0x965  :   26 - 0x1a
    "00000001", -- 2406 - 0x966  :    1 - 0x1
    "00001111", -- 2407 - 0x967  :   15 - 0xf
    "00000000", -- 2408 - 0x968  :    0 - 0x0 -- plane 1
    "11000000", -- 2409 - 0x969  :  192 - 0xc0
    "11110000", -- 2410 - 0x96a  :  240 - 0xf0
    "01101000", -- 2411 - 0x96b  :  104 - 0x68
    "01100100", -- 2412 - 0x96c  :  100 - 0x64
    "11111100", -- 2413 - 0x96d  :  252 - 0xfc
    "11111110", -- 2414 - 0x96e  :  254 - 0xfe
    "11110000", -- 2415 - 0x96f  :  240 - 0xf0
    "01000101", -- 2416 - 0x970  :   69 - 0x45 -- Background 0x97
    "11100001", -- 2417 - 0x971  :  225 - 0xe1
    "11111110", -- 2418 - 0x972  :  254 - 0xfe
    "01111100", -- 2419 - 0x973  :  124 - 0x7c
    "00110000", -- 2420 - 0x974  :   48 - 0x30
    "00110000", -- 2421 - 0x975  :   48 - 0x30
    "10001000", -- 2422 - 0x976  :  136 - 0x88
    "01111000", -- 2423 - 0x977  :  120 - 0x78
    "11111111", -- 2424 - 0x978  :  255 - 0xff -- plane 1
    "11111110", -- 2425 - 0x979  :  254 - 0xfe
    "11111100", -- 2426 - 0x97a  :  252 - 0xfc
    "10110000", -- 2427 - 0x97b  :  176 - 0xb0
    "11000000", -- 2428 - 0x97c  :  192 - 0xc0
    "11000000", -- 2429 - 0x97d  :  192 - 0xc0
    "01110000", -- 2430 - 0x97e  :  112 - 0x70
    "00001000", -- 2431 - 0x97f  :    8 - 0x8
    "00000001", -- 2432 - 0x980  :    1 - 0x1 -- Background 0x98
    "00000000", -- 2433 - 0x981  :    0 - 0x0
    "00000000", -- 2434 - 0x982  :    0 - 0x0
    "00000000", -- 2435 - 0x983  :    0 - 0x0
    "00000001", -- 2436 - 0x984  :    1 - 0x1
    "00000001", -- 2437 - 0x985  :    1 - 0x1
    "00000010", -- 2438 - 0x986  :    2 - 0x2
    "00000110", -- 2439 - 0x987  :    6 - 0x6
    "00000000", -- 2440 - 0x988  :    0 - 0x0 -- plane 1
    "00000001", -- 2441 - 0x989  :    1 - 0x1
    "00000000", -- 2442 - 0x98a  :    0 - 0x0
    "00000000", -- 2443 - 0x98b  :    0 - 0x0
    "00000000", -- 2444 - 0x98c  :    0 - 0x0
    "00000000", -- 2445 - 0x98d  :    0 - 0x0
    "00000001", -- 2446 - 0x98e  :    1 - 0x1
    "00000011", -- 2447 - 0x98f  :    3 - 0x3
    "01111000", -- 2448 - 0x990  :  120 - 0x78 -- Background 0x99
    "00101010", -- 2449 - 0x991  :   42 - 0x2a
    "01010100", -- 2450 - 0x992  :   84 - 0x54
    "00101001", -- 2451 - 0x993  :   41 - 0x29
    "00101111", -- 2452 - 0x994  :   47 - 0x2f
    "00110111", -- 2453 - 0x995  :   55 - 0x37
    "00000011", -- 2454 - 0x996  :    3 - 0x3
    "00000111", -- 2455 - 0x997  :    7 - 0x7
    "00000111", -- 2456 - 0x998  :    7 - 0x7 -- plane 1
    "00010111", -- 2457 - 0x999  :   23 - 0x17
    "00101111", -- 2458 - 0x99a  :   47 - 0x2f
    "00011110", -- 2459 - 0x99b  :   30 - 0x1e
    "00010001", -- 2460 - 0x99c  :   17 - 0x11
    "00000000", -- 2461 - 0x99d  :    0 - 0x0
    "00000001", -- 2462 - 0x99e  :    1 - 0x1
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "10110000", -- 2464 - 0x9a0  :  176 - 0xb0 -- Background 0x9a
    "11101000", -- 2465 - 0x9a1  :  232 - 0xe8
    "10001100", -- 2466 - 0x9a2  :  140 - 0x8c
    "10011110", -- 2467 - 0x9a3  :  158 - 0x9e
    "00011111", -- 2468 - 0x9a4  :   31 - 0x1f
    "00001111", -- 2469 - 0x9a5  :   15 - 0xf
    "10010110", -- 2470 - 0x9a6  :  150 - 0x96
    "00011100", -- 2471 - 0x9a7  :   28 - 0x1c
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0 -- plane 1
    "00010000", -- 2473 - 0x9a9  :   16 - 0x10
    "01111000", -- 2474 - 0x9aa  :  120 - 0x78
    "01110100", -- 2475 - 0x9ab  :  116 - 0x74
    "11111110", -- 2476 - 0x9ac  :  254 - 0xfe
    "11111000", -- 2477 - 0x9ad  :  248 - 0xf8
    "11111100", -- 2478 - 0x9ae  :  252 - 0xfc
    "11111000", -- 2479 - 0x9af  :  248 - 0xf8
    "00001100", -- 2480 - 0x9b0  :   12 - 0xc -- Background 0x9b
    "00111000", -- 2481 - 0x9b1  :   56 - 0x38
    "11101000", -- 2482 - 0x9b2  :  232 - 0xe8
    "11010000", -- 2483 - 0x9b3  :  208 - 0xd0
    "11100000", -- 2484 - 0x9b4  :  224 - 0xe0
    "10000000", -- 2485 - 0x9b5  :  128 - 0x80
    "00000000", -- 2486 - 0x9b6  :    0 - 0x0
    "10000000", -- 2487 - 0x9b7  :  128 - 0x80
    "11111000", -- 2488 - 0x9b8  :  248 - 0xf8 -- plane 1
    "11010000", -- 2489 - 0x9b9  :  208 - 0xd0
    "00110000", -- 2490 - 0x9ba  :   48 - 0x30
    "01100000", -- 2491 - 0x9bb  :   96 - 0x60
    "10000000", -- 2492 - 0x9bc  :  128 - 0x80
    "00000000", -- 2493 - 0x9bd  :    0 - 0x0
    "00000000", -- 2494 - 0x9be  :    0 - 0x0
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00000001", -- 2496 - 0x9c0  :    1 - 0x1 -- Background 0x9c
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000000", -- 2498 - 0x9c2  :    0 - 0x0
    "00000000", -- 2499 - 0x9c3  :    0 - 0x0
    "00000001", -- 2500 - 0x9c4  :    1 - 0x1
    "00000001", -- 2501 - 0x9c5  :    1 - 0x1
    "00000010", -- 2502 - 0x9c6  :    2 - 0x2
    "00000110", -- 2503 - 0x9c7  :    6 - 0x6
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0 -- plane 1
    "00000001", -- 2505 - 0x9c9  :    1 - 0x1
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000001", -- 2510 - 0x9ce  :    1 - 0x1
    "00000011", -- 2511 - 0x9cf  :    3 - 0x3
    "01111000", -- 2512 - 0x9d0  :  120 - 0x78 -- Background 0x9d
    "00101010", -- 2513 - 0x9d1  :   42 - 0x2a
    "01010100", -- 2514 - 0x9d2  :   84 - 0x54
    "00101001", -- 2515 - 0x9d3  :   41 - 0x29
    "00101111", -- 2516 - 0x9d4  :   47 - 0x2f
    "00111100", -- 2517 - 0x9d5  :   60 - 0x3c
    "00011110", -- 2518 - 0x9d6  :   30 - 0x1e
    "00000000", -- 2519 - 0x9d7  :    0 - 0x0
    "00000111", -- 2520 - 0x9d8  :    7 - 0x7 -- plane 1
    "00010111", -- 2521 - 0x9d9  :   23 - 0x17
    "00101111", -- 2522 - 0x9da  :   47 - 0x2f
    "00011110", -- 2523 - 0x9db  :   30 - 0x1e
    "00010000", -- 2524 - 0x9dc  :   16 - 0x10
    "00000100", -- 2525 - 0x9dd  :    4 - 0x4
    "00000000", -- 2526 - 0x9de  :    0 - 0x0
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "10110000", -- 2528 - 0x9e0  :  176 - 0xb0 -- Background 0x9e
    "11101000", -- 2529 - 0x9e1  :  232 - 0xe8
    "10001100", -- 2530 - 0x9e2  :  140 - 0x8c
    "10011110", -- 2531 - 0x9e3  :  158 - 0x9e
    "00011111", -- 2532 - 0x9e4  :   31 - 0x1f
    "00001111", -- 2533 - 0x9e5  :   15 - 0xf
    "10010110", -- 2534 - 0x9e6  :  150 - 0x96
    "00011100", -- 2535 - 0x9e7  :   28 - 0x1c
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0 -- plane 1
    "00010000", -- 2537 - 0x9e9  :   16 - 0x10
    "01111000", -- 2538 - 0x9ea  :  120 - 0x78
    "01110100", -- 2539 - 0x9eb  :  116 - 0x74
    "11111110", -- 2540 - 0x9ec  :  254 - 0xfe
    "11111000", -- 2541 - 0x9ed  :  248 - 0xf8
    "11111100", -- 2542 - 0x9ee  :  252 - 0xfc
    "11111000", -- 2543 - 0x9ef  :  248 - 0xf8
    "00001100", -- 2544 - 0x9f0  :   12 - 0xc -- Background 0x9f
    "00111000", -- 2545 - 0x9f1  :   56 - 0x38
    "11101000", -- 2546 - 0x9f2  :  232 - 0xe8
    "11110000", -- 2547 - 0x9f3  :  240 - 0xf0
    "11000000", -- 2548 - 0x9f4  :  192 - 0xc0
    "01110000", -- 2549 - 0x9f5  :  112 - 0x70
    "11000000", -- 2550 - 0x9f6  :  192 - 0xc0
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "11111000", -- 2552 - 0x9f8  :  248 - 0xf8 -- plane 1
    "11010000", -- 2553 - 0x9f9  :  208 - 0xd0
    "00110000", -- 2554 - 0x9fa  :   48 - 0x30
    "11000000", -- 2555 - 0x9fb  :  192 - 0xc0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00000011", -- 2560 - 0xa00  :    3 - 0x3 -- Background 0xa0
    "00001111", -- 2561 - 0xa01  :   15 - 0xf
    "00011100", -- 2562 - 0xa02  :   28 - 0x1c
    "00110000", -- 2563 - 0xa03  :   48 - 0x30
    "01100000", -- 2564 - 0xa04  :   96 - 0x60
    "01100000", -- 2565 - 0xa05  :   96 - 0x60
    "11000000", -- 2566 - 0xa06  :  192 - 0xc0
    "11000000", -- 2567 - 0xa07  :  192 - 0xc0
    "00000000", -- 2568 - 0xa08  :    0 - 0x0 -- plane 1
    "00000011", -- 2569 - 0xa09  :    3 - 0x3
    "00001111", -- 2570 - 0xa0a  :   15 - 0xf
    "00011111", -- 2571 - 0xa0b  :   31 - 0x1f
    "00111111", -- 2572 - 0xa0c  :   63 - 0x3f
    "00111111", -- 2573 - 0xa0d  :   63 - 0x3f
    "01111111", -- 2574 - 0xa0e  :  127 - 0x7f
    "01111111", -- 2575 - 0xa0f  :  127 - 0x7f
    "11000000", -- 2576 - 0xa10  :  192 - 0xc0 -- Background 0xa1
    "11000000", -- 2577 - 0xa11  :  192 - 0xc0
    "01100000", -- 2578 - 0xa12  :   96 - 0x60
    "01100000", -- 2579 - 0xa13  :   96 - 0x60
    "00110000", -- 2580 - 0xa14  :   48 - 0x30
    "00011010", -- 2581 - 0xa15  :   26 - 0x1a
    "00001101", -- 2582 - 0xa16  :   13 - 0xd
    "00000011", -- 2583 - 0xa17  :    3 - 0x3
    "01111111", -- 2584 - 0xa18  :  127 - 0x7f -- plane 1
    "01111111", -- 2585 - 0xa19  :  127 - 0x7f
    "00111111", -- 2586 - 0xa1a  :   63 - 0x3f
    "00111111", -- 2587 - 0xa1b  :   63 - 0x3f
    "00011111", -- 2588 - 0xa1c  :   31 - 0x1f
    "00000101", -- 2589 - 0xa1d  :    5 - 0x5
    "00000010", -- 2590 - 0xa1e  :    2 - 0x2
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "11000000", -- 2592 - 0xa20  :  192 - 0xc0 -- Background 0xa2
    "11110000", -- 2593 - 0xa21  :  240 - 0xf0
    "00111000", -- 2594 - 0xa22  :   56 - 0x38
    "00001100", -- 2595 - 0xa23  :   12 - 0xc
    "00000110", -- 2596 - 0xa24  :    6 - 0x6
    "00000010", -- 2597 - 0xa25  :    2 - 0x2
    "00000101", -- 2598 - 0xa26  :    5 - 0x5
    "00000011", -- 2599 - 0xa27  :    3 - 0x3
    "00000000", -- 2600 - 0xa28  :    0 - 0x0 -- plane 1
    "11000000", -- 2601 - 0xa29  :  192 - 0xc0
    "11110000", -- 2602 - 0xa2a  :  240 - 0xf0
    "11111000", -- 2603 - 0xa2b  :  248 - 0xf8
    "11111000", -- 2604 - 0xa2c  :  248 - 0xf8
    "11111100", -- 2605 - 0xa2d  :  252 - 0xfc
    "11111010", -- 2606 - 0xa2e  :  250 - 0xfa
    "11111100", -- 2607 - 0xa2f  :  252 - 0xfc
    "00000101", -- 2608 - 0xa30  :    5 - 0x5 -- Background 0xa3
    "00001011", -- 2609 - 0xa31  :   11 - 0xb
    "00010110", -- 2610 - 0xa32  :   22 - 0x16
    "00101010", -- 2611 - 0xa33  :   42 - 0x2a
    "01010100", -- 2612 - 0xa34  :   84 - 0x54
    "10101000", -- 2613 - 0xa35  :  168 - 0xa8
    "01110000", -- 2614 - 0xa36  :  112 - 0x70
    "11000000", -- 2615 - 0xa37  :  192 - 0xc0
    "11111010", -- 2616 - 0xa38  :  250 - 0xfa -- plane 1
    "11110100", -- 2617 - 0xa39  :  244 - 0xf4
    "11101000", -- 2618 - 0xa3a  :  232 - 0xe8
    "11010100", -- 2619 - 0xa3b  :  212 - 0xd4
    "10101000", -- 2620 - 0xa3c  :  168 - 0xa8
    "01010000", -- 2621 - 0xa3d  :   80 - 0x50
    "10000000", -- 2622 - 0xa3e  :  128 - 0x80
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "00000000", -- 2624 - 0xa40  :    0 - 0x0 -- Background 0xa4
    "00001111", -- 2625 - 0xa41  :   15 - 0xf
    "00011111", -- 2626 - 0xa42  :   31 - 0x1f
    "00110001", -- 2627 - 0xa43  :   49 - 0x31
    "00111111", -- 2628 - 0xa44  :   63 - 0x3f
    "01111111", -- 2629 - 0xa45  :  127 - 0x7f
    "11111111", -- 2630 - 0xa46  :  255 - 0xff
    "11011111", -- 2631 - 0xa47  :  223 - 0xdf
    "00000000", -- 2632 - 0xa48  :    0 - 0x0 -- plane 1
    "00000000", -- 2633 - 0xa49  :    0 - 0x0
    "00000000", -- 2634 - 0xa4a  :    0 - 0x0
    "00001110", -- 2635 - 0xa4b  :   14 - 0xe
    "00000000", -- 2636 - 0xa4c  :    0 - 0x0
    "00001010", -- 2637 - 0xa4d  :   10 - 0xa
    "01001010", -- 2638 - 0xa4e  :   74 - 0x4a
    "01100000", -- 2639 - 0xa4f  :   96 - 0x60
    "11000000", -- 2640 - 0xa50  :  192 - 0xc0 -- Background 0xa5
    "11000111", -- 2641 - 0xa51  :  199 - 0xc7
    "01101111", -- 2642 - 0xa52  :  111 - 0x6f
    "01100111", -- 2643 - 0xa53  :  103 - 0x67
    "01100011", -- 2644 - 0xa54  :   99 - 0x63
    "00110000", -- 2645 - 0xa55  :   48 - 0x30
    "00011000", -- 2646 - 0xa56  :   24 - 0x18
    "00000111", -- 2647 - 0xa57  :    7 - 0x7
    "01111111", -- 2648 - 0xa58  :  127 - 0x7f -- plane 1
    "01111000", -- 2649 - 0xa59  :  120 - 0x78
    "00110111", -- 2650 - 0xa5a  :   55 - 0x37
    "00111011", -- 2651 - 0xa5b  :   59 - 0x3b
    "00111100", -- 2652 - 0xa5c  :   60 - 0x3c
    "00011111", -- 2653 - 0xa5d  :   31 - 0x1f
    "00000111", -- 2654 - 0xa5e  :    7 - 0x7
    "00000000", -- 2655 - 0xa5f  :    0 - 0x0
    "00000000", -- 2656 - 0xa60  :    0 - 0x0 -- Background 0xa6
    "11110000", -- 2657 - 0xa61  :  240 - 0xf0
    "11111000", -- 2658 - 0xa62  :  248 - 0xf8
    "10001100", -- 2659 - 0xa63  :  140 - 0x8c
    "11111100", -- 2660 - 0xa64  :  252 - 0xfc
    "11111110", -- 2661 - 0xa65  :  254 - 0xfe
    "11111101", -- 2662 - 0xa66  :  253 - 0xfd
    "11111001", -- 2663 - 0xa67  :  249 - 0xf9
    "00000000", -- 2664 - 0xa68  :    0 - 0x0 -- plane 1
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "00000000", -- 2666 - 0xa6a  :    0 - 0x0
    "01110000", -- 2667 - 0xa6b  :  112 - 0x70
    "00000000", -- 2668 - 0xa6c  :    0 - 0x0
    "01010000", -- 2669 - 0xa6d  :   80 - 0x50
    "01010010", -- 2670 - 0xa6e  :   82 - 0x52
    "00000110", -- 2671 - 0xa6f  :    6 - 0x6
    "00000011", -- 2672 - 0xa70  :    3 - 0x3 -- Background 0xa7
    "11100101", -- 2673 - 0xa71  :  229 - 0xe5
    "11110010", -- 2674 - 0xa72  :  242 - 0xf2
    "11100110", -- 2675 - 0xa73  :  230 - 0xe6
    "11001010", -- 2676 - 0xa74  :  202 - 0xca
    "00010100", -- 2677 - 0xa75  :   20 - 0x14
    "00111000", -- 2678 - 0xa76  :   56 - 0x38
    "11100000", -- 2679 - 0xa77  :  224 - 0xe0
    "11111100", -- 2680 - 0xa78  :  252 - 0xfc -- plane 1
    "00011010", -- 2681 - 0xa79  :   26 - 0x1a
    "11101100", -- 2682 - 0xa7a  :  236 - 0xec
    "11011000", -- 2683 - 0xa7b  :  216 - 0xd8
    "00110100", -- 2684 - 0xa7c  :   52 - 0x34
    "11101000", -- 2685 - 0xa7d  :  232 - 0xe8
    "11000000", -- 2686 - 0xa7e  :  192 - 0xc0
    "00000000", -- 2687 - 0xa7f  :    0 - 0x0
    "00000000", -- 2688 - 0xa80  :    0 - 0x0 -- Background 0xa8
    "00001111", -- 2689 - 0xa81  :   15 - 0xf
    "00011111", -- 2690 - 0xa82  :   31 - 0x1f
    "00110001", -- 2691 - 0xa83  :   49 - 0x31
    "00111111", -- 2692 - 0xa84  :   63 - 0x3f
    "01111111", -- 2693 - 0xa85  :  127 - 0x7f
    "11111111", -- 2694 - 0xa86  :  255 - 0xff
    "11011111", -- 2695 - 0xa87  :  223 - 0xdf
    "00000000", -- 2696 - 0xa88  :    0 - 0x0 -- plane 1
    "00000000", -- 2697 - 0xa89  :    0 - 0x0
    "00000000", -- 2698 - 0xa8a  :    0 - 0x0
    "00001110", -- 2699 - 0xa8b  :   14 - 0xe
    "00000000", -- 2700 - 0xa8c  :    0 - 0x0
    "00001110", -- 2701 - 0xa8d  :   14 - 0xe
    "01001010", -- 2702 - 0xa8e  :   74 - 0x4a
    "01100000", -- 2703 - 0xa8f  :   96 - 0x60
    "11000000", -- 2704 - 0xa90  :  192 - 0xc0 -- Background 0xa9
    "11000011", -- 2705 - 0xa91  :  195 - 0xc3
    "11000111", -- 2706 - 0xa92  :  199 - 0xc7
    "11001111", -- 2707 - 0xa93  :  207 - 0xcf
    "11000111", -- 2708 - 0xa94  :  199 - 0xc7
    "11000000", -- 2709 - 0xa95  :  192 - 0xc0
    "11100000", -- 2710 - 0xa96  :  224 - 0xe0
    "11111111", -- 2711 - 0xa97  :  255 - 0xff
    "01111111", -- 2712 - 0xa98  :  127 - 0x7f -- plane 1
    "01111100", -- 2713 - 0xa99  :  124 - 0x7c
    "01111011", -- 2714 - 0xa9a  :  123 - 0x7b
    "01110111", -- 2715 - 0xa9b  :  119 - 0x77
    "01111000", -- 2716 - 0xa9c  :  120 - 0x78
    "01111111", -- 2717 - 0xa9d  :  127 - 0x7f
    "01111111", -- 2718 - 0xa9e  :  127 - 0x7f
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "00000000", -- 2720 - 0xaa0  :    0 - 0x0 -- Background 0xaa
    "11110000", -- 2721 - 0xaa1  :  240 - 0xf0
    "11111000", -- 2722 - 0xaa2  :  248 - 0xf8
    "10001100", -- 2723 - 0xaa3  :  140 - 0x8c
    "11111100", -- 2724 - 0xaa4  :  252 - 0xfc
    "11111110", -- 2725 - 0xaa5  :  254 - 0xfe
    "11111101", -- 2726 - 0xaa6  :  253 - 0xfd
    "11111001", -- 2727 - 0xaa7  :  249 - 0xf9
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0 -- plane 1
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "00000000", -- 2730 - 0xaaa  :    0 - 0x0
    "01110000", -- 2731 - 0xaab  :  112 - 0x70
    "00000000", -- 2732 - 0xaac  :    0 - 0x0
    "01110000", -- 2733 - 0xaad  :  112 - 0x70
    "01010010", -- 2734 - 0xaae  :   82 - 0x52
    "00000110", -- 2735 - 0xaaf  :    6 - 0x6
    "00000011", -- 2736 - 0xab0  :    3 - 0x3 -- Background 0xab
    "11000101", -- 2737 - 0xab1  :  197 - 0xc5
    "11100011", -- 2738 - 0xab2  :  227 - 0xe3
    "11110101", -- 2739 - 0xab3  :  245 - 0xf5
    "11100011", -- 2740 - 0xab4  :  227 - 0xe3
    "00000101", -- 2741 - 0xab5  :    5 - 0x5
    "00001011", -- 2742 - 0xab6  :   11 - 0xb
    "11111111", -- 2743 - 0xab7  :  255 - 0xff
    "11111100", -- 2744 - 0xab8  :  252 - 0xfc -- plane 1
    "00111010", -- 2745 - 0xab9  :   58 - 0x3a
    "11011100", -- 2746 - 0xaba  :  220 - 0xdc
    "11101010", -- 2747 - 0xabb  :  234 - 0xea
    "00011100", -- 2748 - 0xabc  :   28 - 0x1c
    "11111010", -- 2749 - 0xabd  :  250 - 0xfa
    "11110100", -- 2750 - 0xabe  :  244 - 0xf4
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "10000011", -- 2752 - 0xac0  :  131 - 0x83 -- Background 0xac
    "10001100", -- 2753 - 0xac1  :  140 - 0x8c
    "10010000", -- 2754 - 0xac2  :  144 - 0x90
    "10010000", -- 2755 - 0xac3  :  144 - 0x90
    "11100000", -- 2756 - 0xac4  :  224 - 0xe0
    "10100000", -- 2757 - 0xac5  :  160 - 0xa0
    "10101111", -- 2758 - 0xac6  :  175 - 0xaf
    "01101111", -- 2759 - 0xac7  :  111 - 0x6f
    "00000000", -- 2760 - 0xac8  :    0 - 0x0 -- plane 1
    "00000011", -- 2761 - 0xac9  :    3 - 0x3
    "00001111", -- 2762 - 0xaca  :   15 - 0xf
    "00001111", -- 2763 - 0xacb  :   15 - 0xf
    "00011111", -- 2764 - 0xacc  :   31 - 0x1f
    "01011111", -- 2765 - 0xacd  :   95 - 0x5f
    "01010000", -- 2766 - 0xace  :   80 - 0x50
    "00010000", -- 2767 - 0xacf  :   16 - 0x10
    "11111011", -- 2768 - 0xad0  :  251 - 0xfb -- Background 0xad
    "00000101", -- 2769 - 0xad1  :    5 - 0x5
    "00000101", -- 2770 - 0xad2  :    5 - 0x5
    "00000101", -- 2771 - 0xad3  :    5 - 0x5
    "01000101", -- 2772 - 0xad4  :   69 - 0x45
    "01100101", -- 2773 - 0xad5  :  101 - 0x65
    "11110101", -- 2774 - 0xad6  :  245 - 0xf5
    "11111101", -- 2775 - 0xad7  :  253 - 0xfd
    "00000000", -- 2776 - 0xad8  :    0 - 0x0 -- plane 1
    "11111010", -- 2777 - 0xad9  :  250 - 0xfa
    "11111010", -- 2778 - 0xada  :  250 - 0xfa
    "11111010", -- 2779 - 0xadb  :  250 - 0xfa
    "10111010", -- 2780 - 0xadc  :  186 - 0xba
    "10011010", -- 2781 - 0xadd  :  154 - 0x9a
    "00001010", -- 2782 - 0xade  :   10 - 0xa
    "00000010", -- 2783 - 0xadf  :    2 - 0x2
    "10000011", -- 2784 - 0xae0  :  131 - 0x83 -- Background 0xae
    "10001100", -- 2785 - 0xae1  :  140 - 0x8c
    "10010000", -- 2786 - 0xae2  :  144 - 0x90
    "10010000", -- 2787 - 0xae3  :  144 - 0x90
    "11100000", -- 2788 - 0xae4  :  224 - 0xe0
    "10100000", -- 2789 - 0xae5  :  160 - 0xa0
    "10101111", -- 2790 - 0xae6  :  175 - 0xaf
    "01101111", -- 2791 - 0xae7  :  111 - 0x6f
    "00000000", -- 2792 - 0xae8  :    0 - 0x0 -- plane 1
    "00000011", -- 2793 - 0xae9  :    3 - 0x3
    "00001111", -- 2794 - 0xaea  :   15 - 0xf
    "00001111", -- 2795 - 0xaeb  :   15 - 0xf
    "00011111", -- 2796 - 0xaec  :   31 - 0x1f
    "01011111", -- 2797 - 0xaed  :   95 - 0x5f
    "01010000", -- 2798 - 0xaee  :   80 - 0x50
    "00010111", -- 2799 - 0xaef  :   23 - 0x17
    "11111011", -- 2800 - 0xaf0  :  251 - 0xfb -- Background 0xaf
    "00000101", -- 2801 - 0xaf1  :    5 - 0x5
    "00000101", -- 2802 - 0xaf2  :    5 - 0x5
    "00000101", -- 2803 - 0xaf3  :    5 - 0x5
    "11000101", -- 2804 - 0xaf4  :  197 - 0xc5
    "11100101", -- 2805 - 0xaf5  :  229 - 0xe5
    "11110101", -- 2806 - 0xaf6  :  245 - 0xf5
    "11111101", -- 2807 - 0xaf7  :  253 - 0xfd
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0 -- plane 1
    "11111010", -- 2809 - 0xaf9  :  250 - 0xfa
    "11111010", -- 2810 - 0xafa  :  250 - 0xfa
    "11111010", -- 2811 - 0xafb  :  250 - 0xfa
    "00111010", -- 2812 - 0xafc  :   58 - 0x3a
    "01011010", -- 2813 - 0xafd  :   90 - 0x5a
    "01101010", -- 2814 - 0xafe  :  106 - 0x6a
    "11110010", -- 2815 - 0xaff  :  242 - 0xf2
    "00000000", -- 2816 - 0xb00  :    0 - 0x0 -- Background 0xb0
    "00000011", -- 2817 - 0xb01  :    3 - 0x3
    "00001111", -- 2818 - 0xb02  :   15 - 0xf
    "00111111", -- 2819 - 0xb03  :   63 - 0x3f
    "01111111", -- 2820 - 0xb04  :  127 - 0x7f
    "01111111", -- 2821 - 0xb05  :  127 - 0x7f
    "11111111", -- 2822 - 0xb06  :  255 - 0xff
    "11111111", -- 2823 - 0xb07  :  255 - 0xff
    "00000000", -- 2824 - 0xb08  :    0 - 0x0 -- plane 1
    "00000000", -- 2825 - 0xb09  :    0 - 0x0
    "00000011", -- 2826 - 0xb0a  :    3 - 0x3
    "00001111", -- 2827 - 0xb0b  :   15 - 0xf
    "00111011", -- 2828 - 0xb0c  :   59 - 0x3b
    "00111111", -- 2829 - 0xb0d  :   63 - 0x3f
    "01101111", -- 2830 - 0xb0e  :  111 - 0x6f
    "01111101", -- 2831 - 0xb0f  :  125 - 0x7d
    "11111111", -- 2832 - 0xb10  :  255 - 0xff -- Background 0xb1
    "10001111", -- 2833 - 0xb11  :  143 - 0x8f
    "10000000", -- 2834 - 0xb12  :  128 - 0x80
    "11110000", -- 2835 - 0xb13  :  240 - 0xf0
    "11111111", -- 2836 - 0xb14  :  255 - 0xff
    "11111111", -- 2837 - 0xb15  :  255 - 0xff
    "01111111", -- 2838 - 0xb16  :  127 - 0x7f
    "00001111", -- 2839 - 0xb17  :   15 - 0xf
    "00001111", -- 2840 - 0xb18  :   15 - 0xf -- plane 1
    "01110000", -- 2841 - 0xb19  :  112 - 0x70
    "01111111", -- 2842 - 0xb1a  :  127 - 0x7f
    "00001111", -- 2843 - 0xb1b  :   15 - 0xf
    "01110000", -- 2844 - 0xb1c  :  112 - 0x70
    "01111111", -- 2845 - 0xb1d  :  127 - 0x7f
    "00001111", -- 2846 - 0xb1e  :   15 - 0xf
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "00000000", -- 2848 - 0xb20  :    0 - 0x0 -- Background 0xb2
    "11000000", -- 2849 - 0xb21  :  192 - 0xc0
    "11110000", -- 2850 - 0xb22  :  240 - 0xf0
    "11111100", -- 2851 - 0xb23  :  252 - 0xfc
    "11111110", -- 2852 - 0xb24  :  254 - 0xfe
    "11111110", -- 2853 - 0xb25  :  254 - 0xfe
    "11111111", -- 2854 - 0xb26  :  255 - 0xff
    "11111111", -- 2855 - 0xb27  :  255 - 0xff
    "00000000", -- 2856 - 0xb28  :    0 - 0x0 -- plane 1
    "00000000", -- 2857 - 0xb29  :    0 - 0x0
    "11000000", -- 2858 - 0xb2a  :  192 - 0xc0
    "11110000", -- 2859 - 0xb2b  :  240 - 0xf0
    "10111100", -- 2860 - 0xb2c  :  188 - 0xbc
    "11110100", -- 2861 - 0xb2d  :  244 - 0xf4
    "11111110", -- 2862 - 0xb2e  :  254 - 0xfe
    "11011110", -- 2863 - 0xb2f  :  222 - 0xde
    "11111111", -- 2864 - 0xb30  :  255 - 0xff -- Background 0xb3
    "11110001", -- 2865 - 0xb31  :  241 - 0xf1
    "00000001", -- 2866 - 0xb32  :    1 - 0x1
    "00001111", -- 2867 - 0xb33  :   15 - 0xf
    "11111111", -- 2868 - 0xb34  :  255 - 0xff
    "11111111", -- 2869 - 0xb35  :  255 - 0xff
    "11111110", -- 2870 - 0xb36  :  254 - 0xfe
    "11110000", -- 2871 - 0xb37  :  240 - 0xf0
    "11110000", -- 2872 - 0xb38  :  240 - 0xf0 -- plane 1
    "00001110", -- 2873 - 0xb39  :   14 - 0xe
    "11111110", -- 2874 - 0xb3a  :  254 - 0xfe
    "11110000", -- 2875 - 0xb3b  :  240 - 0xf0
    "00001110", -- 2876 - 0xb3c  :   14 - 0xe
    "11111110", -- 2877 - 0xb3d  :  254 - 0xfe
    "11110000", -- 2878 - 0xb3e  :  240 - 0xf0
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "00000000", -- 2880 - 0xb40  :    0 - 0x0 -- Background 0xb4
    "00000011", -- 2881 - 0xb41  :    3 - 0x3
    "00001110", -- 2882 - 0xb42  :   14 - 0xe
    "00110101", -- 2883 - 0xb43  :   53 - 0x35
    "01101110", -- 2884 - 0xb44  :  110 - 0x6e
    "01010101", -- 2885 - 0xb45  :   85 - 0x55
    "10111010", -- 2886 - 0xb46  :  186 - 0xba
    "11010111", -- 2887 - 0xb47  :  215 - 0xd7
    "00000000", -- 2888 - 0xb48  :    0 - 0x0 -- plane 1
    "00000000", -- 2889 - 0xb49  :    0 - 0x0
    "00000011", -- 2890 - 0xb4a  :    3 - 0x3
    "00001111", -- 2891 - 0xb4b  :   15 - 0xf
    "00111011", -- 2892 - 0xb4c  :   59 - 0x3b
    "00111111", -- 2893 - 0xb4d  :   63 - 0x3f
    "01101111", -- 2894 - 0xb4e  :  111 - 0x6f
    "01111101", -- 2895 - 0xb4f  :  125 - 0x7d
    "11111010", -- 2896 - 0xb50  :  250 - 0xfa -- Background 0xb5
    "10001111", -- 2897 - 0xb51  :  143 - 0x8f
    "10000000", -- 2898 - 0xb52  :  128 - 0x80
    "11110000", -- 2899 - 0xb53  :  240 - 0xf0
    "10101111", -- 2900 - 0xb54  :  175 - 0xaf
    "11010101", -- 2901 - 0xb55  :  213 - 0xd5
    "01111010", -- 2902 - 0xb56  :  122 - 0x7a
    "00001111", -- 2903 - 0xb57  :   15 - 0xf
    "00001111", -- 2904 - 0xb58  :   15 - 0xf -- plane 1
    "01110000", -- 2905 - 0xb59  :  112 - 0x70
    "01111111", -- 2906 - 0xb5a  :  127 - 0x7f
    "00001111", -- 2907 - 0xb5b  :   15 - 0xf
    "01110000", -- 2908 - 0xb5c  :  112 - 0x70
    "01111111", -- 2909 - 0xb5d  :  127 - 0x7f
    "00001111", -- 2910 - 0xb5e  :   15 - 0xf
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "00000000", -- 2912 - 0xb60  :    0 - 0x0 -- Background 0xb6
    "11000000", -- 2913 - 0xb61  :  192 - 0xc0
    "10110000", -- 2914 - 0xb62  :  176 - 0xb0
    "01011100", -- 2915 - 0xb63  :   92 - 0x5c
    "11101010", -- 2916 - 0xb64  :  234 - 0xea
    "01011110", -- 2917 - 0xb65  :   94 - 0x5e
    "10101011", -- 2918 - 0xb66  :  171 - 0xab
    "01110101", -- 2919 - 0xb67  :  117 - 0x75
    "00000000", -- 2920 - 0xb68  :    0 - 0x0 -- plane 1
    "00000000", -- 2921 - 0xb69  :    0 - 0x0
    "11000000", -- 2922 - 0xb6a  :  192 - 0xc0
    "11110000", -- 2923 - 0xb6b  :  240 - 0xf0
    "10111100", -- 2924 - 0xb6c  :  188 - 0xbc
    "11110100", -- 2925 - 0xb6d  :  244 - 0xf4
    "11111110", -- 2926 - 0xb6e  :  254 - 0xfe
    "11011110", -- 2927 - 0xb6f  :  222 - 0xde
    "10101111", -- 2928 - 0xb70  :  175 - 0xaf -- Background 0xb7
    "11110001", -- 2929 - 0xb71  :  241 - 0xf1
    "00000001", -- 2930 - 0xb72  :    1 - 0x1
    "00001111", -- 2931 - 0xb73  :   15 - 0xf
    "11111011", -- 2932 - 0xb74  :  251 - 0xfb
    "01010101", -- 2933 - 0xb75  :   85 - 0x55
    "10101110", -- 2934 - 0xb76  :  174 - 0xae
    "11110000", -- 2935 - 0xb77  :  240 - 0xf0
    "11110000", -- 2936 - 0xb78  :  240 - 0xf0 -- plane 1
    "00001110", -- 2937 - 0xb79  :   14 - 0xe
    "11111110", -- 2938 - 0xb7a  :  254 - 0xfe
    "11110000", -- 2939 - 0xb7b  :  240 - 0xf0
    "00001110", -- 2940 - 0xb7c  :   14 - 0xe
    "11111110", -- 2941 - 0xb7d  :  254 - 0xfe
    "11110000", -- 2942 - 0xb7e  :  240 - 0xf0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "00000000", -- 2944 - 0xb80  :    0 - 0x0 -- Background 0xb8
    "00000011", -- 2945 - 0xb81  :    3 - 0x3
    "00001100", -- 2946 - 0xb82  :   12 - 0xc
    "00110000", -- 2947 - 0xb83  :   48 - 0x30
    "01000100", -- 2948 - 0xb84  :   68 - 0x44
    "01000000", -- 2949 - 0xb85  :   64 - 0x40
    "10010000", -- 2950 - 0xb86  :  144 - 0x90
    "10000010", -- 2951 - 0xb87  :  130 - 0x82
    "00000000", -- 2952 - 0xb88  :    0 - 0x0 -- plane 1
    "00000000", -- 2953 - 0xb89  :    0 - 0x0
    "00000011", -- 2954 - 0xb8a  :    3 - 0x3
    "00001111", -- 2955 - 0xb8b  :   15 - 0xf
    "00111011", -- 2956 - 0xb8c  :   59 - 0x3b
    "00111111", -- 2957 - 0xb8d  :   63 - 0x3f
    "01101111", -- 2958 - 0xb8e  :  111 - 0x6f
    "01111101", -- 2959 - 0xb8f  :  125 - 0x7d
    "11110000", -- 2960 - 0xb90  :  240 - 0xf0 -- Background 0xb9
    "11111111", -- 2961 - 0xb91  :  255 - 0xff
    "11111111", -- 2962 - 0xb92  :  255 - 0xff
    "11111111", -- 2963 - 0xb93  :  255 - 0xff
    "10001111", -- 2964 - 0xb94  :  143 - 0x8f
    "10000000", -- 2965 - 0xb95  :  128 - 0x80
    "01110000", -- 2966 - 0xb96  :  112 - 0x70
    "00001111", -- 2967 - 0xb97  :   15 - 0xf
    "00001111", -- 2968 - 0xb98  :   15 - 0xf -- plane 1
    "00100000", -- 2969 - 0xb99  :   32 - 0x20
    "01010101", -- 2970 - 0xb9a  :   85 - 0x55
    "00001010", -- 2971 - 0xb9b  :   10 - 0xa
    "01110000", -- 2972 - 0xb9c  :  112 - 0x70
    "01111111", -- 2973 - 0xb9d  :  127 - 0x7f
    "00001111", -- 2974 - 0xb9e  :   15 - 0xf
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "00000000", -- 2976 - 0xba0  :    0 - 0x0 -- Background 0xba
    "11000000", -- 2977 - 0xba1  :  192 - 0xc0
    "00110000", -- 2978 - 0xba2  :   48 - 0x30
    "00001100", -- 2979 - 0xba3  :   12 - 0xc
    "01000010", -- 2980 - 0xba4  :   66 - 0x42
    "00001010", -- 2981 - 0xba5  :   10 - 0xa
    "00000001", -- 2982 - 0xba6  :    1 - 0x1
    "00100001", -- 2983 - 0xba7  :   33 - 0x21
    "00000000", -- 2984 - 0xba8  :    0 - 0x0 -- plane 1
    "00000000", -- 2985 - 0xba9  :    0 - 0x0
    "11000000", -- 2986 - 0xbaa  :  192 - 0xc0
    "11110000", -- 2987 - 0xbab  :  240 - 0xf0
    "10111100", -- 2988 - 0xbac  :  188 - 0xbc
    "11110100", -- 2989 - 0xbad  :  244 - 0xf4
    "11111110", -- 2990 - 0xbae  :  254 - 0xfe
    "11011110", -- 2991 - 0xbaf  :  222 - 0xde
    "00001111", -- 2992 - 0xbb0  :   15 - 0xf -- Background 0xbb
    "11111111", -- 2993 - 0xbb1  :  255 - 0xff
    "11111111", -- 2994 - 0xbb2  :  255 - 0xff
    "11111111", -- 2995 - 0xbb3  :  255 - 0xff
    "11110001", -- 2996 - 0xbb4  :  241 - 0xf1
    "00000001", -- 2997 - 0xbb5  :    1 - 0x1
    "00001110", -- 2998 - 0xbb6  :   14 - 0xe
    "11110000", -- 2999 - 0xbb7  :  240 - 0xf0
    "11110000", -- 3000 - 0xbb8  :  240 - 0xf0 -- plane 1
    "00001010", -- 3001 - 0xbb9  :   10 - 0xa
    "01010100", -- 3002 - 0xbba  :   84 - 0x54
    "10100000", -- 3003 - 0xbbb  :  160 - 0xa0
    "00001110", -- 3004 - 0xbbc  :   14 - 0xe
    "11111110", -- 3005 - 0xbbd  :  254 - 0xfe
    "11110000", -- 3006 - 0xbbe  :  240 - 0xf0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "11110011", -- 3008 - 0xbc0  :  243 - 0xf3 -- Background 0xbc
    "11111111", -- 3009 - 0xbc1  :  255 - 0xff
    "11000100", -- 3010 - 0xbc2  :  196 - 0xc4
    "11000000", -- 3011 - 0xbc3  :  192 - 0xc0
    "01000000", -- 3012 - 0xbc4  :   64 - 0x40
    "01100011", -- 3013 - 0xbc5  :   99 - 0x63
    "11000111", -- 3014 - 0xbc6  :  199 - 0xc7
    "11000110", -- 3015 - 0xbc7  :  198 - 0xc6
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0 -- plane 1
    "01110011", -- 3017 - 0xbc9  :  115 - 0x73
    "01111011", -- 3018 - 0xbca  :  123 - 0x7b
    "01111111", -- 3019 - 0xbcb  :  127 - 0x7f
    "00111111", -- 3020 - 0xbcc  :   63 - 0x3f
    "00011100", -- 3021 - 0xbcd  :   28 - 0x1c
    "01111011", -- 3022 - 0xbce  :  123 - 0x7b
    "01111011", -- 3023 - 0xbcf  :  123 - 0x7b
    "11000110", -- 3024 - 0xbd0  :  198 - 0xc6 -- Background 0xbd
    "11000110", -- 3025 - 0xbd1  :  198 - 0xc6
    "01100011", -- 3026 - 0xbd2  :   99 - 0x63
    "01000000", -- 3027 - 0xbd3  :   64 - 0x40
    "11000000", -- 3028 - 0xbd4  :  192 - 0xc0
    "11000100", -- 3029 - 0xbd5  :  196 - 0xc4
    "11001100", -- 3030 - 0xbd6  :  204 - 0xcc
    "11110011", -- 3031 - 0xbd7  :  243 - 0xf3
    "01111011", -- 3032 - 0xbd8  :  123 - 0x7b -- plane 1
    "01111011", -- 3033 - 0xbd9  :  123 - 0x7b
    "00011100", -- 3034 - 0xbda  :   28 - 0x1c
    "00111111", -- 3035 - 0xbdb  :   63 - 0x3f
    "01111111", -- 3036 - 0xbdc  :  127 - 0x7f
    "01111011", -- 3037 - 0xbdd  :  123 - 0x7b
    "01110011", -- 3038 - 0xbde  :  115 - 0x73
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "11001111", -- 3040 - 0xbe0  :  207 - 0xcf -- Background 0xbe
    "11111111", -- 3041 - 0xbe1  :  255 - 0xff
    "00100001", -- 3042 - 0xbe2  :   33 - 0x21
    "00000001", -- 3043 - 0xbe3  :    1 - 0x1
    "00000010", -- 3044 - 0xbe4  :    2 - 0x2
    "11000110", -- 3045 - 0xbe5  :  198 - 0xc6
    "11100001", -- 3046 - 0xbe6  :  225 - 0xe1
    "00100001", -- 3047 - 0xbe7  :   33 - 0x21
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0 -- plane 1
    "11001110", -- 3049 - 0xbe9  :  206 - 0xce
    "11011110", -- 3050 - 0xbea  :  222 - 0xde
    "11111110", -- 3051 - 0xbeb  :  254 - 0xfe
    "11111100", -- 3052 - 0xbec  :  252 - 0xfc
    "00111000", -- 3053 - 0xbed  :   56 - 0x38
    "11011110", -- 3054 - 0xbee  :  222 - 0xde
    "11011110", -- 3055 - 0xbef  :  222 - 0xde
    "00100001", -- 3056 - 0xbf0  :   33 - 0x21 -- Background 0xbf
    "00100001", -- 3057 - 0xbf1  :   33 - 0x21
    "11000110", -- 3058 - 0xbf2  :  198 - 0xc6
    "00000010", -- 3059 - 0xbf3  :    2 - 0x2
    "00000001", -- 3060 - 0xbf4  :    1 - 0x1
    "00100001", -- 3061 - 0xbf5  :   33 - 0x21
    "00110001", -- 3062 - 0xbf6  :   49 - 0x31
    "11001111", -- 3063 - 0xbf7  :  207 - 0xcf
    "11011110", -- 3064 - 0xbf8  :  222 - 0xde -- plane 1
    "11011110", -- 3065 - 0xbf9  :  222 - 0xde
    "00111000", -- 3066 - 0xbfa  :   56 - 0x38
    "11111100", -- 3067 - 0xbfb  :  252 - 0xfc
    "11111110", -- 3068 - 0xbfc  :  254 - 0xfe
    "11011110", -- 3069 - 0xbfd  :  222 - 0xde
    "11001110", -- 3070 - 0xbfe  :  206 - 0xce
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00000000", -- 3072 - 0xc00  :    0 - 0x0 -- Background 0xc0
    "01010000", -- 3073 - 0xc01  :   80 - 0x50
    "10110011", -- 3074 - 0xc02  :  179 - 0xb3
    "10010111", -- 3075 - 0xc03  :  151 - 0x97
    "10011111", -- 3076 - 0xc04  :  159 - 0x9f
    "01101111", -- 3077 - 0xc05  :  111 - 0x6f
    "00011111", -- 3078 - 0xc06  :   31 - 0x1f
    "00011111", -- 3079 - 0xc07  :   31 - 0x1f
    "00000000", -- 3080 - 0xc08  :    0 - 0x0 -- plane 1
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "01000000", -- 3082 - 0xc0a  :   64 - 0x40
    "01100000", -- 3083 - 0xc0b  :   96 - 0x60
    "01100001", -- 3084 - 0xc0c  :   97 - 0x61
    "00000010", -- 3085 - 0xc0d  :    2 - 0x2
    "00000010", -- 3086 - 0xc0e  :    2 - 0x2
    "00000111", -- 3087 - 0xc0f  :    7 - 0x7
    "00011111", -- 3088 - 0xc10  :   31 - 0x1f -- Background 0xc1
    "00011111", -- 3089 - 0xc11  :   31 - 0x1f
    "00001111", -- 3090 - 0xc12  :   15 - 0xf
    "00000111", -- 3091 - 0xc13  :    7 - 0x7
    "00011101", -- 3092 - 0xc14  :   29 - 0x1d
    "00101100", -- 3093 - 0xc15  :   44 - 0x2c
    "01010100", -- 3094 - 0xc16  :   84 - 0x54
    "01111100", -- 3095 - 0xc17  :  124 - 0x7c
    "00000111", -- 3096 - 0xc18  :    7 - 0x7 -- plane 1
    "00000100", -- 3097 - 0xc19  :    4 - 0x4
    "00000111", -- 3098 - 0xc1a  :    7 - 0x7
    "00000001", -- 3099 - 0xc1b  :    1 - 0x1
    "00000000", -- 3100 - 0xc1c  :    0 - 0x0
    "00010000", -- 3101 - 0xc1d  :   16 - 0x10
    "00101000", -- 3102 - 0xc1e  :   40 - 0x28
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00000000", -- 3104 - 0xc20  :    0 - 0x0 -- Background 0xc2
    "00001010", -- 3105 - 0xc21  :   10 - 0xa
    "11001101", -- 3106 - 0xc22  :  205 - 0xcd
    "11101001", -- 3107 - 0xc23  :  233 - 0xe9
    "11111001", -- 3108 - 0xc24  :  249 - 0xf9
    "11110110", -- 3109 - 0xc25  :  246 - 0xf6
    "11110000", -- 3110 - 0xc26  :  240 - 0xf0
    "11111000", -- 3111 - 0xc27  :  248 - 0xf8
    "00000000", -- 3112 - 0xc28  :    0 - 0x0 -- plane 1
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000010", -- 3114 - 0xc2a  :    2 - 0x2
    "00000110", -- 3115 - 0xc2b  :    6 - 0x6
    "11100110", -- 3116 - 0xc2c  :  230 - 0xe6
    "10100000", -- 3117 - 0xc2d  :  160 - 0xa0
    "10100000", -- 3118 - 0xc2e  :  160 - 0xa0
    "11110000", -- 3119 - 0xc2f  :  240 - 0xf0
    "11111000", -- 3120 - 0xc30  :  248 - 0xf8 -- Background 0xc3
    "11111000", -- 3121 - 0xc31  :  248 - 0xf8
    "11110000", -- 3122 - 0xc32  :  240 - 0xf0
    "11000000", -- 3123 - 0xc33  :  192 - 0xc0
    "10111000", -- 3124 - 0xc34  :  184 - 0xb8
    "00110100", -- 3125 - 0xc35  :   52 - 0x34
    "00101010", -- 3126 - 0xc36  :   42 - 0x2a
    "00111110", -- 3127 - 0xc37  :   62 - 0x3e
    "11110000", -- 3128 - 0xc38  :  240 - 0xf0 -- plane 1
    "00110000", -- 3129 - 0xc39  :   48 - 0x30
    "11000000", -- 3130 - 0xc3a  :  192 - 0xc0
    "10000000", -- 3131 - 0xc3b  :  128 - 0x80
    "00000000", -- 3132 - 0xc3c  :    0 - 0x0
    "00001000", -- 3133 - 0xc3d  :    8 - 0x8
    "00010100", -- 3134 - 0xc3e  :   20 - 0x14
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00000101", -- 3136 - 0xc40  :    5 - 0x5 -- Background 0xc4
    "00001010", -- 3137 - 0xc41  :   10 - 0xa
    "00001000", -- 3138 - 0xc42  :    8 - 0x8
    "00001111", -- 3139 - 0xc43  :   15 - 0xf
    "00000001", -- 3140 - 0xc44  :    1 - 0x1
    "00000011", -- 3141 - 0xc45  :    3 - 0x3
    "00000111", -- 3142 - 0xc46  :    7 - 0x7
    "00001111", -- 3143 - 0xc47  :   15 - 0xf
    "00000000", -- 3144 - 0xc48  :    0 - 0x0 -- plane 1
    "00000101", -- 3145 - 0xc49  :    5 - 0x5
    "00000111", -- 3146 - 0xc4a  :    7 - 0x7
    "00000000", -- 3147 - 0xc4b  :    0 - 0x0
    "00000000", -- 3148 - 0xc4c  :    0 - 0x0
    "00000000", -- 3149 - 0xc4d  :    0 - 0x0
    "00000000", -- 3150 - 0xc4e  :    0 - 0x0
    "00000001", -- 3151 - 0xc4f  :    1 - 0x1
    "00001111", -- 3152 - 0xc50  :   15 - 0xf -- Background 0xc5
    "11101111", -- 3153 - 0xc51  :  239 - 0xef
    "11011111", -- 3154 - 0xc52  :  223 - 0xdf
    "10101111", -- 3155 - 0xc53  :  175 - 0xaf
    "01100111", -- 3156 - 0xc54  :  103 - 0x67
    "00001101", -- 3157 - 0xc55  :   13 - 0xd
    "00001010", -- 3158 - 0xc56  :   10 - 0xa
    "00000111", -- 3159 - 0xc57  :    7 - 0x7
    "00000010", -- 3160 - 0xc58  :    2 - 0x2 -- plane 1
    "00000111", -- 3161 - 0xc59  :    7 - 0x7
    "00100111", -- 3162 - 0xc5a  :   39 - 0x27
    "01010011", -- 3163 - 0xc5b  :   83 - 0x53
    "00000000", -- 3164 - 0xc5c  :    0 - 0x0
    "00000010", -- 3165 - 0xc5d  :    2 - 0x2
    "00000101", -- 3166 - 0xc5e  :    5 - 0x5
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "00000000", -- 3168 - 0xc60  :    0 - 0x0 -- Background 0xc6
    "10000000", -- 3169 - 0xc61  :  128 - 0x80
    "10000000", -- 3170 - 0xc62  :  128 - 0x80
    "11110000", -- 3171 - 0xc63  :  240 - 0xf0
    "11111000", -- 3172 - 0xc64  :  248 - 0xf8
    "11111100", -- 3173 - 0xc65  :  252 - 0xfc
    "11111100", -- 3174 - 0xc66  :  252 - 0xfc
    "11111100", -- 3175 - 0xc67  :  252 - 0xfc
    "00000000", -- 3176 - 0xc68  :    0 - 0x0 -- plane 1
    "00000000", -- 3177 - 0xc69  :    0 - 0x0
    "00000000", -- 3178 - 0xc6a  :    0 - 0x0
    "00000000", -- 3179 - 0xc6b  :    0 - 0x0
    "00000000", -- 3180 - 0xc6c  :    0 - 0x0
    "01100000", -- 3181 - 0xc6d  :   96 - 0x60
    "11011000", -- 3182 - 0xc6e  :  216 - 0xd8
    "10110000", -- 3183 - 0xc6f  :  176 - 0xb0
    "11111100", -- 3184 - 0xc70  :  252 - 0xfc -- Background 0xc7
    "11111110", -- 3185 - 0xc71  :  254 - 0xfe
    "11111001", -- 3186 - 0xc72  :  249 - 0xf9
    "11111010", -- 3187 - 0xc73  :  250 - 0xfa
    "11101001", -- 3188 - 0xc74  :  233 - 0xe9
    "00001110", -- 3189 - 0xc75  :   14 - 0xe
    "10000000", -- 3190 - 0xc76  :  128 - 0x80
    "00000000", -- 3191 - 0xc77  :    0 - 0x0
    "11101000", -- 3192 - 0xc78  :  232 - 0xe8 -- plane 1
    "01111000", -- 3193 - 0xc79  :  120 - 0x78
    "10110110", -- 3194 - 0xc7a  :  182 - 0xb6
    "11100100", -- 3195 - 0xc7b  :  228 - 0xe4
    "00000110", -- 3196 - 0xc7c  :    6 - 0x6
    "00000000", -- 3197 - 0xc7d  :    0 - 0x0
    "00000000", -- 3198 - 0xc7e  :    0 - 0x0
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Background 0xc8
    "11000000", -- 3201 - 0xc81  :  192 - 0xc0
    "10100000", -- 3202 - 0xc82  :  160 - 0xa0
    "11010011", -- 3203 - 0xc83  :  211 - 0xd3
    "10110111", -- 3204 - 0xc84  :  183 - 0xb7
    "11111111", -- 3205 - 0xc85  :  255 - 0xff
    "00001111", -- 3206 - 0xc86  :   15 - 0xf
    "00011111", -- 3207 - 0xc87  :   31 - 0x1f
    "00000000", -- 3208 - 0xc88  :    0 - 0x0 -- plane 1
    "00000000", -- 3209 - 0xc89  :    0 - 0x0
    "01000000", -- 3210 - 0xc8a  :   64 - 0x40
    "00100000", -- 3211 - 0xc8b  :   32 - 0x20
    "01000000", -- 3212 - 0xc8c  :   64 - 0x40
    "00000111", -- 3213 - 0xc8d  :    7 - 0x7
    "00000101", -- 3214 - 0xc8e  :    5 - 0x5
    "00001101", -- 3215 - 0xc8f  :   13 - 0xd
    "00011111", -- 3216 - 0xc90  :   31 - 0x1f -- Background 0xc9
    "00001111", -- 3217 - 0xc91  :   15 - 0xf
    "11110111", -- 3218 - 0xc92  :  247 - 0xf7
    "10110111", -- 3219 - 0xc93  :  183 - 0xb7
    "11010011", -- 3220 - 0xc94  :  211 - 0xd3
    "10100000", -- 3221 - 0xc95  :  160 - 0xa0
    "11000000", -- 3222 - 0xc96  :  192 - 0xc0
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "00001101", -- 3224 - 0xc98  :   13 - 0xd -- plane 1
    "00000101", -- 3225 - 0xc99  :    5 - 0x5
    "00000011", -- 3226 - 0xc9a  :    3 - 0x3
    "01000011", -- 3227 - 0xc9b  :   67 - 0x43
    "00100000", -- 3228 - 0xc9c  :   32 - 0x20
    "01000000", -- 3229 - 0xc9d  :   64 - 0x40
    "00000000", -- 3230 - 0xc9e  :    0 - 0x0
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00011100", -- 3232 - 0xca0  :   28 - 0x1c -- Background 0xca
    "00100010", -- 3233 - 0xca1  :   34 - 0x22
    "00100100", -- 3234 - 0xca2  :   36 - 0x24
    "11011110", -- 3235 - 0xca3  :  222 - 0xde
    "11110000", -- 3236 - 0xca4  :  240 - 0xf0
    "11111000", -- 3237 - 0xca5  :  248 - 0xf8
    "11111100", -- 3238 - 0xca6  :  252 - 0xfc
    "11111100", -- 3239 - 0xca7  :  252 - 0xfc
    "00000000", -- 3240 - 0xca8  :    0 - 0x0 -- plane 1
    "00011100", -- 3241 - 0xca9  :   28 - 0x1c
    "00011000", -- 3242 - 0xcaa  :   24 - 0x18
    "00000000", -- 3243 - 0xcab  :    0 - 0x0
    "00000000", -- 3244 - 0xcac  :    0 - 0x0
    "10000000", -- 3245 - 0xcad  :  128 - 0x80
    "11100000", -- 3246 - 0xcae  :  224 - 0xe0
    "10010000", -- 3247 - 0xcaf  :  144 - 0x90
    "11111100", -- 3248 - 0xcb0  :  252 - 0xfc -- Background 0xcb
    "11111100", -- 3249 - 0xcb1  :  252 - 0xfc
    "11111000", -- 3250 - 0xcb2  :  248 - 0xf8
    "11110000", -- 3251 - 0xcb3  :  240 - 0xf0
    "10011110", -- 3252 - 0xcb4  :  158 - 0x9e
    "00100100", -- 3253 - 0xcb5  :   36 - 0x24
    "00100010", -- 3254 - 0xcb6  :   34 - 0x22
    "00011100", -- 3255 - 0xcb7  :   28 - 0x1c
    "11110000", -- 3256 - 0xcb8  :  240 - 0xf0 -- plane 1
    "10010000", -- 3257 - 0xcb9  :  144 - 0x90
    "11110000", -- 3258 - 0xcba  :  240 - 0xf0
    "10000000", -- 3259 - 0xcbb  :  128 - 0x80
    "00000000", -- 3260 - 0xcbc  :    0 - 0x0
    "00011000", -- 3261 - 0xcbd  :   24 - 0x18
    "00011100", -- 3262 - 0xcbe  :   28 - 0x1c
    "00000000", -- 3263 - 0xcbf  :    0 - 0x0
    "00001110", -- 3264 - 0xcc0  :   14 - 0xe -- Background 0xcc
    "00010110", -- 3265 - 0xcc1  :   22 - 0x16
    "00011010", -- 3266 - 0xcc2  :   26 - 0x1a
    "00000100", -- 3267 - 0xcc3  :    4 - 0x4
    "01101111", -- 3268 - 0xcc4  :  111 - 0x6f
    "10111111", -- 3269 - 0xcc5  :  191 - 0xbf
    "11011111", -- 3270 - 0xcc6  :  223 - 0xdf
    "10111111", -- 3271 - 0xcc7  :  191 - 0xbf
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0 -- plane 1
    "00001000", -- 3273 - 0xcc9  :    8 - 0x8
    "00000100", -- 3274 - 0xcca  :    4 - 0x4
    "00001000", -- 3275 - 0xccb  :    8 - 0x8
    "00000000", -- 3276 - 0xccc  :    0 - 0x0
    "01000110", -- 3277 - 0xccd  :   70 - 0x46
    "00101111", -- 3278 - 0xcce  :   47 - 0x2f
    "01001110", -- 3279 - 0xccf  :   78 - 0x4e
    "01011111", -- 3280 - 0xcd0  :   95 - 0x5f -- Background 0xcd
    "00011111", -- 3281 - 0xcd1  :   31 - 0x1f
    "00011111", -- 3282 - 0xcd2  :   31 - 0x1f
    "00001111", -- 3283 - 0xcd3  :   15 - 0xf
    "00111111", -- 3284 - 0xcd4  :   63 - 0x3f
    "00100011", -- 3285 - 0xcd5  :   35 - 0x23
    "00101010", -- 3286 - 0xcd6  :   42 - 0x2a
    "00010100", -- 3287 - 0xcd7  :   20 - 0x14
    "00001101", -- 3288 - 0xcd8  :   13 - 0xd -- plane 1
    "00001011", -- 3289 - 0xcd9  :   11 - 0xb
    "00001111", -- 3290 - 0xcda  :   15 - 0xf
    "00000110", -- 3291 - 0xcdb  :    6 - 0x6
    "00000011", -- 3292 - 0xcdc  :    3 - 0x3
    "00011100", -- 3293 - 0xcdd  :   28 - 0x1c
    "00010100", -- 3294 - 0xcde  :   20 - 0x14
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Background 0xce
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "00000000", -- 3299 - 0xce3  :    0 - 0x0
    "10001110", -- 3300 - 0xce4  :  142 - 0x8e
    "11001001", -- 3301 - 0xce5  :  201 - 0xc9
    "11101010", -- 3302 - 0xce6  :  234 - 0xea
    "11111001", -- 3303 - 0xce7  :  249 - 0xf9
    "00000000", -- 3304 - 0xce8  :    0 - 0x0 -- plane 1
    "00000000", -- 3305 - 0xce9  :    0 - 0x0
    "00000000", -- 3306 - 0xcea  :    0 - 0x0
    "00000000", -- 3307 - 0xceb  :    0 - 0x0
    "00000000", -- 3308 - 0xcec  :    0 - 0x0
    "00000110", -- 3309 - 0xced  :    6 - 0x6
    "00000100", -- 3310 - 0xcee  :    4 - 0x4
    "10000110", -- 3311 - 0xcef  :  134 - 0x86
    "11111110", -- 3312 - 0xcf0  :  254 - 0xfe -- Background 0xcf
    "11111000", -- 3313 - 0xcf1  :  248 - 0xf8
    "11111000", -- 3314 - 0xcf2  :  248 - 0xf8
    "11111000", -- 3315 - 0xcf3  :  248 - 0xf8
    "11110000", -- 3316 - 0xcf4  :  240 - 0xf0
    "11100000", -- 3317 - 0xcf5  :  224 - 0xe0
    "00000000", -- 3318 - 0xcf6  :    0 - 0x0
    "00000000", -- 3319 - 0xcf7  :    0 - 0x0
    "11000000", -- 3320 - 0xcf8  :  192 - 0xc0 -- plane 1
    "01100000", -- 3321 - 0xcf9  :   96 - 0x60
    "10100000", -- 3322 - 0xcfa  :  160 - 0xa0
    "11000000", -- 3323 - 0xcfb  :  192 - 0xc0
    "01000000", -- 3324 - 0xcfc  :   64 - 0x40
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00000000", -- 3328 - 0xd00  :    0 - 0x0 -- Background 0xd0
    "00000000", -- 3329 - 0xd01  :    0 - 0x0
    "00000100", -- 3330 - 0xd02  :    4 - 0x4
    "00100110", -- 3331 - 0xd03  :   38 - 0x26
    "00101011", -- 3332 - 0xd04  :   43 - 0x2b
    "01110001", -- 3333 - 0xd05  :  113 - 0x71
    "01000000", -- 3334 - 0xd06  :   64 - 0x40
    "01000111", -- 3335 - 0xd07  :   71 - 0x47
    "00000000", -- 3336 - 0xd08  :    0 - 0x0 -- plane 1
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "00000000", -- 3338 - 0xd0a  :    0 - 0x0
    "00000000", -- 3339 - 0xd0b  :    0 - 0x0
    "00000100", -- 3340 - 0xd0c  :    4 - 0x4
    "00001110", -- 3341 - 0xd0d  :   14 - 0xe
    "00111111", -- 3342 - 0xd0e  :   63 - 0x3f
    "00111001", -- 3343 - 0xd0f  :   57 - 0x39
    "10001111", -- 3344 - 0xd10  :  143 - 0x8f -- Background 0xd1
    "10001111", -- 3345 - 0xd11  :  143 - 0x8f
    "01001111", -- 3346 - 0xd12  :   79 - 0x4f
    "01001111", -- 3347 - 0xd13  :   79 - 0x4f
    "00111111", -- 3348 - 0xd14  :   63 - 0x3f
    "00010011", -- 3349 - 0xd15  :   19 - 0x13
    "00010001", -- 3350 - 0xd16  :   17 - 0x11
    "00011111", -- 3351 - 0xd17  :   31 - 0x1f
    "01110000", -- 3352 - 0xd18  :  112 - 0x70 -- plane 1
    "01111000", -- 3353 - 0xd19  :  120 - 0x78
    "00111111", -- 3354 - 0xd1a  :   63 - 0x3f
    "00111111", -- 3355 - 0xd1b  :   63 - 0x3f
    "00000011", -- 3356 - 0xd1c  :    3 - 0x3
    "00001100", -- 3357 - 0xd1d  :   12 - 0xc
    "00001110", -- 3358 - 0xd1e  :   14 - 0xe
    "00000000", -- 3359 - 0xd1f  :    0 - 0x0
    "00000000", -- 3360 - 0xd20  :    0 - 0x0 -- Background 0xd2
    "10000000", -- 3361 - 0xd21  :  128 - 0x80
    "11001000", -- 3362 - 0xd22  :  200 - 0xc8
    "11010100", -- 3363 - 0xd23  :  212 - 0xd4
    "00100100", -- 3364 - 0xd24  :   36 - 0x24
    "00000010", -- 3365 - 0xd25  :    2 - 0x2
    "00000010", -- 3366 - 0xd26  :    2 - 0x2
    "11110010", -- 3367 - 0xd27  :  242 - 0xf2
    "00000000", -- 3368 - 0xd28  :    0 - 0x0 -- plane 1
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "00000000", -- 3370 - 0xd2a  :    0 - 0x0
    "00001000", -- 3371 - 0xd2b  :    8 - 0x8
    "11011000", -- 3372 - 0xd2c  :  216 - 0xd8
    "11111100", -- 3373 - 0xd2d  :  252 - 0xfc
    "11111100", -- 3374 - 0xd2e  :  252 - 0xfc
    "10011100", -- 3375 - 0xd2f  :  156 - 0x9c
    "11110010", -- 3376 - 0xd30  :  242 - 0xf2 -- Background 0xd3
    "11110010", -- 3377 - 0xd31  :  242 - 0xf2
    "11110100", -- 3378 - 0xd32  :  244 - 0xf4
    "11110100", -- 3379 - 0xd33  :  244 - 0xf4
    "11110100", -- 3380 - 0xd34  :  244 - 0xf4
    "11001000", -- 3381 - 0xd35  :  200 - 0xc8
    "01000100", -- 3382 - 0xd36  :   68 - 0x44
    "01111100", -- 3383 - 0xd37  :  124 - 0x7c
    "00001100", -- 3384 - 0xd38  :   12 - 0xc -- plane 1
    "10011100", -- 3385 - 0xd39  :  156 - 0x9c
    "11111000", -- 3386 - 0xd3a  :  248 - 0xf8
    "01111000", -- 3387 - 0xd3b  :  120 - 0x78
    "10001000", -- 3388 - 0xd3c  :  136 - 0x88
    "00110000", -- 3389 - 0xd3d  :   48 - 0x30
    "00111000", -- 3390 - 0xd3e  :   56 - 0x38
    "00000000", -- 3391 - 0xd3f  :    0 - 0x0
    "00000000", -- 3392 - 0xd40  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 3393 - 0xd41  :    0 - 0x0
    "00000000", -- 3394 - 0xd42  :    0 - 0x0
    "00001001", -- 3395 - 0xd43  :    9 - 0x9
    "00011010", -- 3396 - 0xd44  :   26 - 0x1a
    "00010100", -- 3397 - 0xd45  :   20 - 0x14
    "00100000", -- 3398 - 0xd46  :   32 - 0x20
    "01000111", -- 3399 - 0xd47  :   71 - 0x47
    "00000000", -- 3400 - 0xd48  :    0 - 0x0 -- plane 1
    "00000000", -- 3401 - 0xd49  :    0 - 0x0
    "00000000", -- 3402 - 0xd4a  :    0 - 0x0
    "00000000", -- 3403 - 0xd4b  :    0 - 0x0
    "00000001", -- 3404 - 0xd4c  :    1 - 0x1
    "00001011", -- 3405 - 0xd4d  :   11 - 0xb
    "00011111", -- 3406 - 0xd4e  :   31 - 0x1f
    "00111001", -- 3407 - 0xd4f  :   57 - 0x39
    "10001111", -- 3408 - 0xd50  :  143 - 0x8f -- Background 0xd5
    "10001111", -- 3409 - 0xd51  :  143 - 0x8f
    "01001111", -- 3410 - 0xd52  :   79 - 0x4f
    "01001111", -- 3411 - 0xd53  :   79 - 0x4f
    "00111111", -- 3412 - 0xd54  :   63 - 0x3f
    "01000111", -- 3413 - 0xd55  :   71 - 0x47
    "00100010", -- 3414 - 0xd56  :   34 - 0x22
    "00011100", -- 3415 - 0xd57  :   28 - 0x1c
    "01110000", -- 3416 - 0xd58  :  112 - 0x70 -- plane 1
    "01111000", -- 3417 - 0xd59  :  120 - 0x78
    "00111111", -- 3418 - 0xd5a  :   63 - 0x3f
    "00111111", -- 3419 - 0xd5b  :   63 - 0x3f
    "00000011", -- 3420 - 0xd5c  :    3 - 0x3
    "00111000", -- 3421 - 0xd5d  :   56 - 0x38
    "00011100", -- 3422 - 0xd5e  :   28 - 0x1c
    "00000000", -- 3423 - 0xd5f  :    0 - 0x0
    "00000000", -- 3424 - 0xd60  :    0 - 0x0 -- Background 0xd6
    "01000000", -- 3425 - 0xd61  :   64 - 0x40
    "11000000", -- 3426 - 0xd62  :  192 - 0xc0
    "00101100", -- 3427 - 0xd63  :   44 - 0x2c
    "00110100", -- 3428 - 0xd64  :   52 - 0x34
    "00000100", -- 3429 - 0xd65  :    4 - 0x4
    "00000010", -- 3430 - 0xd66  :    2 - 0x2
    "11110010", -- 3431 - 0xd67  :  242 - 0xf2
    "00000000", -- 3432 - 0xd68  :    0 - 0x0 -- plane 1
    "00000000", -- 3433 - 0xd69  :    0 - 0x0
    "00000000", -- 3434 - 0xd6a  :    0 - 0x0
    "11000000", -- 3435 - 0xd6b  :  192 - 0xc0
    "11001000", -- 3436 - 0xd6c  :  200 - 0xc8
    "11111000", -- 3437 - 0xd6d  :  248 - 0xf8
    "11111100", -- 3438 - 0xd6e  :  252 - 0xfc
    "10011100", -- 3439 - 0xd6f  :  156 - 0x9c
    "11110010", -- 3440 - 0xd70  :  242 - 0xf2 -- Background 0xd7
    "11110010", -- 3441 - 0xd71  :  242 - 0xf2
    "11110100", -- 3442 - 0xd72  :  244 - 0xf4
    "11110111", -- 3443 - 0xd73  :  247 - 0xf7
    "11111101", -- 3444 - 0xd74  :  253 - 0xfd
    "11100001", -- 3445 - 0xd75  :  225 - 0xe1
    "00010010", -- 3446 - 0xd76  :   18 - 0x12
    "00001100", -- 3447 - 0xd77  :   12 - 0xc
    "00001100", -- 3448 - 0xd78  :   12 - 0xc -- plane 1
    "10011100", -- 3449 - 0xd79  :  156 - 0x9c
    "11111000", -- 3450 - 0xd7a  :  248 - 0xf8
    "01111000", -- 3451 - 0xd7b  :  120 - 0x78
    "11100010", -- 3452 - 0xd7c  :  226 - 0xe2
    "00011110", -- 3453 - 0xd7d  :   30 - 0x1e
    "00001100", -- 3454 - 0xd7e  :   12 - 0xc
    "00000000", -- 3455 - 0xd7f  :    0 - 0x0
    "01111000", -- 3456 - 0xd80  :  120 - 0x78 -- Background 0xd8
    "01001110", -- 3457 - 0xd81  :   78 - 0x4e
    "11000010", -- 3458 - 0xd82  :  194 - 0xc2
    "10011010", -- 3459 - 0xd83  :  154 - 0x9a
    "10011011", -- 3460 - 0xd84  :  155 - 0x9b
    "11011001", -- 3461 - 0xd85  :  217 - 0xd9
    "01100011", -- 3462 - 0xd86  :   99 - 0x63
    "00111110", -- 3463 - 0xd87  :   62 - 0x3e
    "00000000", -- 3464 - 0xd88  :    0 - 0x0 -- plane 1
    "00110000", -- 3465 - 0xd89  :   48 - 0x30
    "00111100", -- 3466 - 0xd8a  :   60 - 0x3c
    "01111100", -- 3467 - 0xd8b  :  124 - 0x7c
    "01111100", -- 3468 - 0xd8c  :  124 - 0x7c
    "00111110", -- 3469 - 0xd8d  :   62 - 0x3e
    "00011100", -- 3470 - 0xd8e  :   28 - 0x1c
    "00000000", -- 3471 - 0xd8f  :    0 - 0x0
    "00011110", -- 3472 - 0xd90  :   30 - 0x1e -- Background 0xd9
    "01110001", -- 3473 - 0xd91  :  113 - 0x71
    "01001001", -- 3474 - 0xd92  :   73 - 0x49
    "10111001", -- 3475 - 0xd93  :  185 - 0xb9
    "10011101", -- 3476 - 0xd94  :  157 - 0x9d
    "01010010", -- 3477 - 0xd95  :   82 - 0x52
    "01110010", -- 3478 - 0xd96  :  114 - 0x72
    "00011110", -- 3479 - 0xd97  :   30 - 0x1e
    "00000000", -- 3480 - 0xd98  :    0 - 0x0 -- plane 1
    "00001110", -- 3481 - 0xd99  :   14 - 0xe
    "00111110", -- 3482 - 0xd9a  :   62 - 0x3e
    "01111110", -- 3483 - 0xd9b  :  126 - 0x7e
    "01111110", -- 3484 - 0xd9c  :  126 - 0x7e
    "00111100", -- 3485 - 0xd9d  :   60 - 0x3c
    "00001100", -- 3486 - 0xd9e  :   12 - 0xc
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "01100000", -- 3488 - 0xda0  :   96 - 0x60 -- Background 0xda
    "01011110", -- 3489 - 0xda1  :   94 - 0x5e
    "10001001", -- 3490 - 0xda2  :  137 - 0x89
    "10111101", -- 3491 - 0xda3  :  189 - 0xbd
    "10011101", -- 3492 - 0xda4  :  157 - 0x9d
    "11010011", -- 3493 - 0xda5  :  211 - 0xd3
    "01000110", -- 3494 - 0xda6  :   70 - 0x46
    "01111100", -- 3495 - 0xda7  :  124 - 0x7c
    "00000000", -- 3496 - 0xda8  :    0 - 0x0 -- plane 1
    "00100000", -- 3497 - 0xda9  :   32 - 0x20
    "01111110", -- 3498 - 0xdaa  :  126 - 0x7e
    "01111110", -- 3499 - 0xdab  :  126 - 0x7e
    "01111110", -- 3500 - 0xdac  :  126 - 0x7e
    "00111100", -- 3501 - 0xdad  :   60 - 0x3c
    "00111000", -- 3502 - 0xdae  :   56 - 0x38
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00011110", -- 3504 - 0xdb0  :   30 - 0x1e -- Background 0xdb
    "00100011", -- 3505 - 0xdb1  :   35 - 0x23
    "01001001", -- 3506 - 0xdb2  :   73 - 0x49
    "10111101", -- 3507 - 0xdb3  :  189 - 0xbd
    "10011001", -- 3508 - 0xdb4  :  153 - 0x99
    "01000011", -- 3509 - 0xdb5  :   67 - 0x43
    "01101110", -- 3510 - 0xdb6  :  110 - 0x6e
    "00011000", -- 3511 - 0xdb7  :   24 - 0x18
    "00000000", -- 3512 - 0xdb8  :    0 - 0x0 -- plane 1
    "00011100", -- 3513 - 0xdb9  :   28 - 0x1c
    "00111110", -- 3514 - 0xdba  :   62 - 0x3e
    "01111110", -- 3515 - 0xdbb  :  126 - 0x7e
    "01111110", -- 3516 - 0xdbc  :  126 - 0x7e
    "00111100", -- 3517 - 0xdbd  :   60 - 0x3c
    "00010000", -- 3518 - 0xdbe  :   16 - 0x10
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 3521 - 0xdc1  :    0 - 0x0
    "00000001", -- 3522 - 0xdc2  :    1 - 0x1
    "00000010", -- 3523 - 0xdc3  :    2 - 0x2
    "00000100", -- 3524 - 0xdc4  :    4 - 0x4
    "00000010", -- 3525 - 0xdc5  :    2 - 0x2
    "00011110", -- 3526 - 0xdc6  :   30 - 0x1e
    "00010000", -- 3527 - 0xdc7  :   16 - 0x10
    "00000000", -- 3528 - 0xdc8  :    0 - 0x0 -- plane 1
    "00000000", -- 3529 - 0xdc9  :    0 - 0x0
    "00000000", -- 3530 - 0xdca  :    0 - 0x0
    "00000001", -- 3531 - 0xdcb  :    1 - 0x1
    "00000011", -- 3532 - 0xdcc  :    3 - 0x3
    "00000001", -- 3533 - 0xdcd  :    1 - 0x1
    "00000001", -- 3534 - 0xdce  :    1 - 0x1
    "00001111", -- 3535 - 0xdcf  :   15 - 0xf
    "00001000", -- 3536 - 0xdd0  :    8 - 0x8 -- Background 0xdd
    "00001101", -- 3537 - 0xdd1  :   13 - 0xd
    "00111010", -- 3538 - 0xdd2  :   58 - 0x3a
    "00100101", -- 3539 - 0xdd3  :   37 - 0x25
    "00011011", -- 3540 - 0xdd4  :   27 - 0x1b
    "00001111", -- 3541 - 0xdd5  :   15 - 0xf
    "00000111", -- 3542 - 0xdd6  :    7 - 0x7
    "00000011", -- 3543 - 0xdd7  :    3 - 0x3
    "00000111", -- 3544 - 0xdd8  :    7 - 0x7 -- plane 1
    "00000111", -- 3545 - 0xdd9  :    7 - 0x7
    "00000111", -- 3546 - 0xdda  :    7 - 0x7
    "00011111", -- 3547 - 0xddb  :   31 - 0x1f
    "00001111", -- 3548 - 0xddc  :   15 - 0xf
    "00000111", -- 3549 - 0xddd  :    7 - 0x7
    "00000011", -- 3550 - 0xdde  :    3 - 0x3
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "00000000", -- 3552 - 0xde0  :    0 - 0x0 -- Background 0xde
    "00000000", -- 3553 - 0xde1  :    0 - 0x0
    "00000000", -- 3554 - 0xde2  :    0 - 0x0
    "11000000", -- 3555 - 0xde3  :  192 - 0xc0
    "01000000", -- 3556 - 0xde4  :   64 - 0x40
    "01011000", -- 3557 - 0xde5  :   88 - 0x58
    "01101000", -- 3558 - 0xde6  :  104 - 0x68
    "00001000", -- 3559 - 0xde7  :    8 - 0x8
    "00000000", -- 3560 - 0xde8  :    0 - 0x0 -- plane 1
    "00000000", -- 3561 - 0xde9  :    0 - 0x0
    "00000000", -- 3562 - 0xdea  :    0 - 0x0
    "00000000", -- 3563 - 0xdeb  :    0 - 0x0
    "10000000", -- 3564 - 0xdec  :  128 - 0x80
    "10000000", -- 3565 - 0xded  :  128 - 0x80
    "10010000", -- 3566 - 0xdee  :  144 - 0x90
    "11110000", -- 3567 - 0xdef  :  240 - 0xf0
    "00010000", -- 3568 - 0xdf0  :   16 - 0x10 -- Background 0xdf
    "01011100", -- 3569 - 0xdf1  :   92 - 0x5c
    "10101000", -- 3570 - 0xdf2  :  168 - 0xa8
    "11011000", -- 3571 - 0xdf3  :  216 - 0xd8
    "10111000", -- 3572 - 0xdf4  :  184 - 0xb8
    "11110000", -- 3573 - 0xdf5  :  240 - 0xf0
    "11100000", -- 3574 - 0xdf6  :  224 - 0xe0
    "11000000", -- 3575 - 0xdf7  :  192 - 0xc0
    "11100000", -- 3576 - 0xdf8  :  224 - 0xe0 -- plane 1
    "11100000", -- 3577 - 0xdf9  :  224 - 0xe0
    "11110000", -- 3578 - 0xdfa  :  240 - 0xf0
    "11110000", -- 3579 - 0xdfb  :  240 - 0xf0
    "11100000", -- 3580 - 0xdfc  :  224 - 0xe0
    "11000000", -- 3581 - 0xdfd  :  192 - 0xc0
    "11000000", -- 3582 - 0xdfe  :  192 - 0xc0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "00000000", -- 3584 - 0xe00  :    0 - 0x0 -- Background 0xe0
    "00000000", -- 3585 - 0xe01  :    0 - 0x0
    "00000000", -- 3586 - 0xe02  :    0 - 0x0
    "00010011", -- 3587 - 0xe03  :   19 - 0x13
    "00010011", -- 3588 - 0xe04  :   19 - 0x13
    "00110111", -- 3589 - 0xe05  :   55 - 0x37
    "00110111", -- 3590 - 0xe06  :   55 - 0x37
    "00000111", -- 3591 - 0xe07  :    7 - 0x7
    "00001111", -- 3592 - 0xe08  :   15 - 0xf -- plane 1
    "00011111", -- 3593 - 0xe09  :   31 - 0x1f
    "00011111", -- 3594 - 0xe0a  :   31 - 0x1f
    "00111111", -- 3595 - 0xe0b  :   63 - 0x3f
    "01111111", -- 3596 - 0xe0c  :  127 - 0x7f
    "11111111", -- 3597 - 0xe0d  :  255 - 0xff
    "11111111", -- 3598 - 0xe0e  :  255 - 0xff
    "11111111", -- 3599 - 0xe0f  :  255 - 0xff
    "00000111", -- 3600 - 0xe10  :    7 - 0x7 -- Background 0xe1
    "00000100", -- 3601 - 0xe11  :    4 - 0x4
    "00000000", -- 3602 - 0xe12  :    0 - 0x0
    "00000000", -- 3603 - 0xe13  :    0 - 0x0
    "00000000", -- 3604 - 0xe14  :    0 - 0x0
    "00100000", -- 3605 - 0xe15  :   32 - 0x20
    "01110000", -- 3606 - 0xe16  :  112 - 0x70
    "11111000", -- 3607 - 0xe17  :  248 - 0xf8
    "11111111", -- 3608 - 0xe18  :  255 - 0xff -- plane 1
    "11111111", -- 3609 - 0xe19  :  255 - 0xff
    "01111111", -- 3610 - 0xe1a  :  127 - 0x7f
    "00111111", -- 3611 - 0xe1b  :   63 - 0x3f
    "00111111", -- 3612 - 0xe1c  :   63 - 0x3f
    "00011111", -- 3613 - 0xe1d  :   31 - 0x1f
    "00001111", -- 3614 - 0xe1e  :   15 - 0xf
    "00000111", -- 3615 - 0xe1f  :    7 - 0x7
    "00000000", -- 3616 - 0xe20  :    0 - 0x0 -- Background 0xe2
    "00000000", -- 3617 - 0xe21  :    0 - 0x0
    "00000000", -- 3618 - 0xe22  :    0 - 0x0
    "11111000", -- 3619 - 0xe23  :  248 - 0xf8
    "11111100", -- 3620 - 0xe24  :  252 - 0xfc
    "11111100", -- 3621 - 0xe25  :  252 - 0xfc
    "11111100", -- 3622 - 0xe26  :  252 - 0xfc
    "11111101", -- 3623 - 0xe27  :  253 - 0xfd
    "11111110", -- 3624 - 0xe28  :  254 - 0xfe -- plane 1
    "11111111", -- 3625 - 0xe29  :  255 - 0xff
    "11111111", -- 3626 - 0xe2a  :  255 - 0xff
    "00001111", -- 3627 - 0xe2b  :   15 - 0xf
    "10111111", -- 3628 - 0xe2c  :  191 - 0xbf
    "10100011", -- 3629 - 0xe2d  :  163 - 0xa3
    "11110111", -- 3630 - 0xe2e  :  247 - 0xf7
    "11110111", -- 3631 - 0xe2f  :  247 - 0xf7
    "11111100", -- 3632 - 0xe30  :  252 - 0xfc -- Background 0xe3
    "00011100", -- 3633 - 0xe31  :   28 - 0x1c
    "11000000", -- 3634 - 0xe32  :  192 - 0xc0
    "11100000", -- 3635 - 0xe33  :  224 - 0xe0
    "00000000", -- 3636 - 0xe34  :    0 - 0x0
    "00000000", -- 3637 - 0xe35  :    0 - 0x0
    "00000110", -- 3638 - 0xe36  :    6 - 0x6
    "00001111", -- 3639 - 0xe37  :   15 - 0xf
    "11111111", -- 3640 - 0xe38  :  255 - 0xff -- plane 1
    "11111111", -- 3641 - 0xe39  :  255 - 0xff
    "00111111", -- 3642 - 0xe3a  :   63 - 0x3f
    "00011111", -- 3643 - 0xe3b  :   31 - 0x1f
    "11111110", -- 3644 - 0xe3c  :  254 - 0xfe
    "11111100", -- 3645 - 0xe3d  :  252 - 0xfc
    "11111000", -- 3646 - 0xe3e  :  248 - 0xf8
    "11110000", -- 3647 - 0xe3f  :  240 - 0xf0
    "00000000", -- 3648 - 0xe40  :    0 - 0x0 -- Background 0xe4
    "00000000", -- 3649 - 0xe41  :    0 - 0x0
    "00000000", -- 3650 - 0xe42  :    0 - 0x0
    "00010011", -- 3651 - 0xe43  :   19 - 0x13
    "00010011", -- 3652 - 0xe44  :   19 - 0x13
    "00110111", -- 3653 - 0xe45  :   55 - 0x37
    "00110111", -- 3654 - 0xe46  :   55 - 0x37
    "00000111", -- 3655 - 0xe47  :    7 - 0x7
    "00001111", -- 3656 - 0xe48  :   15 - 0xf -- plane 1
    "00011111", -- 3657 - 0xe49  :   31 - 0x1f
    "00011111", -- 3658 - 0xe4a  :   31 - 0x1f
    "00111111", -- 3659 - 0xe4b  :   63 - 0x3f
    "01111111", -- 3660 - 0xe4c  :  127 - 0x7f
    "11111111", -- 3661 - 0xe4d  :  255 - 0xff
    "11111111", -- 3662 - 0xe4e  :  255 - 0xff
    "11111111", -- 3663 - 0xe4f  :  255 - 0xff
    "00000111", -- 3664 - 0xe50  :    7 - 0x7 -- Background 0xe5
    "00000100", -- 3665 - 0xe51  :    4 - 0x4
    "00000001", -- 3666 - 0xe52  :    1 - 0x1
    "00000000", -- 3667 - 0xe53  :    0 - 0x0
    "00000000", -- 3668 - 0xe54  :    0 - 0x0
    "00100000", -- 3669 - 0xe55  :   32 - 0x20
    "01110000", -- 3670 - 0xe56  :  112 - 0x70
    "11111000", -- 3671 - 0xe57  :  248 - 0xf8
    "11111111", -- 3672 - 0xe58  :  255 - 0xff -- plane 1
    "11111111", -- 3673 - 0xe59  :  255 - 0xff
    "01111110", -- 3674 - 0xe5a  :  126 - 0x7e
    "00111111", -- 3675 - 0xe5b  :   63 - 0x3f
    "00111111", -- 3676 - 0xe5c  :   63 - 0x3f
    "00011111", -- 3677 - 0xe5d  :   31 - 0x1f
    "00001111", -- 3678 - 0xe5e  :   15 - 0xf
    "00000111", -- 3679 - 0xe5f  :    7 - 0x7
    "00000000", -- 3680 - 0xe60  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 3681 - 0xe61  :    0 - 0x0
    "00000000", -- 3682 - 0xe62  :    0 - 0x0
    "11111100", -- 3683 - 0xe63  :  252 - 0xfc
    "11111100", -- 3684 - 0xe64  :  252 - 0xfc
    "11111100", -- 3685 - 0xe65  :  252 - 0xfc
    "11111100", -- 3686 - 0xe66  :  252 - 0xfc
    "11111101", -- 3687 - 0xe67  :  253 - 0xfd
    "11111110", -- 3688 - 0xe68  :  254 - 0xfe -- plane 1
    "11111111", -- 3689 - 0xe69  :  255 - 0xff
    "11111111", -- 3690 - 0xe6a  :  255 - 0xff
    "11100011", -- 3691 - 0xe6b  :  227 - 0xe3
    "00010111", -- 3692 - 0xe6c  :   23 - 0x17
    "10110111", -- 3693 - 0xe6d  :  183 - 0xb7
    "10111111", -- 3694 - 0xe6e  :  191 - 0xbf
    "11111111", -- 3695 - 0xe6f  :  255 - 0xff
    "11111100", -- 3696 - 0xe70  :  252 - 0xfc -- Background 0xe7
    "00001100", -- 3697 - 0xe71  :   12 - 0xc
    "11000000", -- 3698 - 0xe72  :  192 - 0xc0
    "11110000", -- 3699 - 0xe73  :  240 - 0xf0
    "11110000", -- 3700 - 0xe74  :  240 - 0xf0
    "00000000", -- 3701 - 0xe75  :    0 - 0x0
    "00000110", -- 3702 - 0xe76  :    6 - 0x6
    "00001111", -- 3703 - 0xe77  :   15 - 0xf
    "11111111", -- 3704 - 0xe78  :  255 - 0xff -- plane 1
    "11111111", -- 3705 - 0xe79  :  255 - 0xff
    "00111111", -- 3706 - 0xe7a  :   63 - 0x3f
    "00001111", -- 3707 - 0xe7b  :   15 - 0xf
    "00001110", -- 3708 - 0xe7c  :   14 - 0xe
    "11111100", -- 3709 - 0xe7d  :  252 - 0xfc
    "11111000", -- 3710 - 0xe7e  :  248 - 0xf8
    "11110000", -- 3711 - 0xe7f  :  240 - 0xf0
    "11111111", -- 3712 - 0xe80  :  255 - 0xff -- Background 0xe8
    "11111111", -- 3713 - 0xe81  :  255 - 0xff
    "01111111", -- 3714 - 0xe82  :  127 - 0x7f
    "01111111", -- 3715 - 0xe83  :  127 - 0x7f
    "01111111", -- 3716 - 0xe84  :  127 - 0x7f
    "00111111", -- 3717 - 0xe85  :   63 - 0x3f
    "00111111", -- 3718 - 0xe86  :   63 - 0x3f
    "00111111", -- 3719 - 0xe87  :   63 - 0x3f
    "00000000", -- 3720 - 0xe88  :    0 - 0x0 -- plane 1
    "00000101", -- 3721 - 0xe89  :    5 - 0x5
    "00000111", -- 3722 - 0xe8a  :    7 - 0x7
    "00000011", -- 3723 - 0xe8b  :    3 - 0x3
    "00000000", -- 3724 - 0xe8c  :    0 - 0x0
    "00000000", -- 3725 - 0xe8d  :    0 - 0x0
    "00000000", -- 3726 - 0xe8e  :    0 - 0x0
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "00111100", -- 3728 - 0xe90  :   60 - 0x3c -- Background 0xe9
    "00111110", -- 3729 - 0xe91  :   62 - 0x3e
    "00011111", -- 3730 - 0xe92  :   31 - 0x1f
    "00001111", -- 3731 - 0xe93  :   15 - 0xf
    "00000111", -- 3732 - 0xe94  :    7 - 0x7
    "00000000", -- 3733 - 0xe95  :    0 - 0x0
    "00000000", -- 3734 - 0xe96  :    0 - 0x0
    "00000000", -- 3735 - 0xe97  :    0 - 0x0
    "00000000", -- 3736 - 0xe98  :    0 - 0x0 -- plane 1
    "00000000", -- 3737 - 0xe99  :    0 - 0x0
    "00000000", -- 3738 - 0xe9a  :    0 - 0x0
    "00000000", -- 3739 - 0xe9b  :    0 - 0x0
    "00000000", -- 3740 - 0xe9c  :    0 - 0x0
    "00000000", -- 3741 - 0xe9d  :    0 - 0x0
    "00000000", -- 3742 - 0xe9e  :    0 - 0x0
    "00000000", -- 3743 - 0xe9f  :    0 - 0x0
    "11111111", -- 3744 - 0xea0  :  255 - 0xff -- Background 0xea
    "11111110", -- 3745 - 0xea1  :  254 - 0xfe
    "11111110", -- 3746 - 0xea2  :  254 - 0xfe
    "11111100", -- 3747 - 0xea3  :  252 - 0xfc
    "11111000", -- 3748 - 0xea4  :  248 - 0xf8
    "11110000", -- 3749 - 0xea5  :  240 - 0xf0
    "10110000", -- 3750 - 0xea6  :  176 - 0xb0
    "00111001", -- 3751 - 0xea7  :   57 - 0x39
    "00000011", -- 3752 - 0xea8  :    3 - 0x3 -- plane 1
    "10011110", -- 3753 - 0xea9  :  158 - 0x9e
    "00001110", -- 3754 - 0xeaa  :   14 - 0xe
    "00000000", -- 3755 - 0xeab  :    0 - 0x0
    "00000000", -- 3756 - 0xeac  :    0 - 0x0
    "00000000", -- 3757 - 0xead  :    0 - 0x0
    "00000000", -- 3758 - 0xeae  :    0 - 0x0
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "00011111", -- 3760 - 0xeb0  :   31 - 0x1f -- Background 0xeb
    "11001111", -- 3761 - 0xeb1  :  207 - 0xcf
    "11000110", -- 3762 - 0xeb2  :  198 - 0xc6
    "10000000", -- 3763 - 0xeb3  :  128 - 0x80
    "00000000", -- 3764 - 0xeb4  :    0 - 0x0
    "00000000", -- 3765 - 0xeb5  :    0 - 0x0
    "00000000", -- 3766 - 0xeb6  :    0 - 0x0
    "00000000", -- 3767 - 0xeb7  :    0 - 0x0
    "00000000", -- 3768 - 0xeb8  :    0 - 0x0 -- plane 1
    "00000000", -- 3769 - 0xeb9  :    0 - 0x0
    "00000000", -- 3770 - 0xeba  :    0 - 0x0
    "00000000", -- 3771 - 0xebb  :    0 - 0x0
    "00000000", -- 3772 - 0xebc  :    0 - 0x0
    "00000000", -- 3773 - 0xebd  :    0 - 0x0
    "00000000", -- 3774 - 0xebe  :    0 - 0x0
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Background 0xec
    "00000000", -- 3777 - 0xec1  :    0 - 0x0
    "00000000", -- 3778 - 0xec2  :    0 - 0x0
    "00000000", -- 3779 - 0xec3  :    0 - 0x0
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00000000", -- 3781 - 0xec5  :    0 - 0x0
    "00001100", -- 3782 - 0xec6  :   12 - 0xc
    "00001100", -- 3783 - 0xec7  :   12 - 0xc
    "00000000", -- 3784 - 0xec8  :    0 - 0x0 -- plane 1
    "00000000", -- 3785 - 0xec9  :    0 - 0x0
    "00000000", -- 3786 - 0xeca  :    0 - 0x0
    "00000000", -- 3787 - 0xecb  :    0 - 0x0
    "00000100", -- 3788 - 0xecc  :    4 - 0x4
    "00001110", -- 3789 - 0xecd  :   14 - 0xe
    "00001111", -- 3790 - 0xece  :   15 - 0xf
    "00001011", -- 3791 - 0xecf  :   11 - 0xb
    "00110000", -- 3792 - 0xed0  :   48 - 0x30 -- Background 0xed
    "01000011", -- 3793 - 0xed1  :   67 - 0x43
    "01000000", -- 3794 - 0xed2  :   64 - 0x40
    "01100000", -- 3795 - 0xed3  :   96 - 0x60
    "00000011", -- 3796 - 0xed4  :    3 - 0x3
    "00000000", -- 3797 - 0xed5  :    0 - 0x0
    "01111111", -- 3798 - 0xed6  :  127 - 0x7f
    "00000000", -- 3799 - 0xed7  :    0 - 0x0
    "00001111", -- 3800 - 0xed8  :   15 - 0xf -- plane 1
    "00001100", -- 3801 - 0xed9  :   12 - 0xc
    "00001111", -- 3802 - 0xeda  :   15 - 0xf
    "00001111", -- 3803 - 0xedb  :   15 - 0xf
    "00000000", -- 3804 - 0xedc  :    0 - 0x0
    "01111111", -- 3805 - 0xedd  :  127 - 0x7f
    "11010101", -- 3806 - 0xede  :  213 - 0xd5
    "01111111", -- 3807 - 0xedf  :  127 - 0x7f
    "00000000", -- 3808 - 0xee0  :    0 - 0x0 -- Background 0xee
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000000", -- 3811 - 0xee3  :    0 - 0x0
    "00000000", -- 3812 - 0xee4  :    0 - 0x0
    "00000000", -- 3813 - 0xee5  :    0 - 0x0
    "00110000", -- 3814 - 0xee6  :   48 - 0x30
    "00110000", -- 3815 - 0xee7  :   48 - 0x30
    "00000000", -- 3816 - 0xee8  :    0 - 0x0 -- plane 1
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "00000000", -- 3818 - 0xeea  :    0 - 0x0
    "00000000", -- 3819 - 0xeeb  :    0 - 0x0
    "00100000", -- 3820 - 0xeec  :   32 - 0x20
    "01110000", -- 3821 - 0xeed  :  112 - 0x70
    "11110000", -- 3822 - 0xeee  :  240 - 0xf0
    "11100000", -- 3823 - 0xeef  :  224 - 0xe0
    "00001110", -- 3824 - 0xef0  :   14 - 0xe -- Background 0xef
    "11001011", -- 3825 - 0xef1  :  203 - 0xcb
    "00000000", -- 3826 - 0xef2  :    0 - 0x0
    "00000000", -- 3827 - 0xef3  :    0 - 0x0
    "11000000", -- 3828 - 0xef4  :  192 - 0xc0
    "00000000", -- 3829 - 0xef5  :    0 - 0x0
    "11111110", -- 3830 - 0xef6  :  254 - 0xfe
    "00000000", -- 3831 - 0xef7  :    0 - 0x0
    "11110000", -- 3832 - 0xef8  :  240 - 0xf0 -- plane 1
    "00110000", -- 3833 - 0xef9  :   48 - 0x30
    "11110000", -- 3834 - 0xefa  :  240 - 0xf0
    "11110000", -- 3835 - 0xefb  :  240 - 0xf0
    "00000000", -- 3836 - 0xefc  :    0 - 0x0
    "11111110", -- 3837 - 0xefd  :  254 - 0xfe
    "01010101", -- 3838 - 0xefe  :   85 - 0x55
    "11111110", -- 3839 - 0xeff  :  254 - 0xfe
    "00000000", -- 3840 - 0xf00  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 3841 - 0xf01  :    0 - 0x0
    "00000000", -- 3842 - 0xf02  :    0 - 0x0
    "00000000", -- 3843 - 0xf03  :    0 - 0x0
    "00000000", -- 3844 - 0xf04  :    0 - 0x0
    "00000000", -- 3845 - 0xf05  :    0 - 0x0
    "00001100", -- 3846 - 0xf06  :   12 - 0xc
    "00001100", -- 3847 - 0xf07  :   12 - 0xc
    "00000000", -- 3848 - 0xf08  :    0 - 0x0 -- plane 1
    "00000000", -- 3849 - 0xf09  :    0 - 0x0
    "00000000", -- 3850 - 0xf0a  :    0 - 0x0
    "00000000", -- 3851 - 0xf0b  :    0 - 0x0
    "00000100", -- 3852 - 0xf0c  :    4 - 0x4
    "00001110", -- 3853 - 0xf0d  :   14 - 0xe
    "00001111", -- 3854 - 0xf0e  :   15 - 0xf
    "00001011", -- 3855 - 0xf0f  :   11 - 0xb
    "00110000", -- 3856 - 0xf10  :   48 - 0x30 -- Background 0xf1
    "00100011", -- 3857 - 0xf11  :   35 - 0x23
    "00100000", -- 3858 - 0xf12  :   32 - 0x20
    "01100000", -- 3859 - 0xf13  :   96 - 0x60
    "00000011", -- 3860 - 0xf14  :    3 - 0x3
    "00000000", -- 3861 - 0xf15  :    0 - 0x0
    "01111111", -- 3862 - 0xf16  :  127 - 0x7f
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "00001111", -- 3864 - 0xf18  :   15 - 0xf -- plane 1
    "00001100", -- 3865 - 0xf19  :   12 - 0xc
    "00001111", -- 3866 - 0xf1a  :   15 - 0xf
    "00001111", -- 3867 - 0xf1b  :   15 - 0xf
    "00000000", -- 3868 - 0xf1c  :    0 - 0x0
    "01111111", -- 3869 - 0xf1d  :  127 - 0x7f
    "10101010", -- 3870 - 0xf1e  :  170 - 0xaa
    "01111111", -- 3871 - 0xf1f  :  127 - 0x7f
    "00000000", -- 3872 - 0xf20  :    0 - 0x0 -- Background 0xf2
    "00000000", -- 3873 - 0xf21  :    0 - 0x0
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000000", -- 3876 - 0xf24  :    0 - 0x0
    "00000000", -- 3877 - 0xf25  :    0 - 0x0
    "00110000", -- 3878 - 0xf26  :   48 - 0x30
    "00110000", -- 3879 - 0xf27  :   48 - 0x30
    "00000000", -- 3880 - 0xf28  :    0 - 0x0 -- plane 1
    "00000000", -- 3881 - 0xf29  :    0 - 0x0
    "00000000", -- 3882 - 0xf2a  :    0 - 0x0
    "00000000", -- 3883 - 0xf2b  :    0 - 0x0
    "00100000", -- 3884 - 0xf2c  :   32 - 0x20
    "01110000", -- 3885 - 0xf2d  :  112 - 0x70
    "11110000", -- 3886 - 0xf2e  :  240 - 0xf0
    "11100000", -- 3887 - 0xf2f  :  224 - 0xe0
    "00001001", -- 3888 - 0xf30  :    9 - 0x9 -- Background 0xf3
    "11001111", -- 3889 - 0xf31  :  207 - 0xcf
    "00000000", -- 3890 - 0xf32  :    0 - 0x0
    "00000000", -- 3891 - 0xf33  :    0 - 0x0
    "11000000", -- 3892 - 0xf34  :  192 - 0xc0
    "00000000", -- 3893 - 0xf35  :    0 - 0x0
    "11111110", -- 3894 - 0xf36  :  254 - 0xfe
    "00000000", -- 3895 - 0xf37  :    0 - 0x0
    "11110000", -- 3896 - 0xf38  :  240 - 0xf0 -- plane 1
    "00110000", -- 3897 - 0xf39  :   48 - 0x30
    "11110000", -- 3898 - 0xf3a  :  240 - 0xf0
    "11110000", -- 3899 - 0xf3b  :  240 - 0xf0
    "00000000", -- 3900 - 0xf3c  :    0 - 0x0
    "11111110", -- 3901 - 0xf3d  :  254 - 0xfe
    "10101011", -- 3902 - 0xf3e  :  171 - 0xab
    "11111110", -- 3903 - 0xf3f  :  254 - 0xfe
    "00111111", -- 3904 - 0xf40  :   63 - 0x3f -- Background 0xf4
    "00110101", -- 3905 - 0xf41  :   53 - 0x35
    "00011010", -- 3906 - 0xf42  :   26 - 0x1a
    "00001101", -- 3907 - 0xf43  :   13 - 0xd
    "00001010", -- 3908 - 0xf44  :   10 - 0xa
    "00001101", -- 3909 - 0xf45  :   13 - 0xd
    "00001000", -- 3910 - 0xf46  :    8 - 0x8
    "00111000", -- 3911 - 0xf47  :   56 - 0x38
    "00000000", -- 3912 - 0xf48  :    0 - 0x0 -- plane 1
    "00010101", -- 3913 - 0xf49  :   21 - 0x15
    "00001010", -- 3914 - 0xf4a  :   10 - 0xa
    "00000101", -- 3915 - 0xf4b  :    5 - 0x5
    "00000010", -- 3916 - 0xf4c  :    2 - 0x2
    "00000101", -- 3917 - 0xf4d  :    5 - 0x5
    "00000111", -- 3918 - 0xf4e  :    7 - 0x7
    "00000111", -- 3919 - 0xf4f  :    7 - 0x7
    "01110011", -- 3920 - 0xf50  :  115 - 0x73 -- Background 0xf5
    "11000100", -- 3921 - 0xf51  :  196 - 0xc4
    "11000100", -- 3922 - 0xf52  :  196 - 0xc4
    "11000000", -- 3923 - 0xf53  :  192 - 0xc0
    "11000001", -- 3924 - 0xf54  :  193 - 0xc1
    "11000000", -- 3925 - 0xf55  :  192 - 0xc0
    "01100001", -- 3926 - 0xf56  :   97 - 0x61
    "00111111", -- 3927 - 0xf57  :   63 - 0x3f
    "00111100", -- 3928 - 0xf58  :   60 - 0x3c -- plane 1
    "01111011", -- 3929 - 0xf59  :  123 - 0x7b
    "01111011", -- 3930 - 0xf5a  :  123 - 0x7b
    "01111111", -- 3931 - 0xf5b  :  127 - 0x7f
    "01111110", -- 3932 - 0xf5c  :  126 - 0x7e
    "01111111", -- 3933 - 0xf5d  :  127 - 0x7f
    "00111110", -- 3934 - 0xf5e  :   62 - 0x3e
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "11111100", -- 3936 - 0xf60  :  252 - 0xfc -- Background 0xf6
    "01010100", -- 3937 - 0xf61  :   84 - 0x54
    "10101000", -- 3938 - 0xf62  :  168 - 0xa8
    "01010000", -- 3939 - 0xf63  :   80 - 0x50
    "10110000", -- 3940 - 0xf64  :  176 - 0xb0
    "01010000", -- 3941 - 0xf65  :   80 - 0x50
    "10010000", -- 3942 - 0xf66  :  144 - 0x90
    "00011100", -- 3943 - 0xf67  :   28 - 0x1c
    "00000000", -- 3944 - 0xf68  :    0 - 0x0 -- plane 1
    "01010000", -- 3945 - 0xf69  :   80 - 0x50
    "10100000", -- 3946 - 0xf6a  :  160 - 0xa0
    "01000000", -- 3947 - 0xf6b  :   64 - 0x40
    "10100000", -- 3948 - 0xf6c  :  160 - 0xa0
    "01000000", -- 3949 - 0xf6d  :   64 - 0x40
    "11100000", -- 3950 - 0xf6e  :  224 - 0xe0
    "11100000", -- 3951 - 0xf6f  :  224 - 0xe0
    "10000110", -- 3952 - 0xf70  :  134 - 0x86 -- Background 0xf7
    "01000010", -- 3953 - 0xf71  :   66 - 0x42
    "01000111", -- 3954 - 0xf72  :   71 - 0x47
    "01000001", -- 3955 - 0xf73  :   65 - 0x41
    "10000011", -- 3956 - 0xf74  :  131 - 0x83
    "00000001", -- 3957 - 0xf75  :    1 - 0x1
    "10000110", -- 3958 - 0xf76  :  134 - 0x86
    "11111100", -- 3959 - 0xf77  :  252 - 0xfc
    "01111000", -- 3960 - 0xf78  :  120 - 0x78 -- plane 1
    "10111100", -- 3961 - 0xf79  :  188 - 0xbc
    "10111000", -- 3962 - 0xf7a  :  184 - 0xb8
    "10111110", -- 3963 - 0xf7b  :  190 - 0xbe
    "01111100", -- 3964 - 0xf7c  :  124 - 0x7c
    "11111110", -- 3965 - 0xf7d  :  254 - 0xfe
    "01111000", -- 3966 - 0xf7e  :  120 - 0x78
    "00000000", -- 3967 - 0xf7f  :    0 - 0x0
    "11100100", -- 3968 - 0xf80  :  228 - 0xe4 -- Background 0xf8
    "11100100", -- 3969 - 0xf81  :  228 - 0xe4
    "11101111", -- 3970 - 0xf82  :  239 - 0xef
    "11101111", -- 3971 - 0xf83  :  239 - 0xef
    "11111111", -- 3972 - 0xf84  :  255 - 0xff
    "11111111", -- 3973 - 0xf85  :  255 - 0xff
    "01111111", -- 3974 - 0xf86  :  127 - 0x7f
    "01111111", -- 3975 - 0xf87  :  127 - 0x7f
    "00000011", -- 3976 - 0xf88  :    3 - 0x3 -- plane 1
    "00000011", -- 3977 - 0xf89  :    3 - 0x3
    "00000000", -- 3978 - 0xf8a  :    0 - 0x0
    "00000011", -- 3979 - 0xf8b  :    3 - 0x3
    "00000111", -- 3980 - 0xf8c  :    7 - 0x7
    "00000110", -- 3981 - 0xf8d  :    6 - 0x6
    "00000111", -- 3982 - 0xf8e  :    7 - 0x7
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "00111111", -- 3984 - 0xf90  :   63 - 0x3f -- Background 0xf9
    "01111111", -- 3985 - 0xf91  :  127 - 0x7f
    "01111111", -- 3986 - 0xf92  :  127 - 0x7f
    "11111111", -- 3987 - 0xf93  :  255 - 0xff
    "11111111", -- 3988 - 0xf94  :  255 - 0xff
    "11111111", -- 3989 - 0xf95  :  255 - 0xff
    "11111111", -- 3990 - 0xf96  :  255 - 0xff
    "11111111", -- 3991 - 0xf97  :  255 - 0xff
    "00000000", -- 3992 - 0xf98  :    0 - 0x0 -- plane 1
    "00011111", -- 3993 - 0xf99  :   31 - 0x1f
    "00011111", -- 3994 - 0xf9a  :   31 - 0x1f
    "00001111", -- 3995 - 0xf9b  :   15 - 0xf
    "00000011", -- 3996 - 0xf9c  :    3 - 0x3
    "00000000", -- 3997 - 0xf9d  :    0 - 0x0
    "00000000", -- 3998 - 0xf9e  :    0 - 0x0
    "00000000", -- 3999 - 0xf9f  :    0 - 0x0
    "00010011", -- 4000 - 0xfa0  :   19 - 0x13 -- Background 0xfa
    "00010011", -- 4001 - 0xfa1  :   19 - 0x13
    "11111011", -- 4002 - 0xfa2  :  251 - 0xfb
    "11111011", -- 4003 - 0xfa3  :  251 - 0xfb
    "11111111", -- 4004 - 0xfa4  :  255 - 0xff
    "11111111", -- 4005 - 0xfa5  :  255 - 0xff
    "11111110", -- 4006 - 0xfa6  :  254 - 0xfe
    "11111110", -- 4007 - 0xfa7  :  254 - 0xfe
    "11100000", -- 4008 - 0xfa8  :  224 - 0xe0 -- plane 1
    "11100000", -- 4009 - 0xfa9  :  224 - 0xe0
    "00000000", -- 4010 - 0xfaa  :    0 - 0x0
    "00110000", -- 4011 - 0xfab  :   48 - 0x30
    "01110000", -- 4012 - 0xfac  :  112 - 0x70
    "01100000", -- 4013 - 0xfad  :   96 - 0x60
    "01110000", -- 4014 - 0xfae  :  112 - 0x70
    "00000000", -- 4015 - 0xfaf  :    0 - 0x0
    "11111110", -- 4016 - 0xfb0  :  254 - 0xfe -- Background 0xfb
    "11111111", -- 4017 - 0xfb1  :  255 - 0xff
    "11111111", -- 4018 - 0xfb2  :  255 - 0xff
    "11111111", -- 4019 - 0xfb3  :  255 - 0xff
    "11111111", -- 4020 - 0xfb4  :  255 - 0xff
    "11111111", -- 4021 - 0xfb5  :  255 - 0xff
    "11111111", -- 4022 - 0xfb6  :  255 - 0xff
    "11111111", -- 4023 - 0xfb7  :  255 - 0xff
    "00000000", -- 4024 - 0xfb8  :    0 - 0x0 -- plane 1
    "11111000", -- 4025 - 0xfb9  :  248 - 0xf8
    "11111000", -- 4026 - 0xfba  :  248 - 0xf8
    "11110000", -- 4027 - 0xfbb  :  240 - 0xf0
    "11000000", -- 4028 - 0xfbc  :  192 - 0xc0
    "00000000", -- 4029 - 0xfbd  :    0 - 0x0
    "00000000", -- 4030 - 0xfbe  :    0 - 0x0
    "00000000", -- 4031 - 0xfbf  :    0 - 0x0
    "00000000", -- 4032 - 0xfc0  :    0 - 0x0 -- Background 0xfc
    "00000000", -- 4033 - 0xfc1  :    0 - 0x0
    "01111100", -- 4034 - 0xfc2  :  124 - 0x7c
    "11111110", -- 4035 - 0xfc3  :  254 - 0xfe
    "11111110", -- 4036 - 0xfc4  :  254 - 0xfe
    "01111100", -- 4037 - 0xfc5  :  124 - 0x7c
    "01000100", -- 4038 - 0xfc6  :   68 - 0x44
    "10000010", -- 4039 - 0xfc7  :  130 - 0x82
    "00111000", -- 4040 - 0xfc8  :   56 - 0x38 -- plane 1
    "00111000", -- 4041 - 0xfc9  :   56 - 0x38
    "00000000", -- 4042 - 0xfca  :    0 - 0x0
    "01111100", -- 4043 - 0xfcb  :  124 - 0x7c
    "00000000", -- 4044 - 0xfcc  :    0 - 0x0
    "00111000", -- 4045 - 0xfcd  :   56 - 0x38
    "00111000", -- 4046 - 0xfce  :   56 - 0x38
    "01111100", -- 4047 - 0xfcf  :  124 - 0x7c
    "10000010", -- 4048 - 0xfd0  :  130 - 0x82 -- Background 0xfd
    "10000010", -- 4049 - 0xfd1  :  130 - 0x82
    "10000010", -- 4050 - 0xfd2  :  130 - 0x82
    "11000110", -- 4051 - 0xfd3  :  198 - 0xc6
    "11111110", -- 4052 - 0xfd4  :  254 - 0xfe
    "11111110", -- 4053 - 0xfd5  :  254 - 0xfe
    "10111010", -- 4054 - 0xfd6  :  186 - 0xba
    "01111100", -- 4055 - 0xfd7  :  124 - 0x7c
    "01111100", -- 4056 - 0xfd8  :  124 - 0x7c -- plane 1
    "01111100", -- 4057 - 0xfd9  :  124 - 0x7c
    "01111100", -- 4058 - 0xfda  :  124 - 0x7c
    "00111000", -- 4059 - 0xfdb  :   56 - 0x38
    "00000000", -- 4060 - 0xfdc  :    0 - 0x0
    "01111100", -- 4061 - 0xfdd  :  124 - 0x7c
    "01111100", -- 4062 - 0xfde  :  124 - 0x7c
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00000000", -- 4064 - 0xfe0  :    0 - 0x0 -- Background 0xfe
    "00011001", -- 4065 - 0xfe1  :   25 - 0x19
    "00111110", -- 4066 - 0xfe2  :   62 - 0x3e
    "00111100", -- 4067 - 0xfe3  :   60 - 0x3c
    "00111100", -- 4068 - 0xfe4  :   60 - 0x3c
    "00111100", -- 4069 - 0xfe5  :   60 - 0x3c
    "00111110", -- 4070 - 0xfe6  :   62 - 0x3e
    "00011001", -- 4071 - 0xfe7  :   25 - 0x19
    "00000000", -- 4072 - 0xfe8  :    0 - 0x0 -- plane 1
    "00000000", -- 4073 - 0xfe9  :    0 - 0x0
    "00010001", -- 4074 - 0xfea  :   17 - 0x11
    "11010111", -- 4075 - 0xfeb  :  215 - 0xd7
    "11010111", -- 4076 - 0xfec  :  215 - 0xd7
    "11010111", -- 4077 - 0xfed  :  215 - 0xd7
    "00010001", -- 4078 - 0xfee  :   17 - 0x11
    "00000000", -- 4079 - 0xfef  :    0 - 0x0
    "00000000", -- 4080 - 0xff0  :    0 - 0x0 -- Background 0xff
    "11111110", -- 4081 - 0xff1  :  254 - 0xfe
    "00011101", -- 4082 - 0xff2  :   29 - 0x1d
    "00001111", -- 4083 - 0xff3  :   15 - 0xf
    "00001111", -- 4084 - 0xff4  :   15 - 0xf
    "00001111", -- 4085 - 0xff5  :   15 - 0xf
    "00011101", -- 4086 - 0xff6  :   29 - 0x1d
    "11111110", -- 4087 - 0xff7  :  254 - 0xfe
    "00000000", -- 4088 - 0xff8  :    0 - 0x0 -- plane 1
    "00000000", -- 4089 - 0xff9  :    0 - 0x0
    "11100110", -- 4090 - 0xffa  :  230 - 0xe6
    "11110110", -- 4091 - 0xffb  :  246 - 0xf6
    "11110110", -- 4092 - 0xffc  :  246 - 0xf6
    "11110110", -- 4093 - 0xffd  :  246 - 0xf6
    "11100110", -- 4094 - 0xffe  :  230 - 0xe6
    "00000000"  -- 4095 - 0xfff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
