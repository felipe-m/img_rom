//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: lawnmower_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_LAWN_color0
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout <= 8'b11111111; //    0 : 255 - 0xff -- Sprite 0x0
      12'h1: dout <= 8'b11111111; //    1 : 255 - 0xff
      12'h2: dout <= 8'b11111111; //    2 : 255 - 0xff
      12'h3: dout <= 8'b11111111; //    3 : 255 - 0xff
      12'h4: dout <= 8'b11111111; //    4 : 255 - 0xff
      12'h5: dout <= 8'b11111111; //    5 : 255 - 0xff
      12'h6: dout <= 8'b11111111; //    6 : 255 - 0xff
      12'h7: dout <= 8'b11111111; //    7 : 255 - 0xff
      12'h8: dout <= 8'b11111111; //    8 : 255 - 0xff -- Sprite 0x1
      12'h9: dout <= 8'b11111111; //    9 : 255 - 0xff
      12'hA: dout <= 8'b11111111; //   10 : 255 - 0xff
      12'hB: dout <= 8'b11111111; //   11 : 255 - 0xff
      12'hC: dout <= 8'b11111111; //   12 : 255 - 0xff
      12'hD: dout <= 8'b11111111; //   13 : 255 - 0xff
      12'hE: dout <= 8'b11111100; //   14 : 252 - 0xfc
      12'hF: dout <= 8'b11111100; //   15 : 252 - 0xfc
      12'h10: dout <= 8'b11111111; //   16 : 255 - 0xff -- Sprite 0x2
      12'h11: dout <= 8'b11111111; //   17 : 255 - 0xff
      12'h12: dout <= 8'b11111111; //   18 : 255 - 0xff
      12'h13: dout <= 8'b11111111; //   19 : 255 - 0xff
      12'h14: dout <= 8'b11111111; //   20 : 255 - 0xff
      12'h15: dout <= 8'b11111111; //   21 : 255 - 0xff
      12'h16: dout <= 8'b00000000; //   22 :   0 - 0x0
      12'h17: dout <= 8'b00000000; //   23 :   0 - 0x0
      12'h18: dout <= 8'b11111111; //   24 : 255 - 0xff -- Sprite 0x3
      12'h19: dout <= 8'b11111111; //   25 : 255 - 0xff
      12'h1A: dout <= 8'b11111111; //   26 : 255 - 0xff
      12'h1B: dout <= 8'b11111111; //   27 : 255 - 0xff
      12'h1C: dout <= 8'b11111111; //   28 : 255 - 0xff
      12'h1D: dout <= 8'b11111111; //   29 : 255 - 0xff
      12'h1E: dout <= 8'b00011111; //   30 :  31 - 0x1f
      12'h1F: dout <= 8'b01000111; //   31 :  71 - 0x47
      12'h20: dout <= 8'b11111111; //   32 : 255 - 0xff -- Sprite 0x4
      12'h21: dout <= 8'b11111111; //   33 : 255 - 0xff
      12'h22: dout <= 8'b11111111; //   34 : 255 - 0xff
      12'h23: dout <= 8'b11111111; //   35 : 255 - 0xff
      12'h24: dout <= 8'b11111111; //   36 : 255 - 0xff
      12'h25: dout <= 8'b11111111; //   37 : 255 - 0xff
      12'h26: dout <= 8'b11100000; //   38 : 224 - 0xe0
      12'h27: dout <= 8'b10000000; //   39 : 128 - 0x80
      12'h28: dout <= 8'b11111111; //   40 : 255 - 0xff -- Sprite 0x5
      12'h29: dout <= 8'b11111111; //   41 : 255 - 0xff
      12'h2A: dout <= 8'b11111111; //   42 : 255 - 0xff
      12'h2B: dout <= 8'b11111111; //   43 : 255 - 0xff
      12'h2C: dout <= 8'b11111111; //   44 : 255 - 0xff
      12'h2D: dout <= 8'b11110111; //   45 : 247 - 0xf7
      12'h2E: dout <= 8'b00000001; //   46 :   1 - 0x1
      12'h2F: dout <= 8'b00000100; //   47 :   4 - 0x4
      12'h30: dout <= 8'b11111111; //   48 : 255 - 0xff -- Sprite 0x6
      12'h31: dout <= 8'b11111111; //   49 : 255 - 0xff
      12'h32: dout <= 8'b11111111; //   50 : 255 - 0xff
      12'h33: dout <= 8'b11111111; //   51 : 255 - 0xff
      12'h34: dout <= 8'b11111111; //   52 : 255 - 0xff
      12'h35: dout <= 8'b11011111; //   53 : 223 - 0xdf
      12'h36: dout <= 8'b00011100; //   54 :  28 - 0x1c
      12'h37: dout <= 8'b01000100; //   55 :  68 - 0x44
      12'h38: dout <= 8'b11111111; //   56 : 255 - 0xff -- Sprite 0x7
      12'h39: dout <= 8'b11111111; //   57 : 255 - 0xff
      12'h3A: dout <= 8'b11111111; //   58 : 255 - 0xff
      12'h3B: dout <= 8'b11111111; //   59 : 255 - 0xff
      12'h3C: dout <= 8'b11111111; //   60 : 255 - 0xff
      12'h3D: dout <= 8'b10111111; //   61 : 191 - 0xbf
      12'h3E: dout <= 8'b00111100; //   62 :  60 - 0x3c
      12'h3F: dout <= 8'b01001100; //   63 :  76 - 0x4c
      12'h40: dout <= 8'b11111100; //   64 : 252 - 0xfc -- Sprite 0x8
      12'h41: dout <= 8'b11111100; //   65 : 252 - 0xfc
      12'h42: dout <= 8'b11111100; //   66 : 252 - 0xfc
      12'h43: dout <= 8'b11111100; //   67 : 252 - 0xfc
      12'h44: dout <= 8'b11111100; //   68 : 252 - 0xfc
      12'h45: dout <= 8'b11111100; //   69 : 252 - 0xfc
      12'h46: dout <= 8'b11111100; //   70 : 252 - 0xfc
      12'h47: dout <= 8'b11111100; //   71 : 252 - 0xfc
      12'h48: dout <= 8'b00010000; //   72 :  16 - 0x10 -- Sprite 0x9
      12'h49: dout <= 8'b00111000; //   73 :  56 - 0x38
      12'h4A: dout <= 8'b01111100; //   74 : 124 - 0x7c
      12'h4B: dout <= 8'b11111000; //   75 : 248 - 0xf8
      12'h4C: dout <= 8'b01110000; //   76 : 112 - 0x70
      12'h4D: dout <= 8'b00100010; //   77 :  34 - 0x22
      12'h4E: dout <= 8'b00000101; //   78 :   5 - 0x5
      12'h4F: dout <= 8'b00000010; //   79 :   2 - 0x2
      12'h50: dout <= 8'b01000111; //   80 :  71 - 0x47 -- Sprite 0xa
      12'h51: dout <= 8'b01000111; //   81 :  71 - 0x47
      12'h52: dout <= 8'b01000111; //   82 :  71 - 0x47
      12'h53: dout <= 8'b01000111; //   83 :  71 - 0x47
      12'h54: dout <= 8'b01000111; //   84 :  71 - 0x47
      12'h55: dout <= 8'b01000111; //   85 :  71 - 0x47
      12'h56: dout <= 8'b01000111; //   86 :  71 - 0x47
      12'h57: dout <= 8'b01000111; //   87 :  71 - 0x47
      12'h58: dout <= 8'b11111111; //   88 : 255 - 0xff -- Sprite 0xb
      12'h59: dout <= 8'b11111110; //   89 : 254 - 0xfe
      12'h5A: dout <= 8'b11111110; //   90 : 254 - 0xfe
      12'h5B: dout <= 8'b11111100; //   91 : 252 - 0xfc
      12'h5C: dout <= 8'b11111100; //   92 : 252 - 0xfc
      12'h5D: dout <= 8'b11111100; //   93 : 252 - 0xfc
      12'h5E: dout <= 8'b11111100; //   94 : 252 - 0xfc
      12'h5F: dout <= 8'b11111100; //   95 : 252 - 0xfc
      12'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0xc
      12'h61: dout <= 8'b00001000; //   97 :   8 - 0x8
      12'h62: dout <= 8'b00011100; //   98 :  28 - 0x1c
      12'h63: dout <= 8'b00111000; //   99 :  56 - 0x38
      12'h64: dout <= 8'b01110000; //  100 : 112 - 0x70
      12'h65: dout <= 8'b00100010; //  101 :  34 - 0x22
      12'h66: dout <= 8'b00000101; //  102 :   5 - 0x5
      12'h67: dout <= 8'b00000010; //  103 :   2 - 0x2
      12'h68: dout <= 8'b00000010; //  104 :   2 - 0x2 -- Sprite 0xd
      12'h69: dout <= 8'b00110001; //  105 :  49 - 0x31
      12'h6A: dout <= 8'b01111000; //  106 : 120 - 0x78
      12'h6B: dout <= 8'b11111000; //  107 : 248 - 0xf8
      12'h6C: dout <= 8'b01110000; //  108 : 112 - 0x70
      12'h6D: dout <= 8'b00100010; //  109 :  34 - 0x22
      12'h6E: dout <= 8'b00000101; //  110 :   5 - 0x5
      12'h6F: dout <= 8'b00000010; //  111 :   2 - 0x2
      12'h70: dout <= 8'b01111100; //  112 : 124 - 0x7c -- Sprite 0xe
      12'h71: dout <= 8'b00111100; //  113 :  60 - 0x3c
      12'h72: dout <= 8'b10011100; //  114 : 156 - 0x9c
      12'h73: dout <= 8'b10001100; //  115 : 140 - 0x8c
      12'h74: dout <= 8'b01001100; //  116 :  76 - 0x4c
      12'h75: dout <= 8'b01000100; //  117 :  68 - 0x44
      12'h76: dout <= 8'b01000100; //  118 :  68 - 0x44
      12'h77: dout <= 8'b01000100; //  119 :  68 - 0x44
      12'h78: dout <= 8'b01000100; //  120 :  68 - 0x44 -- Sprite 0xf
      12'h79: dout <= 8'b01000100; //  121 :  68 - 0x44
      12'h7A: dout <= 8'b01000100; //  122 :  68 - 0x44
      12'h7B: dout <= 8'b01000100; //  123 :  68 - 0x44
      12'h7C: dout <= 8'b01000100; //  124 :  68 - 0x44
      12'h7D: dout <= 8'b01000100; //  125 :  68 - 0x44
      12'h7E: dout <= 8'b01000100; //  126 :  68 - 0x44
      12'h7F: dout <= 8'b01000100; //  127 :  68 - 0x44
      12'h80: dout <= 8'b01001100; //  128 :  76 - 0x4c -- Sprite 0x10
      12'h81: dout <= 8'b00100100; //  129 :  36 - 0x24
      12'h82: dout <= 8'b00100100; //  130 :  36 - 0x24
      12'h83: dout <= 8'b10010100; //  131 : 148 - 0x94
      12'h84: dout <= 8'b00010000; //  132 :  16 - 0x10
      12'h85: dout <= 8'b00001000; //  133 :   8 - 0x8
      12'h86: dout <= 8'b00001000; //  134 :   8 - 0x8
      12'h87: dout <= 8'b00000100; //  135 :   4 - 0x4
      12'h88: dout <= 8'b00000000; //  136 :   0 - 0x0 -- Sprite 0x11
      12'h89: dout <= 8'b00111100; //  137 :  60 - 0x3c
      12'h8A: dout <= 8'b01000000; //  138 :  64 - 0x40
      12'h8B: dout <= 8'b01000100; //  139 :  68 - 0x44
      12'h8C: dout <= 8'b01000100; //  140 :  68 - 0x44
      12'h8D: dout <= 8'b01000100; //  141 :  68 - 0x44
      12'h8E: dout <= 8'b01000100; //  142 :  68 - 0x44
      12'h8F: dout <= 8'b01000100; //  143 :  68 - 0x44
      12'h90: dout <= 8'b00000100; //  144 :   4 - 0x4 -- Sprite 0x12
      12'h91: dout <= 8'b00010010; //  145 :  18 - 0x12
      12'h92: dout <= 8'b00110010; //  146 :  50 - 0x32
      12'h93: dout <= 8'b01111000; //  147 : 120 - 0x78
      12'h94: dout <= 8'b11111000; //  148 : 248 - 0xf8
      12'h95: dout <= 8'b01110000; //  149 : 112 - 0x70
      12'h96: dout <= 8'b00100100; //  150 :  36 - 0x24
      12'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      12'h98: dout <= 8'b01000100; //  152 :  68 - 0x44 -- Sprite 0x13
      12'h99: dout <= 8'b01000100; //  153 :  68 - 0x44
      12'h9A: dout <= 8'b01000100; //  154 :  68 - 0x44
      12'h9B: dout <= 8'b01000100; //  155 :  68 - 0x44
      12'h9C: dout <= 8'b01000100; //  156 :  68 - 0x44
      12'h9D: dout <= 8'b01000100; //  157 :  68 - 0x44
      12'h9E: dout <= 8'b01000100; //  158 :  68 - 0x44
      12'h9F: dout <= 8'b01011100; //  159 :  92 - 0x5c
      12'hA0: dout <= 8'b00010000; //  160 :  16 - 0x10 -- Sprite 0x14
      12'hA1: dout <= 8'b00111000; //  161 :  56 - 0x38
      12'hA2: dout <= 8'b00111100; //  162 :  60 - 0x3c
      12'hA3: dout <= 8'b00111000; //  163 :  56 - 0x38
      12'hA4: dout <= 8'b00010000; //  164 :  16 - 0x10
      12'hA5: dout <= 8'b00000010; //  165 :   2 - 0x2
      12'hA6: dout <= 8'b01000101; //  166 :  69 - 0x45
      12'hA7: dout <= 8'b01000010; //  167 :  66 - 0x42
      12'hA8: dout <= 8'b01000100; //  168 :  68 - 0x44 -- Sprite 0x15
      12'hA9: dout <= 8'b01000100; //  169 :  68 - 0x44
      12'hAA: dout <= 8'b01000100; //  170 :  68 - 0x44
      12'hAB: dout <= 8'b01000100; //  171 :  68 - 0x44
      12'hAC: dout <= 8'b01000100; //  172 :  68 - 0x44
      12'hAD: dout <= 8'b01011100; //  173 :  92 - 0x5c
      12'hAE: dout <= 8'b01000000; //  174 :  64 - 0x40
      12'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      12'hB0: dout <= 8'b01000000; //  176 :  64 - 0x40 -- Sprite 0x16
      12'hB1: dout <= 8'b01000000; //  177 :  64 - 0x40
      12'hB2: dout <= 8'b00000000; //  178 :   0 - 0x0
      12'hB3: dout <= 8'b00000000; //  179 :   0 - 0x0
      12'hB4: dout <= 8'b00011000; //  180 :  24 - 0x18
      12'hB5: dout <= 8'b00111000; //  181 :  56 - 0x38
      12'hB6: dout <= 8'b00010000; //  182 :  16 - 0x10
      12'hB7: dout <= 8'b00000000; //  183 :   0 - 0x0
      12'hB8: dout <= 8'b01000000; //  184 :  64 - 0x40 -- Sprite 0x17
      12'hB9: dout <= 8'b01000000; //  185 :  64 - 0x40
      12'hBA: dout <= 8'b01000000; //  186 :  64 - 0x40
      12'hBB: dout <= 8'b01000000; //  187 :  64 - 0x40
      12'hBC: dout <= 8'b01010000; //  188 :  80 - 0x50
      12'hBD: dout <= 8'b01010000; //  189 :  80 - 0x50
      12'hBE: dout <= 8'b01001000; //  190 :  72 - 0x48
      12'hBF: dout <= 8'b01001000; //  191 :  72 - 0x48
      12'hC0: dout <= 8'b01000111; //  192 :  71 - 0x47 -- Sprite 0x18
      12'hC1: dout <= 8'b01000111; //  193 :  71 - 0x47
      12'hC2: dout <= 8'b01000111; //  194 :  71 - 0x47
      12'hC3: dout <= 8'b01000111; //  195 :  71 - 0x47
      12'hC4: dout <= 8'b01000111; //  196 :  71 - 0x47
      12'hC5: dout <= 8'b01011111; //  197 :  95 - 0x5f
      12'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      12'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      12'hC8: dout <= 8'b11111100; //  200 : 252 - 0xfc -- Sprite 0x19
      12'hC9: dout <= 8'b11111100; //  201 : 252 - 0xfc
      12'hCA: dout <= 8'b11111100; //  202 : 252 - 0xfc
      12'hCB: dout <= 8'b11111100; //  203 : 252 - 0xfc
      12'hCC: dout <= 8'b11111100; //  204 : 252 - 0xfc
      12'hCD: dout <= 8'b11011100; //  205 : 220 - 0xdc
      12'hCE: dout <= 8'b00011100; //  206 :  28 - 0x1c
      12'hCF: dout <= 8'b01000100; //  207 :  68 - 0x44
      12'hD0: dout <= 8'b00010000; //  208 :  16 - 0x10 -- Sprite 0x1a
      12'hD1: dout <= 8'b00111000; //  209 :  56 - 0x38
      12'hD2: dout <= 8'b01111100; //  210 : 124 - 0x7c
      12'hD3: dout <= 8'b11100000; //  211 : 224 - 0xe0
      12'hD4: dout <= 8'b01000000; //  212 :  64 - 0x40
      12'hD5: dout <= 8'b00000000; //  213 :   0 - 0x0
      12'hD6: dout <= 8'b00010000; //  214 :  16 - 0x10
      12'hD7: dout <= 8'b00100000; //  215 :  32 - 0x20
      12'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x1b
      12'hD9: dout <= 8'b01111100; //  217 : 124 - 0x7c
      12'hDA: dout <= 8'b01000000; //  218 :  64 - 0x40
      12'hDB: dout <= 8'b01000100; //  219 :  68 - 0x44
      12'hDC: dout <= 8'b01000100; //  220 :  68 - 0x44
      12'hDD: dout <= 8'b01000100; //  221 :  68 - 0x44
      12'hDE: dout <= 8'b01000100; //  222 :  68 - 0x44
      12'hDF: dout <= 8'b01000100; //  223 :  68 - 0x44
      12'hE0: dout <= 8'b00010000; //  224 :  16 - 0x10 -- Sprite 0x1c
      12'hE1: dout <= 8'b00111000; //  225 :  56 - 0x38
      12'hE2: dout <= 8'b01110001; //  226 : 113 - 0x71
      12'hE3: dout <= 8'b11100010; //  227 : 226 - 0xe2
      12'hE4: dout <= 8'b01000100; //  228 :  68 - 0x44
      12'hE5: dout <= 8'b00001000; //  229 :   8 - 0x8
      12'hE6: dout <= 8'b00010000; //  230 :  16 - 0x10
      12'hE7: dout <= 8'b00100000; //  231 :  32 - 0x20
      12'hE8: dout <= 8'b01000000; //  232 :  64 - 0x40 -- Sprite 0x1d
      12'hE9: dout <= 8'b10000100; //  233 : 132 - 0x84
      12'hEA: dout <= 8'b00000010; //  234 :   2 - 0x2
      12'hEB: dout <= 8'b00000111; //  235 :   7 - 0x7
      12'hEC: dout <= 8'b00001111; //  236 :  15 - 0xf
      12'hED: dout <= 8'b00011111; //  237 :  31 - 0x1f
      12'hEE: dout <= 8'b00111111; //  238 :  63 - 0x3f
      12'hEF: dout <= 8'b01111111; //  239 : 127 - 0x7f
      12'hF0: dout <= 8'b00010000; //  240 :  16 - 0x10 -- Sprite 0x1e
      12'hF1: dout <= 8'b00011000; //  241 :  24 - 0x18
      12'hF2: dout <= 8'b00001100; //  242 :  12 - 0xc
      12'hF3: dout <= 8'b00000110; //  243 :   6 - 0x6
      12'hF4: dout <= 8'b10000000; //  244 : 128 - 0x80
      12'hF5: dout <= 8'b11000000; //  245 : 192 - 0xc0
      12'hF6: dout <= 8'b11100000; //  246 : 224 - 0xe0
      12'hF7: dout <= 8'b11110000; //  247 : 240 - 0xf0
      12'hF8: dout <= 8'b11111100; //  248 : 252 - 0xfc -- Sprite 0x1f
      12'hF9: dout <= 8'b11111101; //  249 : 253 - 0xfd
      12'hFA: dout <= 8'b11111100; //  250 : 252 - 0xfc
      12'hFB: dout <= 8'b11111110; //  251 : 254 - 0xfe
      12'hFC: dout <= 8'b11111110; //  252 : 254 - 0xfe
      12'hFD: dout <= 8'b11111111; //  253 : 255 - 0xff
      12'hFE: dout <= 8'b11111111; //  254 : 255 - 0xff
      12'hFF: dout <= 8'b11111111; //  255 : 255 - 0xff
      12'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      12'h101: dout <= 8'b11111111; //  257 : 255 - 0xff
      12'h102: dout <= 8'b00000000; //  258 :   0 - 0x0
      12'h103: dout <= 8'b00000000; //  259 :   0 - 0x0
      12'h104: dout <= 8'b00000000; //  260 :   0 - 0x0
      12'h105: dout <= 8'b11111111; //  261 : 255 - 0xff
      12'h106: dout <= 8'b11111111; //  262 : 255 - 0xff
      12'h107: dout <= 8'b11111111; //  263 : 255 - 0xff
      12'h108: dout <= 8'b01000100; //  264 :  68 - 0x44 -- Sprite 0x21
      12'h109: dout <= 8'b11000101; //  265 : 197 - 0xc5
      12'h10A: dout <= 8'b00000000; //  266 :   0 - 0x0
      12'h10B: dout <= 8'b00000110; //  267 :   6 - 0x6
      12'h10C: dout <= 8'b00000110; //  268 :   6 - 0x6
      12'h10D: dout <= 8'b11111111; //  269 : 255 - 0xff
      12'h10E: dout <= 8'b11111111; //  270 : 255 - 0xff
      12'h10F: dout <= 8'b11111111; //  271 : 255 - 0xff
      12'h110: dout <= 8'b01000000; //  272 :  64 - 0x40 -- Sprite 0x22
      12'h111: dout <= 8'b10000001; //  273 : 129 - 0x81
      12'h112: dout <= 8'b00000011; //  274 :   3 - 0x3
      12'h113: dout <= 8'b00000111; //  275 :   7 - 0x7
      12'h114: dout <= 8'b00001111; //  276 :  15 - 0xf
      12'h115: dout <= 8'b11111111; //  277 : 255 - 0xff
      12'h116: dout <= 8'b11111111; //  278 : 255 - 0xff
      12'h117: dout <= 8'b11111111; //  279 : 255 - 0xff
      12'h118: dout <= 8'b11111000; //  280 : 248 - 0xf8 -- Sprite 0x23
      12'h119: dout <= 8'b11111100; //  281 : 252 - 0xfc
      12'h11A: dout <= 8'b11111110; //  282 : 254 - 0xfe
      12'h11B: dout <= 8'b11111110; //  283 : 254 - 0xfe
      12'h11C: dout <= 8'b11111111; //  284 : 255 - 0xff
      12'h11D: dout <= 8'b11111111; //  285 : 255 - 0xff
      12'h11E: dout <= 8'b11111111; //  286 : 255 - 0xff
      12'h11F: dout <= 8'b11111111; //  287 : 255 - 0xff
      12'h120: dout <= 8'b01000111; //  288 :  71 - 0x47 -- Sprite 0x24
      12'h121: dout <= 8'b11000111; //  289 : 199 - 0xc7
      12'h122: dout <= 8'b00000111; //  290 :   7 - 0x7
      12'h123: dout <= 8'b00000111; //  291 :   7 - 0x7
      12'h124: dout <= 8'b00000111; //  292 :   7 - 0x7
      12'h125: dout <= 8'b11111111; //  293 : 255 - 0xff
      12'h126: dout <= 8'b11111111; //  294 : 255 - 0xff
      12'h127: dout <= 8'b11111111; //  295 : 255 - 0xff
      12'h128: dout <= 8'b11111111; //  296 : 255 - 0xff -- Sprite 0x25
      12'h129: dout <= 8'b11111111; //  297 : 255 - 0xff
      12'h12A: dout <= 8'b11111111; //  298 : 255 - 0xff
      12'h12B: dout <= 8'b11111111; //  299 : 255 - 0xff
      12'h12C: dout <= 8'b11111111; //  300 : 255 - 0xff
      12'h12D: dout <= 8'b11111111; //  301 : 255 - 0xff
      12'h12E: dout <= 8'b00011111; //  302 :  31 - 0x1f
      12'h12F: dout <= 8'b00001111; //  303 :  15 - 0xf
      12'h130: dout <= 8'b11111111; //  304 : 255 - 0xff -- Sprite 0x26
      12'h131: dout <= 8'b11111111; //  305 : 255 - 0xff
      12'h132: dout <= 8'b11111111; //  306 : 255 - 0xff
      12'h133: dout <= 8'b11111111; //  307 : 255 - 0xff
      12'h134: dout <= 8'b11111111; //  308 : 255 - 0xff
      12'h135: dout <= 8'b11111111; //  309 : 255 - 0xff
      12'h136: dout <= 8'b11111100; //  310 : 252 - 0xfc
      12'h137: dout <= 8'b11111000; //  311 : 248 - 0xf8
      12'h138: dout <= 8'b00100111; //  312 :  39 - 0x27 -- Sprite 0x27
      12'h139: dout <= 8'b00010011; //  313 :  19 - 0x13
      12'h13A: dout <= 8'b00001001; //  314 :   9 - 0x9
      12'h13B: dout <= 8'b11000100; //  315 : 196 - 0xc4
      12'h13C: dout <= 8'b01100010; //  316 :  98 - 0x62
      12'h13D: dout <= 8'b00100001; //  317 :  33 - 0x21
      12'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout <= 8'b11111111; //  320 : 255 - 0xff -- Sprite 0x28
      12'h141: dout <= 8'b11111111; //  321 : 255 - 0xff
      12'h142: dout <= 8'b11111111; //  322 : 255 - 0xff
      12'h143: dout <= 8'b11111111; //  323 : 255 - 0xff
      12'h144: dout <= 8'b01111111; //  324 : 127 - 0x7f
      12'h145: dout <= 8'b00111110; //  325 :  62 - 0x3e
      12'h146: dout <= 8'b10011100; //  326 : 156 - 0x9c
      12'h147: dout <= 8'b01001000; //  327 :  72 - 0x48
      12'h148: dout <= 8'b11110000; //  328 : 240 - 0xf0 -- Sprite 0x29
      12'h149: dout <= 8'b11100000; //  329 : 224 - 0xe0
      12'h14A: dout <= 8'b11000000; //  330 : 192 - 0xc0
      12'h14B: dout <= 8'b10000000; //  331 : 128 - 0x80
      12'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      12'h14D: dout <= 8'b00000010; //  333 :   2 - 0x2
      12'h14E: dout <= 8'b00000101; //  334 :   5 - 0x5
      12'h14F: dout <= 8'b00000010; //  335 :   2 - 0x2
      12'h150: dout <= 8'b01000111; //  336 :  71 - 0x47 -- Sprite 0x2a
      12'h151: dout <= 8'b01000110; //  337 :  70 - 0x46
      12'h152: dout <= 8'b01000110; //  338 :  70 - 0x46
      12'h153: dout <= 8'b01000100; //  339 :  68 - 0x44
      12'h154: dout <= 8'b01000100; //  340 :  68 - 0x44
      12'h155: dout <= 8'b01000100; //  341 :  68 - 0x44
      12'h156: dout <= 8'b01000100; //  342 :  68 - 0x44
      12'h157: dout <= 8'b01000100; //  343 :  68 - 0x44
      12'h158: dout <= 8'b01111111; //  344 : 127 - 0x7f -- Sprite 0x2b
      12'h159: dout <= 8'b00111111; //  345 :  63 - 0x3f
      12'h15A: dout <= 8'b10011111; //  346 : 159 - 0x9f
      12'h15B: dout <= 8'b10001111; //  347 : 143 - 0x8f
      12'h15C: dout <= 8'b01001111; //  348 :  79 - 0x4f
      12'h15D: dout <= 8'b01000111; //  349 :  71 - 0x47
      12'h15E: dout <= 8'b01000111; //  350 :  71 - 0x47
      12'h15F: dout <= 8'b01000111; //  351 :  71 - 0x47
      12'h160: dout <= 8'b00100000; //  352 :  32 - 0x20 -- Sprite 0x2c
      12'h161: dout <= 8'b00010000; //  353 :  16 - 0x10
      12'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      12'h163: dout <= 8'b11000000; //  355 : 192 - 0xc0
      12'h164: dout <= 8'b01100000; //  356 :  96 - 0x60
      12'h165: dout <= 8'b00100010; //  357 :  34 - 0x22
      12'h166: dout <= 8'b00000101; //  358 :   5 - 0x5
      12'h167: dout <= 8'b00000010; //  359 :   2 - 0x2
      12'h168: dout <= 8'b00000000; //  360 :   0 - 0x0 -- Sprite 0x2d
      12'h169: dout <= 8'b01111111; //  361 : 127 - 0x7f
      12'h16A: dout <= 8'b01000000; //  362 :  64 - 0x40
      12'h16B: dout <= 8'b01000000; //  363 :  64 - 0x40
      12'h16C: dout <= 8'b01000000; //  364 :  64 - 0x40
      12'h16D: dout <= 8'b01000111; //  365 :  71 - 0x47
      12'h16E: dout <= 8'b01000111; //  366 :  71 - 0x47
      12'h16F: dout <= 8'b01000111; //  367 :  71 - 0x47
      12'h170: dout <= 8'b01000100; //  368 :  68 - 0x44 -- Sprite 0x2e
      12'h171: dout <= 8'b11000100; //  369 : 196 - 0xc4
      12'h172: dout <= 8'b00000100; //  370 :   4 - 0x4
      12'h173: dout <= 8'b00000100; //  371 :   4 - 0x4
      12'h174: dout <= 8'b00000100; //  372 :   4 - 0x4
      12'h175: dout <= 8'b11111100; //  373 : 252 - 0xfc
      12'h176: dout <= 8'b11111100; //  374 : 252 - 0xfc
      12'h177: dout <= 8'b11111100; //  375 : 252 - 0xfc
      12'h178: dout <= 8'b00000001; //  376 :   1 - 0x1 -- Sprite 0x2f
      12'h179: dout <= 8'b01111100; //  377 : 124 - 0x7c
      12'h17A: dout <= 8'b01000000; //  378 :  64 - 0x40
      12'h17B: dout <= 8'b01000100; //  379 :  68 - 0x44
      12'h17C: dout <= 8'b01000100; //  380 :  68 - 0x44
      12'h17D: dout <= 8'b01000100; //  381 :  68 - 0x44
      12'h17E: dout <= 8'b01000100; //  382 :  68 - 0x44
      12'h17F: dout <= 8'b01000100; //  383 :  68 - 0x44
      12'h180: dout <= 8'b00010000; //  384 :  16 - 0x10 -- Sprite 0x30
      12'h181: dout <= 8'b00111000; //  385 :  56 - 0x38
      12'h182: dout <= 8'b00111100; //  386 :  60 - 0x3c
      12'h183: dout <= 8'b00011000; //  387 :  24 - 0x18
      12'h184: dout <= 8'b00000000; //  388 :   0 - 0x0
      12'h185: dout <= 8'b01000010; //  389 :  66 - 0x42
      12'h186: dout <= 8'b01000100; //  390 :  68 - 0x44
      12'h187: dout <= 8'b01001000; //  391 :  72 - 0x48
      12'h188: dout <= 8'b01000111; //  392 :  71 - 0x47 -- Sprite 0x31
      12'h189: dout <= 8'b01011111; //  393 :  95 - 0x5f
      12'h18A: dout <= 8'b00000000; //  394 :   0 - 0x0
      12'h18B: dout <= 8'b00000000; //  395 :   0 - 0x0
      12'h18C: dout <= 8'b01110000; //  396 : 112 - 0x70
      12'h18D: dout <= 8'b00100010; //  397 :  34 - 0x22
      12'h18E: dout <= 8'b00000101; //  398 :   5 - 0x5
      12'h18F: dout <= 8'b00000010; //  399 :   2 - 0x2
      12'h190: dout <= 8'b11111111; //  400 : 255 - 0xff -- Sprite 0x32
      12'h191: dout <= 8'b11111111; //  401 : 255 - 0xff
      12'h192: dout <= 8'b00000000; //  402 :   0 - 0x0
      12'h193: dout <= 8'b00000000; //  403 :   0 - 0x0
      12'h194: dout <= 8'b01110000; //  404 : 112 - 0x70
      12'h195: dout <= 8'b00100010; //  405 :  34 - 0x22
      12'h196: dout <= 8'b00000101; //  406 :   5 - 0x5
      12'h197: dout <= 8'b00000010; //  407 :   2 - 0x2
      12'h198: dout <= 8'b11111111; //  408 : 255 - 0xff -- Sprite 0x33
      12'h199: dout <= 8'b11011111; //  409 : 223 - 0xdf
      12'h19A: dout <= 8'b00011111; //  410 :  31 - 0x1f
      12'h19B: dout <= 8'b01000111; //  411 :  71 - 0x47
      12'h19C: dout <= 8'b01000111; //  412 :  71 - 0x47
      12'h19D: dout <= 8'b01000111; //  413 :  71 - 0x47
      12'h19E: dout <= 8'b01000111; //  414 :  71 - 0x47
      12'h19F: dout <= 8'b01000111; //  415 :  71 - 0x47
      12'h1A0: dout <= 8'b01000100; //  416 :  68 - 0x44 -- Sprite 0x34
      12'h1A1: dout <= 8'b01000100; //  417 :  68 - 0x44
      12'h1A2: dout <= 8'b01000100; //  418 :  68 - 0x44
      12'h1A3: dout <= 8'b01000100; //  419 :  68 - 0x44
      12'h1A4: dout <= 8'b01000100; //  420 :  68 - 0x44
      12'h1A5: dout <= 8'b01000100; //  421 :  68 - 0x44
      12'h1A6: dout <= 8'b01000100; //  422 :  68 - 0x44
      12'h1A7: dout <= 8'b01000100; //  423 :  68 - 0x44
      12'h1A8: dout <= 8'b00010000; //  424 :  16 - 0x10 -- Sprite 0x35
      12'h1A9: dout <= 8'b00111000; //  425 :  56 - 0x38
      12'h1AA: dout <= 8'b01111100; //  426 : 124 - 0x7c
      12'h1AB: dout <= 8'b11111000; //  427 : 248 - 0xf8
      12'h1AC: dout <= 8'b00000000; //  428 :   0 - 0x0
      12'h1AD: dout <= 8'b01111111; //  429 : 127 - 0x7f
      12'h1AE: dout <= 8'b01000000; //  430 :  64 - 0x40
      12'h1AF: dout <= 8'b01000000; //  431 :  64 - 0x40
      12'h1B0: dout <= 8'b00010000; //  432 :  16 - 0x10 -- Sprite 0x36
      12'h1B1: dout <= 8'b00111000; //  433 :  56 - 0x38
      12'h1B2: dout <= 8'b01111100; //  434 : 124 - 0x7c
      12'h1B3: dout <= 8'b11111000; //  435 : 248 - 0xf8
      12'h1B4: dout <= 8'b00000000; //  436 :   0 - 0x0
      12'h1B5: dout <= 8'b11111111; //  437 : 255 - 0xff
      12'h1B6: dout <= 8'b00000000; //  438 :   0 - 0x0
      12'h1B7: dout <= 8'b00000000; //  439 :   0 - 0x0
      12'h1B8: dout <= 8'b01000111; //  440 :  71 - 0x47 -- Sprite 0x37
      12'h1B9: dout <= 8'b01000111; //  441 :  71 - 0x47
      12'h1BA: dout <= 8'b01000111; //  442 :  71 - 0x47
      12'h1BB: dout <= 8'b01000111; //  443 :  71 - 0x47
      12'h1BC: dout <= 8'b01000111; //  444 :  71 - 0x47
      12'h1BD: dout <= 8'b11000111; //  445 : 199 - 0xc7
      12'h1BE: dout <= 8'b00000111; //  446 :   7 - 0x7
      12'h1BF: dout <= 8'b00000111; //  447 :   7 - 0x7
      12'h1C0: dout <= 8'b01000100; //  448 :  68 - 0x44 -- Sprite 0x38
      12'h1C1: dout <= 8'b01000100; //  449 :  68 - 0x44
      12'h1C2: dout <= 8'b01000100; //  450 :  68 - 0x44
      12'h1C3: dout <= 8'b01000100; //  451 :  68 - 0x44
      12'h1C4: dout <= 8'b01000100; //  452 :  68 - 0x44
      12'h1C5: dout <= 8'b01011000; //  453 :  88 - 0x58
      12'h1C6: dout <= 8'b00000000; //  454 :   0 - 0x0
      12'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      12'h1C8: dout <= 8'b00010000; //  456 :  16 - 0x10 -- Sprite 0x39
      12'h1C9: dout <= 8'b00111000; //  457 :  56 - 0x38
      12'h1CA: dout <= 8'b01111100; //  458 : 124 - 0x7c
      12'h1CB: dout <= 8'b11111000; //  459 : 248 - 0xf8
      12'h1CC: dout <= 8'b01110000; //  460 : 112 - 0x70
      12'h1CD: dout <= 8'b00100010; //  461 :  34 - 0x22
      12'h1CE: dout <= 8'b00000100; //  462 :   4 - 0x4
      12'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout <= 8'b01000100; //  464 :  68 - 0x44 -- Sprite 0x3a
      12'h1D1: dout <= 8'b01000100; //  465 :  68 - 0x44
      12'h1D2: dout <= 8'b01000100; //  466 :  68 - 0x44
      12'h1D3: dout <= 8'b01000100; //  467 :  68 - 0x44
      12'h1D4: dout <= 8'b01000100; //  468 :  68 - 0x44
      12'h1D5: dout <= 8'b01011000; //  469 :  88 - 0x58
      12'h1D6: dout <= 8'b00000000; //  470 :   0 - 0x0
      12'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      12'h1D8: dout <= 8'b01000000; //  472 :  64 - 0x40 -- Sprite 0x3b
      12'h1D9: dout <= 8'b01000111; //  473 :  71 - 0x47
      12'h1DA: dout <= 8'b01000111; //  474 :  71 - 0x47
      12'h1DB: dout <= 8'b01000111; //  475 :  71 - 0x47
      12'h1DC: dout <= 8'b01000111; //  476 :  71 - 0x47
      12'h1DD: dout <= 8'b01011111; //  477 :  95 - 0x5f
      12'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      12'h1E1: dout <= 8'b11111111; //  481 : 255 - 0xff
      12'h1E2: dout <= 8'b11111111; //  482 : 255 - 0xff
      12'h1E3: dout <= 8'b11111111; //  483 : 255 - 0xff
      12'h1E4: dout <= 8'b11111111; //  484 : 255 - 0xff
      12'h1E5: dout <= 8'b11111111; //  485 : 255 - 0xff
      12'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      12'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout <= 8'b00000111; //  488 :   7 - 0x7 -- Sprite 0x3d
      12'h1E9: dout <= 8'b11111111; //  489 : 255 - 0xff
      12'h1EA: dout <= 8'b11111111; //  490 : 255 - 0xff
      12'h1EB: dout <= 8'b11111111; //  491 : 255 - 0xff
      12'h1EC: dout <= 8'b11111111; //  492 : 255 - 0xff
      12'h1ED: dout <= 8'b11111111; //  493 : 255 - 0xff
      12'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      12'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout <= 8'b00010000; //  496 :  16 - 0x10 -- Sprite 0x3e
      12'h1F1: dout <= 8'b00111000; //  497 :  56 - 0x38
      12'h1F2: dout <= 8'b01110001; //  498 : 113 - 0x71
      12'h1F3: dout <= 8'b11100010; //  499 : 226 - 0xe2
      12'h1F4: dout <= 8'b01100010; //  500 :  98 - 0x62
      12'h1F5: dout <= 8'b00100001; //  501 :  33 - 0x21
      12'h1F6: dout <= 8'b00000000; //  502 :   0 - 0x0
      12'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      12'h1F8: dout <= 8'b10000111; //  504 : 135 - 0x87 -- Sprite 0x3f
      12'h1F9: dout <= 8'b10000111; //  505 : 135 - 0x87
      12'h1FA: dout <= 8'b00000111; //  506 :   7 - 0x7
      12'h1FB: dout <= 8'b00001111; //  507 :  15 - 0xf
      12'h1FC: dout <= 8'b00001111; //  508 :  15 - 0xf
      12'h1FD: dout <= 8'b00011111; //  509 :  31 - 0x1f
      12'h1FE: dout <= 8'b10011111; //  510 : 159 - 0x9f
      12'h1FF: dout <= 8'b10001111; //  511 : 143 - 0x8f
      12'h200: dout <= 8'b01000100; //  512 :  68 - 0x44 -- Sprite 0x40
      12'h201: dout <= 8'b01000100; //  513 :  68 - 0x44
      12'h202: dout <= 8'b01000100; //  514 :  68 - 0x44
      12'h203: dout <= 8'b01000100; //  515 :  68 - 0x44
      12'h204: dout <= 8'b01000100; //  516 :  68 - 0x44
      12'h205: dout <= 8'b01000110; //  517 :  70 - 0x46
      12'h206: dout <= 8'b01000110; //  518 :  70 - 0x46
      12'h207: dout <= 8'b01000111; //  519 :  71 - 0x47
      12'h208: dout <= 8'b00010000; //  520 :  16 - 0x10 -- Sprite 0x41
      12'h209: dout <= 8'b00111000; //  521 :  56 - 0x38
      12'h20A: dout <= 8'b01111100; //  522 : 124 - 0x7c
      12'h20B: dout <= 8'b01111000; //  523 : 120 - 0x78
      12'h20C: dout <= 8'b00110000; //  524 :  48 - 0x30
      12'h20D: dout <= 8'b00000010; //  525 :   2 - 0x2
      12'h20E: dout <= 8'b00000101; //  526 :   5 - 0x5
      12'h20F: dout <= 8'b00000010; //  527 :   2 - 0x2
      12'h210: dout <= 8'b00010000; //  528 :  16 - 0x10 -- Sprite 0x42
      12'h211: dout <= 8'b00111000; //  529 :  56 - 0x38
      12'h212: dout <= 8'b01111100; //  530 : 124 - 0x7c
      12'h213: dout <= 8'b11111000; //  531 : 248 - 0xf8
      12'h214: dout <= 8'b01110000; //  532 : 112 - 0x70
      12'h215: dout <= 8'b00100000; //  533 :  32 - 0x20
      12'h216: dout <= 8'b00000001; //  534 :   1 - 0x1
      12'h217: dout <= 8'b00000010; //  535 :   2 - 0x2
      12'h218: dout <= 8'b01000100; //  536 :  68 - 0x44 -- Sprite 0x43
      12'h219: dout <= 8'b01000100; //  537 :  68 - 0x44
      12'h21A: dout <= 8'b01000100; //  538 :  68 - 0x44
      12'h21B: dout <= 8'b01000100; //  539 :  68 - 0x44
      12'h21C: dout <= 8'b10000100; //  540 : 132 - 0x84
      12'h21D: dout <= 8'b10000100; //  541 : 132 - 0x84
      12'h21E: dout <= 8'b00000100; //  542 :   4 - 0x4
      12'h21F: dout <= 8'b00001100; //  543 :  12 - 0xc
      12'h220: dout <= 8'b00010000; //  544 :  16 - 0x10 -- Sprite 0x44
      12'h221: dout <= 8'b00111000; //  545 :  56 - 0x38
      12'h222: dout <= 8'b01111100; //  546 : 124 - 0x7c
      12'h223: dout <= 8'b11111000; //  547 : 248 - 0xf8
      12'h224: dout <= 8'b01110000; //  548 : 112 - 0x70
      12'h225: dout <= 8'b00100010; //  549 :  34 - 0x22
      12'h226: dout <= 8'b00000101; //  550 :   5 - 0x5
      12'h227: dout <= 8'b00000010; //  551 :   2 - 0x2
      12'h228: dout <= 8'b01001111; //  552 :  79 - 0x4f -- Sprite 0x45
      12'h229: dout <= 8'b01000111; //  553 :  71 - 0x47
      12'h22A: dout <= 8'b01000111; //  554 :  71 - 0x47
      12'h22B: dout <= 8'b01000111; //  555 :  71 - 0x47
      12'h22C: dout <= 8'b01000111; //  556 :  71 - 0x47
      12'h22D: dout <= 8'b01000111; //  557 :  71 - 0x47
      12'h22E: dout <= 8'b01000111; //  558 :  71 - 0x47
      12'h22F: dout <= 8'b01000111; //  559 :  71 - 0x47
      12'h230: dout <= 8'b10100000; //  560 : 160 - 0xa0 -- Sprite 0x46
      12'h231: dout <= 8'b10011111; //  561 : 159 - 0x9f
      12'h232: dout <= 8'b11000000; //  562 : 192 - 0xc0
      12'h233: dout <= 8'b11100000; //  563 : 224 - 0xe0
      12'h234: dout <= 8'b11111000; //  564 : 248 - 0xf8
      12'h235: dout <= 8'b11111111; //  565 : 255 - 0xff
      12'h236: dout <= 8'b11111111; //  566 : 255 - 0xff
      12'h237: dout <= 8'b11111111; //  567 : 255 - 0xff
      12'h238: dout <= 8'b00001100; //  568 :  12 - 0xc -- Sprite 0x47
      12'h239: dout <= 8'b11110000; //  569 : 240 - 0xf0
      12'h23A: dout <= 8'b00000000; //  570 :   0 - 0x0
      12'h23B: dout <= 8'b00000000; //  571 :   0 - 0x0
      12'h23C: dout <= 8'b00000001; //  572 :   1 - 0x1
      12'h23D: dout <= 8'b11111111; //  573 : 255 - 0xff
      12'h23E: dout <= 8'b11111111; //  574 : 255 - 0xff
      12'h23F: dout <= 8'b11111111; //  575 : 255 - 0xff
      12'h240: dout <= 8'b00001100; //  576 :  12 - 0xc -- Sprite 0x48
      12'h241: dout <= 8'b00011101; //  577 :  29 - 0x1d
      12'h242: dout <= 8'b00111000; //  578 :  56 - 0x38
      12'h243: dout <= 8'b01111110; //  579 : 126 - 0x7e
      12'h244: dout <= 8'b11111110; //  580 : 254 - 0xfe
      12'h245: dout <= 8'b11111111; //  581 : 255 - 0xff
      12'h246: dout <= 8'b11111111; //  582 : 255 - 0xff
      12'h247: dout <= 8'b11111111; //  583 : 255 - 0xff
      12'h248: dout <= 8'b11111111; //  584 : 255 - 0xff -- Sprite 0x49
      12'h249: dout <= 8'b11111111; //  585 : 255 - 0xff
      12'h24A: dout <= 8'b11111111; //  586 : 255 - 0xff
      12'h24B: dout <= 8'b11111111; //  587 : 255 - 0xff
      12'h24C: dout <= 8'b11111111; //  588 : 255 - 0xff
      12'h24D: dout <= 8'b11111111; //  589 : 255 - 0xff
      12'h24E: dout <= 8'b11111111; //  590 : 255 - 0xff
      12'h24F: dout <= 8'b11111111; //  591 : 255 - 0xff
      12'h250: dout <= 8'b11111111; //  592 : 255 - 0xff -- Sprite 0x4a
      12'h251: dout <= 8'b11101111; //  593 : 239 - 0xef
      12'h252: dout <= 8'b11111101; //  594 : 253 - 0xfd
      12'h253: dout <= 8'b11111111; //  595 : 255 - 0xff
      12'h254: dout <= 8'b11111111; //  596 : 255 - 0xff
      12'h255: dout <= 8'b11101111; //  597 : 239 - 0xef
      12'h256: dout <= 8'b11111110; //  598 : 254 - 0xfe
      12'h257: dout <= 8'b11111111; //  599 : 255 - 0xff
      12'h258: dout <= 8'b11111111; //  600 : 255 - 0xff -- Sprite 0x4b
      12'h259: dout <= 8'b11101010; //  601 : 234 - 0xea
      12'h25A: dout <= 8'b11111111; //  602 : 255 - 0xff
      12'h25B: dout <= 8'b10101111; //  603 : 175 - 0xaf
      12'h25C: dout <= 8'b11111111; //  604 : 255 - 0xff
      12'h25D: dout <= 8'b11111111; //  605 : 255 - 0xff
      12'h25E: dout <= 8'b11111010; //  606 : 250 - 0xfa
      12'h25F: dout <= 8'b11111111; //  607 : 255 - 0xff
      12'h260: dout <= 8'b11111111; //  608 : 255 - 0xff -- Sprite 0x4c
      12'h261: dout <= 8'b11111111; //  609 : 255 - 0xff
      12'h262: dout <= 8'b11111111; //  610 : 255 - 0xff
      12'h263: dout <= 8'b11111111; //  611 : 255 - 0xff
      12'h264: dout <= 8'b11111111; //  612 : 255 - 0xff
      12'h265: dout <= 8'b11111111; //  613 : 255 - 0xff
      12'h266: dout <= 8'b11111110; //  614 : 254 - 0xfe
      12'h267: dout <= 8'b11111111; //  615 : 255 - 0xff
      12'h268: dout <= 8'b11111111; //  616 : 255 - 0xff -- Sprite 0x4d
      12'h269: dout <= 8'b10111111; //  617 : 191 - 0xbf
      12'h26A: dout <= 8'b11111110; //  618 : 254 - 0xfe
      12'h26B: dout <= 8'b10101111; //  619 : 175 - 0xaf
      12'h26C: dout <= 8'b11111111; //  620 : 255 - 0xff
      12'h26D: dout <= 8'b11111111; //  621 : 255 - 0xff
      12'h26E: dout <= 8'b11101111; //  622 : 239 - 0xef
      12'h26F: dout <= 8'b11111111; //  623 : 255 - 0xff
      12'h270: dout <= 8'b11111111; //  624 : 255 - 0xff -- Sprite 0x4e
      12'h271: dout <= 8'b11111111; //  625 : 255 - 0xff
      12'h272: dout <= 8'b11111011; //  626 : 251 - 0xfb
      12'h273: dout <= 8'b11111111; //  627 : 255 - 0xff
      12'h274: dout <= 8'b11111111; //  628 : 255 - 0xff
      12'h275: dout <= 8'b11111111; //  629 : 255 - 0xff
      12'h276: dout <= 8'b11111110; //  630 : 254 - 0xfe
      12'h277: dout <= 8'b11111111; //  631 : 255 - 0xff
      12'h278: dout <= 8'b11111111; //  632 : 255 - 0xff -- Sprite 0x4f
      12'h279: dout <= 8'b11111111; //  633 : 255 - 0xff
      12'h27A: dout <= 8'b11110111; //  634 : 247 - 0xf7
      12'h27B: dout <= 8'b11111110; //  635 : 254 - 0xfe
      12'h27C: dout <= 8'b11111011; //  636 : 251 - 0xfb
      12'h27D: dout <= 8'b11111111; //  637 : 255 - 0xff
      12'h27E: dout <= 8'b11101111; //  638 : 239 - 0xef
      12'h27F: dout <= 8'b11111101; //  639 : 253 - 0xfd
      12'h280: dout <= 8'b11111111; //  640 : 255 - 0xff -- Sprite 0x50
      12'h281: dout <= 8'b11111111; //  641 : 255 - 0xff
      12'h282: dout <= 8'b00000011; //  642 :   3 - 0x3
      12'h283: dout <= 8'b00000001; //  643 :   1 - 0x1
      12'h284: dout <= 8'b11101110; //  644 : 238 - 0xee
      12'h285: dout <= 8'b00000000; //  645 :   0 - 0x0
      12'h286: dout <= 8'b11101110; //  646 : 238 - 0xee
      12'h287: dout <= 8'b11101110; //  647 : 238 - 0xee
      12'h288: dout <= 8'b11111111; //  648 : 255 - 0xff -- Sprite 0x51
      12'h289: dout <= 8'b11111111; //  649 : 255 - 0xff
      12'h28A: dout <= 8'b00000011; //  650 :   3 - 0x3
      12'h28B: dout <= 8'b00000001; //  651 :   1 - 0x1
      12'h28C: dout <= 8'b11101110; //  652 : 238 - 0xee
      12'h28D: dout <= 8'b00000000; //  653 :   0 - 0x0
      12'h28E: dout <= 8'b11101110; //  654 : 238 - 0xee
      12'h28F: dout <= 8'b11101110; //  655 : 238 - 0xee
      12'h290: dout <= 8'b11111111; //  656 : 255 - 0xff -- Sprite 0x52
      12'h291: dout <= 8'b11111111; //  657 : 255 - 0xff
      12'h292: dout <= 8'b00000001; //  658 :   1 - 0x1
      12'h293: dout <= 8'b00000000; //  659 :   0 - 0x0
      12'h294: dout <= 8'b11100000; //  660 : 224 - 0xe0
      12'h295: dout <= 8'b00001111; //  661 :  15 - 0xf
      12'h296: dout <= 8'b11111111; //  662 : 255 - 0xff
      12'h297: dout <= 8'b11111011; //  663 : 251 - 0xfb
      12'h298: dout <= 8'b11111111; //  664 : 255 - 0xff -- Sprite 0x53
      12'h299: dout <= 8'b11111111; //  665 : 255 - 0xff
      12'h29A: dout <= 8'b10000011; //  666 : 131 - 0x83
      12'h29B: dout <= 8'b00000001; //  667 :   1 - 0x1
      12'h29C: dout <= 8'b11101110; //  668 : 238 - 0xee
      12'h29D: dout <= 8'b00000000; //  669 :   0 - 0x0
      12'h29E: dout <= 8'b11111111; //  670 : 255 - 0xff
      12'h29F: dout <= 8'b11111111; //  671 : 255 - 0xff
      12'h2A0: dout <= 8'b11111111; //  672 : 255 - 0xff -- Sprite 0x54
      12'h2A1: dout <= 8'b11111111; //  673 : 255 - 0xff
      12'h2A2: dout <= 8'b00000001; //  674 :   1 - 0x1
      12'h2A3: dout <= 8'b00000000; //  675 :   0 - 0x0
      12'h2A4: dout <= 8'b10111000; //  676 : 184 - 0xb8
      12'h2A5: dout <= 8'b11000011; //  677 : 195 - 0xc3
      12'h2A6: dout <= 8'b11111011; //  678 : 251 - 0xfb
      12'h2A7: dout <= 8'b11111011; //  679 : 251 - 0xfb
      12'h2A8: dout <= 8'b11111111; //  680 : 255 - 0xff -- Sprite 0x55
      12'h2A9: dout <= 8'b11111111; //  681 : 255 - 0xff
      12'h2AA: dout <= 8'b10000011; //  682 : 131 - 0x83
      12'h2AB: dout <= 8'b00000001; //  683 :   1 - 0x1
      12'h2AC: dout <= 8'b11101110; //  684 : 238 - 0xee
      12'h2AD: dout <= 8'b00000000; //  685 :   0 - 0x0
      12'h2AE: dout <= 8'b11101110; //  686 : 238 - 0xee
      12'h2AF: dout <= 8'b11101110; //  687 : 238 - 0xee
      12'h2B0: dout <= 8'b11111111; //  688 : 255 - 0xff -- Sprite 0x56
      12'h2B1: dout <= 8'b11111111; //  689 : 255 - 0xff
      12'h2B2: dout <= 8'b00011111; //  690 :  31 - 0x1f
      12'h2B3: dout <= 8'b00001111; //  691 :  15 - 0xf
      12'h2B4: dout <= 8'b11101111; //  692 : 239 - 0xef
      12'h2B5: dout <= 8'b00001111; //  693 :  15 - 0xf
      12'h2B6: dout <= 8'b11101111; //  694 : 239 - 0xef
      12'h2B7: dout <= 8'b11101111; //  695 : 239 - 0xef
      12'h2B8: dout <= 8'b11111111; //  696 : 255 - 0xff -- Sprite 0x57
      12'h2B9: dout <= 8'b11111111; //  697 : 255 - 0xff
      12'h2BA: dout <= 8'b00010001; //  698 :  17 - 0x11
      12'h2BB: dout <= 8'b00000000; //  699 :   0 - 0x0
      12'h2BC: dout <= 8'b11101110; //  700 : 238 - 0xee
      12'h2BD: dout <= 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout <= 8'b11101110; //  702 : 238 - 0xee
      12'h2BF: dout <= 8'b11101110; //  703 : 238 - 0xee
      12'h2C0: dout <= 8'b11111111; //  704 : 255 - 0xff -- Sprite 0x58
      12'h2C1: dout <= 8'b11111111; //  705 : 255 - 0xff
      12'h2C2: dout <= 8'b01110001; //  706 : 113 - 0x71
      12'h2C3: dout <= 8'b00110000; //  707 :  48 - 0x30
      12'h2C4: dout <= 8'b11111110; //  708 : 254 - 0xfe
      12'h2C5: dout <= 8'b00000000; //  709 :   0 - 0x0
      12'h2C6: dout <= 8'b11111110; //  710 : 254 - 0xfe
      12'h2C7: dout <= 8'b11101110; //  711 : 238 - 0xee
      12'h2C8: dout <= 8'b11111111; //  712 : 255 - 0xff -- Sprite 0x59
      12'h2C9: dout <= 8'b11111111; //  713 : 255 - 0xff
      12'h2CA: dout <= 8'b00000011; //  714 :   3 - 0x3
      12'h2CB: dout <= 8'b00000001; //  715 :   1 - 0x1
      12'h2CC: dout <= 8'b11101110; //  716 : 238 - 0xee
      12'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      12'h2CE: dout <= 8'b11101110; //  718 : 238 - 0xee
      12'h2CF: dout <= 8'b11101110; //  719 : 238 - 0xee
      12'h2D0: dout <= 8'b11111111; //  720 : 255 - 0xff -- Sprite 0x5a
      12'h2D1: dout <= 8'b11111111; //  721 : 255 - 0xff
      12'h2D2: dout <= 8'b10000011; //  722 : 131 - 0x83
      12'h2D3: dout <= 8'b00000001; //  723 :   1 - 0x1
      12'h2D4: dout <= 8'b11101110; //  724 : 238 - 0xee
      12'h2D5: dout <= 8'b00000000; //  725 :   0 - 0x0
      12'h2D6: dout <= 8'b11101110; //  726 : 238 - 0xee
      12'h2D7: dout <= 8'b11101110; //  727 : 238 - 0xee
      12'h2D8: dout <= 8'b11111111; //  728 : 255 - 0xff -- Sprite 0x5b
      12'h2D9: dout <= 8'b11111111; //  729 : 255 - 0xff
      12'h2DA: dout <= 8'b00000001; //  730 :   1 - 0x1
      12'h2DB: dout <= 8'b00000000; //  731 :   0 - 0x0
      12'h2DC: dout <= 8'b11100000; //  732 : 224 - 0xe0
      12'h2DD: dout <= 8'b00001111; //  733 :  15 - 0xf
      12'h2DE: dout <= 8'b11111111; //  734 : 255 - 0xff
      12'h2DF: dout <= 8'b11111011; //  735 : 251 - 0xfb
      12'h2E0: dout <= 8'b11111111; //  736 : 255 - 0xff -- Sprite 0x5c
      12'h2E1: dout <= 8'b11111111; //  737 : 255 - 0xff
      12'h2E2: dout <= 8'b11111111; //  738 : 255 - 0xff
      12'h2E3: dout <= 8'b11111111; //  739 : 255 - 0xff
      12'h2E4: dout <= 8'b11111111; //  740 : 255 - 0xff
      12'h2E5: dout <= 8'b11111111; //  741 : 255 - 0xff
      12'h2E6: dout <= 8'b11111111; //  742 : 255 - 0xff
      12'h2E7: dout <= 8'b11011101; //  743 : 221 - 0xdd
      12'h2E8: dout <= 8'b11111111; //  744 : 255 - 0xff -- Sprite 0x5d
      12'h2E9: dout <= 8'b11111111; //  745 : 255 - 0xff
      12'h2EA: dout <= 8'b00000001; //  746 :   1 - 0x1
      12'h2EB: dout <= 8'b00000000; //  747 :   0 - 0x0
      12'h2EC: dout <= 8'b11100000; //  748 : 224 - 0xe0
      12'h2ED: dout <= 8'b00001111; //  749 :  15 - 0xf
      12'h2EE: dout <= 8'b11111111; //  750 : 255 - 0xff
      12'h2EF: dout <= 8'b11111011; //  751 : 251 - 0xfb
      12'h2F0: dout <= 8'b11111111; //  752 : 255 - 0xff -- Sprite 0x5e
      12'h2F1: dout <= 8'b11111111; //  753 : 255 - 0xff
      12'h2F2: dout <= 8'b00010001; //  754 :  17 - 0x11
      12'h2F3: dout <= 8'b00000000; //  755 :   0 - 0x0
      12'h2F4: dout <= 8'b11101110; //  756 : 238 - 0xee
      12'h2F5: dout <= 8'b00000000; //  757 :   0 - 0x0
      12'h2F6: dout <= 8'b11101110; //  758 : 238 - 0xee
      12'h2F7: dout <= 8'b11101110; //  759 : 238 - 0xee
      12'h2F8: dout <= 8'b10111101; //  760 : 189 - 0xbd -- Sprite 0x5f
      12'h2F9: dout <= 8'b11111111; //  761 : 255 - 0xff
      12'h2FA: dout <= 8'b11111111; //  762 : 255 - 0xff
      12'h2FB: dout <= 8'b11111111; //  763 : 255 - 0xff
      12'h2FC: dout <= 8'b11111111; //  764 : 255 - 0xff
      12'h2FD: dout <= 8'b11111111; //  765 : 255 - 0xff
      12'h2FE: dout <= 8'b11111111; //  766 : 255 - 0xff
      12'h2FF: dout <= 8'b11111111; //  767 : 255 - 0xff
      12'h300: dout <= 8'b11101110; //  768 : 238 - 0xee -- Sprite 0x60
      12'h301: dout <= 8'b00000000; //  769 :   0 - 0x0
      12'h302: dout <= 8'b11111110; //  770 : 254 - 0xfe
      12'h303: dout <= 8'b00000000; //  771 :   0 - 0x0
      12'h304: dout <= 8'b00000001; //  772 :   1 - 0x1
      12'h305: dout <= 8'b00001111; //  773 :  15 - 0xf
      12'h306: dout <= 8'b10001111; //  774 : 143 - 0x8f
      12'h307: dout <= 8'b11111111; //  775 : 255 - 0xff
      12'h308: dout <= 8'b11101110; //  776 : 238 - 0xee -- Sprite 0x61
      12'h309: dout <= 8'b00000000; //  777 :   0 - 0x0
      12'h30A: dout <= 8'b11111100; //  778 : 252 - 0xfc
      12'h30B: dout <= 8'b00000001; //  779 :   1 - 0x1
      12'h30C: dout <= 8'b00000001; //  780 :   1 - 0x1
      12'h30D: dout <= 8'b00000000; //  781 :   0 - 0x0
      12'h30E: dout <= 8'b10001000; //  782 : 136 - 0x88
      12'h30F: dout <= 8'b11111111; //  783 : 255 - 0xff
      12'h310: dout <= 8'b11100011; //  784 : 227 - 0xe3 -- Sprite 0x62
      12'h311: dout <= 8'b00001111; //  785 :  15 - 0xf
      12'h312: dout <= 8'b11101111; //  786 : 239 - 0xef
      12'h313: dout <= 8'b00001111; //  787 :  15 - 0xf
      12'h314: dout <= 8'b00000001; //  788 :   1 - 0x1
      12'h315: dout <= 8'b00000000; //  789 :   0 - 0x0
      12'h316: dout <= 8'b10000000; //  790 : 128 - 0x80
      12'h317: dout <= 8'b11111111; //  791 : 255 - 0xff
      12'h318: dout <= 8'b11001110; //  792 : 206 - 0xce -- Sprite 0x63
      12'h319: dout <= 8'b11110000; //  793 : 240 - 0xf0
      12'h31A: dout <= 8'b11111110; //  794 : 254 - 0xfe
      12'h31B: dout <= 8'b00010000; //  795 :  16 - 0x10
      12'h31C: dout <= 8'b00000000; //  796 :   0 - 0x0
      12'h31D: dout <= 8'b10000000; //  797 : 128 - 0x80
      12'h31E: dout <= 8'b11000001; //  798 : 193 - 0xc1
      12'h31F: dout <= 8'b11111111; //  799 : 255 - 0xff
      12'h320: dout <= 8'b11111011; //  800 : 251 - 0xfb -- Sprite 0x64
      12'h321: dout <= 8'b11000011; //  801 : 195 - 0xc3
      12'h322: dout <= 8'b11111011; //  802 : 251 - 0xfb
      12'h323: dout <= 8'b11000011; //  803 : 195 - 0xc3
      12'h324: dout <= 8'b11000011; //  804 : 195 - 0xc3
      12'h325: dout <= 8'b11000011; //  805 : 195 - 0xc3
      12'h326: dout <= 8'b11100011; //  806 : 227 - 0xe3
      12'h327: dout <= 8'b11111111; //  807 : 255 - 0xff
      12'h328: dout <= 8'b11101110; //  808 : 238 - 0xee -- Sprite 0x65
      12'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout <= 8'b11111110; //  810 : 254 - 0xfe
      12'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      12'h32C: dout <= 8'b00000000; //  812 :   0 - 0x0
      12'h32D: dout <= 8'b00000000; //  813 :   0 - 0x0
      12'h32E: dout <= 8'b10001000; //  814 : 136 - 0x88
      12'h32F: dout <= 8'b11111111; //  815 : 255 - 0xff
      12'h330: dout <= 8'b11101111; //  816 : 239 - 0xef -- Sprite 0x66
      12'h331: dout <= 8'b00001111; //  817 :  15 - 0xf
      12'h332: dout <= 8'b11101111; //  818 : 239 - 0xef
      12'h333: dout <= 8'b00000001; //  819 :   1 - 0x1
      12'h334: dout <= 8'b00000000; //  820 :   0 - 0x0
      12'h335: dout <= 8'b00000000; //  821 :   0 - 0x0
      12'h336: dout <= 8'b10000000; //  822 : 128 - 0x80
      12'h337: dout <= 8'b11111111; //  823 : 255 - 0xff
      12'h338: dout <= 8'b11101110; //  824 : 238 - 0xee -- Sprite 0x67
      12'h339: dout <= 8'b00000000; //  825 :   0 - 0x0
      12'h33A: dout <= 8'b11111110; //  826 : 254 - 0xfe
      12'h33B: dout <= 8'b00000000; //  827 :   0 - 0x0
      12'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      12'h33D: dout <= 8'b00001000; //  829 :   8 - 0x8
      12'h33E: dout <= 8'b10011100; //  830 : 156 - 0x9c
      12'h33F: dout <= 8'b11111111; //  831 : 255 - 0xff
      12'h340: dout <= 8'b11101110; //  832 : 238 - 0xee -- Sprite 0x68
      12'h341: dout <= 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout <= 8'b11101110; //  834 : 238 - 0xee
      12'h343: dout <= 8'b00000000; //  835 :   0 - 0x0
      12'h344: dout <= 8'b00000000; //  836 :   0 - 0x0
      12'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout <= 8'b10001000; //  838 : 136 - 0x88
      12'h347: dout <= 8'b11111111; //  839 : 255 - 0xff
      12'h348: dout <= 8'b11101110; //  840 : 238 - 0xee -- Sprite 0x69
      12'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout <= 8'b11101110; //  842 : 238 - 0xee
      12'h34B: dout <= 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout <= 8'b00000000; //  844 :   0 - 0x0
      12'h34D: dout <= 8'b00000000; //  845 :   0 - 0x0
      12'h34E: dout <= 8'b10000001; //  846 : 129 - 0x81
      12'h34F: dout <= 8'b11111111; //  847 : 255 - 0xff
      12'h350: dout <= 8'b11101110; //  848 : 238 - 0xee -- Sprite 0x6a
      12'h351: dout <= 8'b00000000; //  849 :   0 - 0x0
      12'h352: dout <= 8'b11101110; //  850 : 238 - 0xee
      12'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      12'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout <= 8'b10000000; //  853 : 128 - 0x80
      12'h356: dout <= 8'b11000001; //  854 : 193 - 0xc1
      12'h357: dout <= 8'b11111111; //  855 : 255 - 0xff
      12'h358: dout <= 8'b11100011; //  856 : 227 - 0xe3 -- Sprite 0x6b
      12'h359: dout <= 8'b00001111; //  857 :  15 - 0xf
      12'h35A: dout <= 8'b11101111; //  858 : 239 - 0xef
      12'h35B: dout <= 8'b00001111; //  859 :  15 - 0xf
      12'h35C: dout <= 8'b00000001; //  860 :   1 - 0x1
      12'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout <= 8'b10000000; //  862 : 128 - 0x80
      12'h35F: dout <= 8'b11111111; //  863 : 255 - 0xff
      12'h360: dout <= 8'b10011001; //  864 : 153 - 0x99 -- Sprite 0x6c
      12'h361: dout <= 8'b11100011; //  865 : 227 - 0xe3
      12'h362: dout <= 8'b11110011; //  866 : 243 - 0xf3
      12'h363: dout <= 8'b11000111; //  867 : 199 - 0xc7
      12'h364: dout <= 8'b10000001; //  868 : 129 - 0x81
      12'h365: dout <= 8'b10001000; //  869 : 136 - 0x88
      12'h366: dout <= 8'b11001100; //  870 : 204 - 0xcc
      12'h367: dout <= 8'b11111111; //  871 : 255 - 0xff
      12'h368: dout <= 8'b11100011; //  872 : 227 - 0xe3 -- Sprite 0x6d
      12'h369: dout <= 8'b00001111; //  873 :  15 - 0xf
      12'h36A: dout <= 8'b11101111; //  874 : 239 - 0xef
      12'h36B: dout <= 8'b00001111; //  875 :  15 - 0xf
      12'h36C: dout <= 8'b00001111; //  876 :  15 - 0xf
      12'h36D: dout <= 8'b00001111; //  877 :  15 - 0xf
      12'h36E: dout <= 8'b10001111; //  878 : 143 - 0x8f
      12'h36F: dout <= 8'b11111111; //  879 : 255 - 0xff
      12'h370: dout <= 8'b11101110; //  880 : 238 - 0xee -- Sprite 0x6e
      12'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout <= 8'b11101110; //  882 : 238 - 0xee
      12'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      12'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      12'h375: dout <= 8'b10000000; //  885 : 128 - 0x80
      12'h376: dout <= 8'b11000001; //  886 : 193 - 0xc1
      12'h377: dout <= 8'b11111111; //  887 : 255 - 0xff
      12'h378: dout <= 8'b11111111; //  888 : 255 - 0xff -- Sprite 0x6f
      12'h379: dout <= 8'b11111111; //  889 : 255 - 0xff
      12'h37A: dout <= 8'b11111111; //  890 : 255 - 0xff
      12'h37B: dout <= 8'b10111101; //  891 : 189 - 0xbd
      12'h37C: dout <= 8'b11111111; //  892 : 255 - 0xff
      12'h37D: dout <= 8'b11011011; //  893 : 219 - 0xdb
      12'h37E: dout <= 8'b11111111; //  894 : 255 - 0xff
      12'h37F: dout <= 8'b11111111; //  895 : 255 - 0xff
      12'h380: dout <= 8'b11111011; //  896 : 251 - 0xfb -- Sprite 0x70
      12'h381: dout <= 8'b11101111; //  897 : 239 - 0xef
      12'h382: dout <= 8'b11011111; //  898 : 223 - 0xdf
      12'h383: dout <= 8'b11111111; //  899 : 255 - 0xff
      12'h384: dout <= 8'b10111111; //  900 : 191 - 0xbf
      12'h385: dout <= 8'b10111111; //  901 : 191 - 0xbf
      12'h386: dout <= 8'b11111110; //  902 : 254 - 0xfe
      12'h387: dout <= 8'b11111111; //  903 : 255 - 0xff
      12'h388: dout <= 8'b11011111; //  904 : 223 - 0xdf -- Sprite 0x71
      12'h389: dout <= 8'b11110111; //  905 : 247 - 0xf7
      12'h38A: dout <= 8'b11111011; //  906 : 251 - 0xfb
      12'h38B: dout <= 8'b11111111; //  907 : 255 - 0xff
      12'h38C: dout <= 8'b11111101; //  908 : 253 - 0xfd
      12'h38D: dout <= 8'b11111101; //  909 : 253 - 0xfd
      12'h38E: dout <= 8'b01111111; //  910 : 127 - 0x7f
      12'h38F: dout <= 8'b11111111; //  911 : 255 - 0xff
      12'h390: dout <= 8'b11111111; //  912 : 255 - 0xff -- Sprite 0x72
      12'h391: dout <= 8'b11111111; //  913 : 255 - 0xff
      12'h392: dout <= 8'b11111111; //  914 : 255 - 0xff
      12'h393: dout <= 8'b11111111; //  915 : 255 - 0xff
      12'h394: dout <= 8'b11111111; //  916 : 255 - 0xff
      12'h395: dout <= 8'b11111111; //  917 : 255 - 0xff
      12'h396: dout <= 8'b11111111; //  918 : 255 - 0xff
      12'h397: dout <= 8'b11111111; //  919 : 255 - 0xff
      12'h398: dout <= 8'b11111111; //  920 : 255 - 0xff -- Sprite 0x73
      12'h399: dout <= 8'b11111110; //  921 : 254 - 0xfe
      12'h39A: dout <= 8'b10111111; //  922 : 191 - 0xbf
      12'h39B: dout <= 8'b10111111; //  923 : 191 - 0xbf
      12'h39C: dout <= 8'b11111111; //  924 : 255 - 0xff
      12'h39D: dout <= 8'b11011111; //  925 : 223 - 0xdf
      12'h39E: dout <= 8'b11101111; //  926 : 239 - 0xef
      12'h39F: dout <= 8'b11111011; //  927 : 251 - 0xfb
      12'h3A0: dout <= 8'b11111111; //  928 : 255 - 0xff -- Sprite 0x74
      12'h3A1: dout <= 8'b01111111; //  929 : 127 - 0x7f
      12'h3A2: dout <= 8'b11111101; //  930 : 253 - 0xfd
      12'h3A3: dout <= 8'b11111101; //  931 : 253 - 0xfd
      12'h3A4: dout <= 8'b11111111; //  932 : 255 - 0xff
      12'h3A5: dout <= 8'b11111011; //  933 : 251 - 0xfb
      12'h3A6: dout <= 8'b11110111; //  934 : 247 - 0xf7
      12'h3A7: dout <= 8'b11011111; //  935 : 223 - 0xdf
      12'h3A8: dout <= 8'b11111111; //  936 : 255 - 0xff -- Sprite 0x75
      12'h3A9: dout <= 8'b11111111; //  937 : 255 - 0xff
      12'h3AA: dout <= 8'b11111111; //  938 : 255 - 0xff
      12'h3AB: dout <= 8'b11111111; //  939 : 255 - 0xff
      12'h3AC: dout <= 8'b11111111; //  940 : 255 - 0xff
      12'h3AD: dout <= 8'b11111111; //  941 : 255 - 0xff
      12'h3AE: dout <= 8'b11111111; //  942 : 255 - 0xff
      12'h3AF: dout <= 8'b11111111; //  943 : 255 - 0xff
      12'h3B0: dout <= 8'b11111111; //  944 : 255 - 0xff -- Sprite 0x76
      12'h3B1: dout <= 8'b11111111; //  945 : 255 - 0xff
      12'h3B2: dout <= 8'b11111111; //  946 : 255 - 0xff
      12'h3B3: dout <= 8'b11111111; //  947 : 255 - 0xff
      12'h3B4: dout <= 8'b11111111; //  948 : 255 - 0xff
      12'h3B5: dout <= 8'b11111111; //  949 : 255 - 0xff
      12'h3B6: dout <= 8'b11111111; //  950 : 255 - 0xff
      12'h3B7: dout <= 8'b11111111; //  951 : 255 - 0xff
      12'h3B8: dout <= 8'b11111111; //  952 : 255 - 0xff -- Sprite 0x77
      12'h3B9: dout <= 8'b11111111; //  953 : 255 - 0xff
      12'h3BA: dout <= 8'b11111111; //  954 : 255 - 0xff
      12'h3BB: dout <= 8'b11111111; //  955 : 255 - 0xff
      12'h3BC: dout <= 8'b11111111; //  956 : 255 - 0xff
      12'h3BD: dout <= 8'b11111111; //  957 : 255 - 0xff
      12'h3BE: dout <= 8'b11111111; //  958 : 255 - 0xff
      12'h3BF: dout <= 8'b11111111; //  959 : 255 - 0xff
      12'h3C0: dout <= 8'b11111111; //  960 : 255 - 0xff -- Sprite 0x78
      12'h3C1: dout <= 8'b11111111; //  961 : 255 - 0xff
      12'h3C2: dout <= 8'b11111111; //  962 : 255 - 0xff
      12'h3C3: dout <= 8'b11111111; //  963 : 255 - 0xff
      12'h3C4: dout <= 8'b11111111; //  964 : 255 - 0xff
      12'h3C5: dout <= 8'b11111111; //  965 : 255 - 0xff
      12'h3C6: dout <= 8'b11111111; //  966 : 255 - 0xff
      12'h3C7: dout <= 8'b11111111; //  967 : 255 - 0xff
      12'h3C8: dout <= 8'b11111111; //  968 : 255 - 0xff -- Sprite 0x79
      12'h3C9: dout <= 8'b11111111; //  969 : 255 - 0xff
      12'h3CA: dout <= 8'b11111111; //  970 : 255 - 0xff
      12'h3CB: dout <= 8'b11111111; //  971 : 255 - 0xff
      12'h3CC: dout <= 8'b11111111; //  972 : 255 - 0xff
      12'h3CD: dout <= 8'b11111111; //  973 : 255 - 0xff
      12'h3CE: dout <= 8'b11111111; //  974 : 255 - 0xff
      12'h3CF: dout <= 8'b11111111; //  975 : 255 - 0xff
      12'h3D0: dout <= 8'b11111111; //  976 : 255 - 0xff -- Sprite 0x7a
      12'h3D1: dout <= 8'b11111111; //  977 : 255 - 0xff
      12'h3D2: dout <= 8'b11111111; //  978 : 255 - 0xff
      12'h3D3: dout <= 8'b11111111; //  979 : 255 - 0xff
      12'h3D4: dout <= 8'b11111111; //  980 : 255 - 0xff
      12'h3D5: dout <= 8'b11111111; //  981 : 255 - 0xff
      12'h3D6: dout <= 8'b11111111; //  982 : 255 - 0xff
      12'h3D7: dout <= 8'b11111111; //  983 : 255 - 0xff
      12'h3D8: dout <= 8'b11111111; //  984 : 255 - 0xff -- Sprite 0x7b
      12'h3D9: dout <= 8'b11111111; //  985 : 255 - 0xff
      12'h3DA: dout <= 8'b11111111; //  986 : 255 - 0xff
      12'h3DB: dout <= 8'b11111111; //  987 : 255 - 0xff
      12'h3DC: dout <= 8'b11111111; //  988 : 255 - 0xff
      12'h3DD: dout <= 8'b11111111; //  989 : 255 - 0xff
      12'h3DE: dout <= 8'b11111111; //  990 : 255 - 0xff
      12'h3DF: dout <= 8'b11111111; //  991 : 255 - 0xff
      12'h3E0: dout <= 8'b11111111; //  992 : 255 - 0xff -- Sprite 0x7c
      12'h3E1: dout <= 8'b11111111; //  993 : 255 - 0xff
      12'h3E2: dout <= 8'b11111111; //  994 : 255 - 0xff
      12'h3E3: dout <= 8'b11111111; //  995 : 255 - 0xff
      12'h3E4: dout <= 8'b11111111; //  996 : 255 - 0xff
      12'h3E5: dout <= 8'b11111111; //  997 : 255 - 0xff
      12'h3E6: dout <= 8'b11111111; //  998 : 255 - 0xff
      12'h3E7: dout <= 8'b11111111; //  999 : 255 - 0xff
      12'h3E8: dout <= 8'b11111111; // 1000 : 255 - 0xff -- Sprite 0x7d
      12'h3E9: dout <= 8'b11111111; // 1001 : 255 - 0xff
      12'h3EA: dout <= 8'b11111111; // 1002 : 255 - 0xff
      12'h3EB: dout <= 8'b11111111; // 1003 : 255 - 0xff
      12'h3EC: dout <= 8'b11111111; // 1004 : 255 - 0xff
      12'h3ED: dout <= 8'b11111111; // 1005 : 255 - 0xff
      12'h3EE: dout <= 8'b11111111; // 1006 : 255 - 0xff
      12'h3EF: dout <= 8'b11111111; // 1007 : 255 - 0xff
      12'h3F0: dout <= 8'b11111111; // 1008 : 255 - 0xff -- Sprite 0x7e
      12'h3F1: dout <= 8'b11111111; // 1009 : 255 - 0xff
      12'h3F2: dout <= 8'b11111111; // 1010 : 255 - 0xff
      12'h3F3: dout <= 8'b11111111; // 1011 : 255 - 0xff
      12'h3F4: dout <= 8'b11111111; // 1012 : 255 - 0xff
      12'h3F5: dout <= 8'b11111111; // 1013 : 255 - 0xff
      12'h3F6: dout <= 8'b11111111; // 1014 : 255 - 0xff
      12'h3F7: dout <= 8'b11111111; // 1015 : 255 - 0xff
      12'h3F8: dout <= 8'b11111111; // 1016 : 255 - 0xff -- Sprite 0x7f
      12'h3F9: dout <= 8'b11111111; // 1017 : 255 - 0xff
      12'h3FA: dout <= 8'b11111111; // 1018 : 255 - 0xff
      12'h3FB: dout <= 8'b11111111; // 1019 : 255 - 0xff
      12'h3FC: dout <= 8'b11111111; // 1020 : 255 - 0xff
      12'h3FD: dout <= 8'b11111111; // 1021 : 255 - 0xff
      12'h3FE: dout <= 8'b11111111; // 1022 : 255 - 0xff
      12'h3FF: dout <= 8'b11111111; // 1023 : 255 - 0xff
      12'h400: dout <= 8'b10111111; // 1024 : 191 - 0xbf -- Sprite 0x80
      12'h401: dout <= 8'b11110111; // 1025 : 247 - 0xf7
      12'h402: dout <= 8'b11111101; // 1026 : 253 - 0xfd
      12'h403: dout <= 8'b11011111; // 1027 : 223 - 0xdf
      12'h404: dout <= 8'b11111011; // 1028 : 251 - 0xfb
      12'h405: dout <= 8'b10111111; // 1029 : 191 - 0xbf
      12'h406: dout <= 8'b11111110; // 1030 : 254 - 0xfe
      12'h407: dout <= 8'b11101111; // 1031 : 239 - 0xef
      12'h408: dout <= 8'b11111111; // 1032 : 255 - 0xff -- Sprite 0x81
      12'h409: dout <= 8'b11101110; // 1033 : 238 - 0xee
      12'h40A: dout <= 8'b11111111; // 1034 : 255 - 0xff
      12'h40B: dout <= 8'b11011111; // 1035 : 223 - 0xdf
      12'h40C: dout <= 8'b01110111; // 1036 : 119 - 0x77
      12'h40D: dout <= 8'b11111101; // 1037 : 253 - 0xfd
      12'h40E: dout <= 8'b11011111; // 1038 : 223 - 0xdf
      12'h40F: dout <= 8'b10111111; // 1039 : 191 - 0xbf
      12'h410: dout <= 8'b11111110; // 1040 : 254 - 0xfe -- Sprite 0x82
      12'h411: dout <= 8'b11101111; // 1041 : 239 - 0xef
      12'h412: dout <= 8'b10111111; // 1042 : 191 - 0xbf
      12'h413: dout <= 8'b11110111; // 1043 : 247 - 0xf7
      12'h414: dout <= 8'b11111101; // 1044 : 253 - 0xfd
      12'h415: dout <= 8'b11011111; // 1045 : 223 - 0xdf
      12'h416: dout <= 8'b11111011; // 1046 : 251 - 0xfb
      12'h417: dout <= 8'b10111111; // 1047 : 191 - 0xbf
      12'h418: dout <= 8'b11101111; // 1048 : 239 - 0xef -- Sprite 0x83
      12'h419: dout <= 8'b11111111; // 1049 : 255 - 0xff
      12'h41A: dout <= 8'b10111011; // 1050 : 187 - 0xbb
      12'h41B: dout <= 8'b11111111; // 1051 : 255 - 0xff
      12'h41C: dout <= 8'b11110111; // 1052 : 247 - 0xf7
      12'h41D: dout <= 8'b11011101; // 1053 : 221 - 0xdd
      12'h41E: dout <= 8'b01111111; // 1054 : 127 - 0x7f
      12'h41F: dout <= 8'b11110111; // 1055 : 247 - 0xf7
      12'h420: dout <= 8'b11111111; // 1056 : 255 - 0xff -- Sprite 0x84
      12'h421: dout <= 8'b11101110; // 1057 : 238 - 0xee
      12'h422: dout <= 8'b11111011; // 1058 : 251 - 0xfb
      12'h423: dout <= 8'b10111111; // 1059 : 191 - 0xbf
      12'h424: dout <= 8'b01111111; // 1060 : 127 - 0x7f
      12'h425: dout <= 8'b11101101; // 1061 : 237 - 0xed
      12'h426: dout <= 8'b11111111; // 1062 : 255 - 0xff
      12'h427: dout <= 8'b10111111; // 1063 : 191 - 0xbf
      12'h428: dout <= 8'b11111111; // 1064 : 255 - 0xff -- Sprite 0x85
      12'h429: dout <= 8'b10111111; // 1065 : 191 - 0xbf
      12'h42A: dout <= 8'b01111101; // 1066 : 125 - 0x7d
      12'h42B: dout <= 8'b11110111; // 1067 : 247 - 0xf7
      12'h42C: dout <= 8'b11011011; // 1068 : 219 - 0xdb
      12'h42D: dout <= 8'b11111101; // 1069 : 253 - 0xfd
      12'h42E: dout <= 8'b01111110; // 1070 : 126 - 0x7e
      12'h42F: dout <= 8'b11111011; // 1071 : 251 - 0xfb
      12'h430: dout <= 8'b11111111; // 1072 : 255 - 0xff -- Sprite 0x86
      12'h431: dout <= 8'b11110111; // 1073 : 247 - 0xf7
      12'h432: dout <= 8'b11111111; // 1074 : 255 - 0xff
      12'h433: dout <= 8'b11011101; // 1075 : 221 - 0xdd
      12'h434: dout <= 8'b01111111; // 1076 : 127 - 0x7f
      12'h435: dout <= 8'b11110111; // 1077 : 247 - 0xf7
      12'h436: dout <= 8'b11101111; // 1078 : 239 - 0xef
      12'h437: dout <= 8'b10111101; // 1079 : 189 - 0xbd
      12'h438: dout <= 8'b01011111; // 1080 :  95 - 0x5f -- Sprite 0x87
      12'h439: dout <= 8'b11111101; // 1081 : 253 - 0xfd
      12'h43A: dout <= 8'b11110110; // 1082 : 246 - 0xf6
      12'h43B: dout <= 8'b01111111; // 1083 : 127 - 0x7f
      12'h43C: dout <= 8'b10011111; // 1084 : 159 - 0x9f
      12'h43D: dout <= 8'b11111110; // 1085 : 254 - 0xfe
      12'h43E: dout <= 8'b11111111; // 1086 : 255 - 0xff
      12'h43F: dout <= 8'b11101111; // 1087 : 239 - 0xef
      12'h440: dout <= 8'b11111111; // 1088 : 255 - 0xff -- Sprite 0x88
      12'h441: dout <= 8'b11111111; // 1089 : 255 - 0xff
      12'h442: dout <= 8'b10011111; // 1090 : 159 - 0x9f
      12'h443: dout <= 8'b10110011; // 1091 : 179 - 0xb3
      12'h444: dout <= 8'b11110011; // 1092 : 243 - 0xf3
      12'h445: dout <= 8'b11111111; // 1093 : 255 - 0xff
      12'h446: dout <= 8'b11111111; // 1094 : 255 - 0xff
      12'h447: dout <= 8'b11111111; // 1095 : 255 - 0xff
      12'h448: dout <= 8'b11111111; // 1096 : 255 - 0xff -- Sprite 0x89
      12'h449: dout <= 8'b11001111; // 1097 : 207 - 0xcf
      12'h44A: dout <= 8'b11011111; // 1098 : 223 - 0xdf
      12'h44B: dout <= 8'b11111111; // 1099 : 255 - 0xff
      12'h44C: dout <= 8'b11110011; // 1100 : 243 - 0xf3
      12'h44D: dout <= 8'b11110011; // 1101 : 243 - 0xf3
      12'h44E: dout <= 8'b11111111; // 1102 : 255 - 0xff
      12'h44F: dout <= 8'b11111111; // 1103 : 255 - 0xff
      12'h450: dout <= 8'b10111111; // 1104 : 191 - 0xbf -- Sprite 0x8a
      12'h451: dout <= 8'b11110111; // 1105 : 247 - 0xf7
      12'h452: dout <= 8'b11111101; // 1106 : 253 - 0xfd
      12'h453: dout <= 8'b11111111; // 1107 : 255 - 0xff
      12'h454: dout <= 8'b11111011; // 1108 : 251 - 0xfb
      12'h455: dout <= 8'b10111111; // 1109 : 191 - 0xbf
      12'h456: dout <= 8'b11111110; // 1110 : 254 - 0xfe
      12'h457: dout <= 8'b11101111; // 1111 : 239 - 0xef
      12'h458: dout <= 8'b10111111; // 1112 : 191 - 0xbf -- Sprite 0x8b
      12'h459: dout <= 8'b11111111; // 1113 : 255 - 0xff
      12'h45A: dout <= 8'b11101110; // 1114 : 238 - 0xee
      12'h45B: dout <= 8'b11111111; // 1115 : 255 - 0xff
      12'h45C: dout <= 8'b11011111; // 1116 : 223 - 0xdf
      12'h45D: dout <= 8'b01111101; // 1117 : 125 - 0x7d
      12'h45E: dout <= 8'b11111111; // 1118 : 255 - 0xff
      12'h45F: dout <= 8'b11011111; // 1119 : 223 - 0xdf
      12'h460: dout <= 8'b11111111; // 1120 : 255 - 0xff -- Sprite 0x8c
      12'h461: dout <= 8'b11111000; // 1121 : 248 - 0xf8
      12'h462: dout <= 8'b11100010; // 1122 : 226 - 0xe2
      12'h463: dout <= 8'b11010111; // 1123 : 215 - 0xd7
      12'h464: dout <= 8'b11001111; // 1124 : 207 - 0xcf
      12'h465: dout <= 8'b10011111; // 1125 : 159 - 0x9f
      12'h466: dout <= 8'b10111110; // 1126 : 190 - 0xbe
      12'h467: dout <= 8'b10011101; // 1127 : 157 - 0x9d
      12'h468: dout <= 8'b11111111; // 1128 : 255 - 0xff -- Sprite 0x8d
      12'h469: dout <= 8'b00011111; // 1129 :  31 - 0x1f
      12'h46A: dout <= 8'b10100111; // 1130 : 167 - 0xa7
      12'h46B: dout <= 8'b11000011; // 1131 : 195 - 0xc3
      12'h46C: dout <= 8'b11100011; // 1132 : 227 - 0xe3
      12'h46D: dout <= 8'b01000001; // 1133 :  65 - 0x41
      12'h46E: dout <= 8'b10100001; // 1134 : 161 - 0xa1
      12'h46F: dout <= 8'b00000001; // 1135 :   1 - 0x1
      12'h470: dout <= 8'b10111110; // 1136 : 190 - 0xbe -- Sprite 0x8e
      12'h471: dout <= 8'b11111111; // 1137 : 255 - 0xff
      12'h472: dout <= 8'b11011111; // 1138 : 223 - 0xdf
      12'h473: dout <= 8'b11111111; // 1139 : 255 - 0xff
      12'h474: dout <= 8'b11101111; // 1140 : 239 - 0xef
      12'h475: dout <= 8'b11111111; // 1141 : 255 - 0xff
      12'h476: dout <= 8'b11110111; // 1142 : 247 - 0xf7
      12'h477: dout <= 8'b11111111; // 1143 : 255 - 0xff
      12'h478: dout <= 8'b01111101; // 1144 : 125 - 0x7d -- Sprite 0x8f
      12'h479: dout <= 8'b11111111; // 1145 : 255 - 0xff
      12'h47A: dout <= 8'b11111011; // 1146 : 251 - 0xfb
      12'h47B: dout <= 8'b11111111; // 1147 : 255 - 0xff
      12'h47C: dout <= 8'b11110111; // 1148 : 247 - 0xf7
      12'h47D: dout <= 8'b11111111; // 1149 : 255 - 0xff
      12'h47E: dout <= 8'b11101111; // 1150 : 239 - 0xef
      12'h47F: dout <= 8'b11111111; // 1151 : 255 - 0xff
      12'h480: dout <= 8'b10111110; // 1152 : 190 - 0xbe -- Sprite 0x90
      12'h481: dout <= 8'b11110111; // 1153 : 247 - 0xf7
      12'h482: dout <= 8'b11111111; // 1154 : 255 - 0xff
      12'h483: dout <= 8'b11011111; // 1155 : 223 - 0xdf
      12'h484: dout <= 8'b11111011; // 1156 : 251 - 0xfb
      12'h485: dout <= 8'b11111110; // 1157 : 254 - 0xfe
      12'h486: dout <= 8'b10111111; // 1158 : 191 - 0xbf
      12'h487: dout <= 8'b11110111; // 1159 : 247 - 0xf7
      12'h488: dout <= 8'b11101110; // 1160 : 238 - 0xee -- Sprite 0x91
      12'h489: dout <= 8'b11111111; // 1161 : 255 - 0xff
      12'h48A: dout <= 8'b01111011; // 1162 : 123 - 0x7b
      12'h48B: dout <= 8'b11111101; // 1163 : 253 - 0xfd
      12'h48C: dout <= 8'b11101111; // 1164 : 239 - 0xef
      12'h48D: dout <= 8'b11111111; // 1165 : 255 - 0xff
      12'h48E: dout <= 8'b10111101; // 1166 : 189 - 0xbd
      12'h48F: dout <= 8'b11111111; // 1167 : 255 - 0xff
      12'h490: dout <= 8'b11111011; // 1168 : 251 - 0xfb -- Sprite 0x92
      12'h491: dout <= 8'b10111111; // 1169 : 191 - 0xbf
      12'h492: dout <= 8'b11101111; // 1170 : 239 - 0xef
      12'h493: dout <= 8'b11111101; // 1171 : 253 - 0xfd
      12'h494: dout <= 8'b11111111; // 1172 : 255 - 0xff
      12'h495: dout <= 8'b10111111; // 1173 : 191 - 0xbf
      12'h496: dout <= 8'b11111011; // 1174 : 251 - 0xfb
      12'h497: dout <= 8'b11011111; // 1175 : 223 - 0xdf
      12'h498: dout <= 8'b10111101; // 1176 : 189 - 0xbd -- Sprite 0x93
      12'h499: dout <= 8'b11111111; // 1177 : 255 - 0xff
      12'h49A: dout <= 8'b01110111; // 1178 : 119 - 0x77
      12'h49B: dout <= 8'b11111110; // 1179 : 254 - 0xfe
      12'h49C: dout <= 8'b11011111; // 1180 : 223 - 0xdf
      12'h49D: dout <= 8'b11111011; // 1181 : 251 - 0xfb
      12'h49E: dout <= 8'b11101111; // 1182 : 239 - 0xef
      12'h49F: dout <= 8'b01111111; // 1183 : 127 - 0x7f
      12'h4A0: dout <= 8'b01111111; // 1184 : 127 - 0x7f -- Sprite 0x94
      12'h4A1: dout <= 8'b11110111; // 1185 : 247 - 0xf7
      12'h4A2: dout <= 8'b11011101; // 1186 : 221 - 0xdd
      12'h4A3: dout <= 8'b01111011; // 1187 : 123 - 0x7b
      12'h4A4: dout <= 8'b11111111; // 1188 : 255 - 0xff
      12'h4A5: dout <= 8'b11101110; // 1189 : 238 - 0xee
      12'h4A6: dout <= 8'b10111011; // 1190 : 187 - 0xbb
      12'h4A7: dout <= 8'b11111101; // 1191 : 253 - 0xfd
      12'h4A8: dout <= 8'b11010111; // 1192 : 215 - 0xd7 -- Sprite 0x95
      12'h4A9: dout <= 8'b01111111; // 1193 : 127 - 0x7f
      12'h4AA: dout <= 8'b11111101; // 1194 : 253 - 0xfd
      12'h4AB: dout <= 8'b11101110; // 1195 : 238 - 0xee
      12'h4AC: dout <= 8'b11110111; // 1196 : 247 - 0xf7
      12'h4AD: dout <= 8'b10111011; // 1197 : 187 - 0xbb
      12'h4AE: dout <= 8'b11101111; // 1198 : 239 - 0xef
      12'h4AF: dout <= 8'b11110111; // 1199 : 247 - 0xf7
      12'h4B0: dout <= 8'b10111111; // 1200 : 191 - 0xbf -- Sprite 0x96
      12'h4B1: dout <= 8'b11101110; // 1201 : 238 - 0xee
      12'h4B2: dout <= 8'b11011011; // 1202 : 219 - 0xdb
      12'h4B3: dout <= 8'b11111111; // 1203 : 255 - 0xff
      12'h4B4: dout <= 8'b01110111; // 1204 : 119 - 0x77
      12'h4B5: dout <= 8'b11011101; // 1205 : 221 - 0xdd
      12'h4B6: dout <= 8'b11101111; // 1206 : 239 - 0xef
      12'h4B7: dout <= 8'b11111011; // 1207 : 251 - 0xfb
      12'h4B8: dout <= 8'b11111101; // 1208 : 253 - 0xfd -- Sprite 0x97
      12'h4B9: dout <= 8'b11101110; // 1209 : 238 - 0xee
      12'h4BA: dout <= 8'b11111011; // 1210 : 251 - 0xfb
      12'h4BB: dout <= 8'b11111101; // 1211 : 253 - 0xfd
      12'h4BC: dout <= 8'b11110101; // 1212 : 245 - 0xf5
      12'h4BD: dout <= 8'b11011111; // 1213 : 223 - 0xdf
      12'h4BE: dout <= 8'b01111111; // 1214 : 127 - 0x7f
      12'h4BF: dout <= 8'b10111011; // 1215 : 187 - 0xbb
      12'h4C0: dout <= 8'b11111111; // 1216 : 255 - 0xff -- Sprite 0x98
      12'h4C1: dout <= 8'b11001111; // 1217 : 207 - 0xcf
      12'h4C2: dout <= 8'b11011111; // 1218 : 223 - 0xdf
      12'h4C3: dout <= 8'b11111111; // 1219 : 255 - 0xff
      12'h4C4: dout <= 8'b11110011; // 1220 : 243 - 0xf3
      12'h4C5: dout <= 8'b11110011; // 1221 : 243 - 0xf3
      12'h4C6: dout <= 8'b11111111; // 1222 : 255 - 0xff
      12'h4C7: dout <= 8'b11111111; // 1223 : 255 - 0xff
      12'h4C8: dout <= 8'b11111111; // 1224 : 255 - 0xff -- Sprite 0x99
      12'h4C9: dout <= 8'b11111111; // 1225 : 255 - 0xff
      12'h4CA: dout <= 8'b10011111; // 1226 : 159 - 0x9f
      12'h4CB: dout <= 8'b10110011; // 1227 : 179 - 0xb3
      12'h4CC: dout <= 8'b11110011; // 1228 : 243 - 0xf3
      12'h4CD: dout <= 8'b11111111; // 1229 : 255 - 0xff
      12'h4CE: dout <= 8'b11111111; // 1230 : 255 - 0xff
      12'h4CF: dout <= 8'b11111111; // 1231 : 255 - 0xff
      12'h4D0: dout <= 8'b10111111; // 1232 : 191 - 0xbf -- Sprite 0x9a
      12'h4D1: dout <= 8'b11110111; // 1233 : 247 - 0xf7
      12'h4D2: dout <= 8'b11111111; // 1234 : 255 - 0xff
      12'h4D3: dout <= 8'b11011111; // 1235 : 223 - 0xdf
      12'h4D4: dout <= 8'b11111011; // 1236 : 251 - 0xfb
      12'h4D5: dout <= 8'b11111111; // 1237 : 255 - 0xff
      12'h4D6: dout <= 8'b10111111; // 1238 : 191 - 0xbf
      12'h4D7: dout <= 8'b11110111; // 1239 : 247 - 0xf7
      12'h4D8: dout <= 8'b11011111; // 1240 : 223 - 0xdf -- Sprite 0x9b
      12'h4D9: dout <= 8'b11111111; // 1241 : 255 - 0xff
      12'h4DA: dout <= 8'b01111011; // 1242 : 123 - 0x7b
      12'h4DB: dout <= 8'b11111111; // 1243 : 255 - 0xff
      12'h4DC: dout <= 8'b11101111; // 1244 : 239 - 0xef
      12'h4DD: dout <= 8'b11111101; // 1245 : 253 - 0xfd
      12'h4DE: dout <= 8'b10111111; // 1246 : 191 - 0xbf
      12'h4DF: dout <= 8'b11111111; // 1247 : 255 - 0xff
      12'h4E0: dout <= 8'b10111010; // 1248 : 186 - 0xba -- Sprite 0x9c
      12'h4E1: dout <= 8'b10011100; // 1249 : 156 - 0x9c
      12'h4E2: dout <= 8'b10101010; // 1250 : 170 - 0xaa
      12'h4E3: dout <= 8'b11000000; // 1251 : 192 - 0xc0
      12'h4E4: dout <= 8'b11000000; // 1252 : 192 - 0xc0
      12'h4E5: dout <= 8'b11100000; // 1253 : 224 - 0xe0
      12'h4E6: dout <= 8'b11111000; // 1254 : 248 - 0xf8
      12'h4E7: dout <= 8'b11111111; // 1255 : 255 - 0xff
      12'h4E8: dout <= 8'b00000001; // 1256 :   1 - 0x1 -- Sprite 0x9d
      12'h4E9: dout <= 8'b00000001; // 1257 :   1 - 0x1
      12'h4EA: dout <= 8'b00000001; // 1258 :   1 - 0x1
      12'h4EB: dout <= 8'b00000011; // 1259 :   3 - 0x3
      12'h4EC: dout <= 8'b00000011; // 1260 :   3 - 0x3
      12'h4ED: dout <= 8'b00000111; // 1261 :   7 - 0x7
      12'h4EE: dout <= 8'b00011111; // 1262 :  31 - 0x1f
      12'h4EF: dout <= 8'b11111111; // 1263 : 255 - 0xff
      12'h4F0: dout <= 8'b01111101; // 1264 : 125 - 0x7d -- Sprite 0x9e
      12'h4F1: dout <= 8'b11111111; // 1265 : 255 - 0xff
      12'h4F2: dout <= 8'b11111011; // 1266 : 251 - 0xfb
      12'h4F3: dout <= 8'b11111111; // 1267 : 255 - 0xff
      12'h4F4: dout <= 8'b11111111; // 1268 : 255 - 0xff
      12'h4F5: dout <= 8'b11111011; // 1269 : 251 - 0xfb
      12'h4F6: dout <= 8'b11111111; // 1270 : 255 - 0xff
      12'h4F7: dout <= 8'b01111101; // 1271 : 125 - 0x7d
      12'h4F8: dout <= 8'b11111111; // 1272 : 255 - 0xff -- Sprite 0x9f
      12'h4F9: dout <= 8'b11111111; // 1273 : 255 - 0xff
      12'h4FA: dout <= 8'b10111101; // 1274 : 189 - 0xbd
      12'h4FB: dout <= 8'b11111111; // 1275 : 255 - 0xff
      12'h4FC: dout <= 8'b11111111; // 1276 : 255 - 0xff
      12'h4FD: dout <= 8'b11111111; // 1277 : 255 - 0xff
      12'h4FE: dout <= 8'b11111111; // 1278 : 255 - 0xff
      12'h4FF: dout <= 8'b10111101; // 1279 : 189 - 0xbd
      12'h500: dout <= 8'b11101111; // 1280 : 239 - 0xef -- Sprite 0xa0
      12'h501: dout <= 8'b11000111; // 1281 : 199 - 0xc7
      12'h502: dout <= 8'b10000011; // 1282 : 131 - 0x83
      12'h503: dout <= 8'b00000111; // 1283 :   7 - 0x7
      12'h504: dout <= 8'b10001111; // 1284 : 143 - 0x8f
      12'h505: dout <= 8'b11011101; // 1285 : 221 - 0xdd
      12'h506: dout <= 8'b11111010; // 1286 : 250 - 0xfa
      12'h507: dout <= 8'b11111101; // 1287 : 253 - 0xfd
      12'h508: dout <= 8'b11101111; // 1288 : 239 - 0xef -- Sprite 0xa1
      12'h509: dout <= 8'b11000111; // 1289 : 199 - 0xc7
      12'h50A: dout <= 8'b10000011; // 1290 : 131 - 0x83
      12'h50B: dout <= 8'b00011111; // 1291 :  31 - 0x1f
      12'h50C: dout <= 8'b10010000; // 1292 : 144 - 0x90
      12'h50D: dout <= 8'b11010100; // 1293 : 212 - 0xd4
      12'h50E: dout <= 8'b11110011; // 1294 : 243 - 0xf3
      12'h50F: dout <= 8'b11110010; // 1295 : 242 - 0xf2
      12'h510: dout <= 8'b11101111; // 1296 : 239 - 0xef -- Sprite 0xa2
      12'h511: dout <= 8'b11000111; // 1297 : 199 - 0xc7
      12'h512: dout <= 8'b10000011; // 1298 : 131 - 0x83
      12'h513: dout <= 8'b11111111; // 1299 : 255 - 0xff
      12'h514: dout <= 8'b00000000; // 1300 :   0 - 0x0
      12'h515: dout <= 8'b00000000; // 1301 :   0 - 0x0
      12'h516: dout <= 8'b01010101; // 1302 :  85 - 0x55
      12'h517: dout <= 8'b00000000; // 1303 :   0 - 0x0
      12'h518: dout <= 8'b11110000; // 1304 : 240 - 0xf0 -- Sprite 0xa3
      12'h519: dout <= 8'b11010010; // 1305 : 210 - 0xd2
      12'h51A: dout <= 8'b10010000; // 1306 : 144 - 0x90
      12'h51B: dout <= 8'b00010010; // 1307 :  18 - 0x12
      12'h51C: dout <= 8'b10010000; // 1308 : 144 - 0x90
      12'h51D: dout <= 8'b11010010; // 1309 : 210 - 0xd2
      12'h51E: dout <= 8'b11110000; // 1310 : 240 - 0xf0
      12'h51F: dout <= 8'b11110010; // 1311 : 242 - 0xf2
      12'h520: dout <= 8'b11110000; // 1312 : 240 - 0xf0 -- Sprite 0xa4
      12'h521: dout <= 8'b11010011; // 1313 : 211 - 0xd3
      12'h522: dout <= 8'b10010100; // 1314 : 148 - 0x94
      12'h523: dout <= 8'b00011000; // 1315 :  24 - 0x18
      12'h524: dout <= 8'b10011111; // 1316 : 159 - 0x9f
      12'h525: dout <= 8'b11011101; // 1317 : 221 - 0xdd
      12'h526: dout <= 8'b11111010; // 1318 : 250 - 0xfa
      12'h527: dout <= 8'b11111101; // 1319 : 253 - 0xfd
      12'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0 -- Sprite 0xa5
      12'h529: dout <= 8'b11111111; // 1321 : 255 - 0xff
      12'h52A: dout <= 8'b00000000; // 1322 :   0 - 0x0
      12'h52B: dout <= 8'b00000000; // 1323 :   0 - 0x0
      12'h52C: dout <= 8'b11111111; // 1324 : 255 - 0xff
      12'h52D: dout <= 8'b11011101; // 1325 : 221 - 0xdd
      12'h52E: dout <= 8'b11111010; // 1326 : 250 - 0xfa
      12'h52F: dout <= 8'b11111101; // 1327 : 253 - 0xfd
      12'h530: dout <= 8'b11101111; // 1328 : 239 - 0xef -- Sprite 0xa6
      12'h531: dout <= 8'b11000111; // 1329 : 199 - 0xc7
      12'h532: dout <= 8'b10000011; // 1330 : 131 - 0x83
      12'h533: dout <= 8'b11111111; // 1331 : 255 - 0xff
      12'h534: dout <= 8'b00011111; // 1332 :  31 - 0x1f
      12'h535: dout <= 8'b00101101; // 1333 :  45 - 0x2d
      12'h536: dout <= 8'b01001010; // 1334 :  74 - 0x4a
      12'h537: dout <= 8'b01001101; // 1335 :  77 - 0x4d
      12'h538: dout <= 8'b01001111; // 1336 :  79 - 0x4f -- Sprite 0xa7
      12'h539: dout <= 8'b01001111; // 1337 :  79 - 0x4f
      12'h53A: dout <= 8'b01001011; // 1338 :  75 - 0x4b
      12'h53B: dout <= 8'b01001111; // 1339 :  79 - 0x4f
      12'h53C: dout <= 8'b01001111; // 1340 :  79 - 0x4f
      12'h53D: dout <= 8'b01001101; // 1341 :  77 - 0x4d
      12'h53E: dout <= 8'b01001010; // 1342 :  74 - 0x4a
      12'h53F: dout <= 8'b01001101; // 1343 :  77 - 0x4d
      12'h540: dout <= 8'b01001111; // 1344 :  79 - 0x4f -- Sprite 0xa8
      12'h541: dout <= 8'b11001111; // 1345 : 207 - 0xcf
      12'h542: dout <= 8'b00001011; // 1346 :  11 - 0xb
      12'h543: dout <= 8'b00001111; // 1347 :  15 - 0xf
      12'h544: dout <= 8'b11111111; // 1348 : 255 - 0xff
      12'h545: dout <= 8'b11011101; // 1349 : 221 - 0xdd
      12'h546: dout <= 8'b11111010; // 1350 : 250 - 0xfa
      12'h547: dout <= 8'b11111101; // 1351 : 253 - 0xfd
      12'h548: dout <= 8'b11111111; // 1352 : 255 - 0xff -- Sprite 0xa9
      12'h549: dout <= 8'b11111111; // 1353 : 255 - 0xff
      12'h54A: dout <= 8'b11111111; // 1354 : 255 - 0xff
      12'h54B: dout <= 8'b11111111; // 1355 : 255 - 0xff
      12'h54C: dout <= 8'b11111111; // 1356 : 255 - 0xff
      12'h54D: dout <= 8'b11111111; // 1357 : 255 - 0xff
      12'h54E: dout <= 8'b11111111; // 1358 : 255 - 0xff
      12'h54F: dout <= 8'b11111111; // 1359 : 255 - 0xff
      12'h550: dout <= 8'b11111111; // 1360 : 255 - 0xff -- Sprite 0xaa
      12'h551: dout <= 8'b11111111; // 1361 : 255 - 0xff
      12'h552: dout <= 8'b10101111; // 1362 : 175 - 0xaf
      12'h553: dout <= 8'b01010111; // 1363 :  87 - 0x57
      12'h554: dout <= 8'b10001111; // 1364 : 143 - 0x8f
      12'h555: dout <= 8'b11011101; // 1365 : 221 - 0xdd
      12'h556: dout <= 8'b11111010; // 1366 : 250 - 0xfa
      12'h557: dout <= 8'b11111101; // 1367 : 253 - 0xfd
      12'h558: dout <= 8'b11111111; // 1368 : 255 - 0xff -- Sprite 0xab
      12'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      12'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      12'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      12'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      12'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      12'h560: dout <= 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      12'h561: dout <= 8'b00000000; // 1377 :   0 - 0x0
      12'h562: dout <= 8'b00000000; // 1378 :   0 - 0x0
      12'h563: dout <= 8'b00000000; // 1379 :   0 - 0x0
      12'h564: dout <= 8'b00000000; // 1380 :   0 - 0x0
      12'h565: dout <= 8'b00000000; // 1381 :   0 - 0x0
      12'h566: dout <= 8'b00000000; // 1382 :   0 - 0x0
      12'h567: dout <= 8'b00000000; // 1383 :   0 - 0x0
      12'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0 -- Sprite 0xad
      12'h569: dout <= 8'b11111111; // 1385 : 255 - 0xff
      12'h56A: dout <= 8'b00000000; // 1386 :   0 - 0x0
      12'h56B: dout <= 8'b11111111; // 1387 : 255 - 0xff
      12'h56C: dout <= 8'b11111111; // 1388 : 255 - 0xff
      12'h56D: dout <= 8'b11111111; // 1389 : 255 - 0xff
      12'h56E: dout <= 8'b11111111; // 1390 : 255 - 0xff
      12'h56F: dout <= 8'b11111111; // 1391 : 255 - 0xff
      12'h570: dout <= 8'b11111111; // 1392 : 255 - 0xff -- Sprite 0xae
      12'h571: dout <= 8'b11111111; // 1393 : 255 - 0xff
      12'h572: dout <= 8'b11111111; // 1394 : 255 - 0xff
      12'h573: dout <= 8'b11111111; // 1395 : 255 - 0xff
      12'h574: dout <= 8'b11111111; // 1396 : 255 - 0xff
      12'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      12'h576: dout <= 8'b11111111; // 1398 : 255 - 0xff
      12'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout <= 8'b11111111; // 1400 : 255 - 0xff -- Sprite 0xaf
      12'h579: dout <= 8'b11111111; // 1401 : 255 - 0xff
      12'h57A: dout <= 8'b11111111; // 1402 : 255 - 0xff
      12'h57B: dout <= 8'b11111111; // 1403 : 255 - 0xff
      12'h57C: dout <= 8'b11111111; // 1404 : 255 - 0xff
      12'h57D: dout <= 8'b11111111; // 1405 : 255 - 0xff
      12'h57E: dout <= 8'b11111111; // 1406 : 255 - 0xff
      12'h57F: dout <= 8'b11111111; // 1407 : 255 - 0xff
      12'h580: dout <= 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      12'h581: dout <= 8'b00011111; // 1409 :  31 - 0x1f
      12'h582: dout <= 8'b00010000; // 1410 :  16 - 0x10
      12'h583: dout <= 8'b00010000; // 1411 :  16 - 0x10
      12'h584: dout <= 8'b00010000; // 1412 :  16 - 0x10
      12'h585: dout <= 8'b00010000; // 1413 :  16 - 0x10
      12'h586: dout <= 8'b00010000; // 1414 :  16 - 0x10
      12'h587: dout <= 8'b00010000; // 1415 :  16 - 0x10
      12'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0 -- Sprite 0xb1
      12'h589: dout <= 8'b11111000; // 1417 : 248 - 0xf8
      12'h58A: dout <= 8'b00001000; // 1418 :   8 - 0x8
      12'h58B: dout <= 8'b00001000; // 1419 :   8 - 0x8
      12'h58C: dout <= 8'b00001000; // 1420 :   8 - 0x8
      12'h58D: dout <= 8'b00001000; // 1421 :   8 - 0x8
      12'h58E: dout <= 8'b00001000; // 1422 :   8 - 0x8
      12'h58F: dout <= 8'b00001000; // 1423 :   8 - 0x8
      12'h590: dout <= 8'b00010000; // 1424 :  16 - 0x10 -- Sprite 0xb2
      12'h591: dout <= 8'b00010000; // 1425 :  16 - 0x10
      12'h592: dout <= 8'b00010000; // 1426 :  16 - 0x10
      12'h593: dout <= 8'b00010000; // 1427 :  16 - 0x10
      12'h594: dout <= 8'b00011111; // 1428 :  31 - 0x1f
      12'h595: dout <= 8'b00011111; // 1429 :  31 - 0x1f
      12'h596: dout <= 8'b00001111; // 1430 :  15 - 0xf
      12'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      12'h598: dout <= 8'b00001000; // 1432 :   8 - 0x8 -- Sprite 0xb3
      12'h599: dout <= 8'b00001000; // 1433 :   8 - 0x8
      12'h59A: dout <= 8'b00001000; // 1434 :   8 - 0x8
      12'h59B: dout <= 8'b00001000; // 1435 :   8 - 0x8
      12'h59C: dout <= 8'b11111000; // 1436 : 248 - 0xf8
      12'h59D: dout <= 8'b11111000; // 1437 : 248 - 0xf8
      12'h59E: dout <= 8'b11110000; // 1438 : 240 - 0xf0
      12'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout <= 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0xb4
      12'h5A1: dout <= 8'b00000000; // 1441 :   0 - 0x0
      12'h5A2: dout <= 8'b00111111; // 1442 :  63 - 0x3f
      12'h5A3: dout <= 8'b01100000; // 1443 :  96 - 0x60
      12'h5A4: dout <= 8'b01100000; // 1444 :  96 - 0x60
      12'h5A5: dout <= 8'b01100000; // 1445 :  96 - 0x60
      12'h5A6: dout <= 8'b01100000; // 1446 :  96 - 0x60
      12'h5A7: dout <= 8'b01100000; // 1447 :  96 - 0x60
      12'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0 -- Sprite 0xb5
      12'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      12'h5AA: dout <= 8'b11111100; // 1450 : 252 - 0xfc
      12'h5AB: dout <= 8'b00000110; // 1451 :   6 - 0x6
      12'h5AC: dout <= 8'b00000110; // 1452 :   6 - 0x6
      12'h5AD: dout <= 8'b00000110; // 1453 :   6 - 0x6
      12'h5AE: dout <= 8'b00000110; // 1454 :   6 - 0x6
      12'h5AF: dout <= 8'b00000110; // 1455 :   6 - 0x6
      12'h5B0: dout <= 8'b01100000; // 1456 :  96 - 0x60 -- Sprite 0xb6
      12'h5B1: dout <= 8'b01100000; // 1457 :  96 - 0x60
      12'h5B2: dout <= 8'b01100000; // 1458 :  96 - 0x60
      12'h5B3: dout <= 8'b01111111; // 1459 : 127 - 0x7f
      12'h5B4: dout <= 8'b01111111; // 1460 : 127 - 0x7f
      12'h5B5: dout <= 8'b00111111; // 1461 :  63 - 0x3f
      12'h5B6: dout <= 8'b00000000; // 1462 :   0 - 0x0
      12'h5B7: dout <= 8'b00000000; // 1463 :   0 - 0x0
      12'h5B8: dout <= 8'b00000110; // 1464 :   6 - 0x6 -- Sprite 0xb7
      12'h5B9: dout <= 8'b00000110; // 1465 :   6 - 0x6
      12'h5BA: dout <= 8'b00000110; // 1466 :   6 - 0x6
      12'h5BB: dout <= 8'b11111110; // 1467 : 254 - 0xfe
      12'h5BC: dout <= 8'b11111110; // 1468 : 254 - 0xfe
      12'h5BD: dout <= 8'b11111100; // 1469 : 252 - 0xfc
      12'h5BE: dout <= 8'b00000000; // 1470 :   0 - 0x0
      12'h5BF: dout <= 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout <= 8'b01100000; // 1472 :  96 - 0x60 -- Sprite 0xb8
      12'h5C1: dout <= 8'b11110011; // 1473 : 243 - 0xf3
      12'h5C2: dout <= 8'b11000111; // 1474 : 199 - 0xc7
      12'h5C3: dout <= 8'b10000110; // 1475 : 134 - 0x86
      12'h5C4: dout <= 8'b00000100; // 1476 :   4 - 0x4
      12'h5C5: dout <= 8'b00000100; // 1477 :   4 - 0x4
      12'h5C6: dout <= 8'b00000111; // 1478 :   7 - 0x7
      12'h5C7: dout <= 8'b00000111; // 1479 :   7 - 0x7
      12'h5C8: dout <= 8'b00000110; // 1480 :   6 - 0x6 -- Sprite 0xb9
      12'h5C9: dout <= 8'b10001111; // 1481 : 143 - 0x8f
      12'h5CA: dout <= 8'b11000101; // 1482 : 197 - 0xc5
      12'h5CB: dout <= 8'b00100011; // 1483 :  35 - 0x23
      12'h5CC: dout <= 8'b00101110; // 1484 :  46 - 0x2e
      12'h5CD: dout <= 8'b01100000; // 1485 :  96 - 0x60
      12'h5CE: dout <= 8'b11100001; // 1486 : 225 - 0xe1
      12'h5CF: dout <= 8'b11100001; // 1487 : 225 - 0xe1
      12'h5D0: dout <= 8'b11001000; // 1488 : 200 - 0xc8 -- Sprite 0xba
      12'h5D1: dout <= 8'b11111000; // 1489 : 248 - 0xf8
      12'h5D2: dout <= 8'b10110000; // 1490 : 176 - 0xb0
      12'h5D3: dout <= 8'b00010000; // 1491 :  16 - 0x10
      12'h5D4: dout <= 8'b00110000; // 1492 :  48 - 0x30
      12'h5D5: dout <= 8'b11001000; // 1493 : 200 - 0xc8
      12'h5D6: dout <= 8'b11111000; // 1494 : 248 - 0xf8
      12'h5D7: dout <= 8'b10000000; // 1495 : 128 - 0x80
      12'h5D8: dout <= 8'b00000011; // 1496 :   3 - 0x3 -- Sprite 0xbb
      12'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      12'h5DB: dout <= 8'b01100000; // 1499 :  96 - 0x60
      12'h5DC: dout <= 8'b11110000; // 1500 : 240 - 0xf0
      12'h5DD: dout <= 8'b11010000; // 1501 : 208 - 0xd0
      12'h5DE: dout <= 8'b10010000; // 1502 : 144 - 0x90
      12'h5DF: dout <= 8'b01100000; // 1503 :  96 - 0x60
      12'h5E0: dout <= 8'b11000011; // 1504 : 195 - 0xc3 -- Sprite 0xbc
      12'h5E1: dout <= 8'b00001110; // 1505 :  14 - 0xe
      12'h5E2: dout <= 8'b00000000; // 1506 :   0 - 0x0
      12'h5E3: dout <= 8'b00000110; // 1507 :   6 - 0x6
      12'h5E4: dout <= 8'b00001111; // 1508 :  15 - 0xf
      12'h5E5: dout <= 8'b00001101; // 1509 :  13 - 0xd
      12'h5E6: dout <= 8'b00001001; // 1510 :   9 - 0x9
      12'h5E7: dout <= 8'b00000110; // 1511 :   6 - 0x6
      12'h5E8: dout <= 8'b11100000; // 1512 : 224 - 0xe0 -- Sprite 0xbd
      12'h5E9: dout <= 8'b01100011; // 1513 :  99 - 0x63
      12'h5EA: dout <= 8'b11100111; // 1514 : 231 - 0xe7
      12'h5EB: dout <= 8'b11100110; // 1515 : 230 - 0xe6
      12'h5EC: dout <= 8'b00000100; // 1516 :   4 - 0x4
      12'h5ED: dout <= 8'b00000100; // 1517 :   4 - 0x4
      12'h5EE: dout <= 8'b00000111; // 1518 :   7 - 0x7
      12'h5EF: dout <= 8'b00000111; // 1519 :   7 - 0x7
      12'h5F0: dout <= 8'b00000111; // 1520 :   7 - 0x7 -- Sprite 0xbe
      12'h5F1: dout <= 8'b10000011; // 1521 : 131 - 0x83
      12'h5F2: dout <= 8'b11000111; // 1522 : 199 - 0xc7
      12'h5F3: dout <= 8'b00100111; // 1523 :  39 - 0x27
      12'h5F4: dout <= 8'b00100000; // 1524 :  32 - 0x20
      12'h5F5: dout <= 8'b01100000; // 1525 :  96 - 0x60
      12'h5F6: dout <= 8'b11100000; // 1526 : 224 - 0xe0
      12'h5F7: dout <= 8'b11100000; // 1527 : 224 - 0xe0
      12'h5F8: dout <= 8'b00000011; // 1528 :   3 - 0x3 -- Sprite 0xbf
      12'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout <= 8'b00001100; // 1530 :  12 - 0xc
      12'h5FB: dout <= 8'b00001100; // 1531 :  12 - 0xc
      12'h5FC: dout <= 8'b11100100; // 1532 : 228 - 0xe4
      12'h5FD: dout <= 8'b01101100; // 1533 : 108 - 0x6c
      12'h5FE: dout <= 8'b11101101; // 1534 : 237 - 0xed
      12'h5FF: dout <= 8'b11100111; // 1535 : 231 - 0xe7
      12'h600: dout <= 8'b11000000; // 1536 : 192 - 0xc0 -- Sprite 0xc0
      12'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout <= 8'b00110000; // 1538 :  48 - 0x30
      12'h603: dout <= 8'b00110000; // 1539 :  48 - 0x30
      12'h604: dout <= 8'b00010111; // 1540 :  23 - 0x17
      12'h605: dout <= 8'b00110011; // 1541 :  51 - 0x33
      12'h606: dout <= 8'b01110111; // 1542 : 119 - 0x77
      12'h607: dout <= 8'b11010111; // 1543 : 215 - 0xd7
      12'h608: dout <= 8'b00001100; // 1544 :  12 - 0xc -- Sprite 0xc1
      12'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      12'h60A: dout <= 8'b00000000; // 1546 :   0 - 0x0
      12'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      12'h60C: dout <= 8'b00000000; // 1548 :   0 - 0x0
      12'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      12'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      12'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout <= 8'b00110000; // 1552 :  48 - 0x30 -- Sprite 0xc2
      12'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      12'h612: dout <= 8'b00000000; // 1554 :   0 - 0x0
      12'h613: dout <= 8'b00000000; // 1555 :   0 - 0x0
      12'h614: dout <= 8'b00000000; // 1556 :   0 - 0x0
      12'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      12'h616: dout <= 8'b00000000; // 1558 :   0 - 0x0
      12'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      12'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0 -- Sprite 0xc3
      12'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      12'h61A: dout <= 8'b00000100; // 1562 :   4 - 0x4
      12'h61B: dout <= 8'b00001101; // 1563 :  13 - 0xd
      12'h61C: dout <= 8'b00001111; // 1564 :  15 - 0xf
      12'h61D: dout <= 8'b00001100; // 1565 :  12 - 0xc
      12'h61E: dout <= 8'b00001100; // 1566 :  12 - 0xc
      12'h61F: dout <= 8'b00000100; // 1567 :   4 - 0x4
      12'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      12'h621: dout <= 8'b00000000; // 1569 :   0 - 0x0
      12'h622: dout <= 8'b00010000; // 1570 :  16 - 0x10
      12'h623: dout <= 8'b01110000; // 1571 : 112 - 0x70
      12'h624: dout <= 8'b11110000; // 1572 : 240 - 0xf0
      12'h625: dout <= 8'b00110000; // 1573 :  48 - 0x30
      12'h626: dout <= 8'b00110000; // 1574 :  48 - 0x30
      12'h627: dout <= 8'b00010000; // 1575 :  16 - 0x10
      12'h628: dout <= 8'b11100100; // 1576 : 228 - 0xe4 -- Sprite 0xc5
      12'h629: dout <= 8'b00100100; // 1577 :  36 - 0x24
      12'h62A: dout <= 8'b11101111; // 1578 : 239 - 0xef
      12'h62B: dout <= 8'b11100111; // 1579 : 231 - 0xe7
      12'h62C: dout <= 8'b00000110; // 1580 :   6 - 0x6
      12'h62D: dout <= 8'b00000100; // 1581 :   4 - 0x4
      12'h62E: dout <= 8'b00000100; // 1582 :   4 - 0x4
      12'h62F: dout <= 8'b00000111; // 1583 :   7 - 0x7
      12'h630: dout <= 8'b00010111; // 1584 :  23 - 0x17 -- Sprite 0xc6
      12'h631: dout <= 8'b00010001; // 1585 :  17 - 0x11
      12'h632: dout <= 8'b10110111; // 1586 : 183 - 0xb7
      12'h633: dout <= 8'b11000111; // 1587 : 199 - 0xc7
      12'h634: dout <= 8'b00100000; // 1588 :  32 - 0x20
      12'h635: dout <= 8'b00100000; // 1589 :  32 - 0x20
      12'h636: dout <= 8'b01100000; // 1590 :  96 - 0x60
      12'h637: dout <= 8'b11100000; // 1591 : 224 - 0xe0
      12'h638: dout <= 8'b00000111; // 1592 :   7 - 0x7 -- Sprite 0xc7
      12'h639: dout <= 8'b00000011; // 1593 :   3 - 0x3
      12'h63A: dout <= 8'b00000000; // 1594 :   0 - 0x0
      12'h63B: dout <= 8'b00000000; // 1595 :   0 - 0x0
      12'h63C: dout <= 8'b11100000; // 1596 : 224 - 0xe0
      12'h63D: dout <= 8'b00100000; // 1597 :  32 - 0x20
      12'h63E: dout <= 8'b11100000; // 1598 : 224 - 0xe0
      12'h63F: dout <= 8'b11100000; // 1599 : 224 - 0xe0
      12'h640: dout <= 8'b11100000; // 1600 : 224 - 0xe0 -- Sprite 0xc8
      12'h641: dout <= 8'b11000000; // 1601 : 192 - 0xc0
      12'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      12'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      12'h644: dout <= 8'b00000111; // 1604 :   7 - 0x7
      12'h645: dout <= 8'b00000001; // 1605 :   1 - 0x1
      12'h646: dout <= 8'b00000111; // 1606 :   7 - 0x7
      12'h647: dout <= 8'b00000111; // 1607 :   7 - 0x7
      12'h648: dout <= 8'b00010011; // 1608 :  19 - 0x13 -- Sprite 0xc9
      12'h649: dout <= 8'b00011111; // 1609 :  31 - 0x1f
      12'h64A: dout <= 8'b00001101; // 1610 :  13 - 0xd
      12'h64B: dout <= 8'b00000100; // 1611 :   4 - 0x4
      12'h64C: dout <= 8'b00001100; // 1612 :  12 - 0xc
      12'h64D: dout <= 8'b00010011; // 1613 :  19 - 0x13
      12'h64E: dout <= 8'b00011111; // 1614 :  31 - 0x1f
      12'h64F: dout <= 8'b00000001; // 1615 :   1 - 0x1
      12'h650: dout <= 8'b01100000; // 1616 :  96 - 0x60 -- Sprite 0xca
      12'h651: dout <= 8'b11110011; // 1617 : 243 - 0xf3
      12'h652: dout <= 8'b10100111; // 1618 : 167 - 0xa7
      12'h653: dout <= 8'b11000110; // 1619 : 198 - 0xc6
      12'h654: dout <= 8'b01110100; // 1620 : 116 - 0x74
      12'h655: dout <= 8'b00000100; // 1621 :   4 - 0x4
      12'h656: dout <= 8'b10000111; // 1622 : 135 - 0x87
      12'h657: dout <= 8'b10000111; // 1623 : 135 - 0x87
      12'h658: dout <= 8'b00000110; // 1624 :   6 - 0x6 -- Sprite 0xcb
      12'h659: dout <= 8'b10001111; // 1625 : 143 - 0x8f
      12'h65A: dout <= 8'b11000011; // 1626 : 195 - 0xc3
      12'h65B: dout <= 8'b00100001; // 1627 :  33 - 0x21
      12'h65C: dout <= 8'b00100000; // 1628 :  32 - 0x20
      12'h65D: dout <= 8'b01100000; // 1629 :  96 - 0x60
      12'h65E: dout <= 8'b11100000; // 1630 : 224 - 0xe0
      12'h65F: dout <= 8'b11100000; // 1631 : 224 - 0xe0
      12'h660: dout <= 8'b11000011; // 1632 : 195 - 0xc3 -- Sprite 0xcc
      12'h661: dout <= 8'b01110000; // 1633 : 112 - 0x70
      12'h662: dout <= 8'b00000000; // 1634 :   0 - 0x0
      12'h663: dout <= 8'b01100000; // 1635 :  96 - 0x60
      12'h664: dout <= 8'b11110000; // 1636 : 240 - 0xf0
      12'h665: dout <= 8'b11010000; // 1637 : 208 - 0xd0
      12'h666: dout <= 8'b10010000; // 1638 : 144 - 0x90
      12'h667: dout <= 8'b01100000; // 1639 :  96 - 0x60
      12'h668: dout <= 8'b11000000; // 1640 : 192 - 0xc0 -- Sprite 0xcd
      12'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout <= 8'b00000110; // 1643 :   6 - 0x6
      12'h66C: dout <= 8'b00001111; // 1644 :  15 - 0xf
      12'h66D: dout <= 8'b00001101; // 1645 :  13 - 0xd
      12'h66E: dout <= 8'b00001001; // 1646 :   9 - 0x9
      12'h66F: dout <= 8'b00000110; // 1647 :   6 - 0x6
      12'h670: dout <= 8'b11111100; // 1648 : 252 - 0xfc -- Sprite 0xce
      12'h671: dout <= 8'b11000000; // 1649 : 192 - 0xc0
      12'h672: dout <= 8'b11010001; // 1650 : 209 - 0xd1
      12'h673: dout <= 8'b11000010; // 1651 : 194 - 0xc2
      12'h674: dout <= 8'b10011110; // 1652 : 158 - 0x9e
      12'h675: dout <= 8'b10111111; // 1653 : 191 - 0xbf
      12'h676: dout <= 8'b10110000; // 1654 : 176 - 0xb0
      12'h677: dout <= 8'b10110011; // 1655 : 179 - 0xb3
      12'h678: dout <= 8'b00000111; // 1656 :   7 - 0x7 -- Sprite 0xcf
      12'h679: dout <= 8'b11110011; // 1657 : 243 - 0xf3
      12'h67A: dout <= 8'b00001011; // 1658 :  11 - 0xb
      12'h67B: dout <= 8'b01111011; // 1659 : 123 - 0x7b
      12'h67C: dout <= 8'b01111011; // 1660 : 123 - 0x7b
      12'h67D: dout <= 8'b11111001; // 1661 : 249 - 0xf9
      12'h67E: dout <= 8'b00001101; // 1662 :  13 - 0xd
      12'h67F: dout <= 8'b11101101; // 1663 : 237 - 0xed
      12'h680: dout <= 8'b11111111; // 1664 : 255 - 0xff -- Sprite 0xd0
      12'h681: dout <= 8'b11111111; // 1665 : 255 - 0xff
      12'h682: dout <= 8'b11111111; // 1666 : 255 - 0xff
      12'h683: dout <= 8'b11111111; // 1667 : 255 - 0xff
      12'h684: dout <= 8'b11101110; // 1668 : 238 - 0xee
      12'h685: dout <= 8'b11101110; // 1669 : 238 - 0xee
      12'h686: dout <= 8'b11101110; // 1670 : 238 - 0xee
      12'h687: dout <= 8'b11101110; // 1671 : 238 - 0xee
      12'h688: dout <= 8'b11111111; // 1672 : 255 - 0xff -- Sprite 0xd1
      12'h689: dout <= 8'b11111111; // 1673 : 255 - 0xff
      12'h68A: dout <= 8'b11111111; // 1674 : 255 - 0xff
      12'h68B: dout <= 8'b11111011; // 1675 : 251 - 0xfb
      12'h68C: dout <= 8'b11111011; // 1676 : 251 - 0xfb
      12'h68D: dout <= 8'b11111011; // 1677 : 251 - 0xfb
      12'h68E: dout <= 8'b11111011; // 1678 : 251 - 0xfb
      12'h68F: dout <= 8'b11111011; // 1679 : 251 - 0xfb
      12'h690: dout <= 8'b11111111; // 1680 : 255 - 0xff -- Sprite 0xd2
      12'h691: dout <= 8'b11111111; // 1681 : 255 - 0xff
      12'h692: dout <= 8'b11111111; // 1682 : 255 - 0xff
      12'h693: dout <= 8'b11111111; // 1683 : 255 - 0xff
      12'h694: dout <= 8'b11101110; // 1684 : 238 - 0xee
      12'h695: dout <= 8'b10001110; // 1685 : 142 - 0x8e
      12'h696: dout <= 8'b11111110; // 1686 : 254 - 0xfe
      12'h697: dout <= 8'b11111110; // 1687 : 254 - 0xfe
      12'h698: dout <= 8'b11111111; // 1688 : 255 - 0xff -- Sprite 0xd3
      12'h699: dout <= 8'b11111111; // 1689 : 255 - 0xff
      12'h69A: dout <= 8'b11111111; // 1690 : 255 - 0xff
      12'h69B: dout <= 8'b11111111; // 1691 : 255 - 0xff
      12'h69C: dout <= 8'b11101110; // 1692 : 238 - 0xee
      12'h69D: dout <= 8'b10001110; // 1693 : 142 - 0x8e
      12'h69E: dout <= 8'b11111100; // 1694 : 252 - 0xfc
      12'h69F: dout <= 8'b11111101; // 1695 : 253 - 0xfd
      12'h6A0: dout <= 8'b11111111; // 1696 : 255 - 0xff -- Sprite 0xd4
      12'h6A1: dout <= 8'b11111111; // 1697 : 255 - 0xff
      12'h6A2: dout <= 8'b11111111; // 1698 : 255 - 0xff
      12'h6A3: dout <= 8'b11111110; // 1699 : 254 - 0xfe
      12'h6A4: dout <= 8'b11101110; // 1700 : 238 - 0xee
      12'h6A5: dout <= 8'b11101110; // 1701 : 238 - 0xee
      12'h6A6: dout <= 8'b11101110; // 1702 : 238 - 0xee
      12'h6A7: dout <= 8'b11101110; // 1703 : 238 - 0xee
      12'h6A8: dout <= 8'b11111111; // 1704 : 255 - 0xff -- Sprite 0xd5
      12'h6A9: dout <= 8'b11111111; // 1705 : 255 - 0xff
      12'h6AA: dout <= 8'b11111111; // 1706 : 255 - 0xff
      12'h6AB: dout <= 8'b11111101; // 1707 : 253 - 0xfd
      12'h6AC: dout <= 8'b11100001; // 1708 : 225 - 0xe1
      12'h6AD: dout <= 8'b11101111; // 1709 : 239 - 0xef
      12'h6AE: dout <= 8'b11111111; // 1710 : 255 - 0xff
      12'h6AF: dout <= 8'b11111111; // 1711 : 255 - 0xff
      12'h6B0: dout <= 8'b11111111; // 1712 : 255 - 0xff -- Sprite 0xd6
      12'h6B1: dout <= 8'b11111111; // 1713 : 255 - 0xff
      12'h6B2: dout <= 8'b11111111; // 1714 : 255 - 0xff
      12'h6B3: dout <= 8'b11111101; // 1715 : 253 - 0xfd
      12'h6B4: dout <= 8'b11100001; // 1716 : 225 - 0xe1
      12'h6B5: dout <= 8'b11101111; // 1717 : 239 - 0xef
      12'h6B6: dout <= 8'b11111111; // 1718 : 255 - 0xff
      12'h6B7: dout <= 8'b11111111; // 1719 : 255 - 0xff
      12'h6B8: dout <= 8'b11111111; // 1720 : 255 - 0xff -- Sprite 0xd7
      12'h6B9: dout <= 8'b11111111; // 1721 : 255 - 0xff
      12'h6BA: dout <= 8'b11111111; // 1722 : 255 - 0xff
      12'h6BB: dout <= 8'b11111110; // 1723 : 254 - 0xfe
      12'h6BC: dout <= 8'b11101110; // 1724 : 238 - 0xee
      12'h6BD: dout <= 8'b10001110; // 1725 : 142 - 0x8e
      12'h6BE: dout <= 8'b11111110; // 1726 : 254 - 0xfe
      12'h6BF: dout <= 8'b11111100; // 1727 : 252 - 0xfc
      12'h6C0: dout <= 8'b11111111; // 1728 : 255 - 0xff -- Sprite 0xd8
      12'h6C1: dout <= 8'b11111111; // 1729 : 255 - 0xff
      12'h6C2: dout <= 8'b11111111; // 1730 : 255 - 0xff
      12'h6C3: dout <= 8'b11111111; // 1731 : 255 - 0xff
      12'h6C4: dout <= 8'b11101110; // 1732 : 238 - 0xee
      12'h6C5: dout <= 8'b11101110; // 1733 : 238 - 0xee
      12'h6C6: dout <= 8'b11111100; // 1734 : 252 - 0xfc
      12'h6C7: dout <= 8'b11111111; // 1735 : 255 - 0xff
      12'h6C8: dout <= 8'b11111111; // 1736 : 255 - 0xff -- Sprite 0xd9
      12'h6C9: dout <= 8'b11111111; // 1737 : 255 - 0xff
      12'h6CA: dout <= 8'b11111111; // 1738 : 255 - 0xff
      12'h6CB: dout <= 8'b11111111; // 1739 : 255 - 0xff
      12'h6CC: dout <= 8'b11101110; // 1740 : 238 - 0xee
      12'h6CD: dout <= 8'b11101110; // 1741 : 238 - 0xee
      12'h6CE: dout <= 8'b11101110; // 1742 : 238 - 0xee
      12'h6CF: dout <= 8'b11101110; // 1743 : 238 - 0xee
      12'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0xda
      12'h6D1: dout <= 8'b00000000; // 1745 :   0 - 0x0
      12'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      12'h6D3: dout <= 8'b10000000; // 1747 : 128 - 0x80
      12'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      12'h6D5: dout <= 8'b00000000; // 1749 :   0 - 0x0
      12'h6D6: dout <= 8'b00000100; // 1750 :   4 - 0x4
      12'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      12'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0 -- Sprite 0xdb
      12'h6D9: dout <= 8'b00000100; // 1753 :   4 - 0x4
      12'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      12'h6DB: dout <= 8'b00010001; // 1755 :  17 - 0x11
      12'h6DC: dout <= 8'b00000000; // 1756 :   0 - 0x0
      12'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      12'h6DE: dout <= 8'b00000000; // 1758 :   0 - 0x0
      12'h6DF: dout <= 8'b00100000; // 1759 :  32 - 0x20
      12'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0xdc
      12'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout <= 8'b00100000; // 1763 :  32 - 0x20
      12'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      12'h6E5: dout <= 8'b00000000; // 1765 :   0 - 0x0
      12'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      12'h6E7: dout <= 8'b00000100; // 1767 :   4 - 0x4
      12'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- Sprite 0xdd
      12'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      12'h6EA: dout <= 8'b00010001; // 1770 :  17 - 0x11
      12'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      12'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      12'h6ED: dout <= 8'b10000000; // 1773 : 128 - 0x80
      12'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      12'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      12'h6F0: dout <= 8'b10110011; // 1776 : 179 - 0xb3 -- Sprite 0xde
      12'h6F1: dout <= 8'b10110011; // 1777 : 179 - 0xb3
      12'h6F2: dout <= 8'b10110011; // 1778 : 179 - 0xb3
      12'h6F3: dout <= 8'b10110011; // 1779 : 179 - 0xb3
      12'h6F4: dout <= 8'b10110000; // 1780 : 176 - 0xb0
      12'h6F5: dout <= 8'b10101111; // 1781 : 175 - 0xaf
      12'h6F6: dout <= 8'b10011111; // 1782 : 159 - 0x9f
      12'h6F7: dout <= 8'b11000000; // 1783 : 192 - 0xc0
      12'h6F8: dout <= 8'b11101101; // 1784 : 237 - 0xed -- Sprite 0xdf
      12'h6F9: dout <= 8'b11001101; // 1785 : 205 - 0xcd
      12'h6FA: dout <= 8'b11001101; // 1786 : 205 - 0xcd
      12'h6FB: dout <= 8'b00001101; // 1787 :  13 - 0xd
      12'h6FC: dout <= 8'b00001101; // 1788 :  13 - 0xd
      12'h6FD: dout <= 8'b11111101; // 1789 : 253 - 0xfd
      12'h6FE: dout <= 8'b11111101; // 1790 : 253 - 0xfd
      12'h6FF: dout <= 8'b00000011; // 1791 :   3 - 0x3
      12'h700: dout <= 8'b11101110; // 1792 : 238 - 0xee -- Sprite 0xe0
      12'h701: dout <= 8'b11101110; // 1793 : 238 - 0xee
      12'h702: dout <= 8'b11101110; // 1794 : 238 - 0xee
      12'h703: dout <= 8'b11101110; // 1795 : 238 - 0xee
      12'h704: dout <= 8'b11111110; // 1796 : 254 - 0xfe
      12'h705: dout <= 8'b11111100; // 1797 : 252 - 0xfc
      12'h706: dout <= 8'b11000001; // 1798 : 193 - 0xc1
      12'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      12'h708: dout <= 8'b11111011; // 1800 : 251 - 0xfb -- Sprite 0xe1
      12'h709: dout <= 8'b11111011; // 1801 : 251 - 0xfb
      12'h70A: dout <= 8'b11111011; // 1802 : 251 - 0xfb
      12'h70B: dout <= 8'b11111011; // 1803 : 251 - 0xfb
      12'h70C: dout <= 8'b11111111; // 1804 : 255 - 0xff
      12'h70D: dout <= 8'b11111101; // 1805 : 253 - 0xfd
      12'h70E: dout <= 8'b11000001; // 1806 : 193 - 0xc1
      12'h70F: dout <= 8'b11111111; // 1807 : 255 - 0xff
      12'h710: dout <= 8'b11111100; // 1808 : 252 - 0xfc -- Sprite 0xe2
      12'h711: dout <= 8'b11100001; // 1809 : 225 - 0xe1
      12'h712: dout <= 8'b11101111; // 1810 : 239 - 0xef
      12'h713: dout <= 8'b11101111; // 1811 : 239 - 0xef
      12'h714: dout <= 8'b11111111; // 1812 : 255 - 0xff
      12'h715: dout <= 8'b11111110; // 1813 : 254 - 0xfe
      12'h716: dout <= 8'b10000000; // 1814 : 128 - 0x80
      12'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      12'h718: dout <= 8'b11101110; // 1816 : 238 - 0xee -- Sprite 0xe3
      12'h719: dout <= 8'b11111110; // 1817 : 254 - 0xfe
      12'h71A: dout <= 8'b11111110; // 1818 : 254 - 0xfe
      12'h71B: dout <= 8'b11111110; // 1819 : 254 - 0xfe
      12'h71C: dout <= 8'b11111110; // 1820 : 254 - 0xfe
      12'h71D: dout <= 8'b11111100; // 1821 : 252 - 0xfc
      12'h71E: dout <= 8'b11000001; // 1822 : 193 - 0xc1
      12'h71F: dout <= 8'b11111111; // 1823 : 255 - 0xff
      12'h720: dout <= 8'b11101110; // 1824 : 238 - 0xee -- Sprite 0xe4
      12'h721: dout <= 8'b11101110; // 1825 : 238 - 0xee
      12'h722: dout <= 8'b11111110; // 1826 : 254 - 0xfe
      12'h723: dout <= 8'b11111110; // 1827 : 254 - 0xfe
      12'h724: dout <= 8'b10001110; // 1828 : 142 - 0x8e
      12'h725: dout <= 8'b11111110; // 1829 : 254 - 0xfe
      12'h726: dout <= 8'b11111000; // 1830 : 248 - 0xf8
      12'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      12'h728: dout <= 8'b10001110; // 1832 : 142 - 0x8e -- Sprite 0xe5
      12'h729: dout <= 8'b11111110; // 1833 : 254 - 0xfe
      12'h72A: dout <= 8'b11111110; // 1834 : 254 - 0xfe
      12'h72B: dout <= 8'b11111110; // 1835 : 254 - 0xfe
      12'h72C: dout <= 8'b11111110; // 1836 : 254 - 0xfe
      12'h72D: dout <= 8'b11111100; // 1837 : 252 - 0xfc
      12'h72E: dout <= 8'b11000001; // 1838 : 193 - 0xc1
      12'h72F: dout <= 8'b11111111; // 1839 : 255 - 0xff
      12'h730: dout <= 8'b11101110; // 1840 : 238 - 0xee -- Sprite 0xe6
      12'h731: dout <= 8'b11101110; // 1841 : 238 - 0xee
      12'h732: dout <= 8'b11101110; // 1842 : 238 - 0xee
      12'h733: dout <= 8'b11101110; // 1843 : 238 - 0xee
      12'h734: dout <= 8'b11111110; // 1844 : 254 - 0xfe
      12'h735: dout <= 8'b11111100; // 1845 : 252 - 0xfc
      12'h736: dout <= 8'b11000001; // 1846 : 193 - 0xc1
      12'h737: dout <= 8'b11111111; // 1847 : 255 - 0xff
      12'h738: dout <= 8'b11111101; // 1848 : 253 - 0xfd -- Sprite 0xe7
      12'h739: dout <= 8'b11111101; // 1849 : 253 - 0xfd
      12'h73A: dout <= 8'b11111001; // 1850 : 249 - 0xf9
      12'h73B: dout <= 8'b11111011; // 1851 : 251 - 0xfb
      12'h73C: dout <= 8'b11111011; // 1852 : 251 - 0xfb
      12'h73D: dout <= 8'b11111011; // 1853 : 251 - 0xfb
      12'h73E: dout <= 8'b11100011; // 1854 : 227 - 0xe3
      12'h73F: dout <= 8'b11111111; // 1855 : 255 - 0xff
      12'h740: dout <= 8'b11101110; // 1856 : 238 - 0xee -- Sprite 0xe8
      12'h741: dout <= 8'b11101110; // 1857 : 238 - 0xee
      12'h742: dout <= 8'b11101110; // 1858 : 238 - 0xee
      12'h743: dout <= 8'b11101110; // 1859 : 238 - 0xee
      12'h744: dout <= 8'b11111110; // 1860 : 254 - 0xfe
      12'h745: dout <= 8'b11111100; // 1861 : 252 - 0xfc
      12'h746: dout <= 8'b11000001; // 1862 : 193 - 0xc1
      12'h747: dout <= 8'b11111111; // 1863 : 255 - 0xff
      12'h748: dout <= 8'b11111110; // 1864 : 254 - 0xfe -- Sprite 0xe9
      12'h749: dout <= 8'b11111110; // 1865 : 254 - 0xfe
      12'h74A: dout <= 8'b11001110; // 1866 : 206 - 0xce
      12'h74B: dout <= 8'b11111110; // 1867 : 254 - 0xfe
      12'h74C: dout <= 8'b11111110; // 1868 : 254 - 0xfe
      12'h74D: dout <= 8'b11111100; // 1869 : 252 - 0xfc
      12'h74E: dout <= 8'b11000001; // 1870 : 193 - 0xc1
      12'h74F: dout <= 8'b11111111; // 1871 : 255 - 0xff
      12'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0xea
      12'h751: dout <= 8'b01110000; // 1873 : 112 - 0x70
      12'h752: dout <= 8'b00111000; // 1874 :  56 - 0x38
      12'h753: dout <= 8'b00000000; // 1875 :   0 - 0x0
      12'h754: dout <= 8'b00000010; // 1876 :   2 - 0x2
      12'h755: dout <= 8'b00000111; // 1877 :   7 - 0x7
      12'h756: dout <= 8'b00000011; // 1878 :   3 - 0x3
      12'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout <= 8'b00000000; // 1880 :   0 - 0x0 -- Sprite 0xeb
      12'h759: dout <= 8'b00001100; // 1881 :  12 - 0xc
      12'h75A: dout <= 8'b00000110; // 1882 :   6 - 0x6
      12'h75B: dout <= 8'b00000110; // 1883 :   6 - 0x6
      12'h75C: dout <= 8'b01100000; // 1884 :  96 - 0x60
      12'h75D: dout <= 8'b01110000; // 1885 : 112 - 0x70
      12'h75E: dout <= 8'b00110000; // 1886 :  48 - 0x30
      12'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      12'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      12'h761: dout <= 8'b11000000; // 1889 : 192 - 0xc0
      12'h762: dout <= 8'b11100000; // 1890 : 224 - 0xe0
      12'h763: dout <= 8'b01100000; // 1891 :  96 - 0x60
      12'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      12'h765: dout <= 8'b00001100; // 1893 :  12 - 0xc
      12'h766: dout <= 8'b00001110; // 1894 :  14 - 0xe
      12'h767: dout <= 8'b00000110; // 1895 :   6 - 0x6
      12'h768: dout <= 8'b01100000; // 1896 :  96 - 0x60 -- Sprite 0xed
      12'h769: dout <= 8'b01110000; // 1897 : 112 - 0x70
      12'h76A: dout <= 8'b00110000; // 1898 :  48 - 0x30
      12'h76B: dout <= 8'b00000000; // 1899 :   0 - 0x0
      12'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      12'h76D: dout <= 8'b00001100; // 1901 :  12 - 0xc
      12'h76E: dout <= 8'b00001110; // 1902 :  14 - 0xe
      12'h76F: dout <= 8'b00000110; // 1903 :   6 - 0x6
      12'h770: dout <= 8'b11111111; // 1904 : 255 - 0xff -- Sprite 0xee
      12'h771: dout <= 8'b11111111; // 1905 : 255 - 0xff
      12'h772: dout <= 8'b10111101; // 1906 : 189 - 0xbd
      12'h773: dout <= 8'b11111111; // 1907 : 255 - 0xff
      12'h774: dout <= 8'b11111111; // 1908 : 255 - 0xff
      12'h775: dout <= 8'b11111011; // 1909 : 251 - 0xfb
      12'h776: dout <= 8'b11111111; // 1910 : 255 - 0xff
      12'h777: dout <= 8'b11111111; // 1911 : 255 - 0xff
      12'h778: dout <= 8'b11111111; // 1912 : 255 - 0xff -- Sprite 0xef
      12'h779: dout <= 8'b11111111; // 1913 : 255 - 0xff
      12'h77A: dout <= 8'b11111011; // 1914 : 251 - 0xfb
      12'h77B: dout <= 8'b11111111; // 1915 : 255 - 0xff
      12'h77C: dout <= 8'b11011111; // 1916 : 223 - 0xdf
      12'h77D: dout <= 8'b11111111; // 1917 : 255 - 0xff
      12'h77E: dout <= 8'b11111111; // 1918 : 255 - 0xff
      12'h77F: dout <= 8'b11111111; // 1919 : 255 - 0xff
      12'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      12'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0 -- Sprite 0xf1
      12'h789: dout <= 8'b10000000; // 1929 : 128 - 0x80
      12'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      12'h78B: dout <= 8'b00000000; // 1931 :   0 - 0x0
      12'h78C: dout <= 8'b00000000; // 1932 :   0 - 0x0
      12'h78D: dout <= 8'b00000000; // 1933 :   0 - 0x0
      12'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      12'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0xf2
      12'h791: dout <= 8'b11000000; // 1937 : 192 - 0xc0
      12'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0 -- Sprite 0xf3
      12'h799: dout <= 8'b11100000; // 1945 : 224 - 0xe0
      12'h79A: dout <= 8'b00000000; // 1946 :   0 - 0x0
      12'h79B: dout <= 8'b00000000; // 1947 :   0 - 0x0
      12'h79C: dout <= 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout <= 8'b00000000; // 1949 :   0 - 0x0
      12'h79E: dout <= 8'b00000000; // 1950 :   0 - 0x0
      12'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      12'h7A0: dout <= 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0xf4
      12'h7A1: dout <= 8'b11110000; // 1953 : 240 - 0xf0
      12'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      12'h7A3: dout <= 8'b00000000; // 1955 :   0 - 0x0
      12'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      12'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      12'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout <= 8'b00000000; // 1960 :   0 - 0x0 -- Sprite 0xf5
      12'h7A9: dout <= 8'b11111000; // 1961 : 248 - 0xf8
      12'h7AA: dout <= 8'b00000000; // 1962 :   0 - 0x0
      12'h7AB: dout <= 8'b00000000; // 1963 :   0 - 0x0
      12'h7AC: dout <= 8'b00000000; // 1964 :   0 - 0x0
      12'h7AD: dout <= 8'b00000000; // 1965 :   0 - 0x0
      12'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      12'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      12'h7B1: dout <= 8'b11111100; // 1969 : 252 - 0xfc
      12'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      12'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      12'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      12'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      12'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout <= 8'b00000000; // 1976 :   0 - 0x0 -- Sprite 0xf7
      12'h7B9: dout <= 8'b11111110; // 1977 : 254 - 0xfe
      12'h7BA: dout <= 8'b00000000; // 1978 :   0 - 0x0
      12'h7BB: dout <= 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout <= 8'b00000000; // 1982 :   0 - 0x0
      12'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0xf8
      12'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      12'h7C2: dout <= 8'b00000000; // 1986 :   0 - 0x0
      12'h7C3: dout <= 8'b00000000; // 1987 :   0 - 0x0
      12'h7C4: dout <= 8'b00000000; // 1988 :   0 - 0x0
      12'h7C5: dout <= 8'b00000000; // 1989 :   0 - 0x0
      12'h7C6: dout <= 8'b00000000; // 1990 :   0 - 0x0
      12'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      12'h7C8: dout <= 8'b11111111; // 1992 : 255 - 0xff -- Sprite 0xf9
      12'h7C9: dout <= 8'b11111111; // 1993 : 255 - 0xff
      12'h7CA: dout <= 8'b11111111; // 1994 : 255 - 0xff
      12'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      12'h7CC: dout <= 8'b10000000; // 1996 : 128 - 0x80
      12'h7CD: dout <= 8'b10000000; // 1997 : 128 - 0x80
      12'h7CE: dout <= 8'b11000000; // 1998 : 192 - 0xc0
      12'h7CF: dout <= 8'b11000000; // 1999 : 192 - 0xc0
      12'h7D0: dout <= 8'b11111111; // 2000 : 255 - 0xff -- Sprite 0xfa
      12'h7D1: dout <= 8'b11111111; // 2001 : 255 - 0xff
      12'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      12'h7D3: dout <= 8'b11111111; // 2003 : 255 - 0xff
      12'h7D4: dout <= 8'b00000000; // 2004 :   0 - 0x0
      12'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      12'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      12'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      12'h7D8: dout <= 8'b11111111; // 2008 : 255 - 0xff -- Sprite 0xfb
      12'h7D9: dout <= 8'b11111111; // 2009 : 255 - 0xff
      12'h7DA: dout <= 8'b11111111; // 2010 : 255 - 0xff
      12'h7DB: dout <= 8'b11111111; // 2011 : 255 - 0xff
      12'h7DC: dout <= 8'b00000001; // 2012 :   1 - 0x1
      12'h7DD: dout <= 8'b00000000; // 2013 :   0 - 0x0
      12'h7DE: dout <= 8'b00000010; // 2014 :   2 - 0x2
      12'h7DF: dout <= 8'b00000010; // 2015 :   2 - 0x2
      12'h7E0: dout <= 8'b11000000; // 2016 : 192 - 0xc0 -- Sprite 0xfc
      12'h7E1: dout <= 8'b11000000; // 2017 : 192 - 0xc0
      12'h7E2: dout <= 8'b10000000; // 2018 : 128 - 0x80
      12'h7E3: dout <= 8'b10000000; // 2019 : 128 - 0x80
      12'h7E4: dout <= 8'b11000000; // 2020 : 192 - 0xc0
      12'h7E5: dout <= 8'b11111111; // 2021 : 255 - 0xff
      12'h7E6: dout <= 8'b11111111; // 2022 : 255 - 0xff
      12'h7E7: dout <= 8'b11111111; // 2023 : 255 - 0xff
      12'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0 -- Sprite 0xfd
      12'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout <= 8'b00000000; // 2026 :   0 - 0x0
      12'h7EB: dout <= 8'b00000000; // 2027 :   0 - 0x0
      12'h7EC: dout <= 8'b00000000; // 2028 :   0 - 0x0
      12'h7ED: dout <= 8'b11111111; // 2029 : 255 - 0xff
      12'h7EE: dout <= 8'b11111111; // 2030 : 255 - 0xff
      12'h7EF: dout <= 8'b11111111; // 2031 : 255 - 0xff
      12'h7F0: dout <= 8'b00000010; // 2032 :   2 - 0x2 -- Sprite 0xfe
      12'h7F1: dout <= 8'b00000010; // 2033 :   2 - 0x2
      12'h7F2: dout <= 8'b00000000; // 2034 :   0 - 0x0
      12'h7F3: dout <= 8'b00000000; // 2035 :   0 - 0x0
      12'h7F4: dout <= 8'b00000000; // 2036 :   0 - 0x0
      12'h7F5: dout <= 8'b11111111; // 2037 : 255 - 0xff
      12'h7F6: dout <= 8'b11111111; // 2038 : 255 - 0xff
      12'h7F7: dout <= 8'b11111111; // 2039 : 255 - 0xff
      12'h7F8: dout <= 8'b11111111; // 2040 : 255 - 0xff -- Sprite 0xff
      12'h7F9: dout <= 8'b11111111; // 2041 : 255 - 0xff
      12'h7FA: dout <= 8'b11111111; // 2042 : 255 - 0xff
      12'h7FB: dout <= 8'b11111111; // 2043 : 255 - 0xff
      12'h7FC: dout <= 8'b11111111; // 2044 : 255 - 0xff
      12'h7FD: dout <= 8'b11111111; // 2045 : 255 - 0xff
      12'h7FE: dout <= 8'b11111111; // 2046 : 255 - 0xff
      12'h7FF: dout <= 8'b11111111; // 2047 : 255 - 0xff
          // Background pattern Table
      12'h800: dout <= 8'b00000000; // 2048 :   0 - 0x0 -- Background 0x0
      12'h801: dout <= 8'b00000000; // 2049 :   0 - 0x0
      12'h802: dout <= 8'b00000000; // 2050 :   0 - 0x0
      12'h803: dout <= 8'b00000000; // 2051 :   0 - 0x0
      12'h804: dout <= 8'b00000000; // 2052 :   0 - 0x0
      12'h805: dout <= 8'b00000000; // 2053 :   0 - 0x0
      12'h806: dout <= 8'b00000000; // 2054 :   0 - 0x0
      12'h807: dout <= 8'b00000000; // 2055 :   0 - 0x0
      12'h808: dout <= 8'b00000101; // 2056 :   5 - 0x5 -- Background 0x1
      12'h809: dout <= 8'b01010101; // 2057 :  85 - 0x55
      12'h80A: dout <= 8'b01010101; // 2058 :  85 - 0x55
      12'h80B: dout <= 8'b01010000; // 2059 :  80 - 0x50
      12'h80C: dout <= 8'b00000000; // 2060 :   0 - 0x0
      12'h80D: dout <= 8'b00000000; // 2061 :   0 - 0x0
      12'h80E: dout <= 8'b00000000; // 2062 :   0 - 0x0
      12'h80F: dout <= 8'b00000000; // 2063 :   0 - 0x0
      12'h810: dout <= 8'b00000101; // 2064 :   5 - 0x5 -- Background 0x2
      12'h811: dout <= 8'b01010000; // 2065 :  80 - 0x50
      12'h812: dout <= 8'b00000101; // 2066 :   5 - 0x5
      12'h813: dout <= 8'b01010000; // 2067 :  80 - 0x50
      12'h814: dout <= 8'b00000000; // 2068 :   0 - 0x0
      12'h815: dout <= 8'b00000000; // 2069 :   0 - 0x0
      12'h816: dout <= 8'b00000000; // 2070 :   0 - 0x0
      12'h817: dout <= 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout <= 8'b00000101; // 2072 :   5 - 0x5 -- Background 0x3
      12'h819: dout <= 8'b01010000; // 2073 :  80 - 0x50
      12'h81A: dout <= 8'b00000101; // 2074 :   5 - 0x5
      12'h81B: dout <= 8'b01010000; // 2075 :  80 - 0x50
      12'h81C: dout <= 8'b00000000; // 2076 :   0 - 0x0
      12'h81D: dout <= 8'b00000000; // 2077 :   0 - 0x0
      12'h81E: dout <= 8'b00000000; // 2078 :   0 - 0x0
      12'h81F: dout <= 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout <= 8'b00000101; // 2080 :   5 - 0x5 -- Background 0x4
      12'h821: dout <= 8'b01010101; // 2081 :  85 - 0x55
      12'h822: dout <= 8'b01010101; // 2082 :  85 - 0x55
      12'h823: dout <= 8'b01010000; // 2083 :  80 - 0x50
      12'h824: dout <= 8'b00000000; // 2084 :   0 - 0x0
      12'h825: dout <= 8'b00000000; // 2085 :   0 - 0x0
      12'h826: dout <= 8'b00000000; // 2086 :   0 - 0x0
      12'h827: dout <= 8'b00000000; // 2087 :   0 - 0x0
      12'h828: dout <= 8'b00000000; // 2088 :   0 - 0x0 -- Background 0x5
      12'h829: dout <= 8'b00000000; // 2089 :   0 - 0x0
      12'h82A: dout <= 8'b00000000; // 2090 :   0 - 0x0
      12'h82B: dout <= 8'b00000000; // 2091 :   0 - 0x0
      12'h82C: dout <= 8'b00000000; // 2092 :   0 - 0x0
      12'h82D: dout <= 8'b00000000; // 2093 :   0 - 0x0
      12'h82E: dout <= 8'b00000000; // 2094 :   0 - 0x0
      12'h82F: dout <= 8'b00000000; // 2095 :   0 - 0x0
      12'h830: dout <= 8'b01010101; // 2096 :  85 - 0x55 -- Background 0x6
      12'h831: dout <= 8'b01010101; // 2097 :  85 - 0x55
      12'h832: dout <= 8'b01010100; // 2098 :  84 - 0x54
      12'h833: dout <= 8'b00000000; // 2099 :   0 - 0x0
      12'h834: dout <= 8'b00000000; // 2100 :   0 - 0x0
      12'h835: dout <= 8'b00000000; // 2101 :   0 - 0x0
      12'h836: dout <= 8'b00000000; // 2102 :   0 - 0x0
      12'h837: dout <= 8'b00010101; // 2103 :  21 - 0x15
      12'h838: dout <= 8'b10101010; // 2104 : 170 - 0xaa -- Background 0x7
      12'h839: dout <= 8'b10011010; // 2105 : 154 - 0x9a
      12'h83A: dout <= 8'b10010100; // 2106 : 148 - 0x94
      12'h83B: dout <= 8'b00000000; // 2107 :   0 - 0x0
      12'h83C: dout <= 8'b00000000; // 2108 :   0 - 0x0
      12'h83D: dout <= 8'b00000000; // 2109 :   0 - 0x0
      12'h83E: dout <= 8'b00000000; // 2110 :   0 - 0x0
      12'h83F: dout <= 8'b00010110; // 2111 :  22 - 0x16
      12'h840: dout <= 8'b01010000; // 2112 :  80 - 0x50 -- Background 0x8
      12'h841: dout <= 8'b00000101; // 2113 :   5 - 0x5
      12'h842: dout <= 8'b10010100; // 2114 : 148 - 0x94
      12'h843: dout <= 8'b00000000; // 2115 :   0 - 0x0
      12'h844: dout <= 8'b00000000; // 2116 :   0 - 0x0
      12'h845: dout <= 8'b00000000; // 2117 :   0 - 0x0
      12'h846: dout <= 8'b00000000; // 2118 :   0 - 0x0
      12'h847: dout <= 8'b00010101; // 2119 :  21 - 0x15
      12'h848: dout <= 8'b01010000; // 2120 :  80 - 0x50 -- Background 0x9
      12'h849: dout <= 8'b00000101; // 2121 :   5 - 0x5
      12'h84A: dout <= 8'b10010100; // 2122 : 148 - 0x94
      12'h84B: dout <= 8'b00000000; // 2123 :   0 - 0x0
      12'h84C: dout <= 8'b00000000; // 2124 :   0 - 0x0
      12'h84D: dout <= 8'b00000000; // 2125 :   0 - 0x0
      12'h84E: dout <= 8'b00000000; // 2126 :   0 - 0x0
      12'h84F: dout <= 8'b00010110; // 2127 :  22 - 0x16
      12'h850: dout <= 8'b10100110; // 2128 : 166 - 0xa6 -- Background 0xa
      12'h851: dout <= 8'b10101010; // 2129 : 170 - 0xaa
      12'h852: dout <= 8'b10010100; // 2130 : 148 - 0x94
      12'h853: dout <= 8'b00000000; // 2131 :   0 - 0x0
      12'h854: dout <= 8'b00000000; // 2132 :   0 - 0x0
      12'h855: dout <= 8'b00000000; // 2133 :   0 - 0x0
      12'h856: dout <= 8'b00000000; // 2134 :   0 - 0x0
      12'h857: dout <= 8'b00010101; // 2135 :  21 - 0x15
      12'h858: dout <= 8'b01010101; // 2136 :  85 - 0x55 -- Background 0xb
      12'h859: dout <= 8'b01010101; // 2137 :  85 - 0x55
      12'h85A: dout <= 8'b01010100; // 2138 :  84 - 0x54
      12'h85B: dout <= 8'b00000000; // 2139 :   0 - 0x0
      12'h85C: dout <= 8'b00000000; // 2140 :   0 - 0x0
      12'h85D: dout <= 8'b00000000; // 2141 :   0 - 0x0
      12'h85E: dout <= 8'b00000000; // 2142 :   0 - 0x0
      12'h85F: dout <= 8'b00001110; // 2143 :  14 - 0xe
      12'h860: dout <= 8'b01010101; // 2144 :  85 - 0x55 -- Background 0xc
      12'h861: dout <= 8'b01010100; // 2145 :  84 - 0x54
      12'h862: dout <= 8'b00000000; // 2146 :   0 - 0x0
      12'h863: dout <= 8'b00000000; // 2147 :   0 - 0x0
      12'h864: dout <= 8'b00000000; // 2148 :   0 - 0x0
      12'h865: dout <= 8'b00000000; // 2149 :   0 - 0x0
      12'h866: dout <= 8'b00011010; // 2150 :  26 - 0x1a
      12'h867: dout <= 8'b10011101; // 2151 : 157 - 0x9d
      12'h868: dout <= 8'b01010101; // 2152 :  85 - 0x55 -- Background 0xd
      12'h869: dout <= 8'b01010100; // 2153 :  84 - 0x54
      12'h86A: dout <= 8'b00000000; // 2154 :   0 - 0x0
      12'h86B: dout <= 8'b00000000; // 2155 :   0 - 0x0
      12'h86C: dout <= 8'b00000000; // 2156 :   0 - 0x0
      12'h86D: dout <= 8'b00000000; // 2157 :   0 - 0x0
      12'h86E: dout <= 8'b00010111; // 2158 :  23 - 0x17
      12'h86F: dout <= 8'b01010101; // 2159 :  85 - 0x55
      12'h870: dout <= 8'b00000101; // 2160 :   5 - 0x5 -- Background 0xe
      12'h871: dout <= 8'b01010100; // 2161 :  84 - 0x54
      12'h872: dout <= 8'b00000000; // 2162 :   0 - 0x0
      12'h873: dout <= 8'b00000000; // 2163 :   0 - 0x0
      12'h874: dout <= 8'b00000000; // 2164 :   0 - 0x0
      12'h875: dout <= 8'b00000000; // 2165 :   0 - 0x0
      12'h876: dout <= 8'b00010101; // 2166 :  21 - 0x15
      12'h877: dout <= 8'b01010000; // 2167 :  80 - 0x50
      12'h878: dout <= 8'b00000101; // 2168 :   5 - 0x5 -- Background 0xf
      12'h879: dout <= 8'b01010100; // 2169 :  84 - 0x54
      12'h87A: dout <= 8'b00000000; // 2170 :   0 - 0x0
      12'h87B: dout <= 8'b00000000; // 2171 :   0 - 0x0
      12'h87C: dout <= 8'b00000000; // 2172 :   0 - 0x0
      12'h87D: dout <= 8'b00000000; // 2173 :   0 - 0x0
      12'h87E: dout <= 8'b00010111; // 2174 :  23 - 0x17
      12'h87F: dout <= 8'b01010101; // 2175 :  85 - 0x55
      12'h880: dout <= 8'b01010101; // 2176 :  85 - 0x55 -- Background 0x10
      12'h881: dout <= 8'b01010100; // 2177 :  84 - 0x54
      12'h882: dout <= 8'b00000000; // 2178 :   0 - 0x0
      12'h883: dout <= 8'b00000000; // 2179 :   0 - 0x0
      12'h884: dout <= 8'b00000000; // 2180 :   0 - 0x0
      12'h885: dout <= 8'b00000000; // 2181 :   0 - 0x0
      12'h886: dout <= 8'b00011010; // 2182 :  26 - 0x1a
      12'h887: dout <= 8'b10011101; // 2183 : 157 - 0x9d
      12'h888: dout <= 8'b01010101; // 2184 :  85 - 0x55 -- Background 0x11
      12'h889: dout <= 8'b01010100; // 2185 :  84 - 0x54
      12'h88A: dout <= 8'b00000000; // 2186 :   0 - 0x0
      12'h88B: dout <= 8'b00000000; // 2187 :   0 - 0x0
      12'h88C: dout <= 8'b00000000; // 2188 :   0 - 0x0
      12'h88D: dout <= 8'b00000000; // 2189 :   0 - 0x0
      12'h88E: dout <= 8'b00001110; // 2190 :  14 - 0xe
      12'h88F: dout <= 8'b00000111; // 2191 :   7 - 0x7
      12'h890: dout <= 8'b01010101; // 2192 :  85 - 0x55 -- Background 0x12
      12'h891: dout <= 8'b01010101; // 2193 :  85 - 0x55
      12'h892: dout <= 8'b01000000; // 2194 :  64 - 0x40
      12'h893: dout <= 8'b00000000; // 2195 :   0 - 0x0
      12'h894: dout <= 8'b00000000; // 2196 :   0 - 0x0
      12'h895: dout <= 8'b00010101; // 2197 :  21 - 0x15
      12'h896: dout <= 8'b01010101; // 2198 :  85 - 0x55
      12'h897: dout <= 8'b01010101; // 2199 :  85 - 0x55
      12'h898: dout <= 8'b01010101; // 2200 :  85 - 0x55 -- Background 0x13
      12'h899: dout <= 8'b10101001; // 2201 : 169 - 0xa9
      12'h89A: dout <= 8'b01000000; // 2202 :  64 - 0x40
      12'h89B: dout <= 8'b00000000; // 2203 :   0 - 0x0
      12'h89C: dout <= 8'b00000000; // 2204 :   0 - 0x0
      12'h89D: dout <= 8'b00010110; // 2205 :  22 - 0x16
      12'h89E: dout <= 8'b01010101; // 2206 :  85 - 0x55
      12'h89F: dout <= 8'b01101010; // 2207 : 106 - 0x6a
      12'h8A0: dout <= 8'b01010101; // 2208 :  85 - 0x55 -- Background 0x14
      12'h8A1: dout <= 8'b01011001; // 2209 :  89 - 0x59
      12'h8A2: dout <= 8'b01000000; // 2210 :  64 - 0x40
      12'h8A3: dout <= 8'b00000000; // 2211 :   0 - 0x0
      12'h8A4: dout <= 8'b00000000; // 2212 :   0 - 0x0
      12'h8A5: dout <= 8'b00010101; // 2213 :  21 - 0x15
      12'h8A6: dout <= 8'b01000000; // 2214 :  64 - 0x40
      12'h8A7: dout <= 8'b01010101; // 2215 :  85 - 0x55
      12'h8A8: dout <= 8'b01010101; // 2216 :  85 - 0x55 -- Background 0x15
      12'h8A9: dout <= 8'b01011001; // 2217 :  89 - 0x59
      12'h8AA: dout <= 8'b01000000; // 2218 :  64 - 0x40
      12'h8AB: dout <= 8'b00000000; // 2219 :   0 - 0x0
      12'h8AC: dout <= 8'b00000000; // 2220 :   0 - 0x0
      12'h8AD: dout <= 8'b00010110; // 2221 :  22 - 0x16
      12'h8AE: dout <= 8'b01010101; // 2222 :  85 - 0x55
      12'h8AF: dout <= 8'b01101010; // 2223 : 106 - 0x6a
      12'h8B0: dout <= 8'b01010101; // 2224 :  85 - 0x55 -- Background 0x16
      12'h8B1: dout <= 8'b10101001; // 2225 : 169 - 0xa9
      12'h8B2: dout <= 8'b01000000; // 2226 :  64 - 0x40
      12'h8B3: dout <= 8'b00000000; // 2227 :   0 - 0x0
      12'h8B4: dout <= 8'b00000000; // 2228 :   0 - 0x0
      12'h8B5: dout <= 8'b00010101; // 2229 :  21 - 0x15
      12'h8B6: dout <= 8'b01010101; // 2230 :  85 - 0x55
      12'h8B7: dout <= 8'b01010101; // 2231 :  85 - 0x55
      12'h8B8: dout <= 8'b01010101; // 2232 :  85 - 0x55 -- Background 0x17
      12'h8B9: dout <= 8'b01010101; // 2233 :  85 - 0x55
      12'h8BA: dout <= 8'b01000000; // 2234 :  64 - 0x40
      12'h8BB: dout <= 8'b00000000; // 2235 :   0 - 0x0
      12'h8BC: dout <= 8'b00000000; // 2236 :   0 - 0x0
      12'h8BD: dout <= 8'b00010100; // 2237 :  20 - 0x14
      12'h8BE: dout <= 8'b00000110; // 2238 :   6 - 0x6
      12'h8BF: dout <= 8'b00001000; // 2239 :   8 - 0x8
      12'h8C0: dout <= 8'b01010101; // 2240 :  85 - 0x55 -- Background 0x18
      12'h8C1: dout <= 8'b01000000; // 2241 :  64 - 0x40
      12'h8C2: dout <= 8'b00000000; // 2242 :   0 - 0x0
      12'h8C3: dout <= 8'b00000000; // 2243 :   0 - 0x0
      12'h8C4: dout <= 8'b00011010; // 2244 :  26 - 0x1a
      12'h8C5: dout <= 8'b01010111; // 2245 :  87 - 0x57
      12'h8C6: dout <= 8'b01010101; // 2246 :  85 - 0x55
      12'h8C7: dout <= 8'b01011101; // 2247 :  93 - 0x5d
      12'h8C8: dout <= 8'b01011010; // 2248 :  90 - 0x5a -- Background 0x19
      12'h8C9: dout <= 8'b01000000; // 2249 :  64 - 0x40
      12'h8CA: dout <= 8'b00000000; // 2250 :   0 - 0x0
      12'h8CB: dout <= 8'b00000000; // 2251 :   0 - 0x0
      12'h8CC: dout <= 8'b00010101; // 2252 :  21 - 0x15
      12'h8CD: dout <= 8'b01010111; // 2253 :  87 - 0x57
      12'h8CE: dout <= 8'b01011010; // 2254 :  90 - 0x5a
      12'h8CF: dout <= 8'b01011101; // 2255 :  93 - 0x5d
      12'h8D0: dout <= 8'b01010101; // 2256 :  85 - 0x55 -- Background 0x1a
      12'h8D1: dout <= 8'b01000000; // 2257 :  64 - 0x40
      12'h8D2: dout <= 8'b00000000; // 2258 :   0 - 0x0
      12'h8D3: dout <= 8'b00000000; // 2259 :   0 - 0x0
      12'h8D4: dout <= 8'b00010000; // 2260 :  16 - 0x10
      12'h8D5: dout <= 8'b00010101; // 2261 :  21 - 0x15
      12'h8D6: dout <= 8'b01011010; // 2262 :  90 - 0x5a
      12'h8D7: dout <= 8'b01010101; // 2263 :  85 - 0x55
      12'h8D8: dout <= 8'b01010101; // 2264 :  85 - 0x55 -- Background 0x1b
      12'h8D9: dout <= 8'b01000000; // 2265 :  64 - 0x40
      12'h8DA: dout <= 8'b00000000; // 2266 :   0 - 0x0
      12'h8DB: dout <= 8'b00000000; // 2267 :   0 - 0x0
      12'h8DC: dout <= 8'b00010101; // 2268 :  21 - 0x15
      12'h8DD: dout <= 8'b01010111; // 2269 :  87 - 0x57
      12'h8DE: dout <= 8'b01011010; // 2270 :  90 - 0x5a
      12'h8DF: dout <= 8'b01011101; // 2271 :  93 - 0x5d
      12'h8E0: dout <= 8'b01011010; // 2272 :  90 - 0x5a -- Background 0x1c
      12'h8E1: dout <= 8'b01000000; // 2273 :  64 - 0x40
      12'h8E2: dout <= 8'b00000000; // 2274 :   0 - 0x0
      12'h8E3: dout <= 8'b00000000; // 2275 :   0 - 0x0
      12'h8E4: dout <= 8'b00011010; // 2276 :  26 - 0x1a
      12'h8E5: dout <= 8'b01010111; // 2277 :  87 - 0x57
      12'h8E6: dout <= 8'b01010101; // 2278 :  85 - 0x55
      12'h8E7: dout <= 8'b01011101; // 2279 :  93 - 0x5d
      12'h8E8: dout <= 8'b01010101; // 2280 :  85 - 0x55 -- Background 0x1d
      12'h8E9: dout <= 8'b01000000; // 2281 :  64 - 0x40
      12'h8EA: dout <= 8'b00000000; // 2282 :   0 - 0x0
      12'h8EB: dout <= 8'b00000000; // 2283 :   0 - 0x0
      12'h8EC: dout <= 8'b00010100; // 2284 :  20 - 0x14
      12'h8ED: dout <= 8'b00000011; // 2285 :   3 - 0x3
      12'h8EE: dout <= 8'b00001000; // 2286 :   8 - 0x8
      12'h8EF: dout <= 8'b10101101; // 2287 : 173 - 0xad
      12'h8F0: dout <= 8'b01010101; // 2288 :  85 - 0x55 -- Background 0x1e
      12'h8F1: dout <= 8'b01010000; // 2289 :  80 - 0x50
      12'h8F2: dout <= 8'b00000000; // 2290 :   0 - 0x0
      12'h8F3: dout <= 8'b00010101; // 2291 :  21 - 0x15
      12'h8F4: dout <= 8'b01110101; // 2292 : 117 - 0x75
      12'h8F5: dout <= 8'b01010101; // 2293 :  85 - 0x55
      12'h8F6: dout <= 8'b01010111; // 2294 :  87 - 0x57
      12'h8F7: dout <= 8'b01010101; // 2295 :  85 - 0x55
      12'h8F8: dout <= 8'b01010101; // 2296 :  85 - 0x55 -- Background 0x1f
      12'h8F9: dout <= 8'b01010000; // 2297 :  80 - 0x50
      12'h8FA: dout <= 8'b00000000; // 2298 :   0 - 0x0
      12'h8FB: dout <= 8'b00010101; // 2299 :  21 - 0x15
      12'h8FC: dout <= 8'b01010111; // 2300 :  87 - 0x57
      12'h8FD: dout <= 8'b01010101; // 2301 :  85 - 0x55
      12'h8FE: dout <= 8'b01010101; // 2302 :  85 - 0x55
      12'h8FF: dout <= 8'b01010101; // 2303 :  85 - 0x55
      12'h900: dout <= 8'b01010101; // 2304 :  85 - 0x55 -- Background 0x20
      12'h901: dout <= 8'b11010000; // 2305 : 208 - 0xd0
      12'h902: dout <= 8'b00000000; // 2306 :   0 - 0x0
      12'h903: dout <= 8'b00010111; // 2307 :  23 - 0x17
      12'h904: dout <= 8'b01010101; // 2308 :  85 - 0x55
      12'h905: dout <= 8'b01010101; // 2309 :  85 - 0x55
      12'h906: dout <= 8'b00000001; // 2310 :   1 - 0x1
      12'h907: dout <= 8'b01010111; // 2311 :  87 - 0x57
      12'h908: dout <= 8'b01010101; // 2312 :  85 - 0x55 -- Background 0x21
      12'h909: dout <= 8'b01010000; // 2313 :  80 - 0x50
      12'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout <= 8'b00010101; // 2315 :  21 - 0x15
      12'h90C: dout <= 8'b01010101; // 2316 :  85 - 0x55
      12'h90D: dout <= 8'b01110101; // 2317 : 117 - 0x75
      12'h90E: dout <= 8'b01010101; // 2318 :  85 - 0x55
      12'h90F: dout <= 8'b01010101; // 2319 :  85 - 0x55
      12'h910: dout <= 8'b01010101; // 2320 :  85 - 0x55 -- Background 0x22
      12'h911: dout <= 8'b01010000; // 2321 :  80 - 0x50
      12'h912: dout <= 8'b00000000; // 2322 :   0 - 0x0
      12'h913: dout <= 8'b00010101; // 2323 :  21 - 0x15
      12'h914: dout <= 8'b01110101; // 2324 : 117 - 0x75
      12'h915: dout <= 8'b01010101; // 2325 :  85 - 0x55
      12'h916: dout <= 8'b11010101; // 2326 : 213 - 0xd5
      12'h917: dout <= 8'b01010101; // 2327 :  85 - 0x55
      12'h918: dout <= 8'b01010101; // 2328 :  85 - 0x55 -- Background 0x23
      12'h919: dout <= 8'b01010000; // 2329 :  80 - 0x50
      12'h91A: dout <= 8'b00000000; // 2330 :   0 - 0x0
      12'h91B: dout <= 8'b00011001; // 2331 :  25 - 0x19
      12'h91C: dout <= 8'b00001101; // 2332 :  13 - 0xd
      12'h91D: dout <= 8'b00001000; // 2333 :   8 - 0x8
      12'h91E: dout <= 8'b11110111; // 2334 : 247 - 0xf7
      12'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout <= 8'b01010000; // 2336 :  80 - 0x50 -- Background 0x24
      12'h921: dout <= 8'b00000000; // 2337 :   0 - 0x0
      12'h922: dout <= 8'b00011010; // 2338 :  26 - 0x1a
      12'h923: dout <= 8'b10101001; // 2339 : 169 - 0xa9
      12'h924: dout <= 8'b10101010; // 2340 : 170 - 0xaa
      12'h925: dout <= 8'b10011001; // 2341 : 153 - 0x99
      12'h926: dout <= 8'b01011001; // 2342 :  89 - 0x59
      12'h927: dout <= 8'b10101010; // 2343 : 170 - 0xaa
      12'h928: dout <= 8'b10010000; // 2344 : 144 - 0x90 -- Background 0x25
      12'h929: dout <= 8'b00000000; // 2345 :   0 - 0x0
      12'h92A: dout <= 8'b00010101; // 2346 :  21 - 0x15
      12'h92B: dout <= 8'b01011001; // 2347 :  89 - 0x59
      12'h92C: dout <= 8'b10010101; // 2348 : 149 - 0x95
      12'h92D: dout <= 8'b10011001; // 2349 : 153 - 0x99
      12'h92E: dout <= 8'b01011001; // 2350 :  89 - 0x59
      12'h92F: dout <= 8'b10010101; // 2351 : 149 - 0x95
      12'h930: dout <= 8'b01010000; // 2352 :  80 - 0x50 -- Background 0x26
      12'h931: dout <= 8'b00000000; // 2353 :   0 - 0x0
      12'h932: dout <= 8'b00010000; // 2354 :  16 - 0x10
      12'h933: dout <= 8'b00010101; // 2355 :  21 - 0x15
      12'h934: dout <= 8'b01010101; // 2356 :  85 - 0x55
      12'h935: dout <= 8'b01010101; // 2357 :  85 - 0x55
      12'h936: dout <= 8'b01010101; // 2358 :  85 - 0x55
      12'h937: dout <= 8'b01010101; // 2359 :  85 - 0x55
      12'h938: dout <= 8'b01010000; // 2360 :  80 - 0x50 -- Background 0x27
      12'h939: dout <= 8'b00000000; // 2361 :   0 - 0x0
      12'h93A: dout <= 8'b00010101; // 2362 :  21 - 0x15
      12'h93B: dout <= 8'b01011001; // 2363 :  89 - 0x59
      12'h93C: dout <= 8'b10010101; // 2364 : 149 - 0x95
      12'h93D: dout <= 8'b10011001; // 2365 : 153 - 0x99
      12'h93E: dout <= 8'b01011001; // 2366 :  89 - 0x59
      12'h93F: dout <= 8'b10010101; // 2367 : 149 - 0x95
      12'h940: dout <= 8'b10010000; // 2368 : 144 - 0x90 -- Background 0x28
      12'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout <= 8'b00011010; // 2370 :  26 - 0x1a
      12'h943: dout <= 8'b10101001; // 2371 : 169 - 0xa9
      12'h944: dout <= 8'b10010101; // 2372 : 149 - 0x95
      12'h945: dout <= 8'b10011010; // 2373 : 154 - 0x9a
      12'h946: dout <= 8'b10101001; // 2374 : 169 - 0xa9
      12'h947: dout <= 8'b10101010; // 2375 : 170 - 0xaa
      12'h948: dout <= 8'b01010000; // 2376 :  80 - 0x50 -- Background 0x29
      12'h949: dout <= 8'b00000000; // 2377 :   0 - 0x0
      12'h94A: dout <= 8'b00011001; // 2378 :  25 - 0x19
      12'h94B: dout <= 8'b00000011; // 2379 :   3 - 0x3
      12'h94C: dout <= 8'b00001000; // 2380 :   8 - 0x8
      12'h94D: dout <= 8'b10111110; // 2381 : 190 - 0xbe
      12'h94E: dout <= 8'b00000000; // 2382 :   0 - 0x0
      12'h94F: dout <= 8'b10000110; // 2383 : 134 - 0x86
      12'h950: dout <= 8'b00000000; // 2384 :   0 - 0x0 -- Background 0x2a
      12'h951: dout <= 8'b00010101; // 2385 :  21 - 0x15
      12'h952: dout <= 8'b01010111; // 2386 :  87 - 0x57
      12'h953: dout <= 8'b01101010; // 2387 : 106 - 0x6a
      12'h954: dout <= 8'b01010110; // 2388 :  86 - 0x56
      12'h955: dout <= 8'b10100111; // 2389 : 167 - 0xa7
      12'h956: dout <= 8'b01010101; // 2390 :  85 - 0x55
      12'h957: dout <= 8'b01010000; // 2391 :  80 - 0x50
      12'h958: dout <= 8'b00000000; // 2392 :   0 - 0x0 -- Background 0x2b
      12'h959: dout <= 8'b00010101; // 2393 :  21 - 0x15
      12'h95A: dout <= 8'b01010111; // 2394 :  87 - 0x57
      12'h95B: dout <= 8'b01010101; // 2395 :  85 - 0x55
      12'h95C: dout <= 8'b01110101; // 2396 : 117 - 0x75
      12'h95D: dout <= 8'b01010111; // 2397 :  87 - 0x57
      12'h95E: dout <= 8'b01010101; // 2398 :  85 - 0x55
      12'h95F: dout <= 8'b01010000; // 2399 :  80 - 0x50
      12'h960: dout <= 8'b00000000; // 2400 :   0 - 0x0 -- Background 0x2c
      12'h961: dout <= 8'b00010000; // 2401 :  16 - 0x10
      12'h962: dout <= 8'b00010101; // 2402 :  21 - 0x15
      12'h963: dout <= 8'b01010101; // 2403 :  85 - 0x55
      12'h964: dout <= 8'b01110101; // 2404 : 117 - 0x75
      12'h965: dout <= 8'b01010101; // 2405 :  85 - 0x55
      12'h966: dout <= 8'b01010101; // 2406 :  85 - 0x55
      12'h967: dout <= 8'b01010000; // 2407 :  80 - 0x50
      12'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0 -- Background 0x2d
      12'h969: dout <= 8'b00010101; // 2409 :  21 - 0x15
      12'h96A: dout <= 8'b01010111; // 2410 :  87 - 0x57
      12'h96B: dout <= 8'b01010101; // 2411 :  85 - 0x55
      12'h96C: dout <= 8'b01110101; // 2412 : 117 - 0x75
      12'h96D: dout <= 8'b01010111; // 2413 :  87 - 0x57
      12'h96E: dout <= 8'b01010101; // 2414 :  85 - 0x55
      12'h96F: dout <= 8'b01010000; // 2415 :  80 - 0x50
      12'h970: dout <= 8'b00000000; // 2416 :   0 - 0x0 -- Background 0x2e
      12'h971: dout <= 8'b00010101; // 2417 :  21 - 0x15
      12'h972: dout <= 8'b01010111; // 2418 :  87 - 0x57
      12'h973: dout <= 8'b01101010; // 2419 : 106 - 0x6a
      12'h974: dout <= 8'b01010110; // 2420 :  86 - 0x56
      12'h975: dout <= 8'b10100111; // 2421 : 167 - 0xa7
      12'h976: dout <= 8'b01010101; // 2422 :  85 - 0x55
      12'h977: dout <= 8'b01010000; // 2423 :  80 - 0x50
      12'h978: dout <= 8'b00000000; // 2424 :   0 - 0x0 -- Background 0x2f
      12'h979: dout <= 8'b00011001; // 2425 :  25 - 0x19
      12'h97A: dout <= 8'b00000011; // 2426 :   3 - 0x3
      12'h97B: dout <= 8'b00001000; // 2427 :   8 - 0x8
      12'h97C: dout <= 8'b11011101; // 2428 : 221 - 0xdd
      12'h97D: dout <= 8'b00000000; // 2429 :   0 - 0x0
      12'h97E: dout <= 8'b01110011; // 2430 : 115 - 0x73
      12'h97F: dout <= 8'b00000000; // 2431 :   0 - 0x0
      12'h980: dout <= 8'b00011001; // 2432 :  25 - 0x19 -- Background 0x30
      12'h981: dout <= 8'b01100101; // 2433 : 101 - 0x65
      12'h982: dout <= 8'b10010110; // 2434 : 150 - 0x96
      12'h983: dout <= 8'b10100101; // 2435 : 165 - 0xa5
      12'h984: dout <= 8'b01011010; // 2436 :  90 - 0x5a
      12'h985: dout <= 8'b10010110; // 2437 : 150 - 0x96
      12'h986: dout <= 8'b01011001; // 2438 :  89 - 0x59
      12'h987: dout <= 8'b01100100; // 2439 : 100 - 0x64
      12'h988: dout <= 8'b00011001; // 2440 :  25 - 0x19 -- Background 0x31
      12'h989: dout <= 8'b01100101; // 2441 : 101 - 0x65
      12'h98A: dout <= 8'b10010110; // 2442 : 150 - 0x96
      12'h98B: dout <= 8'b10100101; // 2443 : 165 - 0xa5
      12'h98C: dout <= 8'b01011010; // 2444 :  90 - 0x5a
      12'h98D: dout <= 8'b10010110; // 2445 : 150 - 0x96
      12'h98E: dout <= 8'b01011001; // 2446 :  89 - 0x59
      12'h98F: dout <= 8'b01100100; // 2447 : 100 - 0x64
      12'h990: dout <= 8'b00011111; // 2448 :  31 - 0x1f -- Background 0x32
      12'h991: dout <= 8'b01111101; // 2449 : 125 - 0x7d
      12'h992: dout <= 8'b11010101; // 2450 : 213 - 0xd5
      12'h993: dout <= 8'b01010000; // 2451 :  80 - 0x50
      12'h994: dout <= 8'b00000101; // 2452 :   5 - 0x5
      12'h995: dout <= 8'b01010111; // 2453 :  87 - 0x57
      12'h996: dout <= 8'b11111111; // 2454 : 255 - 0xff
      12'h997: dout <= 8'b01110100; // 2455 : 116 - 0x74
      12'h998: dout <= 8'b00011001; // 2456 :  25 - 0x19 -- Background 0x33
      12'h999: dout <= 8'b01100101; // 2457 : 101 - 0x65
      12'h99A: dout <= 8'b10010110; // 2458 : 150 - 0x96
      12'h99B: dout <= 8'b10100101; // 2459 : 165 - 0xa5
      12'h99C: dout <= 8'b01011010; // 2460 :  90 - 0x5a
      12'h99D: dout <= 8'b10010110; // 2461 : 150 - 0x96
      12'h99E: dout <= 8'b01011001; // 2462 :  89 - 0x59
      12'h99F: dout <= 8'b01100100; // 2463 : 100 - 0x64
      12'h9A0: dout <= 8'b00011001; // 2464 :  25 - 0x19 -- Background 0x34
      12'h9A1: dout <= 8'b01100101; // 2465 : 101 - 0x65
      12'h9A2: dout <= 8'b10010110; // 2466 : 150 - 0x96
      12'h9A3: dout <= 8'b10100101; // 2467 : 165 - 0xa5
      12'h9A4: dout <= 8'b01011010; // 2468 :  90 - 0x5a
      12'h9A5: dout <= 8'b10010110; // 2469 : 150 - 0x96
      12'h9A6: dout <= 8'b01011001; // 2470 :  89 - 0x59
      12'h9A7: dout <= 8'b01100100; // 2471 : 100 - 0x64
      12'h9A8: dout <= 8'b00011110; // 2472 :  30 - 0x1e -- Background 0x35
      12'h9A9: dout <= 8'b00001111; // 2473 :  15 - 0xf
      12'h9AA: dout <= 8'b00001000; // 2474 :   8 - 0x8
      12'h9AB: dout <= 8'b11110111; // 2475 : 247 - 0xf7
      12'h9AC: dout <= 8'b00000000; // 2476 :   0 - 0x0
      12'h9AD: dout <= 8'b01100111; // 2477 : 103 - 0x67
      12'h9AE: dout <= 8'b00000000; // 2478 :   0 - 0x0
      12'h9AF: dout <= 8'b00010101; // 2479 :  21 - 0x15
      12'h9B0: dout <= 8'b01110101; // 2480 : 117 - 0x75 -- Background 0x36
      12'h9B1: dout <= 8'b01010110; // 2481 :  86 - 0x56
      12'h9B2: dout <= 8'b10100101; // 2482 : 165 - 0xa5
      12'h9B3: dout <= 8'b01011010; // 2483 :  90 - 0x5a
      12'h9B4: dout <= 8'b10010101; // 2484 : 149 - 0x95
      12'h9B5: dout <= 8'b01011101; // 2485 :  93 - 0x5d
      12'h9B6: dout <= 8'b11010100; // 2486 : 212 - 0xd4
      12'h9B7: dout <= 8'b00010101; // 2487 :  21 - 0x15
      12'h9B8: dout <= 8'b01010101; // 2488 :  85 - 0x55 -- Background 0x37
      12'h9B9: dout <= 8'b01110101; // 2489 : 117 - 0x75
      12'h9BA: dout <= 8'b01010101; // 2490 :  85 - 0x55
      12'h9BB: dout <= 8'b01010101; // 2491 :  85 - 0x55
      12'h9BC: dout <= 8'b01011101; // 2492 :  93 - 0x5d
      12'h9BD: dout <= 8'b01010101; // 2493 :  85 - 0x55
      12'h9BE: dout <= 8'b11010100; // 2494 : 212 - 0xd4
      12'h9BF: dout <= 8'b00010101; // 2495 :  21 - 0x15
      12'h9C0: dout <= 8'b01101110; // 2496 : 110 - 0x6e -- Background 0x38
      12'h9C1: dout <= 8'b01110101; // 2497 : 117 - 0x75
      12'h9C2: dout <= 8'b01010000; // 2498 :  80 - 0x50
      12'h9C3: dout <= 8'b00000101; // 2499 :   5 - 0x5
      12'h9C4: dout <= 8'b01011101; // 2500 :  93 - 0x5d
      12'h9C5: dout <= 8'b10111001; // 2501 : 185 - 0xb9
      12'h9C6: dout <= 8'b01010100; // 2502 :  84 - 0x54
      12'h9C7: dout <= 8'b00010101; // 2503 :  21 - 0x15
      12'h9C8: dout <= 8'b01010101; // 2504 :  85 - 0x55 -- Background 0x39
      12'h9C9: dout <= 8'b01110101; // 2505 : 117 - 0x75
      12'h9CA: dout <= 8'b01010101; // 2506 :  85 - 0x55
      12'h9CB: dout <= 8'b01010101; // 2507 :  85 - 0x55
      12'h9CC: dout <= 8'b01011101; // 2508 :  93 - 0x5d
      12'h9CD: dout <= 8'b01010101; // 2509 :  85 - 0x55
      12'h9CE: dout <= 8'b11010100; // 2510 : 212 - 0xd4
      12'h9CF: dout <= 8'b00010101; // 2511 :  21 - 0x15
      12'h9D0: dout <= 8'b01110101; // 2512 : 117 - 0x75 -- Background 0x3a
      12'h9D1: dout <= 8'b01010101; // 2513 :  85 - 0x55
      12'h9D2: dout <= 8'b01101010; // 2514 : 106 - 0x6a
      12'h9D3: dout <= 8'b10101001; // 2515 : 169 - 0xa9
      12'h9D4: dout <= 8'b01010101; // 2516 :  85 - 0x55
      12'h9D5: dout <= 8'b01011101; // 2517 :  93 - 0x5d
      12'h9D6: dout <= 8'b11010100; // 2518 : 212 - 0xd4
      12'h9D7: dout <= 8'b00010101; // 2519 :  21 - 0x15
      12'h9D8: dout <= 8'b00001111; // 2520 :  15 - 0xf -- Background 0x3b
      12'h9D9: dout <= 8'b00001000; // 2521 :   8 - 0x8
      12'h9DA: dout <= 8'b11111000; // 2522 : 248 - 0xf8
      12'h9DB: dout <= 8'b00000000; // 2523 :   0 - 0x0
      12'h9DC: dout <= 8'b01100111; // 2524 : 103 - 0x67
      12'h9DD: dout <= 8'b00000000; // 2525 :   0 - 0x0
      12'h9DE: dout <= 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout <= 8'b00000000; // 2528 :   0 - 0x0 -- Background 0x3c
      12'h9E1: dout <= 8'b00000000; // 2529 :   0 - 0x0
      12'h9E2: dout <= 8'b00000000; // 2530 :   0 - 0x0
      12'h9E3: dout <= 8'b00000000; // 2531 :   0 - 0x0
      12'h9E4: dout <= 8'b00000000; // 2532 :   0 - 0x0
      12'h9E5: dout <= 8'b00000000; // 2533 :   0 - 0x0
      12'h9E6: dout <= 8'b00000000; // 2534 :   0 - 0x0
      12'h9E7: dout <= 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0 -- Background 0x3d
      12'h9E9: dout <= 8'b00000000; // 2537 :   0 - 0x0
      12'h9EA: dout <= 8'b00000000; // 2538 :   0 - 0x0
      12'h9EB: dout <= 8'b00000000; // 2539 :   0 - 0x0
      12'h9EC: dout <= 8'b00000000; // 2540 :   0 - 0x0
      12'h9ED: dout <= 8'b00000000; // 2541 :   0 - 0x0
      12'h9EE: dout <= 8'b00000000; // 2542 :   0 - 0x0
      12'h9EF: dout <= 8'b00000000; // 2543 :   0 - 0x0
      12'h9F0: dout <= 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x3e
      12'h9F1: dout <= 8'b00000000; // 2545 :   0 - 0x0
      12'h9F2: dout <= 8'b00000000; // 2546 :   0 - 0x0
      12'h9F3: dout <= 8'b00000000; // 2547 :   0 - 0x0
      12'h9F4: dout <= 8'b00000000; // 2548 :   0 - 0x0
      12'h9F5: dout <= 8'b00000000; // 2549 :   0 - 0x0
      12'h9F6: dout <= 8'b00000000; // 2550 :   0 - 0x0
      12'h9F7: dout <= 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- Background 0x3f
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout <= 8'b00000000; // 2560 :   0 - 0x0 -- Background 0x40
      12'hA01: dout <= 8'b00000000; // 2561 :   0 - 0x0
      12'hA02: dout <= 8'b00000000; // 2562 :   0 - 0x0
      12'hA03: dout <= 8'b00000000; // 2563 :   0 - 0x0
      12'hA04: dout <= 8'b00000000; // 2564 :   0 - 0x0
      12'hA05: dout <= 8'b00000000; // 2565 :   0 - 0x0
      12'hA06: dout <= 8'b00000000; // 2566 :   0 - 0x0
      12'hA07: dout <= 8'b00000000; // 2567 :   0 - 0x0
      12'hA08: dout <= 8'b00000000; // 2568 :   0 - 0x0 -- Background 0x41
      12'hA09: dout <= 8'b00000000; // 2569 :   0 - 0x0
      12'hA0A: dout <= 8'b00000000; // 2570 :   0 - 0x0
      12'hA0B: dout <= 8'b00000000; // 2571 :   0 - 0x0
      12'hA0C: dout <= 8'b00000000; // 2572 :   0 - 0x0
      12'hA0D: dout <= 8'b00000000; // 2573 :   0 - 0x0
      12'hA0E: dout <= 8'b00000000; // 2574 :   0 - 0x0
      12'hA0F: dout <= 8'b00000000; // 2575 :   0 - 0x0
      12'hA10: dout <= 8'b00000000; // 2576 :   0 - 0x0 -- Background 0x42
      12'hA11: dout <= 8'b00000000; // 2577 :   0 - 0x0
      12'hA12: dout <= 8'b00000000; // 2578 :   0 - 0x0
      12'hA13: dout <= 8'b00000000; // 2579 :   0 - 0x0
      12'hA14: dout <= 8'b00000000; // 2580 :   0 - 0x0
      12'hA15: dout <= 8'b00000000; // 2581 :   0 - 0x0
      12'hA16: dout <= 8'b00000000; // 2582 :   0 - 0x0
      12'hA17: dout <= 8'b00000000; // 2583 :   0 - 0x0
      12'hA18: dout <= 8'b00000000; // 2584 :   0 - 0x0 -- Background 0x43
      12'hA19: dout <= 8'b00000000; // 2585 :   0 - 0x0
      12'hA1A: dout <= 8'b00000000; // 2586 :   0 - 0x0
      12'hA1B: dout <= 8'b00000000; // 2587 :   0 - 0x0
      12'hA1C: dout <= 8'b00000000; // 2588 :   0 - 0x0
      12'hA1D: dout <= 8'b00000000; // 2589 :   0 - 0x0
      12'hA1E: dout <= 8'b00000000; // 2590 :   0 - 0x0
      12'hA1F: dout <= 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout <= 8'b00000000; // 2592 :   0 - 0x0 -- Background 0x44
      12'hA21: dout <= 8'b00000000; // 2593 :   0 - 0x0
      12'hA22: dout <= 8'b00000000; // 2594 :   0 - 0x0
      12'hA23: dout <= 8'b00000000; // 2595 :   0 - 0x0
      12'hA24: dout <= 8'b00000000; // 2596 :   0 - 0x0
      12'hA25: dout <= 8'b00000000; // 2597 :   0 - 0x0
      12'hA26: dout <= 8'b00000000; // 2598 :   0 - 0x0
      12'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0 -- Background 0x45
      12'hA29: dout <= 8'b00000000; // 2601 :   0 - 0x0
      12'hA2A: dout <= 8'b00000000; // 2602 :   0 - 0x0
      12'hA2B: dout <= 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout <= 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout <= 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout <= 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout <= 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout <= 8'b00000000; // 2608 :   0 - 0x0 -- Background 0x46
      12'hA31: dout <= 8'b00000000; // 2609 :   0 - 0x0
      12'hA32: dout <= 8'b00000000; // 2610 :   0 - 0x0
      12'hA33: dout <= 8'b00000000; // 2611 :   0 - 0x0
      12'hA34: dout <= 8'b00000000; // 2612 :   0 - 0x0
      12'hA35: dout <= 8'b00000000; // 2613 :   0 - 0x0
      12'hA36: dout <= 8'b00000000; // 2614 :   0 - 0x0
      12'hA37: dout <= 8'b00000000; // 2615 :   0 - 0x0
      12'hA38: dout <= 8'b00000000; // 2616 :   0 - 0x0 -- Background 0x47
      12'hA39: dout <= 8'b00000000; // 2617 :   0 - 0x0
      12'hA3A: dout <= 8'b00000000; // 2618 :   0 - 0x0
      12'hA3B: dout <= 8'b00000000; // 2619 :   0 - 0x0
      12'hA3C: dout <= 8'b00000000; // 2620 :   0 - 0x0
      12'hA3D: dout <= 8'b00000000; // 2621 :   0 - 0x0
      12'hA3E: dout <= 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout <= 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout <= 8'b00000000; // 2624 :   0 - 0x0 -- Background 0x48
      12'hA41: dout <= 8'b00000000; // 2625 :   0 - 0x0
      12'hA42: dout <= 8'b00000000; // 2626 :   0 - 0x0
      12'hA43: dout <= 8'b00000000; // 2627 :   0 - 0x0
      12'hA44: dout <= 8'b00000000; // 2628 :   0 - 0x0
      12'hA45: dout <= 8'b00000000; // 2629 :   0 - 0x0
      12'hA46: dout <= 8'b00000000; // 2630 :   0 - 0x0
      12'hA47: dout <= 8'b00000000; // 2631 :   0 - 0x0
      12'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0 -- Background 0x49
      12'hA49: dout <= 8'b00000000; // 2633 :   0 - 0x0
      12'hA4A: dout <= 8'b00000000; // 2634 :   0 - 0x0
      12'hA4B: dout <= 8'b00000000; // 2635 :   0 - 0x0
      12'hA4C: dout <= 8'b00000000; // 2636 :   0 - 0x0
      12'hA4D: dout <= 8'b00000000; // 2637 :   0 - 0x0
      12'hA4E: dout <= 8'b00000000; // 2638 :   0 - 0x0
      12'hA4F: dout <= 8'b00000000; // 2639 :   0 - 0x0
      12'hA50: dout <= 8'b00000000; // 2640 :   0 - 0x0 -- Background 0x4a
      12'hA51: dout <= 8'b00000000; // 2641 :   0 - 0x0
      12'hA52: dout <= 8'b00000000; // 2642 :   0 - 0x0
      12'hA53: dout <= 8'b00000000; // 2643 :   0 - 0x0
      12'hA54: dout <= 8'b00000000; // 2644 :   0 - 0x0
      12'hA55: dout <= 8'b00000000; // 2645 :   0 - 0x0
      12'hA56: dout <= 8'b00000000; // 2646 :   0 - 0x0
      12'hA57: dout <= 8'b00000000; // 2647 :   0 - 0x0
      12'hA58: dout <= 8'b00000000; // 2648 :   0 - 0x0 -- Background 0x4b
      12'hA59: dout <= 8'b00000000; // 2649 :   0 - 0x0
      12'hA5A: dout <= 8'b00000000; // 2650 :   0 - 0x0
      12'hA5B: dout <= 8'b00000000; // 2651 :   0 - 0x0
      12'hA5C: dout <= 8'b00000000; // 2652 :   0 - 0x0
      12'hA5D: dout <= 8'b00000000; // 2653 :   0 - 0x0
      12'hA5E: dout <= 8'b00000000; // 2654 :   0 - 0x0
      12'hA5F: dout <= 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout <= 8'b00000000; // 2656 :   0 - 0x0 -- Background 0x4c
      12'hA61: dout <= 8'b00000000; // 2657 :   0 - 0x0
      12'hA62: dout <= 8'b00000000; // 2658 :   0 - 0x0
      12'hA63: dout <= 8'b00000000; // 2659 :   0 - 0x0
      12'hA64: dout <= 8'b00000000; // 2660 :   0 - 0x0
      12'hA65: dout <= 8'b00000000; // 2661 :   0 - 0x0
      12'hA66: dout <= 8'b00000000; // 2662 :   0 - 0x0
      12'hA67: dout <= 8'b00000000; // 2663 :   0 - 0x0
      12'hA68: dout <= 8'b00000000; // 2664 :   0 - 0x0 -- Background 0x4d
      12'hA69: dout <= 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout <= 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout <= 8'b00000000; // 2667 :   0 - 0x0
      12'hA6C: dout <= 8'b00000000; // 2668 :   0 - 0x0
      12'hA6D: dout <= 8'b00000000; // 2669 :   0 - 0x0
      12'hA6E: dout <= 8'b00000000; // 2670 :   0 - 0x0
      12'hA6F: dout <= 8'b00000000; // 2671 :   0 - 0x0
      12'hA70: dout <= 8'b00000000; // 2672 :   0 - 0x0 -- Background 0x4e
      12'hA71: dout <= 8'b00000000; // 2673 :   0 - 0x0
      12'hA72: dout <= 8'b00000000; // 2674 :   0 - 0x0
      12'hA73: dout <= 8'b00000000; // 2675 :   0 - 0x0
      12'hA74: dout <= 8'b00000000; // 2676 :   0 - 0x0
      12'hA75: dout <= 8'b00000000; // 2677 :   0 - 0x0
      12'hA76: dout <= 8'b00000000; // 2678 :   0 - 0x0
      12'hA77: dout <= 8'b00000000; // 2679 :   0 - 0x0
      12'hA78: dout <= 8'b00000000; // 2680 :   0 - 0x0 -- Background 0x4f
      12'hA79: dout <= 8'b00000000; // 2681 :   0 - 0x0
      12'hA7A: dout <= 8'b00000000; // 2682 :   0 - 0x0
      12'hA7B: dout <= 8'b00000000; // 2683 :   0 - 0x0
      12'hA7C: dout <= 8'b00000000; // 2684 :   0 - 0x0
      12'hA7D: dout <= 8'b00000000; // 2685 :   0 - 0x0
      12'hA7E: dout <= 8'b00000000; // 2686 :   0 - 0x0
      12'hA7F: dout <= 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout <= 8'b00000000; // 2688 :   0 - 0x0 -- Background 0x50
      12'hA81: dout <= 8'b00000000; // 2689 :   0 - 0x0
      12'hA82: dout <= 8'b00000000; // 2690 :   0 - 0x0
      12'hA83: dout <= 8'b00000000; // 2691 :   0 - 0x0
      12'hA84: dout <= 8'b00000000; // 2692 :   0 - 0x0
      12'hA85: dout <= 8'b00000000; // 2693 :   0 - 0x0
      12'hA86: dout <= 8'b00000000; // 2694 :   0 - 0x0
      12'hA87: dout <= 8'b00000000; // 2695 :   0 - 0x0
      12'hA88: dout <= 8'b00000000; // 2696 :   0 - 0x0 -- Background 0x51
      12'hA89: dout <= 8'b00000000; // 2697 :   0 - 0x0
      12'hA8A: dout <= 8'b00000000; // 2698 :   0 - 0x0
      12'hA8B: dout <= 8'b00000000; // 2699 :   0 - 0x0
      12'hA8C: dout <= 8'b00000000; // 2700 :   0 - 0x0
      12'hA8D: dout <= 8'b00000000; // 2701 :   0 - 0x0
      12'hA8E: dout <= 8'b00000000; // 2702 :   0 - 0x0
      12'hA8F: dout <= 8'b00000000; // 2703 :   0 - 0x0
      12'hA90: dout <= 8'b00000000; // 2704 :   0 - 0x0 -- Background 0x52
      12'hA91: dout <= 8'b00000000; // 2705 :   0 - 0x0
      12'hA92: dout <= 8'b00000000; // 2706 :   0 - 0x0
      12'hA93: dout <= 8'b00000000; // 2707 :   0 - 0x0
      12'hA94: dout <= 8'b00000000; // 2708 :   0 - 0x0
      12'hA95: dout <= 8'b00000000; // 2709 :   0 - 0x0
      12'hA96: dout <= 8'b00000000; // 2710 :   0 - 0x0
      12'hA97: dout <= 8'b00000000; // 2711 :   0 - 0x0
      12'hA98: dout <= 8'b00000000; // 2712 :   0 - 0x0 -- Background 0x53
      12'hA99: dout <= 8'b00000000; // 2713 :   0 - 0x0
      12'hA9A: dout <= 8'b00000000; // 2714 :   0 - 0x0
      12'hA9B: dout <= 8'b00000000; // 2715 :   0 - 0x0
      12'hA9C: dout <= 8'b00000000; // 2716 :   0 - 0x0
      12'hA9D: dout <= 8'b00000000; // 2717 :   0 - 0x0
      12'hA9E: dout <= 8'b00000000; // 2718 :   0 - 0x0
      12'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout <= 8'b00000000; // 2720 :   0 - 0x0 -- Background 0x54
      12'hAA1: dout <= 8'b00000000; // 2721 :   0 - 0x0
      12'hAA2: dout <= 8'b00000000; // 2722 :   0 - 0x0
      12'hAA3: dout <= 8'b00000000; // 2723 :   0 - 0x0
      12'hAA4: dout <= 8'b00000000; // 2724 :   0 - 0x0
      12'hAA5: dout <= 8'b00000000; // 2725 :   0 - 0x0
      12'hAA6: dout <= 8'b00000000; // 2726 :   0 - 0x0
      12'hAA7: dout <= 8'b00000000; // 2727 :   0 - 0x0
      12'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0 -- Background 0x55
      12'hAA9: dout <= 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout <= 8'b00000000; // 2730 :   0 - 0x0
      12'hAAB: dout <= 8'b00000000; // 2731 :   0 - 0x0
      12'hAAC: dout <= 8'b00000000; // 2732 :   0 - 0x0
      12'hAAD: dout <= 8'b00000000; // 2733 :   0 - 0x0
      12'hAAE: dout <= 8'b00000000; // 2734 :   0 - 0x0
      12'hAAF: dout <= 8'b00000000; // 2735 :   0 - 0x0
      12'hAB0: dout <= 8'b00000000; // 2736 :   0 - 0x0 -- Background 0x56
      12'hAB1: dout <= 8'b00000000; // 2737 :   0 - 0x0
      12'hAB2: dout <= 8'b00000000; // 2738 :   0 - 0x0
      12'hAB3: dout <= 8'b00000000; // 2739 :   0 - 0x0
      12'hAB4: dout <= 8'b00000000; // 2740 :   0 - 0x0
      12'hAB5: dout <= 8'b00000000; // 2741 :   0 - 0x0
      12'hAB6: dout <= 8'b00000000; // 2742 :   0 - 0x0
      12'hAB7: dout <= 8'b00000000; // 2743 :   0 - 0x0
      12'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0 -- Background 0x57
      12'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout <= 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout <= 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout <= 8'b00000000; // 2752 :   0 - 0x0 -- Background 0x58
      12'hAC1: dout <= 8'b00000000; // 2753 :   0 - 0x0
      12'hAC2: dout <= 8'b00000000; // 2754 :   0 - 0x0
      12'hAC3: dout <= 8'b00000000; // 2755 :   0 - 0x0
      12'hAC4: dout <= 8'b00000000; // 2756 :   0 - 0x0
      12'hAC5: dout <= 8'b00000000; // 2757 :   0 - 0x0
      12'hAC6: dout <= 8'b00000000; // 2758 :   0 - 0x0
      12'hAC7: dout <= 8'b00000000; // 2759 :   0 - 0x0
      12'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0 -- Background 0x59
      12'hAC9: dout <= 8'b00000000; // 2761 :   0 - 0x0
      12'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout <= 8'b00000000; // 2763 :   0 - 0x0
      12'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      12'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout <= 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout <= 8'b00000000; // 2768 :   0 - 0x0 -- Background 0x5a
      12'hAD1: dout <= 8'b00000000; // 2769 :   0 - 0x0
      12'hAD2: dout <= 8'b00000000; // 2770 :   0 - 0x0
      12'hAD3: dout <= 8'b00000000; // 2771 :   0 - 0x0
      12'hAD4: dout <= 8'b00000000; // 2772 :   0 - 0x0
      12'hAD5: dout <= 8'b00000000; // 2773 :   0 - 0x0
      12'hAD6: dout <= 8'b00000000; // 2774 :   0 - 0x0
      12'hAD7: dout <= 8'b00000000; // 2775 :   0 - 0x0
      12'hAD8: dout <= 8'b00000000; // 2776 :   0 - 0x0 -- Background 0x5b
      12'hAD9: dout <= 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout <= 8'b00000000; // 2778 :   0 - 0x0
      12'hADB: dout <= 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout <= 8'b00000000; // 2780 :   0 - 0x0
      12'hADD: dout <= 8'b00000000; // 2781 :   0 - 0x0
      12'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      12'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout <= 8'b00000000; // 2784 :   0 - 0x0 -- Background 0x5c
      12'hAE1: dout <= 8'b00000000; // 2785 :   0 - 0x0
      12'hAE2: dout <= 8'b00000000; // 2786 :   0 - 0x0
      12'hAE3: dout <= 8'b00000000; // 2787 :   0 - 0x0
      12'hAE4: dout <= 8'b00000000; // 2788 :   0 - 0x0
      12'hAE5: dout <= 8'b00000000; // 2789 :   0 - 0x0
      12'hAE6: dout <= 8'b00000000; // 2790 :   0 - 0x0
      12'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0 -- Background 0x5d
      12'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout <= 8'b00000000; // 2794 :   0 - 0x0
      12'hAEB: dout <= 8'b00000000; // 2795 :   0 - 0x0
      12'hAEC: dout <= 8'b00000000; // 2796 :   0 - 0x0
      12'hAED: dout <= 8'b00000000; // 2797 :   0 - 0x0
      12'hAEE: dout <= 8'b00000000; // 2798 :   0 - 0x0
      12'hAEF: dout <= 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout <= 8'b00000000; // 2800 :   0 - 0x0 -- Background 0x5e
      12'hAF1: dout <= 8'b00000000; // 2801 :   0 - 0x0
      12'hAF2: dout <= 8'b00000000; // 2802 :   0 - 0x0
      12'hAF3: dout <= 8'b00000000; // 2803 :   0 - 0x0
      12'hAF4: dout <= 8'b00000000; // 2804 :   0 - 0x0
      12'hAF5: dout <= 8'b00000000; // 2805 :   0 - 0x0
      12'hAF6: dout <= 8'b00000000; // 2806 :   0 - 0x0
      12'hAF7: dout <= 8'b00000000; // 2807 :   0 - 0x0
      12'hAF8: dout <= 8'b00000000; // 2808 :   0 - 0x0 -- Background 0x5f
      12'hAF9: dout <= 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout <= 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout <= 8'b00000000; // 2811 :   0 - 0x0
      12'hAFC: dout <= 8'b00000000; // 2812 :   0 - 0x0
      12'hAFD: dout <= 8'b00000000; // 2813 :   0 - 0x0
      12'hAFE: dout <= 8'b00000000; // 2814 :   0 - 0x0
      12'hAFF: dout <= 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout <= 8'b00000000; // 2816 :   0 - 0x0 -- Background 0x60
      12'hB01: dout <= 8'b00000000; // 2817 :   0 - 0x0
      12'hB02: dout <= 8'b00000000; // 2818 :   0 - 0x0
      12'hB03: dout <= 8'b00000000; // 2819 :   0 - 0x0
      12'hB04: dout <= 8'b00000000; // 2820 :   0 - 0x0
      12'hB05: dout <= 8'b00000000; // 2821 :   0 - 0x0
      12'hB06: dout <= 8'b00000000; // 2822 :   0 - 0x0
      12'hB07: dout <= 8'b00000000; // 2823 :   0 - 0x0
      12'hB08: dout <= 8'b00000000; // 2824 :   0 - 0x0 -- Background 0x61
      12'hB09: dout <= 8'b00000000; // 2825 :   0 - 0x0
      12'hB0A: dout <= 8'b00000000; // 2826 :   0 - 0x0
      12'hB0B: dout <= 8'b00000000; // 2827 :   0 - 0x0
      12'hB0C: dout <= 8'b00000000; // 2828 :   0 - 0x0
      12'hB0D: dout <= 8'b00000000; // 2829 :   0 - 0x0
      12'hB0E: dout <= 8'b00000000; // 2830 :   0 - 0x0
      12'hB0F: dout <= 8'b00000000; // 2831 :   0 - 0x0
      12'hB10: dout <= 8'b00000000; // 2832 :   0 - 0x0 -- Background 0x62
      12'hB11: dout <= 8'b00000000; // 2833 :   0 - 0x0
      12'hB12: dout <= 8'b00000000; // 2834 :   0 - 0x0
      12'hB13: dout <= 8'b00000000; // 2835 :   0 - 0x0
      12'hB14: dout <= 8'b00000000; // 2836 :   0 - 0x0
      12'hB15: dout <= 8'b00000000; // 2837 :   0 - 0x0
      12'hB16: dout <= 8'b00000000; // 2838 :   0 - 0x0
      12'hB17: dout <= 8'b00000000; // 2839 :   0 - 0x0
      12'hB18: dout <= 8'b00000000; // 2840 :   0 - 0x0 -- Background 0x63
      12'hB19: dout <= 8'b00000000; // 2841 :   0 - 0x0
      12'hB1A: dout <= 8'b00000000; // 2842 :   0 - 0x0
      12'hB1B: dout <= 8'b00000000; // 2843 :   0 - 0x0
      12'hB1C: dout <= 8'b00000000; // 2844 :   0 - 0x0
      12'hB1D: dout <= 8'b00000000; // 2845 :   0 - 0x0
      12'hB1E: dout <= 8'b00000000; // 2846 :   0 - 0x0
      12'hB1F: dout <= 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout <= 8'b00000000; // 2848 :   0 - 0x0 -- Background 0x64
      12'hB21: dout <= 8'b00000000; // 2849 :   0 - 0x0
      12'hB22: dout <= 8'b00000000; // 2850 :   0 - 0x0
      12'hB23: dout <= 8'b00000000; // 2851 :   0 - 0x0
      12'hB24: dout <= 8'b00000000; // 2852 :   0 - 0x0
      12'hB25: dout <= 8'b00000000; // 2853 :   0 - 0x0
      12'hB26: dout <= 8'b00000000; // 2854 :   0 - 0x0
      12'hB27: dout <= 8'b00000000; // 2855 :   0 - 0x0
      12'hB28: dout <= 8'b00000000; // 2856 :   0 - 0x0 -- Background 0x65
      12'hB29: dout <= 8'b00000000; // 2857 :   0 - 0x0
      12'hB2A: dout <= 8'b00000000; // 2858 :   0 - 0x0
      12'hB2B: dout <= 8'b00000000; // 2859 :   0 - 0x0
      12'hB2C: dout <= 8'b00000000; // 2860 :   0 - 0x0
      12'hB2D: dout <= 8'b00000000; // 2861 :   0 - 0x0
      12'hB2E: dout <= 8'b00000000; // 2862 :   0 - 0x0
      12'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout <= 8'b00000000; // 2864 :   0 - 0x0 -- Background 0x66
      12'hB31: dout <= 8'b00000000; // 2865 :   0 - 0x0
      12'hB32: dout <= 8'b00000000; // 2866 :   0 - 0x0
      12'hB33: dout <= 8'b00000000; // 2867 :   0 - 0x0
      12'hB34: dout <= 8'b00000000; // 2868 :   0 - 0x0
      12'hB35: dout <= 8'b00000000; // 2869 :   0 - 0x0
      12'hB36: dout <= 8'b00000000; // 2870 :   0 - 0x0
      12'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      12'hB38: dout <= 8'b00000000; // 2872 :   0 - 0x0 -- Background 0x67
      12'hB39: dout <= 8'b00000000; // 2873 :   0 - 0x0
      12'hB3A: dout <= 8'b00000000; // 2874 :   0 - 0x0
      12'hB3B: dout <= 8'b00000000; // 2875 :   0 - 0x0
      12'hB3C: dout <= 8'b00000000; // 2876 :   0 - 0x0
      12'hB3D: dout <= 8'b00000000; // 2877 :   0 - 0x0
      12'hB3E: dout <= 8'b00000000; // 2878 :   0 - 0x0
      12'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout <= 8'b00000000; // 2880 :   0 - 0x0 -- Background 0x68
      12'hB41: dout <= 8'b00000000; // 2881 :   0 - 0x0
      12'hB42: dout <= 8'b00000000; // 2882 :   0 - 0x0
      12'hB43: dout <= 8'b00000000; // 2883 :   0 - 0x0
      12'hB44: dout <= 8'b00000000; // 2884 :   0 - 0x0
      12'hB45: dout <= 8'b00000000; // 2885 :   0 - 0x0
      12'hB46: dout <= 8'b00000000; // 2886 :   0 - 0x0
      12'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout <= 8'b00000000; // 2888 :   0 - 0x0 -- Background 0x69
      12'hB49: dout <= 8'b00000000; // 2889 :   0 - 0x0
      12'hB4A: dout <= 8'b00000000; // 2890 :   0 - 0x0
      12'hB4B: dout <= 8'b00000000; // 2891 :   0 - 0x0
      12'hB4C: dout <= 8'b00000000; // 2892 :   0 - 0x0
      12'hB4D: dout <= 8'b00000000; // 2893 :   0 - 0x0
      12'hB4E: dout <= 8'b00000000; // 2894 :   0 - 0x0
      12'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout <= 8'b00000000; // 2896 :   0 - 0x0 -- Background 0x6a
      12'hB51: dout <= 8'b00000000; // 2897 :   0 - 0x0
      12'hB52: dout <= 8'b00000000; // 2898 :   0 - 0x0
      12'hB53: dout <= 8'b00000000; // 2899 :   0 - 0x0
      12'hB54: dout <= 8'b00000000; // 2900 :   0 - 0x0
      12'hB55: dout <= 8'b00000000; // 2901 :   0 - 0x0
      12'hB56: dout <= 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout <= 8'b00000000; // 2904 :   0 - 0x0 -- Background 0x6b
      12'hB59: dout <= 8'b00000000; // 2905 :   0 - 0x0
      12'hB5A: dout <= 8'b00000000; // 2906 :   0 - 0x0
      12'hB5B: dout <= 8'b00000000; // 2907 :   0 - 0x0
      12'hB5C: dout <= 8'b00000000; // 2908 :   0 - 0x0
      12'hB5D: dout <= 8'b00000000; // 2909 :   0 - 0x0
      12'hB5E: dout <= 8'b00000000; // 2910 :   0 - 0x0
      12'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout <= 8'b00000000; // 2912 :   0 - 0x0 -- Background 0x6c
      12'hB61: dout <= 8'b00000000; // 2913 :   0 - 0x0
      12'hB62: dout <= 8'b00000000; // 2914 :   0 - 0x0
      12'hB63: dout <= 8'b00000000; // 2915 :   0 - 0x0
      12'hB64: dout <= 8'b00000000; // 2916 :   0 - 0x0
      12'hB65: dout <= 8'b00000000; // 2917 :   0 - 0x0
      12'hB66: dout <= 8'b00000000; // 2918 :   0 - 0x0
      12'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout <= 8'b00000000; // 2920 :   0 - 0x0 -- Background 0x6d
      12'hB69: dout <= 8'b00000000; // 2921 :   0 - 0x0
      12'hB6A: dout <= 8'b00000000; // 2922 :   0 - 0x0
      12'hB6B: dout <= 8'b00000000; // 2923 :   0 - 0x0
      12'hB6C: dout <= 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout <= 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout <= 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout <= 8'b00000000; // 2928 :   0 - 0x0 -- Background 0x6e
      12'hB71: dout <= 8'b00000000; // 2929 :   0 - 0x0
      12'hB72: dout <= 8'b00000000; // 2930 :   0 - 0x0
      12'hB73: dout <= 8'b00000000; // 2931 :   0 - 0x0
      12'hB74: dout <= 8'b00000000; // 2932 :   0 - 0x0
      12'hB75: dout <= 8'b00000000; // 2933 :   0 - 0x0
      12'hB76: dout <= 8'b00000000; // 2934 :   0 - 0x0
      12'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout <= 8'b00000000; // 2936 :   0 - 0x0 -- Background 0x6f
      12'hB79: dout <= 8'b00000000; // 2937 :   0 - 0x0
      12'hB7A: dout <= 8'b00000000; // 2938 :   0 - 0x0
      12'hB7B: dout <= 8'b00000000; // 2939 :   0 - 0x0
      12'hB7C: dout <= 8'b00000000; // 2940 :   0 - 0x0
      12'hB7D: dout <= 8'b00000000; // 2941 :   0 - 0x0
      12'hB7E: dout <= 8'b00000000; // 2942 :   0 - 0x0
      12'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout <= 8'b00000000; // 2944 :   0 - 0x0 -- Background 0x70
      12'hB81: dout <= 8'b00000000; // 2945 :   0 - 0x0
      12'hB82: dout <= 8'b00000000; // 2946 :   0 - 0x0
      12'hB83: dout <= 8'b00000000; // 2947 :   0 - 0x0
      12'hB84: dout <= 8'b00000000; // 2948 :   0 - 0x0
      12'hB85: dout <= 8'b00000000; // 2949 :   0 - 0x0
      12'hB86: dout <= 8'b00000000; // 2950 :   0 - 0x0
      12'hB87: dout <= 8'b00000000; // 2951 :   0 - 0x0
      12'hB88: dout <= 8'b00000000; // 2952 :   0 - 0x0 -- Background 0x71
      12'hB89: dout <= 8'b00000000; // 2953 :   0 - 0x0
      12'hB8A: dout <= 8'b00000000; // 2954 :   0 - 0x0
      12'hB8B: dout <= 8'b00000000; // 2955 :   0 - 0x0
      12'hB8C: dout <= 8'b00000000; // 2956 :   0 - 0x0
      12'hB8D: dout <= 8'b00000000; // 2957 :   0 - 0x0
      12'hB8E: dout <= 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b00000000; // 2960 :   0 - 0x0 -- Background 0x72
      12'hB91: dout <= 8'b00000000; // 2961 :   0 - 0x0
      12'hB92: dout <= 8'b00000000; // 2962 :   0 - 0x0
      12'hB93: dout <= 8'b00000000; // 2963 :   0 - 0x0
      12'hB94: dout <= 8'b00000000; // 2964 :   0 - 0x0
      12'hB95: dout <= 8'b00000000; // 2965 :   0 - 0x0
      12'hB96: dout <= 8'b00000000; // 2966 :   0 - 0x0
      12'hB97: dout <= 8'b00000000; // 2967 :   0 - 0x0
      12'hB98: dout <= 8'b00000000; // 2968 :   0 - 0x0 -- Background 0x73
      12'hB99: dout <= 8'b00000000; // 2969 :   0 - 0x0
      12'hB9A: dout <= 8'b00000000; // 2970 :   0 - 0x0
      12'hB9B: dout <= 8'b00000000; // 2971 :   0 - 0x0
      12'hB9C: dout <= 8'b00000000; // 2972 :   0 - 0x0
      12'hB9D: dout <= 8'b00000000; // 2973 :   0 - 0x0
      12'hB9E: dout <= 8'b00000000; // 2974 :   0 - 0x0
      12'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout <= 8'b00000000; // 2976 :   0 - 0x0 -- Background 0x74
      12'hBA1: dout <= 8'b00000000; // 2977 :   0 - 0x0
      12'hBA2: dout <= 8'b00000000; // 2978 :   0 - 0x0
      12'hBA3: dout <= 8'b00000000; // 2979 :   0 - 0x0
      12'hBA4: dout <= 8'b00000000; // 2980 :   0 - 0x0
      12'hBA5: dout <= 8'b00000000; // 2981 :   0 - 0x0
      12'hBA6: dout <= 8'b00000000; // 2982 :   0 - 0x0
      12'hBA7: dout <= 8'b00000000; // 2983 :   0 - 0x0
      12'hBA8: dout <= 8'b00000000; // 2984 :   0 - 0x0 -- Background 0x75
      12'hBA9: dout <= 8'b00000000; // 2985 :   0 - 0x0
      12'hBAA: dout <= 8'b00000000; // 2986 :   0 - 0x0
      12'hBAB: dout <= 8'b00000000; // 2987 :   0 - 0x0
      12'hBAC: dout <= 8'b00000000; // 2988 :   0 - 0x0
      12'hBAD: dout <= 8'b00000000; // 2989 :   0 - 0x0
      12'hBAE: dout <= 8'b00000000; // 2990 :   0 - 0x0
      12'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout <= 8'b00000000; // 2992 :   0 - 0x0 -- Background 0x76
      12'hBB1: dout <= 8'b00000000; // 2993 :   0 - 0x0
      12'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      12'hBB3: dout <= 8'b00000000; // 2995 :   0 - 0x0
      12'hBB4: dout <= 8'b00000000; // 2996 :   0 - 0x0
      12'hBB5: dout <= 8'b00000000; // 2997 :   0 - 0x0
      12'hBB6: dout <= 8'b00000000; // 2998 :   0 - 0x0
      12'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0 -- Background 0x77
      12'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      12'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      12'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      12'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      12'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b00000000; // 3008 :   0 - 0x0 -- Background 0x78
      12'hBC1: dout <= 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout <= 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout <= 8'b00000000; // 3011 :   0 - 0x0
      12'hBC4: dout <= 8'b00000000; // 3012 :   0 - 0x0
      12'hBC5: dout <= 8'b00000000; // 3013 :   0 - 0x0
      12'hBC6: dout <= 8'b00000000; // 3014 :   0 - 0x0
      12'hBC7: dout <= 8'b00000000; // 3015 :   0 - 0x0
      12'hBC8: dout <= 8'b00000000; // 3016 :   0 - 0x0 -- Background 0x79
      12'hBC9: dout <= 8'b00000000; // 3017 :   0 - 0x0
      12'hBCA: dout <= 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout <= 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout <= 8'b00000000; // 3021 :   0 - 0x0
      12'hBCE: dout <= 8'b00000000; // 3022 :   0 - 0x0
      12'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout <= 8'b00000000; // 3024 :   0 - 0x0 -- Background 0x7a
      12'hBD1: dout <= 8'b00000000; // 3025 :   0 - 0x0
      12'hBD2: dout <= 8'b00000000; // 3026 :   0 - 0x0
      12'hBD3: dout <= 8'b00000000; // 3027 :   0 - 0x0
      12'hBD4: dout <= 8'b00000000; // 3028 :   0 - 0x0
      12'hBD5: dout <= 8'b00000000; // 3029 :   0 - 0x0
      12'hBD6: dout <= 8'b00000000; // 3030 :   0 - 0x0
      12'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0 -- Background 0x7b
      12'hBD9: dout <= 8'b00000000; // 3033 :   0 - 0x0
      12'hBDA: dout <= 8'b00000000; // 3034 :   0 - 0x0
      12'hBDB: dout <= 8'b00000000; // 3035 :   0 - 0x0
      12'hBDC: dout <= 8'b00000000; // 3036 :   0 - 0x0
      12'hBDD: dout <= 8'b00000000; // 3037 :   0 - 0x0
      12'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout <= 8'b00000000; // 3040 :   0 - 0x0 -- Background 0x7c
      12'hBE1: dout <= 8'b00000000; // 3041 :   0 - 0x0
      12'hBE2: dout <= 8'b00000000; // 3042 :   0 - 0x0
      12'hBE3: dout <= 8'b00000000; // 3043 :   0 - 0x0
      12'hBE4: dout <= 8'b00000000; // 3044 :   0 - 0x0
      12'hBE5: dout <= 8'b00000000; // 3045 :   0 - 0x0
      12'hBE6: dout <= 8'b00000000; // 3046 :   0 - 0x0
      12'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      12'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0 -- Background 0x7d
      12'hBE9: dout <= 8'b00000000; // 3049 :   0 - 0x0
      12'hBEA: dout <= 8'b00000000; // 3050 :   0 - 0x0
      12'hBEB: dout <= 8'b00000000; // 3051 :   0 - 0x0
      12'hBEC: dout <= 8'b00000000; // 3052 :   0 - 0x0
      12'hBED: dout <= 8'b00000000; // 3053 :   0 - 0x0
      12'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      12'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Background 0x7e
      12'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      12'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      12'hBF4: dout <= 8'b00000000; // 3060 :   0 - 0x0
      12'hBF5: dout <= 8'b00000000; // 3061 :   0 - 0x0
      12'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      12'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0 -- Background 0x7f
      12'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      12'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      12'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      12'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout <= 8'b10111111; // 3072 : 191 - 0xbf -- Background 0x80
      12'hC01: dout <= 8'b11110111; // 3073 : 247 - 0xf7
      12'hC02: dout <= 8'b11111101; // 3074 : 253 - 0xfd
      12'hC03: dout <= 8'b11011111; // 3075 : 223 - 0xdf
      12'hC04: dout <= 8'b11111011; // 3076 : 251 - 0xfb
      12'hC05: dout <= 8'b10111111; // 3077 : 191 - 0xbf
      12'hC06: dout <= 8'b11111110; // 3078 : 254 - 0xfe
      12'hC07: dout <= 8'b11101111; // 3079 : 239 - 0xef
      12'hC08: dout <= 8'b11111111; // 3080 : 255 - 0xff -- Background 0x81
      12'hC09: dout <= 8'b11101110; // 3081 : 238 - 0xee
      12'hC0A: dout <= 8'b11111111; // 3082 : 255 - 0xff
      12'hC0B: dout <= 8'b11011111; // 3083 : 223 - 0xdf
      12'hC0C: dout <= 8'b01110111; // 3084 : 119 - 0x77
      12'hC0D: dout <= 8'b11111101; // 3085 : 253 - 0xfd
      12'hC0E: dout <= 8'b11011111; // 3086 : 223 - 0xdf
      12'hC0F: dout <= 8'b10111111; // 3087 : 191 - 0xbf
      12'hC10: dout <= 8'b11111110; // 3088 : 254 - 0xfe -- Background 0x82
      12'hC11: dout <= 8'b11101111; // 3089 : 239 - 0xef
      12'hC12: dout <= 8'b10111111; // 3090 : 191 - 0xbf
      12'hC13: dout <= 8'b11110111; // 3091 : 247 - 0xf7
      12'hC14: dout <= 8'b11111101; // 3092 : 253 - 0xfd
      12'hC15: dout <= 8'b11011111; // 3093 : 223 - 0xdf
      12'hC16: dout <= 8'b11111011; // 3094 : 251 - 0xfb
      12'hC17: dout <= 8'b10111111; // 3095 : 191 - 0xbf
      12'hC18: dout <= 8'b11101111; // 3096 : 239 - 0xef -- Background 0x83
      12'hC19: dout <= 8'b11111111; // 3097 : 255 - 0xff
      12'hC1A: dout <= 8'b10111011; // 3098 : 187 - 0xbb
      12'hC1B: dout <= 8'b11111111; // 3099 : 255 - 0xff
      12'hC1C: dout <= 8'b11110111; // 3100 : 247 - 0xf7
      12'hC1D: dout <= 8'b11011101; // 3101 : 221 - 0xdd
      12'hC1E: dout <= 8'b01111111; // 3102 : 127 - 0x7f
      12'hC1F: dout <= 8'b11110111; // 3103 : 247 - 0xf7
      12'hC20: dout <= 8'b11111111; // 3104 : 255 - 0xff -- Background 0x84
      12'hC21: dout <= 8'b11101110; // 3105 : 238 - 0xee
      12'hC22: dout <= 8'b11111011; // 3106 : 251 - 0xfb
      12'hC23: dout <= 8'b10111111; // 3107 : 191 - 0xbf
      12'hC24: dout <= 8'b01111111; // 3108 : 127 - 0x7f
      12'hC25: dout <= 8'b11101101; // 3109 : 237 - 0xed
      12'hC26: dout <= 8'b11111111; // 3110 : 255 - 0xff
      12'hC27: dout <= 8'b10111111; // 3111 : 191 - 0xbf
      12'hC28: dout <= 8'b11111111; // 3112 : 255 - 0xff -- Background 0x85
      12'hC29: dout <= 8'b10111111; // 3113 : 191 - 0xbf
      12'hC2A: dout <= 8'b01111101; // 3114 : 125 - 0x7d
      12'hC2B: dout <= 8'b11110111; // 3115 : 247 - 0xf7
      12'hC2C: dout <= 8'b11011011; // 3116 : 219 - 0xdb
      12'hC2D: dout <= 8'b11111101; // 3117 : 253 - 0xfd
      12'hC2E: dout <= 8'b01111110; // 3118 : 126 - 0x7e
      12'hC2F: dout <= 8'b11111011; // 3119 : 251 - 0xfb
      12'hC30: dout <= 8'b11111111; // 3120 : 255 - 0xff -- Background 0x86
      12'hC31: dout <= 8'b11110111; // 3121 : 247 - 0xf7
      12'hC32: dout <= 8'b11111111; // 3122 : 255 - 0xff
      12'hC33: dout <= 8'b11011101; // 3123 : 221 - 0xdd
      12'hC34: dout <= 8'b01111111; // 3124 : 127 - 0x7f
      12'hC35: dout <= 8'b11110111; // 3125 : 247 - 0xf7
      12'hC36: dout <= 8'b11101111; // 3126 : 239 - 0xef
      12'hC37: dout <= 8'b10111101; // 3127 : 189 - 0xbd
      12'hC38: dout <= 8'b01011111; // 3128 :  95 - 0x5f -- Background 0x87
      12'hC39: dout <= 8'b11111101; // 3129 : 253 - 0xfd
      12'hC3A: dout <= 8'b11110110; // 3130 : 246 - 0xf6
      12'hC3B: dout <= 8'b01111111; // 3131 : 127 - 0x7f
      12'hC3C: dout <= 8'b10011111; // 3132 : 159 - 0x9f
      12'hC3D: dout <= 8'b11111110; // 3133 : 254 - 0xfe
      12'hC3E: dout <= 8'b11111111; // 3134 : 255 - 0xff
      12'hC3F: dout <= 8'b11101111; // 3135 : 239 - 0xef
      12'hC40: dout <= 8'b11111111; // 3136 : 255 - 0xff -- Background 0x88
      12'hC41: dout <= 8'b10011111; // 3137 : 159 - 0x9f
      12'hC42: dout <= 8'b10111111; // 3138 : 191 - 0xbf
      12'hC43: dout <= 8'b11111111; // 3139 : 255 - 0xff
      12'hC44: dout <= 8'b11110011; // 3140 : 243 - 0xf3
      12'hC45: dout <= 8'b11110011; // 3141 : 243 - 0xf3
      12'hC46: dout <= 8'b11111111; // 3142 : 255 - 0xff
      12'hC47: dout <= 8'b11111111; // 3143 : 255 - 0xff
      12'hC48: dout <= 8'b11111111; // 3144 : 255 - 0xff -- Background 0x89
      12'hC49: dout <= 8'b10011111; // 3145 : 159 - 0x9f
      12'hC4A: dout <= 8'b10111111; // 3146 : 191 - 0xbf
      12'hC4B: dout <= 8'b11110011; // 3147 : 243 - 0xf3
      12'hC4C: dout <= 8'b11110011; // 3148 : 243 - 0xf3
      12'hC4D: dout <= 8'b11111111; // 3149 : 255 - 0xff
      12'hC4E: dout <= 8'b11111111; // 3150 : 255 - 0xff
      12'hC4F: dout <= 8'b11111111; // 3151 : 255 - 0xff
      12'hC50: dout <= 8'b10111111; // 3152 : 191 - 0xbf -- Background 0x8a
      12'hC51: dout <= 8'b11110111; // 3153 : 247 - 0xf7
      12'hC52: dout <= 8'b11111101; // 3154 : 253 - 0xfd
      12'hC53: dout <= 8'b11111111; // 3155 : 255 - 0xff
      12'hC54: dout <= 8'b11111011; // 3156 : 251 - 0xfb
      12'hC55: dout <= 8'b10111111; // 3157 : 191 - 0xbf
      12'hC56: dout <= 8'b11111110; // 3158 : 254 - 0xfe
      12'hC57: dout <= 8'b11101111; // 3159 : 239 - 0xef
      12'hC58: dout <= 8'b10111111; // 3160 : 191 - 0xbf -- Background 0x8b
      12'hC59: dout <= 8'b11111111; // 3161 : 255 - 0xff
      12'hC5A: dout <= 8'b11101110; // 3162 : 238 - 0xee
      12'hC5B: dout <= 8'b11111111; // 3163 : 255 - 0xff
      12'hC5C: dout <= 8'b11011111; // 3164 : 223 - 0xdf
      12'hC5D: dout <= 8'b01111101; // 3165 : 125 - 0x7d
      12'hC5E: dout <= 8'b11111111; // 3166 : 255 - 0xff
      12'hC5F: dout <= 8'b11011111; // 3167 : 223 - 0xdf
      12'hC60: dout <= 8'b11111111; // 3168 : 255 - 0xff -- Background 0x8c
      12'hC61: dout <= 8'b11111000; // 3169 : 248 - 0xf8
      12'hC62: dout <= 8'b11100010; // 3170 : 226 - 0xe2
      12'hC63: dout <= 8'b11010111; // 3171 : 215 - 0xd7
      12'hC64: dout <= 8'b11001111; // 3172 : 207 - 0xcf
      12'hC65: dout <= 8'b10011111; // 3173 : 159 - 0x9f
      12'hC66: dout <= 8'b10111110; // 3174 : 190 - 0xbe
      12'hC67: dout <= 8'b10011101; // 3175 : 157 - 0x9d
      12'hC68: dout <= 8'b11111111; // 3176 : 255 - 0xff -- Background 0x8d
      12'hC69: dout <= 8'b00011111; // 3177 :  31 - 0x1f
      12'hC6A: dout <= 8'b10100111; // 3178 : 167 - 0xa7
      12'hC6B: dout <= 8'b11000011; // 3179 : 195 - 0xc3
      12'hC6C: dout <= 8'b11100011; // 3180 : 227 - 0xe3
      12'hC6D: dout <= 8'b01000001; // 3181 :  65 - 0x41
      12'hC6E: dout <= 8'b10100001; // 3182 : 161 - 0xa1
      12'hC6F: dout <= 8'b00000001; // 3183 :   1 - 0x1
      12'hC70: dout <= 8'b10111110; // 3184 : 190 - 0xbe -- Background 0x8e
      12'hC71: dout <= 8'b11111111; // 3185 : 255 - 0xff
      12'hC72: dout <= 8'b11011111; // 3186 : 223 - 0xdf
      12'hC73: dout <= 8'b11111111; // 3187 : 255 - 0xff
      12'hC74: dout <= 8'b11101111; // 3188 : 239 - 0xef
      12'hC75: dout <= 8'b11111111; // 3189 : 255 - 0xff
      12'hC76: dout <= 8'b11110111; // 3190 : 247 - 0xf7
      12'hC77: dout <= 8'b11111111; // 3191 : 255 - 0xff
      12'hC78: dout <= 8'b01111101; // 3192 : 125 - 0x7d -- Background 0x8f
      12'hC79: dout <= 8'b11111111; // 3193 : 255 - 0xff
      12'hC7A: dout <= 8'b11111011; // 3194 : 251 - 0xfb
      12'hC7B: dout <= 8'b11111111; // 3195 : 255 - 0xff
      12'hC7C: dout <= 8'b11110111; // 3196 : 247 - 0xf7
      12'hC7D: dout <= 8'b11111111; // 3197 : 255 - 0xff
      12'hC7E: dout <= 8'b11101111; // 3198 : 239 - 0xef
      12'hC7F: dout <= 8'b11111111; // 3199 : 255 - 0xff
      12'hC80: dout <= 8'b10111110; // 3200 : 190 - 0xbe -- Background 0x90
      12'hC81: dout <= 8'b11110111; // 3201 : 247 - 0xf7
      12'hC82: dout <= 8'b11111111; // 3202 : 255 - 0xff
      12'hC83: dout <= 8'b11011111; // 3203 : 223 - 0xdf
      12'hC84: dout <= 8'b11111011; // 3204 : 251 - 0xfb
      12'hC85: dout <= 8'b11111110; // 3205 : 254 - 0xfe
      12'hC86: dout <= 8'b10111111; // 3206 : 191 - 0xbf
      12'hC87: dout <= 8'b11110111; // 3207 : 247 - 0xf7
      12'hC88: dout <= 8'b11101110; // 3208 : 238 - 0xee -- Background 0x91
      12'hC89: dout <= 8'b11111111; // 3209 : 255 - 0xff
      12'hC8A: dout <= 8'b01111011; // 3210 : 123 - 0x7b
      12'hC8B: dout <= 8'b11111101; // 3211 : 253 - 0xfd
      12'hC8C: dout <= 8'b11101111; // 3212 : 239 - 0xef
      12'hC8D: dout <= 8'b11111111; // 3213 : 255 - 0xff
      12'hC8E: dout <= 8'b10111101; // 3214 : 189 - 0xbd
      12'hC8F: dout <= 8'b11111111; // 3215 : 255 - 0xff
      12'hC90: dout <= 8'b11111011; // 3216 : 251 - 0xfb -- Background 0x92
      12'hC91: dout <= 8'b10111111; // 3217 : 191 - 0xbf
      12'hC92: dout <= 8'b11101111; // 3218 : 239 - 0xef
      12'hC93: dout <= 8'b11111101; // 3219 : 253 - 0xfd
      12'hC94: dout <= 8'b11111111; // 3220 : 255 - 0xff
      12'hC95: dout <= 8'b10111111; // 3221 : 191 - 0xbf
      12'hC96: dout <= 8'b11111011; // 3222 : 251 - 0xfb
      12'hC97: dout <= 8'b11011111; // 3223 : 223 - 0xdf
      12'hC98: dout <= 8'b10111101; // 3224 : 189 - 0xbd -- Background 0x93
      12'hC99: dout <= 8'b11111111; // 3225 : 255 - 0xff
      12'hC9A: dout <= 8'b01110111; // 3226 : 119 - 0x77
      12'hC9B: dout <= 8'b11111110; // 3227 : 254 - 0xfe
      12'hC9C: dout <= 8'b11011111; // 3228 : 223 - 0xdf
      12'hC9D: dout <= 8'b11111011; // 3229 : 251 - 0xfb
      12'hC9E: dout <= 8'b11101111; // 3230 : 239 - 0xef
      12'hC9F: dout <= 8'b01111111; // 3231 : 127 - 0x7f
      12'hCA0: dout <= 8'b01111111; // 3232 : 127 - 0x7f -- Background 0x94
      12'hCA1: dout <= 8'b11110111; // 3233 : 247 - 0xf7
      12'hCA2: dout <= 8'b11011101; // 3234 : 221 - 0xdd
      12'hCA3: dout <= 8'b01111011; // 3235 : 123 - 0x7b
      12'hCA4: dout <= 8'b11111111; // 3236 : 255 - 0xff
      12'hCA5: dout <= 8'b11101110; // 3237 : 238 - 0xee
      12'hCA6: dout <= 8'b10111011; // 3238 : 187 - 0xbb
      12'hCA7: dout <= 8'b11111101; // 3239 : 253 - 0xfd
      12'hCA8: dout <= 8'b11010111; // 3240 : 215 - 0xd7 -- Background 0x95
      12'hCA9: dout <= 8'b01111111; // 3241 : 127 - 0x7f
      12'hCAA: dout <= 8'b11111101; // 3242 : 253 - 0xfd
      12'hCAB: dout <= 8'b11101110; // 3243 : 238 - 0xee
      12'hCAC: dout <= 8'b11110111; // 3244 : 247 - 0xf7
      12'hCAD: dout <= 8'b10111011; // 3245 : 187 - 0xbb
      12'hCAE: dout <= 8'b11101111; // 3246 : 239 - 0xef
      12'hCAF: dout <= 8'b11110111; // 3247 : 247 - 0xf7
      12'hCB0: dout <= 8'b10111111; // 3248 : 191 - 0xbf -- Background 0x96
      12'hCB1: dout <= 8'b11101110; // 3249 : 238 - 0xee
      12'hCB2: dout <= 8'b11011011; // 3250 : 219 - 0xdb
      12'hCB3: dout <= 8'b11111111; // 3251 : 255 - 0xff
      12'hCB4: dout <= 8'b01110111; // 3252 : 119 - 0x77
      12'hCB5: dout <= 8'b11011101; // 3253 : 221 - 0xdd
      12'hCB6: dout <= 8'b11101111; // 3254 : 239 - 0xef
      12'hCB7: dout <= 8'b11111011; // 3255 : 251 - 0xfb
      12'hCB8: dout <= 8'b11111101; // 3256 : 253 - 0xfd -- Background 0x97
      12'hCB9: dout <= 8'b11101110; // 3257 : 238 - 0xee
      12'hCBA: dout <= 8'b11111011; // 3258 : 251 - 0xfb
      12'hCBB: dout <= 8'b11111101; // 3259 : 253 - 0xfd
      12'hCBC: dout <= 8'b11110101; // 3260 : 245 - 0xf5
      12'hCBD: dout <= 8'b11011111; // 3261 : 223 - 0xdf
      12'hCBE: dout <= 8'b01111111; // 3262 : 127 - 0x7f
      12'hCBF: dout <= 8'b10111011; // 3263 : 187 - 0xbb
      12'hCC0: dout <= 8'b11111111; // 3264 : 255 - 0xff -- Background 0x98
      12'hCC1: dout <= 8'b10011111; // 3265 : 159 - 0x9f
      12'hCC2: dout <= 8'b10111111; // 3266 : 191 - 0xbf
      12'hCC3: dout <= 8'b11110011; // 3267 : 243 - 0xf3
      12'hCC4: dout <= 8'b11110011; // 3268 : 243 - 0xf3
      12'hCC5: dout <= 8'b11111111; // 3269 : 255 - 0xff
      12'hCC6: dout <= 8'b11111111; // 3270 : 255 - 0xff
      12'hCC7: dout <= 8'b11111111; // 3271 : 255 - 0xff
      12'hCC8: dout <= 8'b11111111; // 3272 : 255 - 0xff -- Background 0x99
      12'hCC9: dout <= 8'b10011111; // 3273 : 159 - 0x9f
      12'hCCA: dout <= 8'b10111111; // 3274 : 191 - 0xbf
      12'hCCB: dout <= 8'b11111111; // 3275 : 255 - 0xff
      12'hCCC: dout <= 8'b11110011; // 3276 : 243 - 0xf3
      12'hCCD: dout <= 8'b11110011; // 3277 : 243 - 0xf3
      12'hCCE: dout <= 8'b11111111; // 3278 : 255 - 0xff
      12'hCCF: dout <= 8'b11111111; // 3279 : 255 - 0xff
      12'hCD0: dout <= 8'b10111111; // 3280 : 191 - 0xbf -- Background 0x9a
      12'hCD1: dout <= 8'b11110111; // 3281 : 247 - 0xf7
      12'hCD2: dout <= 8'b11111111; // 3282 : 255 - 0xff
      12'hCD3: dout <= 8'b11011111; // 3283 : 223 - 0xdf
      12'hCD4: dout <= 8'b11111011; // 3284 : 251 - 0xfb
      12'hCD5: dout <= 8'b11111111; // 3285 : 255 - 0xff
      12'hCD6: dout <= 8'b10111111; // 3286 : 191 - 0xbf
      12'hCD7: dout <= 8'b11110111; // 3287 : 247 - 0xf7
      12'hCD8: dout <= 8'b11011111; // 3288 : 223 - 0xdf -- Background 0x9b
      12'hCD9: dout <= 8'b11111111; // 3289 : 255 - 0xff
      12'hCDA: dout <= 8'b01111011; // 3290 : 123 - 0x7b
      12'hCDB: dout <= 8'b11111111; // 3291 : 255 - 0xff
      12'hCDC: dout <= 8'b11101111; // 3292 : 239 - 0xef
      12'hCDD: dout <= 8'b11111101; // 3293 : 253 - 0xfd
      12'hCDE: dout <= 8'b10111111; // 3294 : 191 - 0xbf
      12'hCDF: dout <= 8'b11111111; // 3295 : 255 - 0xff
      12'hCE0: dout <= 8'b10111010; // 3296 : 186 - 0xba -- Background 0x9c
      12'hCE1: dout <= 8'b10011100; // 3297 : 156 - 0x9c
      12'hCE2: dout <= 8'b10101010; // 3298 : 170 - 0xaa
      12'hCE3: dout <= 8'b11000000; // 3299 : 192 - 0xc0
      12'hCE4: dout <= 8'b11000000; // 3300 : 192 - 0xc0
      12'hCE5: dout <= 8'b11100000; // 3301 : 224 - 0xe0
      12'hCE6: dout <= 8'b11111000; // 3302 : 248 - 0xf8
      12'hCE7: dout <= 8'b11111111; // 3303 : 255 - 0xff
      12'hCE8: dout <= 8'b00000001; // 3304 :   1 - 0x1 -- Background 0x9d
      12'hCE9: dout <= 8'b00000001; // 3305 :   1 - 0x1
      12'hCEA: dout <= 8'b00000001; // 3306 :   1 - 0x1
      12'hCEB: dout <= 8'b00000011; // 3307 :   3 - 0x3
      12'hCEC: dout <= 8'b00000011; // 3308 :   3 - 0x3
      12'hCED: dout <= 8'b00000111; // 3309 :   7 - 0x7
      12'hCEE: dout <= 8'b00011111; // 3310 :  31 - 0x1f
      12'hCEF: dout <= 8'b11111111; // 3311 : 255 - 0xff
      12'hCF0: dout <= 8'b01111101; // 3312 : 125 - 0x7d -- Background 0x9e
      12'hCF1: dout <= 8'b11111111; // 3313 : 255 - 0xff
      12'hCF2: dout <= 8'b11111011; // 3314 : 251 - 0xfb
      12'hCF3: dout <= 8'b11111111; // 3315 : 255 - 0xff
      12'hCF4: dout <= 8'b11111111; // 3316 : 255 - 0xff
      12'hCF5: dout <= 8'b11111011; // 3317 : 251 - 0xfb
      12'hCF6: dout <= 8'b11111111; // 3318 : 255 - 0xff
      12'hCF7: dout <= 8'b01111101; // 3319 : 125 - 0x7d
      12'hCF8: dout <= 8'b11111111; // 3320 : 255 - 0xff -- Background 0x9f
      12'hCF9: dout <= 8'b11111111; // 3321 : 255 - 0xff
      12'hCFA: dout <= 8'b10111101; // 3322 : 189 - 0xbd
      12'hCFB: dout <= 8'b11111111; // 3323 : 255 - 0xff
      12'hCFC: dout <= 8'b11111111; // 3324 : 255 - 0xff
      12'hCFD: dout <= 8'b11111111; // 3325 : 255 - 0xff
      12'hCFE: dout <= 8'b11111111; // 3326 : 255 - 0xff
      12'hCFF: dout <= 8'b10111101; // 3327 : 189 - 0xbd
      12'hD00: dout <= 8'b11101111; // 3328 : 239 - 0xef -- Background 0xa0
      12'hD01: dout <= 8'b11000111; // 3329 : 199 - 0xc7
      12'hD02: dout <= 8'b10000011; // 3330 : 131 - 0x83
      12'hD03: dout <= 8'b00000111; // 3331 :   7 - 0x7
      12'hD04: dout <= 8'b10001111; // 3332 : 143 - 0x8f
      12'hD05: dout <= 8'b11011101; // 3333 : 221 - 0xdd
      12'hD06: dout <= 8'b11111010; // 3334 : 250 - 0xfa
      12'hD07: dout <= 8'b11111101; // 3335 : 253 - 0xfd
      12'hD08: dout <= 8'b11101111; // 3336 : 239 - 0xef -- Background 0xa1
      12'hD09: dout <= 8'b11000111; // 3337 : 199 - 0xc7
      12'hD0A: dout <= 8'b10000011; // 3338 : 131 - 0x83
      12'hD0B: dout <= 8'b00011111; // 3339 :  31 - 0x1f
      12'hD0C: dout <= 8'b10010000; // 3340 : 144 - 0x90
      12'hD0D: dout <= 8'b11010100; // 3341 : 212 - 0xd4
      12'hD0E: dout <= 8'b11110011; // 3342 : 243 - 0xf3
      12'hD0F: dout <= 8'b11110010; // 3343 : 242 - 0xf2
      12'hD10: dout <= 8'b11101111; // 3344 : 239 - 0xef -- Background 0xa2
      12'hD11: dout <= 8'b11000111; // 3345 : 199 - 0xc7
      12'hD12: dout <= 8'b10000011; // 3346 : 131 - 0x83
      12'hD13: dout <= 8'b11111111; // 3347 : 255 - 0xff
      12'hD14: dout <= 8'b00000000; // 3348 :   0 - 0x0
      12'hD15: dout <= 8'b00000000; // 3349 :   0 - 0x0
      12'hD16: dout <= 8'b01010101; // 3350 :  85 - 0x55
      12'hD17: dout <= 8'b00000000; // 3351 :   0 - 0x0
      12'hD18: dout <= 8'b11110000; // 3352 : 240 - 0xf0 -- Background 0xa3
      12'hD19: dout <= 8'b11010010; // 3353 : 210 - 0xd2
      12'hD1A: dout <= 8'b10010000; // 3354 : 144 - 0x90
      12'hD1B: dout <= 8'b00010010; // 3355 :  18 - 0x12
      12'hD1C: dout <= 8'b10010000; // 3356 : 144 - 0x90
      12'hD1D: dout <= 8'b11010010; // 3357 : 210 - 0xd2
      12'hD1E: dout <= 8'b11110000; // 3358 : 240 - 0xf0
      12'hD1F: dout <= 8'b11110010; // 3359 : 242 - 0xf2
      12'hD20: dout <= 8'b11110000; // 3360 : 240 - 0xf0 -- Background 0xa4
      12'hD21: dout <= 8'b11010011; // 3361 : 211 - 0xd3
      12'hD22: dout <= 8'b10010100; // 3362 : 148 - 0x94
      12'hD23: dout <= 8'b00011000; // 3363 :  24 - 0x18
      12'hD24: dout <= 8'b10011111; // 3364 : 159 - 0x9f
      12'hD25: dout <= 8'b11011101; // 3365 : 221 - 0xdd
      12'hD26: dout <= 8'b11111010; // 3366 : 250 - 0xfa
      12'hD27: dout <= 8'b11111101; // 3367 : 253 - 0xfd
      12'hD28: dout <= 8'b00000000; // 3368 :   0 - 0x0 -- Background 0xa5
      12'hD29: dout <= 8'b11111111; // 3369 : 255 - 0xff
      12'hD2A: dout <= 8'b00000000; // 3370 :   0 - 0x0
      12'hD2B: dout <= 8'b00000000; // 3371 :   0 - 0x0
      12'hD2C: dout <= 8'b11111111; // 3372 : 255 - 0xff
      12'hD2D: dout <= 8'b11011101; // 3373 : 221 - 0xdd
      12'hD2E: dout <= 8'b11111010; // 3374 : 250 - 0xfa
      12'hD2F: dout <= 8'b11111101; // 3375 : 253 - 0xfd
      12'hD30: dout <= 8'b11101111; // 3376 : 239 - 0xef -- Background 0xa6
      12'hD31: dout <= 8'b11000111; // 3377 : 199 - 0xc7
      12'hD32: dout <= 8'b10000011; // 3378 : 131 - 0x83
      12'hD33: dout <= 8'b11111111; // 3379 : 255 - 0xff
      12'hD34: dout <= 8'b00011111; // 3380 :  31 - 0x1f
      12'hD35: dout <= 8'b00101101; // 3381 :  45 - 0x2d
      12'hD36: dout <= 8'b01001010; // 3382 :  74 - 0x4a
      12'hD37: dout <= 8'b01001101; // 3383 :  77 - 0x4d
      12'hD38: dout <= 8'b01001111; // 3384 :  79 - 0x4f -- Background 0xa7
      12'hD39: dout <= 8'b01001111; // 3385 :  79 - 0x4f
      12'hD3A: dout <= 8'b01001011; // 3386 :  75 - 0x4b
      12'hD3B: dout <= 8'b01001111; // 3387 :  79 - 0x4f
      12'hD3C: dout <= 8'b01001111; // 3388 :  79 - 0x4f
      12'hD3D: dout <= 8'b01001101; // 3389 :  77 - 0x4d
      12'hD3E: dout <= 8'b01001010; // 3390 :  74 - 0x4a
      12'hD3F: dout <= 8'b01001101; // 3391 :  77 - 0x4d
      12'hD40: dout <= 8'b01001111; // 3392 :  79 - 0x4f -- Background 0xa8
      12'hD41: dout <= 8'b11001111; // 3393 : 207 - 0xcf
      12'hD42: dout <= 8'b00001011; // 3394 :  11 - 0xb
      12'hD43: dout <= 8'b00001111; // 3395 :  15 - 0xf
      12'hD44: dout <= 8'b11111111; // 3396 : 255 - 0xff
      12'hD45: dout <= 8'b11011101; // 3397 : 221 - 0xdd
      12'hD46: dout <= 8'b11111010; // 3398 : 250 - 0xfa
      12'hD47: dout <= 8'b11111101; // 3399 : 253 - 0xfd
      12'hD48: dout <= 8'b11111111; // 3400 : 255 - 0xff -- Background 0xa9
      12'hD49: dout <= 8'b11111111; // 3401 : 255 - 0xff
      12'hD4A: dout <= 8'b11111111; // 3402 : 255 - 0xff
      12'hD4B: dout <= 8'b11111111; // 3403 : 255 - 0xff
      12'hD4C: dout <= 8'b11111111; // 3404 : 255 - 0xff
      12'hD4D: dout <= 8'b11111111; // 3405 : 255 - 0xff
      12'hD4E: dout <= 8'b11111111; // 3406 : 255 - 0xff
      12'hD4F: dout <= 8'b11111111; // 3407 : 255 - 0xff
      12'hD50: dout <= 8'b11111111; // 3408 : 255 - 0xff -- Background 0xaa
      12'hD51: dout <= 8'b11111111; // 3409 : 255 - 0xff
      12'hD52: dout <= 8'b10101111; // 3410 : 175 - 0xaf
      12'hD53: dout <= 8'b01010111; // 3411 :  87 - 0x57
      12'hD54: dout <= 8'b10001111; // 3412 : 143 - 0x8f
      12'hD55: dout <= 8'b11011101; // 3413 : 221 - 0xdd
      12'hD56: dout <= 8'b11111010; // 3414 : 250 - 0xfa
      12'hD57: dout <= 8'b11111101; // 3415 : 253 - 0xfd
      12'hD58: dout <= 8'b11111111; // 3416 : 255 - 0xff -- Background 0xab
      12'hD59: dout <= 8'b00000000; // 3417 :   0 - 0x0
      12'hD5A: dout <= 8'b00000000; // 3418 :   0 - 0x0
      12'hD5B: dout <= 8'b00000000; // 3419 :   0 - 0x0
      12'hD5C: dout <= 8'b00000000; // 3420 :   0 - 0x0
      12'hD5D: dout <= 8'b00000000; // 3421 :   0 - 0x0
      12'hD5E: dout <= 8'b00000000; // 3422 :   0 - 0x0
      12'hD5F: dout <= 8'b00000000; // 3423 :   0 - 0x0
      12'hD60: dout <= 8'b00000000; // 3424 :   0 - 0x0 -- Background 0xac
      12'hD61: dout <= 8'b00000000; // 3425 :   0 - 0x0
      12'hD62: dout <= 8'b00000000; // 3426 :   0 - 0x0
      12'hD63: dout <= 8'b00000000; // 3427 :   0 - 0x0
      12'hD64: dout <= 8'b00000000; // 3428 :   0 - 0x0
      12'hD65: dout <= 8'b00000000; // 3429 :   0 - 0x0
      12'hD66: dout <= 8'b00000000; // 3430 :   0 - 0x0
      12'hD67: dout <= 8'b00000000; // 3431 :   0 - 0x0
      12'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0 -- Background 0xad
      12'hD69: dout <= 8'b11111111; // 3433 : 255 - 0xff
      12'hD6A: dout <= 8'b00000000; // 3434 :   0 - 0x0
      12'hD6B: dout <= 8'b11111111; // 3435 : 255 - 0xff
      12'hD6C: dout <= 8'b11111111; // 3436 : 255 - 0xff
      12'hD6D: dout <= 8'b11111111; // 3437 : 255 - 0xff
      12'hD6E: dout <= 8'b11111111; // 3438 : 255 - 0xff
      12'hD6F: dout <= 8'b11111111; // 3439 : 255 - 0xff
      12'hD70: dout <= 8'b11111111; // 3440 : 255 - 0xff -- Background 0xae
      12'hD71: dout <= 8'b11111111; // 3441 : 255 - 0xff
      12'hD72: dout <= 8'b11111111; // 3442 : 255 - 0xff
      12'hD73: dout <= 8'b11111111; // 3443 : 255 - 0xff
      12'hD74: dout <= 8'b11111111; // 3444 : 255 - 0xff
      12'hD75: dout <= 8'b00000000; // 3445 :   0 - 0x0
      12'hD76: dout <= 8'b11111111; // 3446 : 255 - 0xff
      12'hD77: dout <= 8'b00000000; // 3447 :   0 - 0x0
      12'hD78: dout <= 8'b11111111; // 3448 : 255 - 0xff -- Background 0xaf
      12'hD79: dout <= 8'b11111111; // 3449 : 255 - 0xff
      12'hD7A: dout <= 8'b11111111; // 3450 : 255 - 0xff
      12'hD7B: dout <= 8'b11111111; // 3451 : 255 - 0xff
      12'hD7C: dout <= 8'b11111111; // 3452 : 255 - 0xff
      12'hD7D: dout <= 8'b11111111; // 3453 : 255 - 0xff
      12'hD7E: dout <= 8'b11111111; // 3454 : 255 - 0xff
      12'hD7F: dout <= 8'b11111111; // 3455 : 255 - 0xff
      12'hD80: dout <= 8'b00000000; // 3456 :   0 - 0x0 -- Background 0xb0
      12'hD81: dout <= 8'b00000000; // 3457 :   0 - 0x0
      12'hD82: dout <= 8'b00011111; // 3458 :  31 - 0x1f
      12'hD83: dout <= 8'b00010000; // 3459 :  16 - 0x10
      12'hD84: dout <= 8'b00010000; // 3460 :  16 - 0x10
      12'hD85: dout <= 8'b00010000; // 3461 :  16 - 0x10
      12'hD86: dout <= 8'b00010000; // 3462 :  16 - 0x10
      12'hD87: dout <= 8'b00010000; // 3463 :  16 - 0x10
      12'hD88: dout <= 8'b00000000; // 3464 :   0 - 0x0 -- Background 0xb1
      12'hD89: dout <= 8'b00000000; // 3465 :   0 - 0x0
      12'hD8A: dout <= 8'b11111000; // 3466 : 248 - 0xf8
      12'hD8B: dout <= 8'b00001000; // 3467 :   8 - 0x8
      12'hD8C: dout <= 8'b00001000; // 3468 :   8 - 0x8
      12'hD8D: dout <= 8'b00001000; // 3469 :   8 - 0x8
      12'hD8E: dout <= 8'b00001000; // 3470 :   8 - 0x8
      12'hD8F: dout <= 8'b00001000; // 3471 :   8 - 0x8
      12'hD90: dout <= 8'b00010000; // 3472 :  16 - 0x10 -- Background 0xb2
      12'hD91: dout <= 8'b00010000; // 3473 :  16 - 0x10
      12'hD92: dout <= 8'b00010000; // 3474 :  16 - 0x10
      12'hD93: dout <= 8'b00010000; // 3475 :  16 - 0x10
      12'hD94: dout <= 8'b00010000; // 3476 :  16 - 0x10
      12'hD95: dout <= 8'b00011111; // 3477 :  31 - 0x1f
      12'hD96: dout <= 8'b00011111; // 3478 :  31 - 0x1f
      12'hD97: dout <= 8'b00001111; // 3479 :  15 - 0xf
      12'hD98: dout <= 8'b00001000; // 3480 :   8 - 0x8 -- Background 0xb3
      12'hD99: dout <= 8'b00001000; // 3481 :   8 - 0x8
      12'hD9A: dout <= 8'b00001000; // 3482 :   8 - 0x8
      12'hD9B: dout <= 8'b00001000; // 3483 :   8 - 0x8
      12'hD9C: dout <= 8'b00001000; // 3484 :   8 - 0x8
      12'hD9D: dout <= 8'b11111000; // 3485 : 248 - 0xf8
      12'hD9E: dout <= 8'b11111000; // 3486 : 248 - 0xf8
      12'hD9F: dout <= 8'b11110000; // 3487 : 240 - 0xf0
      12'hDA0: dout <= 8'b00000000; // 3488 :   0 - 0x0 -- Background 0xb4
      12'hDA1: dout <= 8'b00000000; // 3489 :   0 - 0x0
      12'hDA2: dout <= 8'b00000000; // 3490 :   0 - 0x0
      12'hDA3: dout <= 8'b00111111; // 3491 :  63 - 0x3f
      12'hDA4: dout <= 8'b01100000; // 3492 :  96 - 0x60
      12'hDA5: dout <= 8'b01100000; // 3493 :  96 - 0x60
      12'hDA6: dout <= 8'b01100000; // 3494 :  96 - 0x60
      12'hDA7: dout <= 8'b01100000; // 3495 :  96 - 0x60
      12'hDA8: dout <= 8'b00000000; // 3496 :   0 - 0x0 -- Background 0xb5
      12'hDA9: dout <= 8'b00000000; // 3497 :   0 - 0x0
      12'hDAA: dout <= 8'b00000000; // 3498 :   0 - 0x0
      12'hDAB: dout <= 8'b11111100; // 3499 : 252 - 0xfc
      12'hDAC: dout <= 8'b00000110; // 3500 :   6 - 0x6
      12'hDAD: dout <= 8'b00000110; // 3501 :   6 - 0x6
      12'hDAE: dout <= 8'b00000110; // 3502 :   6 - 0x6
      12'hDAF: dout <= 8'b00000110; // 3503 :   6 - 0x6
      12'hDB0: dout <= 8'b01100000; // 3504 :  96 - 0x60 -- Background 0xb6
      12'hDB1: dout <= 8'b01100000; // 3505 :  96 - 0x60
      12'hDB2: dout <= 8'b01100000; // 3506 :  96 - 0x60
      12'hDB3: dout <= 8'b01100000; // 3507 :  96 - 0x60
      12'hDB4: dout <= 8'b01111111; // 3508 : 127 - 0x7f
      12'hDB5: dout <= 8'b01111111; // 3509 : 127 - 0x7f
      12'hDB6: dout <= 8'b00111111; // 3510 :  63 - 0x3f
      12'hDB7: dout <= 8'b00000000; // 3511 :   0 - 0x0
      12'hDB8: dout <= 8'b00000110; // 3512 :   6 - 0x6 -- Background 0xb7
      12'hDB9: dout <= 8'b00000110; // 3513 :   6 - 0x6
      12'hDBA: dout <= 8'b00000110; // 3514 :   6 - 0x6
      12'hDBB: dout <= 8'b00000110; // 3515 :   6 - 0x6
      12'hDBC: dout <= 8'b11111110; // 3516 : 254 - 0xfe
      12'hDBD: dout <= 8'b11111110; // 3517 : 254 - 0xfe
      12'hDBE: dout <= 8'b11111100; // 3518 : 252 - 0xfc
      12'hDBF: dout <= 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout <= 8'b01100000; // 3520 :  96 - 0x60 -- Background 0xb8
      12'hDC1: dout <= 8'b11110000; // 3521 : 240 - 0xf0
      12'hDC2: dout <= 8'b11000011; // 3522 : 195 - 0xc3
      12'hDC3: dout <= 8'b10000111; // 3523 : 135 - 0x87
      12'hDC4: dout <= 8'b00000110; // 3524 :   6 - 0x6
      12'hDC5: dout <= 8'b00000100; // 3525 :   4 - 0x4
      12'hDC6: dout <= 8'b00000100; // 3526 :   4 - 0x4
      12'hDC7: dout <= 8'b00000111; // 3527 :   7 - 0x7
      12'hDC8: dout <= 8'b00000110; // 3528 :   6 - 0x6 -- Background 0xb9
      12'hDC9: dout <= 8'b00001111; // 3529 :  15 - 0xf
      12'hDCA: dout <= 8'b10000111; // 3530 : 135 - 0x87
      12'hDCB: dout <= 8'b11000001; // 3531 : 193 - 0xc1
      12'hDCC: dout <= 8'b00100011; // 3532 :  35 - 0x23
      12'hDCD: dout <= 8'b00101110; // 3533 :  46 - 0x2e
      12'hDCE: dout <= 8'b01100000; // 3534 :  96 - 0x60
      12'hDCF: dout <= 8'b11100001; // 3535 : 225 - 0xe1
      12'hDD0: dout <= 8'b00000000; // 3536 :   0 - 0x0 -- Background 0xba
      12'hDD1: dout <= 8'b11001000; // 3537 : 200 - 0xc8
      12'hDD2: dout <= 8'b11111000; // 3538 : 248 - 0xf8
      12'hDD3: dout <= 8'b10110000; // 3539 : 176 - 0xb0
      12'hDD4: dout <= 8'b00010000; // 3540 :  16 - 0x10
      12'hDD5: dout <= 8'b00110000; // 3541 :  48 - 0x30
      12'hDD6: dout <= 8'b11001000; // 3542 : 200 - 0xc8
      12'hDD7: dout <= 8'b11111000; // 3543 : 248 - 0xf8
      12'hDD8: dout <= 8'b00000111; // 3544 :   7 - 0x7 -- Background 0xbb
      12'hDD9: dout <= 8'b00000011; // 3545 :   3 - 0x3
      12'hDDA: dout <= 8'b00000000; // 3546 :   0 - 0x0
      12'hDDB: dout <= 8'b01100000; // 3547 :  96 - 0x60
      12'hDDC: dout <= 8'b11110000; // 3548 : 240 - 0xf0
      12'hDDD: dout <= 8'b11010000; // 3549 : 208 - 0xd0
      12'hDDE: dout <= 8'b10010000; // 3550 : 144 - 0x90
      12'hDDF: dout <= 8'b01100000; // 3551 :  96 - 0x60
      12'hDE0: dout <= 8'b11100001; // 3552 : 225 - 0xe1 -- Background 0xbc
      12'hDE1: dout <= 8'b11000011; // 3553 : 195 - 0xc3
      12'hDE2: dout <= 8'b00001110; // 3554 :  14 - 0xe
      12'hDE3: dout <= 8'b00000110; // 3555 :   6 - 0x6
      12'hDE4: dout <= 8'b00001111; // 3556 :  15 - 0xf
      12'hDE5: dout <= 8'b00001101; // 3557 :  13 - 0xd
      12'hDE6: dout <= 8'b00001001; // 3558 :   9 - 0x9
      12'hDE7: dout <= 8'b00000110; // 3559 :   6 - 0x6
      12'hDE8: dout <= 8'b11100000; // 3560 : 224 - 0xe0 -- Background 0xbd
      12'hDE9: dout <= 8'b01100000; // 3561 :  96 - 0x60
      12'hDEA: dout <= 8'b11100011; // 3562 : 227 - 0xe3
      12'hDEB: dout <= 8'b11100111; // 3563 : 231 - 0xe7
      12'hDEC: dout <= 8'b00000110; // 3564 :   6 - 0x6
      12'hDED: dout <= 8'b00000100; // 3565 :   4 - 0x4
      12'hDEE: dout <= 8'b00000100; // 3566 :   4 - 0x4
      12'hDEF: dout <= 8'b00000111; // 3567 :   7 - 0x7
      12'hDF0: dout <= 8'b00000111; // 3568 :   7 - 0x7 -- Background 0xbe
      12'hDF1: dout <= 8'b00000011; // 3569 :   3 - 0x3
      12'hDF2: dout <= 8'b10000111; // 3570 : 135 - 0x87
      12'hDF3: dout <= 8'b11000111; // 3571 : 199 - 0xc7
      12'hDF4: dout <= 8'b00100000; // 3572 :  32 - 0x20
      12'hDF5: dout <= 8'b00100000; // 3573 :  32 - 0x20
      12'hDF6: dout <= 8'b01100000; // 3574 :  96 - 0x60
      12'hDF7: dout <= 8'b11100000; // 3575 : 224 - 0xe0
      12'hDF8: dout <= 8'b00000111; // 3576 :   7 - 0x7 -- Background 0xbf
      12'hDF9: dout <= 8'b00000011; // 3577 :   3 - 0x3
      12'hDFA: dout <= 8'b00000000; // 3578 :   0 - 0x0
      12'hDFB: dout <= 8'b00001100; // 3579 :  12 - 0xc
      12'hDFC: dout <= 8'b11101100; // 3580 : 236 - 0xec
      12'hDFD: dout <= 8'b01100100; // 3581 : 100 - 0x64
      12'hDFE: dout <= 8'b11101100; // 3582 : 236 - 0xec
      12'hDFF: dout <= 8'b11101101; // 3583 : 237 - 0xed
      12'hE00: dout <= 8'b11100000; // 3584 : 224 - 0xe0 -- Background 0xc0
      12'hE01: dout <= 8'b11000000; // 3585 : 192 - 0xc0
      12'hE02: dout <= 8'b00000000; // 3586 :   0 - 0x0
      12'hE03: dout <= 8'b00110000; // 3587 :  48 - 0x30
      12'hE04: dout <= 8'b00110111; // 3588 :  55 - 0x37
      12'hE05: dout <= 8'b00010011; // 3589 :  19 - 0x13
      12'hE06: dout <= 8'b00110111; // 3590 :  55 - 0x37
      12'hE07: dout <= 8'b01110111; // 3591 : 119 - 0x77
      12'hE08: dout <= 8'b00001111; // 3592 :  15 - 0xf -- Background 0xc1
      12'hE09: dout <= 8'b00001100; // 3593 :  12 - 0xc
      12'hE0A: dout <= 8'b00000000; // 3594 :   0 - 0x0
      12'hE0B: dout <= 8'b00000000; // 3595 :   0 - 0x0
      12'hE0C: dout <= 8'b00000000; // 3596 :   0 - 0x0
      12'hE0D: dout <= 8'b00000000; // 3597 :   0 - 0x0
      12'hE0E: dout <= 8'b00000000; // 3598 :   0 - 0x0
      12'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout <= 8'b11110000; // 3600 : 240 - 0xf0 -- Background 0xc2
      12'hE11: dout <= 8'b00110000; // 3601 :  48 - 0x30
      12'hE12: dout <= 8'b00000000; // 3602 :   0 - 0x0
      12'hE13: dout <= 8'b00000000; // 3603 :   0 - 0x0
      12'hE14: dout <= 8'b00000000; // 3604 :   0 - 0x0
      12'hE15: dout <= 8'b00000000; // 3605 :   0 - 0x0
      12'hE16: dout <= 8'b00000000; // 3606 :   0 - 0x0
      12'hE17: dout <= 8'b00000000; // 3607 :   0 - 0x0
      12'hE18: dout <= 8'b00000000; // 3608 :   0 - 0x0 -- Background 0xc3
      12'hE19: dout <= 8'b00000000; // 3609 :   0 - 0x0
      12'hE1A: dout <= 8'b00000000; // 3610 :   0 - 0x0
      12'hE1B: dout <= 8'b00000100; // 3611 :   4 - 0x4
      12'hE1C: dout <= 8'b00001101; // 3612 :  13 - 0xd
      12'hE1D: dout <= 8'b00001111; // 3613 :  15 - 0xf
      12'hE1E: dout <= 8'b00001100; // 3614 :  12 - 0xc
      12'hE1F: dout <= 8'b00001100; // 3615 :  12 - 0xc
      12'hE20: dout <= 8'b00000000; // 3616 :   0 - 0x0 -- Background 0xc4
      12'hE21: dout <= 8'b00000000; // 3617 :   0 - 0x0
      12'hE22: dout <= 8'b00000000; // 3618 :   0 - 0x0
      12'hE23: dout <= 8'b00010000; // 3619 :  16 - 0x10
      12'hE24: dout <= 8'b01110000; // 3620 : 112 - 0x70
      12'hE25: dout <= 8'b11110000; // 3621 : 240 - 0xf0
      12'hE26: dout <= 8'b00110000; // 3622 :  48 - 0x30
      12'hE27: dout <= 8'b00110000; // 3623 :  48 - 0x30
      12'hE28: dout <= 8'b11100100; // 3624 : 228 - 0xe4 -- Background 0xc5
      12'hE29: dout <= 8'b00100100; // 3625 :  36 - 0x24
      12'hE2A: dout <= 8'b11100100; // 3626 : 228 - 0xe4
      12'hE2B: dout <= 8'b11101111; // 3627 : 239 - 0xef
      12'hE2C: dout <= 8'b00000111; // 3628 :   7 - 0x7
      12'hE2D: dout <= 8'b00000110; // 3629 :   6 - 0x6
      12'hE2E: dout <= 8'b00000100; // 3630 :   4 - 0x4
      12'hE2F: dout <= 8'b00000100; // 3631 :   4 - 0x4
      12'hE30: dout <= 8'b00010111; // 3632 :  23 - 0x17 -- Background 0xc6
      12'hE31: dout <= 8'b00010001; // 3633 :  17 - 0x11
      12'hE32: dout <= 8'b00010111; // 3634 :  23 - 0x17
      12'hE33: dout <= 8'b10110111; // 3635 : 183 - 0xb7
      12'hE34: dout <= 8'b11000000; // 3636 : 192 - 0xc0
      12'hE35: dout <= 8'b00100000; // 3637 :  32 - 0x20
      12'hE36: dout <= 8'b00100000; // 3638 :  32 - 0x20
      12'hE37: dout <= 8'b01100000; // 3639 :  96 - 0x60
      12'hE38: dout <= 8'b00000111; // 3640 :   7 - 0x7 -- Background 0xc7
      12'hE39: dout <= 8'b00000111; // 3641 :   7 - 0x7
      12'hE3A: dout <= 8'b00000011; // 3642 :   3 - 0x3
      12'hE3B: dout <= 8'b00000000; // 3643 :   0 - 0x0
      12'hE3C: dout <= 8'b11100000; // 3644 : 224 - 0xe0
      12'hE3D: dout <= 8'b00100000; // 3645 :  32 - 0x20
      12'hE3E: dout <= 8'b11100000; // 3646 : 224 - 0xe0
      12'hE3F: dout <= 8'b11100000; // 3647 : 224 - 0xe0
      12'hE40: dout <= 8'b11100000; // 3648 : 224 - 0xe0 -- Background 0xc8
      12'hE41: dout <= 8'b11100000; // 3649 : 224 - 0xe0
      12'hE42: dout <= 8'b11000000; // 3650 : 192 - 0xc0
      12'hE43: dout <= 8'b00000000; // 3651 :   0 - 0x0
      12'hE44: dout <= 8'b00000111; // 3652 :   7 - 0x7
      12'hE45: dout <= 8'b00000001; // 3653 :   1 - 0x1
      12'hE46: dout <= 8'b00000111; // 3654 :   7 - 0x7
      12'hE47: dout <= 8'b00000111; // 3655 :   7 - 0x7
      12'hE48: dout <= 8'b00000001; // 3656 :   1 - 0x1 -- Background 0xc9
      12'hE49: dout <= 8'b00010011; // 3657 :  19 - 0x13
      12'hE4A: dout <= 8'b00011111; // 3658 :  31 - 0x1f
      12'hE4B: dout <= 8'b00001101; // 3659 :  13 - 0xd
      12'hE4C: dout <= 8'b00000100; // 3660 :   4 - 0x4
      12'hE4D: dout <= 8'b00001100; // 3661 :  12 - 0xc
      12'hE4E: dout <= 8'b00010011; // 3662 :  19 - 0x13
      12'hE4F: dout <= 8'b00011111; // 3663 :  31 - 0x1f
      12'hE50: dout <= 8'b01100000; // 3664 :  96 - 0x60 -- Background 0xca
      12'hE51: dout <= 8'b01110000; // 3665 : 112 - 0x70
      12'hE52: dout <= 8'b10100011; // 3666 : 163 - 0xa3
      12'hE53: dout <= 8'b10000111; // 3667 : 135 - 0x87
      12'hE54: dout <= 8'b11000110; // 3668 : 198 - 0xc6
      12'hE55: dout <= 8'b01110100; // 3669 : 116 - 0x74
      12'hE56: dout <= 8'b00000100; // 3670 :   4 - 0x4
      12'hE57: dout <= 8'b10000111; // 3671 : 135 - 0x87
      12'hE58: dout <= 8'b00000110; // 3672 :   6 - 0x6 -- Background 0xcb
      12'hE59: dout <= 8'b00001111; // 3673 :  15 - 0xf
      12'hE5A: dout <= 8'b10000011; // 3674 : 131 - 0x83
      12'hE5B: dout <= 8'b11000001; // 3675 : 193 - 0xc1
      12'hE5C: dout <= 8'b00100000; // 3676 :  32 - 0x20
      12'hE5D: dout <= 8'b00100000; // 3677 :  32 - 0x20
      12'hE5E: dout <= 8'b01100000; // 3678 :  96 - 0x60
      12'hE5F: dout <= 8'b11100000; // 3679 : 224 - 0xe0
      12'hE60: dout <= 8'b10000111; // 3680 : 135 - 0x87 -- Background 0xcc
      12'hE61: dout <= 8'b01000011; // 3681 :  67 - 0x43
      12'hE62: dout <= 8'b00110000; // 3682 :  48 - 0x30
      12'hE63: dout <= 8'b01100000; // 3683 :  96 - 0x60
      12'hE64: dout <= 8'b11110000; // 3684 : 240 - 0xf0
      12'hE65: dout <= 8'b11010000; // 3685 : 208 - 0xd0
      12'hE66: dout <= 8'b10010000; // 3686 : 144 - 0x90
      12'hE67: dout <= 8'b01100000; // 3687 :  96 - 0x60
      12'hE68: dout <= 8'b11100000; // 3688 : 224 - 0xe0 -- Background 0xcd
      12'hE69: dout <= 8'b11000000; // 3689 : 192 - 0xc0
      12'hE6A: dout <= 8'b00000000; // 3690 :   0 - 0x0
      12'hE6B: dout <= 8'b00000110; // 3691 :   6 - 0x6
      12'hE6C: dout <= 8'b00001111; // 3692 :  15 - 0xf
      12'hE6D: dout <= 8'b00001101; // 3693 :  13 - 0xd
      12'hE6E: dout <= 8'b00001001; // 3694 :   9 - 0x9
      12'hE6F: dout <= 8'b00000110; // 3695 :   6 - 0x6
      12'hE70: dout <= 8'b11111100; // 3696 : 252 - 0xfc -- Background 0xce
      12'hE71: dout <= 8'b11000000; // 3697 : 192 - 0xc0
      12'hE72: dout <= 8'b11010001; // 3698 : 209 - 0xd1
      12'hE73: dout <= 8'b11000010; // 3699 : 194 - 0xc2
      12'hE74: dout <= 8'b10011110; // 3700 : 158 - 0x9e
      12'hE75: dout <= 8'b10111111; // 3701 : 191 - 0xbf
      12'hE76: dout <= 8'b10110000; // 3702 : 176 - 0xb0
      12'hE77: dout <= 8'b10110011; // 3703 : 179 - 0xb3
      12'hE78: dout <= 8'b00000111; // 3704 :   7 - 0x7 -- Background 0xcf
      12'hE79: dout <= 8'b11110011; // 3705 : 243 - 0xf3
      12'hE7A: dout <= 8'b00001011; // 3706 :  11 - 0xb
      12'hE7B: dout <= 8'b01111011; // 3707 : 123 - 0x7b
      12'hE7C: dout <= 8'b01111011; // 3708 : 123 - 0x7b
      12'hE7D: dout <= 8'b11111001; // 3709 : 249 - 0xf9
      12'hE7E: dout <= 8'b00001101; // 3710 :  13 - 0xd
      12'hE7F: dout <= 8'b11101101; // 3711 : 237 - 0xed
      12'hE80: dout <= 8'b11111111; // 3712 : 255 - 0xff -- Background 0xd0
      12'hE81: dout <= 8'b11111111; // 3713 : 255 - 0xff
      12'hE82: dout <= 8'b11111111; // 3714 : 255 - 0xff
      12'hE83: dout <= 8'b11111111; // 3715 : 255 - 0xff
      12'hE84: dout <= 8'b11101110; // 3716 : 238 - 0xee
      12'hE85: dout <= 8'b11101110; // 3717 : 238 - 0xee
      12'hE86: dout <= 8'b11101110; // 3718 : 238 - 0xee
      12'hE87: dout <= 8'b11101110; // 3719 : 238 - 0xee
      12'hE88: dout <= 8'b11111111; // 3720 : 255 - 0xff -- Background 0xd1
      12'hE89: dout <= 8'b11111111; // 3721 : 255 - 0xff
      12'hE8A: dout <= 8'b11111111; // 3722 : 255 - 0xff
      12'hE8B: dout <= 8'b11111011; // 3723 : 251 - 0xfb
      12'hE8C: dout <= 8'b11111011; // 3724 : 251 - 0xfb
      12'hE8D: dout <= 8'b11111011; // 3725 : 251 - 0xfb
      12'hE8E: dout <= 8'b11111011; // 3726 : 251 - 0xfb
      12'hE8F: dout <= 8'b11111011; // 3727 : 251 - 0xfb
      12'hE90: dout <= 8'b11111111; // 3728 : 255 - 0xff -- Background 0xd2
      12'hE91: dout <= 8'b11111111; // 3729 : 255 - 0xff
      12'hE92: dout <= 8'b11111111; // 3730 : 255 - 0xff
      12'hE93: dout <= 8'b11111111; // 3731 : 255 - 0xff
      12'hE94: dout <= 8'b11101110; // 3732 : 238 - 0xee
      12'hE95: dout <= 8'b10001110; // 3733 : 142 - 0x8e
      12'hE96: dout <= 8'b11111110; // 3734 : 254 - 0xfe
      12'hE97: dout <= 8'b11111110; // 3735 : 254 - 0xfe
      12'hE98: dout <= 8'b11111111; // 3736 : 255 - 0xff -- Background 0xd3
      12'hE99: dout <= 8'b11111111; // 3737 : 255 - 0xff
      12'hE9A: dout <= 8'b11111111; // 3738 : 255 - 0xff
      12'hE9B: dout <= 8'b11111111; // 3739 : 255 - 0xff
      12'hE9C: dout <= 8'b11101110; // 3740 : 238 - 0xee
      12'hE9D: dout <= 8'b10001110; // 3741 : 142 - 0x8e
      12'hE9E: dout <= 8'b11111100; // 3742 : 252 - 0xfc
      12'hE9F: dout <= 8'b11111101; // 3743 : 253 - 0xfd
      12'hEA0: dout <= 8'b11111111; // 3744 : 255 - 0xff -- Background 0xd4
      12'hEA1: dout <= 8'b11111111; // 3745 : 255 - 0xff
      12'hEA2: dout <= 8'b11111111; // 3746 : 255 - 0xff
      12'hEA3: dout <= 8'b11111110; // 3747 : 254 - 0xfe
      12'hEA4: dout <= 8'b11101110; // 3748 : 238 - 0xee
      12'hEA5: dout <= 8'b11101110; // 3749 : 238 - 0xee
      12'hEA6: dout <= 8'b11101110; // 3750 : 238 - 0xee
      12'hEA7: dout <= 8'b11101110; // 3751 : 238 - 0xee
      12'hEA8: dout <= 8'b11111111; // 3752 : 255 - 0xff -- Background 0xd5
      12'hEA9: dout <= 8'b11111111; // 3753 : 255 - 0xff
      12'hEAA: dout <= 8'b11111111; // 3754 : 255 - 0xff
      12'hEAB: dout <= 8'b11111101; // 3755 : 253 - 0xfd
      12'hEAC: dout <= 8'b11100001; // 3756 : 225 - 0xe1
      12'hEAD: dout <= 8'b11101111; // 3757 : 239 - 0xef
      12'hEAE: dout <= 8'b11111111; // 3758 : 255 - 0xff
      12'hEAF: dout <= 8'b11111111; // 3759 : 255 - 0xff
      12'hEB0: dout <= 8'b11111111; // 3760 : 255 - 0xff -- Background 0xd6
      12'hEB1: dout <= 8'b11111111; // 3761 : 255 - 0xff
      12'hEB2: dout <= 8'b11111111; // 3762 : 255 - 0xff
      12'hEB3: dout <= 8'b11111101; // 3763 : 253 - 0xfd
      12'hEB4: dout <= 8'b11100001; // 3764 : 225 - 0xe1
      12'hEB5: dout <= 8'b11101111; // 3765 : 239 - 0xef
      12'hEB6: dout <= 8'b11111111; // 3766 : 255 - 0xff
      12'hEB7: dout <= 8'b11111111; // 3767 : 255 - 0xff
      12'hEB8: dout <= 8'b11111111; // 3768 : 255 - 0xff -- Background 0xd7
      12'hEB9: dout <= 8'b11111111; // 3769 : 255 - 0xff
      12'hEBA: dout <= 8'b11111111; // 3770 : 255 - 0xff
      12'hEBB: dout <= 8'b11111110; // 3771 : 254 - 0xfe
      12'hEBC: dout <= 8'b11101110; // 3772 : 238 - 0xee
      12'hEBD: dout <= 8'b10001110; // 3773 : 142 - 0x8e
      12'hEBE: dout <= 8'b11111110; // 3774 : 254 - 0xfe
      12'hEBF: dout <= 8'b11111100; // 3775 : 252 - 0xfc
      12'hEC0: dout <= 8'b11111111; // 3776 : 255 - 0xff -- Background 0xd8
      12'hEC1: dout <= 8'b11111111; // 3777 : 255 - 0xff
      12'hEC2: dout <= 8'b11111111; // 3778 : 255 - 0xff
      12'hEC3: dout <= 8'b11111111; // 3779 : 255 - 0xff
      12'hEC4: dout <= 8'b11101110; // 3780 : 238 - 0xee
      12'hEC5: dout <= 8'b11101110; // 3781 : 238 - 0xee
      12'hEC6: dout <= 8'b11111100; // 3782 : 252 - 0xfc
      12'hEC7: dout <= 8'b11111111; // 3783 : 255 - 0xff
      12'hEC8: dout <= 8'b11111111; // 3784 : 255 - 0xff -- Background 0xd9
      12'hEC9: dout <= 8'b11111111; // 3785 : 255 - 0xff
      12'hECA: dout <= 8'b11111111; // 3786 : 255 - 0xff
      12'hECB: dout <= 8'b11111111; // 3787 : 255 - 0xff
      12'hECC: dout <= 8'b11101110; // 3788 : 238 - 0xee
      12'hECD: dout <= 8'b11101110; // 3789 : 238 - 0xee
      12'hECE: dout <= 8'b11101110; // 3790 : 238 - 0xee
      12'hECF: dout <= 8'b11101110; // 3791 : 238 - 0xee
      12'hED0: dout <= 8'b00000000; // 3792 :   0 - 0x0 -- Background 0xda
      12'hED1: dout <= 8'b00000000; // 3793 :   0 - 0x0
      12'hED2: dout <= 8'b00000000; // 3794 :   0 - 0x0
      12'hED3: dout <= 8'b10000000; // 3795 : 128 - 0x80
      12'hED4: dout <= 8'b00000000; // 3796 :   0 - 0x0
      12'hED5: dout <= 8'b00000000; // 3797 :   0 - 0x0
      12'hED6: dout <= 8'b00000100; // 3798 :   4 - 0x4
      12'hED7: dout <= 8'b00000000; // 3799 :   0 - 0x0
      12'hED8: dout <= 8'b00000000; // 3800 :   0 - 0x0 -- Background 0xdb
      12'hED9: dout <= 8'b00000100; // 3801 :   4 - 0x4
      12'hEDA: dout <= 8'b00000000; // 3802 :   0 - 0x0
      12'hEDB: dout <= 8'b00010001; // 3803 :  17 - 0x11
      12'hEDC: dout <= 8'b00000000; // 3804 :   0 - 0x0
      12'hEDD: dout <= 8'b00000000; // 3805 :   0 - 0x0
      12'hEDE: dout <= 8'b00000000; // 3806 :   0 - 0x0
      12'hEDF: dout <= 8'b00100000; // 3807 :  32 - 0x20
      12'hEE0: dout <= 8'b00000000; // 3808 :   0 - 0x0 -- Background 0xdc
      12'hEE1: dout <= 8'b00000000; // 3809 :   0 - 0x0
      12'hEE2: dout <= 8'b00000000; // 3810 :   0 - 0x0
      12'hEE3: dout <= 8'b00100000; // 3811 :  32 - 0x20
      12'hEE4: dout <= 8'b00000000; // 3812 :   0 - 0x0
      12'hEE5: dout <= 8'b00000000; // 3813 :   0 - 0x0
      12'hEE6: dout <= 8'b00000000; // 3814 :   0 - 0x0
      12'hEE7: dout <= 8'b00000100; // 3815 :   4 - 0x4
      12'hEE8: dout <= 8'b00000000; // 3816 :   0 - 0x0 -- Background 0xdd
      12'hEE9: dout <= 8'b00000000; // 3817 :   0 - 0x0
      12'hEEA: dout <= 8'b00010001; // 3818 :  17 - 0x11
      12'hEEB: dout <= 8'b00000000; // 3819 :   0 - 0x0
      12'hEEC: dout <= 8'b00000000; // 3820 :   0 - 0x0
      12'hEED: dout <= 8'b10000000; // 3821 : 128 - 0x80
      12'hEEE: dout <= 8'b00000000; // 3822 :   0 - 0x0
      12'hEEF: dout <= 8'b00000000; // 3823 :   0 - 0x0
      12'hEF0: dout <= 8'b10110011; // 3824 : 179 - 0xb3 -- Background 0xde
      12'hEF1: dout <= 8'b10110011; // 3825 : 179 - 0xb3
      12'hEF2: dout <= 8'b10110011; // 3826 : 179 - 0xb3
      12'hEF3: dout <= 8'b10110011; // 3827 : 179 - 0xb3
      12'hEF4: dout <= 8'b10110000; // 3828 : 176 - 0xb0
      12'hEF5: dout <= 8'b10101111; // 3829 : 175 - 0xaf
      12'hEF6: dout <= 8'b10011111; // 3830 : 159 - 0x9f
      12'hEF7: dout <= 8'b11000000; // 3831 : 192 - 0xc0
      12'hEF8: dout <= 8'b11101101; // 3832 : 237 - 0xed -- Background 0xdf
      12'hEF9: dout <= 8'b11001101; // 3833 : 205 - 0xcd
      12'hEFA: dout <= 8'b11001101; // 3834 : 205 - 0xcd
      12'hEFB: dout <= 8'b00001101; // 3835 :  13 - 0xd
      12'hEFC: dout <= 8'b00001101; // 3836 :  13 - 0xd
      12'hEFD: dout <= 8'b11111101; // 3837 : 253 - 0xfd
      12'hEFE: dout <= 8'b11111101; // 3838 : 253 - 0xfd
      12'hEFF: dout <= 8'b00000011; // 3839 :   3 - 0x3
      12'hF00: dout <= 8'b11101110; // 3840 : 238 - 0xee -- Background 0xe0
      12'hF01: dout <= 8'b11101110; // 3841 : 238 - 0xee
      12'hF02: dout <= 8'b11101110; // 3842 : 238 - 0xee
      12'hF03: dout <= 8'b11101110; // 3843 : 238 - 0xee
      12'hF04: dout <= 8'b11111110; // 3844 : 254 - 0xfe
      12'hF05: dout <= 8'b11111100; // 3845 : 252 - 0xfc
      12'hF06: dout <= 8'b11000001; // 3846 : 193 - 0xc1
      12'hF07: dout <= 8'b11111111; // 3847 : 255 - 0xff
      12'hF08: dout <= 8'b11111011; // 3848 : 251 - 0xfb -- Background 0xe1
      12'hF09: dout <= 8'b11111011; // 3849 : 251 - 0xfb
      12'hF0A: dout <= 8'b11111011; // 3850 : 251 - 0xfb
      12'hF0B: dout <= 8'b11111011; // 3851 : 251 - 0xfb
      12'hF0C: dout <= 8'b11111111; // 3852 : 255 - 0xff
      12'hF0D: dout <= 8'b11111101; // 3853 : 253 - 0xfd
      12'hF0E: dout <= 8'b11000001; // 3854 : 193 - 0xc1
      12'hF0F: dout <= 8'b11111111; // 3855 : 255 - 0xff
      12'hF10: dout <= 8'b11111100; // 3856 : 252 - 0xfc -- Background 0xe2
      12'hF11: dout <= 8'b11100001; // 3857 : 225 - 0xe1
      12'hF12: dout <= 8'b11101111; // 3858 : 239 - 0xef
      12'hF13: dout <= 8'b11101111; // 3859 : 239 - 0xef
      12'hF14: dout <= 8'b11111111; // 3860 : 255 - 0xff
      12'hF15: dout <= 8'b11111110; // 3861 : 254 - 0xfe
      12'hF16: dout <= 8'b10000000; // 3862 : 128 - 0x80
      12'hF17: dout <= 8'b11111111; // 3863 : 255 - 0xff
      12'hF18: dout <= 8'b11101110; // 3864 : 238 - 0xee -- Background 0xe3
      12'hF19: dout <= 8'b11111110; // 3865 : 254 - 0xfe
      12'hF1A: dout <= 8'b11111110; // 3866 : 254 - 0xfe
      12'hF1B: dout <= 8'b11111110; // 3867 : 254 - 0xfe
      12'hF1C: dout <= 8'b11111110; // 3868 : 254 - 0xfe
      12'hF1D: dout <= 8'b11111100; // 3869 : 252 - 0xfc
      12'hF1E: dout <= 8'b11000001; // 3870 : 193 - 0xc1
      12'hF1F: dout <= 8'b11111111; // 3871 : 255 - 0xff
      12'hF20: dout <= 8'b11101110; // 3872 : 238 - 0xee -- Background 0xe4
      12'hF21: dout <= 8'b11101110; // 3873 : 238 - 0xee
      12'hF22: dout <= 8'b11111110; // 3874 : 254 - 0xfe
      12'hF23: dout <= 8'b11111110; // 3875 : 254 - 0xfe
      12'hF24: dout <= 8'b10001110; // 3876 : 142 - 0x8e
      12'hF25: dout <= 8'b11111110; // 3877 : 254 - 0xfe
      12'hF26: dout <= 8'b11111000; // 3878 : 248 - 0xf8
      12'hF27: dout <= 8'b11111111; // 3879 : 255 - 0xff
      12'hF28: dout <= 8'b10001110; // 3880 : 142 - 0x8e -- Background 0xe5
      12'hF29: dout <= 8'b11111110; // 3881 : 254 - 0xfe
      12'hF2A: dout <= 8'b11111110; // 3882 : 254 - 0xfe
      12'hF2B: dout <= 8'b11111110; // 3883 : 254 - 0xfe
      12'hF2C: dout <= 8'b11111110; // 3884 : 254 - 0xfe
      12'hF2D: dout <= 8'b11111100; // 3885 : 252 - 0xfc
      12'hF2E: dout <= 8'b11000001; // 3886 : 193 - 0xc1
      12'hF2F: dout <= 8'b11111111; // 3887 : 255 - 0xff
      12'hF30: dout <= 8'b11101110; // 3888 : 238 - 0xee -- Background 0xe6
      12'hF31: dout <= 8'b11101110; // 3889 : 238 - 0xee
      12'hF32: dout <= 8'b11101110; // 3890 : 238 - 0xee
      12'hF33: dout <= 8'b11101110; // 3891 : 238 - 0xee
      12'hF34: dout <= 8'b11111110; // 3892 : 254 - 0xfe
      12'hF35: dout <= 8'b11111100; // 3893 : 252 - 0xfc
      12'hF36: dout <= 8'b11000001; // 3894 : 193 - 0xc1
      12'hF37: dout <= 8'b11111111; // 3895 : 255 - 0xff
      12'hF38: dout <= 8'b11111101; // 3896 : 253 - 0xfd -- Background 0xe7
      12'hF39: dout <= 8'b11111101; // 3897 : 253 - 0xfd
      12'hF3A: dout <= 8'b11111001; // 3898 : 249 - 0xf9
      12'hF3B: dout <= 8'b11111011; // 3899 : 251 - 0xfb
      12'hF3C: dout <= 8'b11111011; // 3900 : 251 - 0xfb
      12'hF3D: dout <= 8'b11111011; // 3901 : 251 - 0xfb
      12'hF3E: dout <= 8'b11100011; // 3902 : 227 - 0xe3
      12'hF3F: dout <= 8'b11111111; // 3903 : 255 - 0xff
      12'hF40: dout <= 8'b11101110; // 3904 : 238 - 0xee -- Background 0xe8
      12'hF41: dout <= 8'b11101110; // 3905 : 238 - 0xee
      12'hF42: dout <= 8'b11101110; // 3906 : 238 - 0xee
      12'hF43: dout <= 8'b11101110; // 3907 : 238 - 0xee
      12'hF44: dout <= 8'b11111110; // 3908 : 254 - 0xfe
      12'hF45: dout <= 8'b11111100; // 3909 : 252 - 0xfc
      12'hF46: dout <= 8'b11000001; // 3910 : 193 - 0xc1
      12'hF47: dout <= 8'b11111111; // 3911 : 255 - 0xff
      12'hF48: dout <= 8'b11111110; // 3912 : 254 - 0xfe -- Background 0xe9
      12'hF49: dout <= 8'b11111110; // 3913 : 254 - 0xfe
      12'hF4A: dout <= 8'b11001110; // 3914 : 206 - 0xce
      12'hF4B: dout <= 8'b11111110; // 3915 : 254 - 0xfe
      12'hF4C: dout <= 8'b11111110; // 3916 : 254 - 0xfe
      12'hF4D: dout <= 8'b11111100; // 3917 : 252 - 0xfc
      12'hF4E: dout <= 8'b11000001; // 3918 : 193 - 0xc1
      12'hF4F: dout <= 8'b11111111; // 3919 : 255 - 0xff
      12'hF50: dout <= 8'b00000000; // 3920 :   0 - 0x0 -- Background 0xea
      12'hF51: dout <= 8'b01110000; // 3921 : 112 - 0x70
      12'hF52: dout <= 8'b00111000; // 3922 :  56 - 0x38
      12'hF53: dout <= 8'b00000000; // 3923 :   0 - 0x0
      12'hF54: dout <= 8'b00000010; // 3924 :   2 - 0x2
      12'hF55: dout <= 8'b00000111; // 3925 :   7 - 0x7
      12'hF56: dout <= 8'b00000011; // 3926 :   3 - 0x3
      12'hF57: dout <= 8'b00000000; // 3927 :   0 - 0x0
      12'hF58: dout <= 8'b00000000; // 3928 :   0 - 0x0 -- Background 0xeb
      12'hF59: dout <= 8'b00001100; // 3929 :  12 - 0xc
      12'hF5A: dout <= 8'b00000110; // 3930 :   6 - 0x6
      12'hF5B: dout <= 8'b00000110; // 3931 :   6 - 0x6
      12'hF5C: dout <= 8'b01100000; // 3932 :  96 - 0x60
      12'hF5D: dout <= 8'b01110000; // 3933 : 112 - 0x70
      12'hF5E: dout <= 8'b00110000; // 3934 :  48 - 0x30
      12'hF5F: dout <= 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Background 0xec
      12'hF61: dout <= 8'b11000000; // 3937 : 192 - 0xc0
      12'hF62: dout <= 8'b11100000; // 3938 : 224 - 0xe0
      12'hF63: dout <= 8'b01100000; // 3939 :  96 - 0x60
      12'hF64: dout <= 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout <= 8'b00001100; // 3941 :  12 - 0xc
      12'hF66: dout <= 8'b00001110; // 3942 :  14 - 0xe
      12'hF67: dout <= 8'b00000110; // 3943 :   6 - 0x6
      12'hF68: dout <= 8'b01100000; // 3944 :  96 - 0x60 -- Background 0xed
      12'hF69: dout <= 8'b01110000; // 3945 : 112 - 0x70
      12'hF6A: dout <= 8'b00110000; // 3946 :  48 - 0x30
      12'hF6B: dout <= 8'b00000000; // 3947 :   0 - 0x0
      12'hF6C: dout <= 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout <= 8'b00001100; // 3949 :  12 - 0xc
      12'hF6E: dout <= 8'b00001110; // 3950 :  14 - 0xe
      12'hF6F: dout <= 8'b00000110; // 3951 :   6 - 0x6
      12'hF70: dout <= 8'b11111111; // 3952 : 255 - 0xff -- Background 0xee
      12'hF71: dout <= 8'b11111111; // 3953 : 255 - 0xff
      12'hF72: dout <= 8'b10111101; // 3954 : 189 - 0xbd
      12'hF73: dout <= 8'b11111111; // 3955 : 255 - 0xff
      12'hF74: dout <= 8'b11111111; // 3956 : 255 - 0xff
      12'hF75: dout <= 8'b11111011; // 3957 : 251 - 0xfb
      12'hF76: dout <= 8'b11111111; // 3958 : 255 - 0xff
      12'hF77: dout <= 8'b11111111; // 3959 : 255 - 0xff
      12'hF78: dout <= 8'b11111111; // 3960 : 255 - 0xff -- Background 0xef
      12'hF79: dout <= 8'b11111111; // 3961 : 255 - 0xff
      12'hF7A: dout <= 8'b11111011; // 3962 : 251 - 0xfb
      12'hF7B: dout <= 8'b11111111; // 3963 : 255 - 0xff
      12'hF7C: dout <= 8'b11011111; // 3964 : 223 - 0xdf
      12'hF7D: dout <= 8'b11111111; // 3965 : 255 - 0xff
      12'hF7E: dout <= 8'b11111111; // 3966 : 255 - 0xff
      12'hF7F: dout <= 8'b11111111; // 3967 : 255 - 0xff
      12'hF80: dout <= 8'b00000000; // 3968 :   0 - 0x0 -- Background 0xf0
      12'hF81: dout <= 8'b00000000; // 3969 :   0 - 0x0
      12'hF82: dout <= 8'b00000000; // 3970 :   0 - 0x0
      12'hF83: dout <= 8'b00000000; // 3971 :   0 - 0x0
      12'hF84: dout <= 8'b00000000; // 3972 :   0 - 0x0
      12'hF85: dout <= 8'b00000000; // 3973 :   0 - 0x0
      12'hF86: dout <= 8'b00000000; // 3974 :   0 - 0x0
      12'hF87: dout <= 8'b00000000; // 3975 :   0 - 0x0
      12'hF88: dout <= 8'b00000000; // 3976 :   0 - 0x0 -- Background 0xf1
      12'hF89: dout <= 8'b10000000; // 3977 : 128 - 0x80
      12'hF8A: dout <= 8'b00000000; // 3978 :   0 - 0x0
      12'hF8B: dout <= 8'b00000000; // 3979 :   0 - 0x0
      12'hF8C: dout <= 8'b00000000; // 3980 :   0 - 0x0
      12'hF8D: dout <= 8'b00000000; // 3981 :   0 - 0x0
      12'hF8E: dout <= 8'b00000000; // 3982 :   0 - 0x0
      12'hF8F: dout <= 8'b00000000; // 3983 :   0 - 0x0
      12'hF90: dout <= 8'b00000000; // 3984 :   0 - 0x0 -- Background 0xf2
      12'hF91: dout <= 8'b11000000; // 3985 : 192 - 0xc0
      12'hF92: dout <= 8'b00000000; // 3986 :   0 - 0x0
      12'hF93: dout <= 8'b00000000; // 3987 :   0 - 0x0
      12'hF94: dout <= 8'b00000000; // 3988 :   0 - 0x0
      12'hF95: dout <= 8'b00000000; // 3989 :   0 - 0x0
      12'hF96: dout <= 8'b00000000; // 3990 :   0 - 0x0
      12'hF97: dout <= 8'b00000000; // 3991 :   0 - 0x0
      12'hF98: dout <= 8'b00000000; // 3992 :   0 - 0x0 -- Background 0xf3
      12'hF99: dout <= 8'b11100000; // 3993 : 224 - 0xe0
      12'hF9A: dout <= 8'b00000000; // 3994 :   0 - 0x0
      12'hF9B: dout <= 8'b00000000; // 3995 :   0 - 0x0
      12'hF9C: dout <= 8'b00000000; // 3996 :   0 - 0x0
      12'hF9D: dout <= 8'b00000000; // 3997 :   0 - 0x0
      12'hF9E: dout <= 8'b00000000; // 3998 :   0 - 0x0
      12'hF9F: dout <= 8'b00000000; // 3999 :   0 - 0x0
      12'hFA0: dout <= 8'b00000000; // 4000 :   0 - 0x0 -- Background 0xf4
      12'hFA1: dout <= 8'b11110000; // 4001 : 240 - 0xf0
      12'hFA2: dout <= 8'b00000000; // 4002 :   0 - 0x0
      12'hFA3: dout <= 8'b00000000; // 4003 :   0 - 0x0
      12'hFA4: dout <= 8'b00000000; // 4004 :   0 - 0x0
      12'hFA5: dout <= 8'b00000000; // 4005 :   0 - 0x0
      12'hFA6: dout <= 8'b00000000; // 4006 :   0 - 0x0
      12'hFA7: dout <= 8'b00000000; // 4007 :   0 - 0x0
      12'hFA8: dout <= 8'b00000000; // 4008 :   0 - 0x0 -- Background 0xf5
      12'hFA9: dout <= 8'b11111000; // 4009 : 248 - 0xf8
      12'hFAA: dout <= 8'b00000000; // 4010 :   0 - 0x0
      12'hFAB: dout <= 8'b00000000; // 4011 :   0 - 0x0
      12'hFAC: dout <= 8'b00000000; // 4012 :   0 - 0x0
      12'hFAD: dout <= 8'b00000000; // 4013 :   0 - 0x0
      12'hFAE: dout <= 8'b00000000; // 4014 :   0 - 0x0
      12'hFAF: dout <= 8'b00000000; // 4015 :   0 - 0x0
      12'hFB0: dout <= 8'b00000000; // 4016 :   0 - 0x0 -- Background 0xf6
      12'hFB1: dout <= 8'b11111100; // 4017 : 252 - 0xfc
      12'hFB2: dout <= 8'b00000000; // 4018 :   0 - 0x0
      12'hFB3: dout <= 8'b00000000; // 4019 :   0 - 0x0
      12'hFB4: dout <= 8'b00000000; // 4020 :   0 - 0x0
      12'hFB5: dout <= 8'b00000000; // 4021 :   0 - 0x0
      12'hFB6: dout <= 8'b00000000; // 4022 :   0 - 0x0
      12'hFB7: dout <= 8'b00000000; // 4023 :   0 - 0x0
      12'hFB8: dout <= 8'b00000000; // 4024 :   0 - 0x0 -- Background 0xf7
      12'hFB9: dout <= 8'b11111110; // 4025 : 254 - 0xfe
      12'hFBA: dout <= 8'b00000000; // 4026 :   0 - 0x0
      12'hFBB: dout <= 8'b00000000; // 4027 :   0 - 0x0
      12'hFBC: dout <= 8'b00000000; // 4028 :   0 - 0x0
      12'hFBD: dout <= 8'b00000000; // 4029 :   0 - 0x0
      12'hFBE: dout <= 8'b00000000; // 4030 :   0 - 0x0
      12'hFBF: dout <= 8'b00000000; // 4031 :   0 - 0x0
      12'hFC0: dout <= 8'b00000000; // 4032 :   0 - 0x0 -- Background 0xf8
      12'hFC1: dout <= 8'b11111111; // 4033 : 255 - 0xff
      12'hFC2: dout <= 8'b00000000; // 4034 :   0 - 0x0
      12'hFC3: dout <= 8'b00000000; // 4035 :   0 - 0x0
      12'hFC4: dout <= 8'b00000000; // 4036 :   0 - 0x0
      12'hFC5: dout <= 8'b00000000; // 4037 :   0 - 0x0
      12'hFC6: dout <= 8'b00000000; // 4038 :   0 - 0x0
      12'hFC7: dout <= 8'b00000000; // 4039 :   0 - 0x0
      12'hFC8: dout <= 8'b11111111; // 4040 : 255 - 0xff -- Background 0xf9
      12'hFC9: dout <= 8'b11111111; // 4041 : 255 - 0xff
      12'hFCA: dout <= 8'b11111111; // 4042 : 255 - 0xff
      12'hFCB: dout <= 8'b11111111; // 4043 : 255 - 0xff
      12'hFCC: dout <= 8'b10000000; // 4044 : 128 - 0x80
      12'hFCD: dout <= 8'b10000000; // 4045 : 128 - 0x80
      12'hFCE: dout <= 8'b11000000; // 4046 : 192 - 0xc0
      12'hFCF: dout <= 8'b11000000; // 4047 : 192 - 0xc0
      12'hFD0: dout <= 8'b11111111; // 4048 : 255 - 0xff -- Background 0xfa
      12'hFD1: dout <= 8'b11111111; // 4049 : 255 - 0xff
      12'hFD2: dout <= 8'b11111111; // 4050 : 255 - 0xff
      12'hFD3: dout <= 8'b11111111; // 4051 : 255 - 0xff
      12'hFD4: dout <= 8'b00000000; // 4052 :   0 - 0x0
      12'hFD5: dout <= 8'b00000000; // 4053 :   0 - 0x0
      12'hFD6: dout <= 8'b00000000; // 4054 :   0 - 0x0
      12'hFD7: dout <= 8'b00000000; // 4055 :   0 - 0x0
      12'hFD8: dout <= 8'b11111111; // 4056 : 255 - 0xff -- Background 0xfb
      12'hFD9: dout <= 8'b11111111; // 4057 : 255 - 0xff
      12'hFDA: dout <= 8'b11111111; // 4058 : 255 - 0xff
      12'hFDB: dout <= 8'b11111111; // 4059 : 255 - 0xff
      12'hFDC: dout <= 8'b00000001; // 4060 :   1 - 0x1
      12'hFDD: dout <= 8'b00000000; // 4061 :   0 - 0x0
      12'hFDE: dout <= 8'b00000010; // 4062 :   2 - 0x2
      12'hFDF: dout <= 8'b00000010; // 4063 :   2 - 0x2
      12'hFE0: dout <= 8'b11000000; // 4064 : 192 - 0xc0 -- Background 0xfc
      12'hFE1: dout <= 8'b11000000; // 4065 : 192 - 0xc0
      12'hFE2: dout <= 8'b10000000; // 4066 : 128 - 0x80
      12'hFE3: dout <= 8'b10000000; // 4067 : 128 - 0x80
      12'hFE4: dout <= 8'b11000000; // 4068 : 192 - 0xc0
      12'hFE5: dout <= 8'b11111111; // 4069 : 255 - 0xff
      12'hFE6: dout <= 8'b11111111; // 4070 : 255 - 0xff
      12'hFE7: dout <= 8'b11111111; // 4071 : 255 - 0xff
      12'hFE8: dout <= 8'b00000000; // 4072 :   0 - 0x0 -- Background 0xfd
      12'hFE9: dout <= 8'b00000000; // 4073 :   0 - 0x0
      12'hFEA: dout <= 8'b00000000; // 4074 :   0 - 0x0
      12'hFEB: dout <= 8'b00000000; // 4075 :   0 - 0x0
      12'hFEC: dout <= 8'b00000000; // 4076 :   0 - 0x0
      12'hFED: dout <= 8'b11111111; // 4077 : 255 - 0xff
      12'hFEE: dout <= 8'b11111111; // 4078 : 255 - 0xff
      12'hFEF: dout <= 8'b11111111; // 4079 : 255 - 0xff
      12'hFF0: dout <= 8'b00000010; // 4080 :   2 - 0x2 -- Background 0xfe
      12'hFF1: dout <= 8'b00000010; // 4081 :   2 - 0x2
      12'hFF2: dout <= 8'b00000000; // 4082 :   0 - 0x0
      12'hFF3: dout <= 8'b00000000; // 4083 :   0 - 0x0
      12'hFF4: dout <= 8'b00000000; // 4084 :   0 - 0x0
      12'hFF5: dout <= 8'b11111111; // 4085 : 255 - 0xff
      12'hFF6: dout <= 8'b11111111; // 4086 : 255 - 0xff
      12'hFF7: dout <= 8'b11111111; // 4087 : 255 - 0xff
      12'hFF8: dout <= 8'b11111111; // 4088 : 255 - 0xff -- Background 0xff
      12'hFF9: dout <= 8'b11111111; // 4089 : 255 - 0xff
      12'hFFA: dout <= 8'b11111111; // 4090 : 255 - 0xff
      12'hFFB: dout <= 8'b11111111; // 4091 : 255 - 0xff
      12'hFFC: dout <= 8'b11111111; // 4092 : 255 - 0xff
      12'hFFD: dout <= 8'b11111111; // 4093 : 255 - 0xff
      12'hFFE: dout <= 8'b11111111; // 4094 : 255 - 0xff
      12'hFFF: dout <= 8'b11111111; // 4095 : 255 - 0xff
    endcase
  end

endmodule
