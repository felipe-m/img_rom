--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: nova_ntable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_NOVA_00 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_NOVA_00;

architecture BEHAVIORAL of ROM_NTABLE_NOVA_00 is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "00110000", --    0 -  0x0  :   48 - 0x30 -- line 0x0
    "00111111", --    1 -  0x1  :   63 - 0x3f
    "00110000", --    2 -  0x2  :   48 - 0x30
    "00111111", --    3 -  0x3  :   63 - 0x3f
    "00110000", --    4 -  0x4  :   48 - 0x30
    "00111111", --    5 -  0x5  :   63 - 0x3f
    "00110000", --    6 -  0x6  :   48 - 0x30
    "00111111", --    7 -  0x7  :   63 - 0x3f
    "00110000", --    8 -  0x8  :   48 - 0x30
    "00111111", --    9 -  0x9  :   63 - 0x3f
    "00110000", --   10 -  0xa  :   48 - 0x30
    "00111111", --   11 -  0xb  :   63 - 0x3f
    "00110000", --   12 -  0xc  :   48 - 0x30
    "00111111", --   13 -  0xd  :   63 - 0x3f
    "00110000", --   14 -  0xe  :   48 - 0x30
    "00111111", --   15 -  0xf  :   63 - 0x3f
    "00110000", --   16 - 0x10  :   48 - 0x30
    "00111111", --   17 - 0x11  :   63 - 0x3f
    "00110000", --   18 - 0x12  :   48 - 0x30
    "00111111", --   19 - 0x13  :   63 - 0x3f
    "01110000", --   20 - 0x14  :  112 - 0x70
    "01110001", --   21 - 0x15  :  113 - 0x71
    "01110001", --   22 - 0x16  :  113 - 0x71
    "01110001", --   23 - 0x17  :  113 - 0x71
    "01110001", --   24 - 0x18  :  113 - 0x71
    "01110001", --   25 - 0x19  :  113 - 0x71
    "01110001", --   26 - 0x1a  :  113 - 0x71
    "01110001", --   27 - 0x1b  :  113 - 0x71
    "01110001", --   28 - 0x1c  :  113 - 0x71
    "01110001", --   29 - 0x1d  :  113 - 0x71
    "01110001", --   30 - 0x1e  :  113 - 0x71
    "01110001", --   31 - 0x1f  :  113 - 0x71
    "00111111", --   32 - 0x20  :   63 - 0x3f -- line 0x1
    "00110000", --   33 - 0x21  :   48 - 0x30
    "00111111", --   34 - 0x22  :   63 - 0x3f
    "00110000", --   35 - 0x23  :   48 - 0x30
    "00111111", --   36 - 0x24  :   63 - 0x3f
    "00110000", --   37 - 0x25  :   48 - 0x30
    "00111111", --   38 - 0x26  :   63 - 0x3f
    "00110000", --   39 - 0x27  :   48 - 0x30
    "00111111", --   40 - 0x28  :   63 - 0x3f
    "00110000", --   41 - 0x29  :   48 - 0x30
    "00111111", --   42 - 0x2a  :   63 - 0x3f
    "00110000", --   43 - 0x2b  :   48 - 0x30
    "00111111", --   44 - 0x2c  :   63 - 0x3f
    "00110000", --   45 - 0x2d  :   48 - 0x30
    "00111111", --   46 - 0x2e  :   63 - 0x3f
    "00110000", --   47 - 0x2f  :   48 - 0x30
    "00111111", --   48 - 0x30  :   63 - 0x3f
    "00110000", --   49 - 0x31  :   48 - 0x30
    "00111111", --   50 - 0x32  :   63 - 0x3f
    "00110000", --   51 - 0x33  :   48 - 0x30
    "01100000", --   52 - 0x34  :   96 - 0x60
    "01110111", --   53 - 0x35  :  119 - 0x77
    "01110111", --   54 - 0x36  :  119 - 0x77
    "01110111", --   55 - 0x37  :  119 - 0x77
    "01110111", --   56 - 0x38  :  119 - 0x77
    "01110111", --   57 - 0x39  :  119 - 0x77
    "01110111", --   58 - 0x3a  :  119 - 0x77
    "01110111", --   59 - 0x3b  :  119 - 0x77
    "01110111", --   60 - 0x3c  :  119 - 0x77
    "01110111", --   61 - 0x3d  :  119 - 0x77
    "01110111", --   62 - 0x3e  :  119 - 0x77
    "01110111", --   63 - 0x3f  :  119 - 0x77
    "00110000", --   64 - 0x40  :   48 - 0x30 -- line 0x2
    "00111111", --   65 - 0x41  :   63 - 0x3f
    "00110000", --   66 - 0x42  :   48 - 0x30
    "00111111", --   67 - 0x43  :   63 - 0x3f
    "00110000", --   68 - 0x44  :   48 - 0x30
    "00111111", --   69 - 0x45  :   63 - 0x3f
    "00110000", --   70 - 0x46  :   48 - 0x30
    "00111111", --   71 - 0x47  :   63 - 0x3f
    "00110000", --   72 - 0x48  :   48 - 0x30
    "00111111", --   73 - 0x49  :   63 - 0x3f
    "00110000", --   74 - 0x4a  :   48 - 0x30
    "00111111", --   75 - 0x4b  :   63 - 0x3f
    "00110000", --   76 - 0x4c  :   48 - 0x30
    "00111111", --   77 - 0x4d  :   63 - 0x3f
    "00110000", --   78 - 0x4e  :   48 - 0x30
    "00111111", --   79 - 0x4f  :   63 - 0x3f
    "00110000", --   80 - 0x50  :   48 - 0x30
    "00111111", --   81 - 0x51  :   63 - 0x3f
    "00110000", --   82 - 0x52  :   48 - 0x30
    "00111111", --   83 - 0x53  :   63 - 0x3f
    "00111001", --   84 - 0x54  :   57 - 0x39
    "00111001", --   85 - 0x55  :   57 - 0x39
    "00111001", --   86 - 0x56  :   57 - 0x39
    "00111001", --   87 - 0x57  :   57 - 0x39
    "00111001", --   88 - 0x58  :   57 - 0x39
    "00111001", --   89 - 0x59  :   57 - 0x39
    "00111001", --   90 - 0x5a  :   57 - 0x39
    "00111001", --   91 - 0x5b  :   57 - 0x39
    "00111001", --   92 - 0x5c  :   57 - 0x39
    "00111001", --   93 - 0x5d  :   57 - 0x39
    "00111001", --   94 - 0x5e  :   57 - 0x39
    "00111001", --   95 - 0x5f  :   57 - 0x39
    "00111111", --   96 - 0x60  :   63 - 0x3f -- line 0x3
    "00110000", --   97 - 0x61  :   48 - 0x30
    "00111111", --   98 - 0x62  :   63 - 0x3f
    "00110000", --   99 - 0x63  :   48 - 0x30
    "00111111", --  100 - 0x64  :   63 - 0x3f
    "00110000", --  101 - 0x65  :   48 - 0x30
    "00111111", --  102 - 0x66  :   63 - 0x3f
    "00110000", --  103 - 0x67  :   48 - 0x30
    "00111111", --  104 - 0x68  :   63 - 0x3f
    "00110000", --  105 - 0x69  :   48 - 0x30
    "00111111", --  106 - 0x6a  :   63 - 0x3f
    "00110000", --  107 - 0x6b  :   48 - 0x30
    "00111111", --  108 - 0x6c  :   63 - 0x3f
    "00110000", --  109 - 0x6d  :   48 - 0x30
    "00111111", --  110 - 0x6e  :   63 - 0x3f
    "00110000", --  111 - 0x6f  :   48 - 0x30
    "00111111", --  112 - 0x70  :   63 - 0x3f
    "00110000", --  113 - 0x71  :   48 - 0x30
    "00111111", --  114 - 0x72  :   63 - 0x3f
    "00110000", --  115 - 0x73  :   48 - 0x30
    "00111111", --  116 - 0x74  :   63 - 0x3f
    "00111111", --  117 - 0x75  :   63 - 0x3f
    "00111111", --  118 - 0x76  :   63 - 0x3f
    "00111111", --  119 - 0x77  :   63 - 0x3f
    "00111111", --  120 - 0x78  :   63 - 0x3f
    "00111111", --  121 - 0x79  :   63 - 0x3f
    "00111111", --  122 - 0x7a  :   63 - 0x3f
    "00111111", --  123 - 0x7b  :   63 - 0x3f
    "00111111", --  124 - 0x7c  :   63 - 0x3f
    "00111111", --  125 - 0x7d  :   63 - 0x3f
    "00111111", --  126 - 0x7e  :   63 - 0x3f
    "00111111", --  127 - 0x7f  :   63 - 0x3f
    "00111111", --  128 - 0x80  :   63 - 0x3f -- line 0x4
    "00111111", --  129 - 0x81  :   63 - 0x3f
    "00111111", --  130 - 0x82  :   63 - 0x3f
    "00111111", --  131 - 0x83  :   63 - 0x3f
    "00111111", --  132 - 0x84  :   63 - 0x3f
    "00111111", --  133 - 0x85  :   63 - 0x3f
    "00111111", --  134 - 0x86  :   63 - 0x3f
    "00111111", --  135 - 0x87  :   63 - 0x3f
    "00111111", --  136 - 0x88  :   63 - 0x3f
    "00111111", --  137 - 0x89  :   63 - 0x3f
    "00111111", --  138 - 0x8a  :   63 - 0x3f
    "00111111", --  139 - 0x8b  :   63 - 0x3f
    "00111111", --  140 - 0x8c  :   63 - 0x3f
    "00111111", --  141 - 0x8d  :   63 - 0x3f
    "00111111", --  142 - 0x8e  :   63 - 0x3f
    "00111111", --  143 - 0x8f  :   63 - 0x3f
    "00111111", --  144 - 0x90  :   63 - 0x3f
    "00111111", --  145 - 0x91  :   63 - 0x3f
    "00111111", --  146 - 0x92  :   63 - 0x3f
    "00111111", --  147 - 0x93  :   63 - 0x3f
    "00111111", --  148 - 0x94  :   63 - 0x3f
    "00111111", --  149 - 0x95  :   63 - 0x3f
    "00111111", --  150 - 0x96  :   63 - 0x3f
    "00111111", --  151 - 0x97  :   63 - 0x3f
    "00111111", --  152 - 0x98  :   63 - 0x3f
    "00111111", --  153 - 0x99  :   63 - 0x3f
    "00000100", --  154 - 0x9a  :    4 - 0x4
    "00000110", --  155 - 0x9b  :    6 - 0x6
    "00111111", --  156 - 0x9c  :   63 - 0x3f
    "00111111", --  157 - 0x9d  :   63 - 0x3f
    "00010100", --  158 - 0x9e  :   20 - 0x14
    "00010110", --  159 - 0x9f  :   22 - 0x16
    "00111111", --  160 - 0xa0  :   63 - 0x3f -- line 0x5
    "00111111", --  161 - 0xa1  :   63 - 0x3f
    "00111111", --  162 - 0xa2  :   63 - 0x3f
    "00111111", --  163 - 0xa3  :   63 - 0x3f
    "00111111", --  164 - 0xa4  :   63 - 0x3f
    "00111111", --  165 - 0xa5  :   63 - 0x3f
    "00111111", --  166 - 0xa6  :   63 - 0x3f
    "00111111", --  167 - 0xa7  :   63 - 0x3f
    "00111111", --  168 - 0xa8  :   63 - 0x3f
    "00111111", --  169 - 0xa9  :   63 - 0x3f
    "00111111", --  170 - 0xaa  :   63 - 0x3f
    "00111111", --  171 - 0xab  :   63 - 0x3f
    "00111111", --  172 - 0xac  :   63 - 0x3f
    "00111111", --  173 - 0xad  :   63 - 0x3f
    "00111111", --  174 - 0xae  :   63 - 0x3f
    "00111111", --  175 - 0xaf  :   63 - 0x3f
    "00111111", --  176 - 0xb0  :   63 - 0x3f
    "00111111", --  177 - 0xb1  :   63 - 0x3f
    "00111111", --  178 - 0xb2  :   63 - 0x3f
    "00111111", --  179 - 0xb3  :   63 - 0x3f
    "00111111", --  180 - 0xb4  :   63 - 0x3f
    "00111111", --  181 - 0xb5  :   63 - 0x3f
    "00111111", --  182 - 0xb6  :   63 - 0x3f
    "00111111", --  183 - 0xb7  :   63 - 0x3f
    "00111111", --  184 - 0xb8  :   63 - 0x3f
    "00111111", --  185 - 0xb9  :   63 - 0x3f
    "00000101", --  186 - 0xba  :    5 - 0x5
    "00000111", --  187 - 0xbb  :    7 - 0x7
    "00111111", --  188 - 0xbc  :   63 - 0x3f
    "00111111", --  189 - 0xbd  :   63 - 0x3f
    "00010101", --  190 - 0xbe  :   21 - 0x15
    "00010111", --  191 - 0xbf  :   23 - 0x17
    "00111111", --  192 - 0xc0  :   63 - 0x3f -- line 0x6
    "00111111", --  193 - 0xc1  :   63 - 0x3f
    "00111111", --  194 - 0xc2  :   63 - 0x3f
    "00111111", --  195 - 0xc3  :   63 - 0x3f
    "00111111", --  196 - 0xc4  :   63 - 0x3f
    "00111111", --  197 - 0xc5  :   63 - 0x3f
    "00111111", --  198 - 0xc6  :   63 - 0x3f
    "00111111", --  199 - 0xc7  :   63 - 0x3f
    "00111111", --  200 - 0xc8  :   63 - 0x3f
    "00111111", --  201 - 0xc9  :   63 - 0x3f
    "00111111", --  202 - 0xca  :   63 - 0x3f
    "00111111", --  203 - 0xcb  :   63 - 0x3f
    "00111111", --  204 - 0xcc  :   63 - 0x3f
    "00111111", --  205 - 0xcd  :   63 - 0x3f
    "00111111", --  206 - 0xce  :   63 - 0x3f
    "00111111", --  207 - 0xcf  :   63 - 0x3f
    "00111111", --  208 - 0xd0  :   63 - 0x3f
    "00111111", --  209 - 0xd1  :   63 - 0x3f
    "00111111", --  210 - 0xd2  :   63 - 0x3f
    "00111111", --  211 - 0xd3  :   63 - 0x3f
    "00111111", --  212 - 0xd4  :   63 - 0x3f
    "00111111", --  213 - 0xd5  :   63 - 0x3f
    "00111111", --  214 - 0xd6  :   63 - 0x3f
    "00111111", --  215 - 0xd7  :   63 - 0x3f
    "00111111", --  216 - 0xd8  :   63 - 0x3f
    "00111111", --  217 - 0xd9  :   63 - 0x3f
    "00111111", --  218 - 0xda  :   63 - 0x3f
    "00111111", --  219 - 0xdb  :   63 - 0x3f
    "00111111", --  220 - 0xdc  :   63 - 0x3f
    "00111111", --  221 - 0xdd  :   63 - 0x3f
    "00111111", --  222 - 0xde  :   63 - 0x3f
    "00111111", --  223 - 0xdf  :   63 - 0x3f
    "00111111", --  224 - 0xe0  :   63 - 0x3f -- line 0x7
    "00111111", --  225 - 0xe1  :   63 - 0x3f
    "00111111", --  226 - 0xe2  :   63 - 0x3f
    "00111111", --  227 - 0xe3  :   63 - 0x3f
    "00111111", --  228 - 0xe4  :   63 - 0x3f
    "00111111", --  229 - 0xe5  :   63 - 0x3f
    "00111111", --  230 - 0xe6  :   63 - 0x3f
    "00111111", --  231 - 0xe7  :   63 - 0x3f
    "00111111", --  232 - 0xe8  :   63 - 0x3f
    "00111111", --  233 - 0xe9  :   63 - 0x3f
    "00111111", --  234 - 0xea  :   63 - 0x3f
    "00111111", --  235 - 0xeb  :   63 - 0x3f
    "00111111", --  236 - 0xec  :   63 - 0x3f
    "00111111", --  237 - 0xed  :   63 - 0x3f
    "00111111", --  238 - 0xee  :   63 - 0x3f
    "00111111", --  239 - 0xef  :   63 - 0x3f
    "00111111", --  240 - 0xf0  :   63 - 0x3f
    "00111111", --  241 - 0xf1  :   63 - 0x3f
    "00111111", --  242 - 0xf2  :   63 - 0x3f
    "00111111", --  243 - 0xf3  :   63 - 0x3f
    "00111111", --  244 - 0xf4  :   63 - 0x3f
    "00111111", --  245 - 0xf5  :   63 - 0x3f
    "00111111", --  246 - 0xf6  :   63 - 0x3f
    "00111111", --  247 - 0xf7  :   63 - 0x3f
    "00111111", --  248 - 0xf8  :   63 - 0x3f
    "00111111", --  249 - 0xf9  :   63 - 0x3f
    "00111111", --  250 - 0xfa  :   63 - 0x3f
    "00111111", --  251 - 0xfb  :   63 - 0x3f
    "00111111", --  252 - 0xfc  :   63 - 0x3f
    "00111111", --  253 - 0xfd  :   63 - 0x3f
    "00111111", --  254 - 0xfe  :   63 - 0x3f
    "00111111", --  255 - 0xff  :   63 - 0x3f
    "00111111", --  256 - 0x100  :   63 - 0x3f -- line 0x8
    "00111111", --  257 - 0x101  :   63 - 0x3f
    "00111111", --  258 - 0x102  :   63 - 0x3f
    "00111111", --  259 - 0x103  :   63 - 0x3f
    "00111111", --  260 - 0x104  :   63 - 0x3f
    "00111111", --  261 - 0x105  :   63 - 0x3f
    "00111111", --  262 - 0x106  :   63 - 0x3f
    "00111111", --  263 - 0x107  :   63 - 0x3f
    "00111111", --  264 - 0x108  :   63 - 0x3f
    "00111111", --  265 - 0x109  :   63 - 0x3f
    "00111111", --  266 - 0x10a  :   63 - 0x3f
    "00111111", --  267 - 0x10b  :   63 - 0x3f
    "00111111", --  268 - 0x10c  :   63 - 0x3f
    "00111111", --  269 - 0x10d  :   63 - 0x3f
    "00111111", --  270 - 0x10e  :   63 - 0x3f
    "00111111", --  271 - 0x10f  :   63 - 0x3f
    "00111111", --  272 - 0x110  :   63 - 0x3f
    "00111111", --  273 - 0x111  :   63 - 0x3f
    "00111111", --  274 - 0x112  :   63 - 0x3f
    "00111111", --  275 - 0x113  :   63 - 0x3f
    "00001100", --  276 - 0x114  :   12 - 0xc
    "00001110", --  277 - 0x115  :   14 - 0xe
    "00111111", --  278 - 0x116  :   63 - 0x3f
    "00111111", --  279 - 0x117  :   63 - 0x3f
    "00111111", --  280 - 0x118  :   63 - 0x3f
    "00111111", --  281 - 0x119  :   63 - 0x3f
    "00111111", --  282 - 0x11a  :   63 - 0x3f
    "00111111", --  283 - 0x11b  :   63 - 0x3f
    "00111111", --  284 - 0x11c  :   63 - 0x3f
    "00111111", --  285 - 0x11d  :   63 - 0x3f
    "00111111", --  286 - 0x11e  :   63 - 0x3f
    "00111111", --  287 - 0x11f  :   63 - 0x3f
    "00111111", --  288 - 0x120  :   63 - 0x3f -- line 0x9
    "00111111", --  289 - 0x121  :   63 - 0x3f
    "00111111", --  290 - 0x122  :   63 - 0x3f
    "00111111", --  291 - 0x123  :   63 - 0x3f
    "00111111", --  292 - 0x124  :   63 - 0x3f
    "00111111", --  293 - 0x125  :   63 - 0x3f
    "00111111", --  294 - 0x126  :   63 - 0x3f
    "00111111", --  295 - 0x127  :   63 - 0x3f
    "00111111", --  296 - 0x128  :   63 - 0x3f
    "00111111", --  297 - 0x129  :   63 - 0x3f
    "00111111", --  298 - 0x12a  :   63 - 0x3f
    "00111111", --  299 - 0x12b  :   63 - 0x3f
    "00111111", --  300 - 0x12c  :   63 - 0x3f
    "00111111", --  301 - 0x12d  :   63 - 0x3f
    "00111111", --  302 - 0x12e  :   63 - 0x3f
    "00111111", --  303 - 0x12f  :   63 - 0x3f
    "00111111", --  304 - 0x130  :   63 - 0x3f
    "00111111", --  305 - 0x131  :   63 - 0x3f
    "00111111", --  306 - 0x132  :   63 - 0x3f
    "00111111", --  307 - 0x133  :   63 - 0x3f
    "00001101", --  308 - 0x134  :   13 - 0xd
    "00001111", --  309 - 0x135  :   15 - 0xf
    "00111111", --  310 - 0x136  :   63 - 0x3f
    "00111111", --  311 - 0x137  :   63 - 0x3f
    "00111111", --  312 - 0x138  :   63 - 0x3f
    "00111111", --  313 - 0x139  :   63 - 0x3f
    "00111111", --  314 - 0x13a  :   63 - 0x3f
    "00111111", --  315 - 0x13b  :   63 - 0x3f
    "00111111", --  316 - 0x13c  :   63 - 0x3f
    "00111111", --  317 - 0x13d  :   63 - 0x3f
    "00111111", --  318 - 0x13e  :   63 - 0x3f
    "00111111", --  319 - 0x13f  :   63 - 0x3f
    "00111111", --  320 - 0x140  :   63 - 0x3f -- line 0xa
    "00111111", --  321 - 0x141  :   63 - 0x3f
    "00111111", --  322 - 0x142  :   63 - 0x3f
    "00111111", --  323 - 0x143  :   63 - 0x3f
    "00111111", --  324 - 0x144  :   63 - 0x3f
    "00111111", --  325 - 0x145  :   63 - 0x3f
    "00111111", --  326 - 0x146  :   63 - 0x3f
    "00111111", --  327 - 0x147  :   63 - 0x3f
    "00111111", --  328 - 0x148  :   63 - 0x3f
    "00111111", --  329 - 0x149  :   63 - 0x3f
    "00111111", --  330 - 0x14a  :   63 - 0x3f
    "00111111", --  331 - 0x14b  :   63 - 0x3f
    "00111111", --  332 - 0x14c  :   63 - 0x3f
    "00111111", --  333 - 0x14d  :   63 - 0x3f
    "00111111", --  334 - 0x14e  :   63 - 0x3f
    "00111111", --  335 - 0x14f  :   63 - 0x3f
    "00111111", --  336 - 0x150  :   63 - 0x3f
    "00111111", --  337 - 0x151  :   63 - 0x3f
    "00111111", --  338 - 0x152  :   63 - 0x3f
    "00111111", --  339 - 0x153  :   63 - 0x3f
    "01010111", --  340 - 0x154  :   87 - 0x57
    "01011000", --  341 - 0x155  :   88 - 0x58
    "01011000", --  342 - 0x156  :   88 - 0x58
    "01011000", --  343 - 0x157  :   88 - 0x58
    "01011000", --  344 - 0x158  :   88 - 0x58
    "01011000", --  345 - 0x159  :   88 - 0x58
    "01011000", --  346 - 0x15a  :   88 - 0x58
    "01011000", --  347 - 0x15b  :   88 - 0x58
    "01011000", --  348 - 0x15c  :   88 - 0x58
    "01011000", --  349 - 0x15d  :   88 - 0x58
    "01011000", --  350 - 0x15e  :   88 - 0x58
    "01011000", --  351 - 0x15f  :   88 - 0x58
    "00111111", --  352 - 0x160  :   63 - 0x3f -- line 0xb
    "00111111", --  353 - 0x161  :   63 - 0x3f
    "00111111", --  354 - 0x162  :   63 - 0x3f
    "00111111", --  355 - 0x163  :   63 - 0x3f
    "00111111", --  356 - 0x164  :   63 - 0x3f
    "00111111", --  357 - 0x165  :   63 - 0x3f
    "00111111", --  358 - 0x166  :   63 - 0x3f
    "00111111", --  359 - 0x167  :   63 - 0x3f
    "00111111", --  360 - 0x168  :   63 - 0x3f
    "00111111", --  361 - 0x169  :   63 - 0x3f
    "00111111", --  362 - 0x16a  :   63 - 0x3f
    "00111111", --  363 - 0x16b  :   63 - 0x3f
    "00111111", --  364 - 0x16c  :   63 - 0x3f
    "00111111", --  365 - 0x16d  :   63 - 0x3f
    "00111111", --  366 - 0x16e  :   63 - 0x3f
    "00111111", --  367 - 0x16f  :   63 - 0x3f
    "00111111", --  368 - 0x170  :   63 - 0x3f
    "00111111", --  369 - 0x171  :   63 - 0x3f
    "00111111", --  370 - 0x172  :   63 - 0x3f
    "00111111", --  371 - 0x173  :   63 - 0x3f
    "00111111", --  372 - 0x174  :   63 - 0x3f
    "00111111", --  373 - 0x175  :   63 - 0x3f
    "00111111", --  374 - 0x176  :   63 - 0x3f
    "00111111", --  375 - 0x177  :   63 - 0x3f
    "00111111", --  376 - 0x178  :   63 - 0x3f
    "00111111", --  377 - 0x179  :   63 - 0x3f
    "00111111", --  378 - 0x17a  :   63 - 0x3f
    "00111111", --  379 - 0x17b  :   63 - 0x3f
    "00111111", --  380 - 0x17c  :   63 - 0x3f
    "00111111", --  381 - 0x17d  :   63 - 0x3f
    "00111111", --  382 - 0x17e  :   63 - 0x3f
    "00111111", --  383 - 0x17f  :   63 - 0x3f
    "00111111", --  384 - 0x180  :   63 - 0x3f -- line 0xc
    "00111111", --  385 - 0x181  :   63 - 0x3f
    "00111111", --  386 - 0x182  :   63 - 0x3f
    "00111111", --  387 - 0x183  :   63 - 0x3f
    "00111111", --  388 - 0x184  :   63 - 0x3f
    "00111111", --  389 - 0x185  :   63 - 0x3f
    "00111111", --  390 - 0x186  :   63 - 0x3f
    "00111111", --  391 - 0x187  :   63 - 0x3f
    "00111111", --  392 - 0x188  :   63 - 0x3f
    "00111111", --  393 - 0x189  :   63 - 0x3f
    "00111111", --  394 - 0x18a  :   63 - 0x3f
    "00111111", --  395 - 0x18b  :   63 - 0x3f
    "00111111", --  396 - 0x18c  :   63 - 0x3f
    "00111111", --  397 - 0x18d  :   63 - 0x3f
    "00111111", --  398 - 0x18e  :   63 - 0x3f
    "00111111", --  399 - 0x18f  :   63 - 0x3f
    "00111111", --  400 - 0x190  :   63 - 0x3f
    "00111111", --  401 - 0x191  :   63 - 0x3f
    "00111111", --  402 - 0x192  :   63 - 0x3f
    "00111111", --  403 - 0x193  :   63 - 0x3f
    "00111111", --  404 - 0x194  :   63 - 0x3f
    "00111111", --  405 - 0x195  :   63 - 0x3f
    "00111111", --  406 - 0x196  :   63 - 0x3f
    "00111111", --  407 - 0x197  :   63 - 0x3f
    "00111111", --  408 - 0x198  :   63 - 0x3f
    "00111111", --  409 - 0x199  :   63 - 0x3f
    "00111111", --  410 - 0x19a  :   63 - 0x3f
    "00111111", --  411 - 0x19b  :   63 - 0x3f
    "00111111", --  412 - 0x19c  :   63 - 0x3f
    "00111111", --  413 - 0x19d  :   63 - 0x3f
    "00111111", --  414 - 0x19e  :   63 - 0x3f
    "00111111", --  415 - 0x19f  :   63 - 0x3f
    "00111111", --  416 - 0x1a0  :   63 - 0x3f -- line 0xd
    "00111111", --  417 - 0x1a1  :   63 - 0x3f
    "00111111", --  418 - 0x1a2  :   63 - 0x3f
    "00111111", --  419 - 0x1a3  :   63 - 0x3f
    "00111111", --  420 - 0x1a4  :   63 - 0x3f
    "00111111", --  421 - 0x1a5  :   63 - 0x3f
    "00111111", --  422 - 0x1a6  :   63 - 0x3f
    "00111111", --  423 - 0x1a7  :   63 - 0x3f
    "00111111", --  424 - 0x1a8  :   63 - 0x3f
    "00111111", --  425 - 0x1a9  :   63 - 0x3f
    "00111111", --  426 - 0x1aa  :   63 - 0x3f
    "00111111", --  427 - 0x1ab  :   63 - 0x3f
    "00111111", --  428 - 0x1ac  :   63 - 0x3f
    "00111111", --  429 - 0x1ad  :   63 - 0x3f
    "00111111", --  430 - 0x1ae  :   63 - 0x3f
    "00111111", --  431 - 0x1af  :   63 - 0x3f
    "00111111", --  432 - 0x1b0  :   63 - 0x3f
    "00111111", --  433 - 0x1b1  :   63 - 0x3f
    "00111111", --  434 - 0x1b2  :   63 - 0x3f
    "00111111", --  435 - 0x1b3  :   63 - 0x3f
    "00111111", --  436 - 0x1b4  :   63 - 0x3f
    "00111111", --  437 - 0x1b5  :   63 - 0x3f
    "00111111", --  438 - 0x1b6  :   63 - 0x3f
    "00111111", --  439 - 0x1b7  :   63 - 0x3f
    "00111111", --  440 - 0x1b8  :   63 - 0x3f
    "00111111", --  441 - 0x1b9  :   63 - 0x3f
    "00111111", --  442 - 0x1ba  :   63 - 0x3f
    "00111111", --  443 - 0x1bb  :   63 - 0x3f
    "00111111", --  444 - 0x1bc  :   63 - 0x3f
    "00111111", --  445 - 0x1bd  :   63 - 0x3f
    "00111111", --  446 - 0x1be  :   63 - 0x3f
    "00111111", --  447 - 0x1bf  :   63 - 0x3f
    "00111111", --  448 - 0x1c0  :   63 - 0x3f -- line 0xe
    "00111111", --  449 - 0x1c1  :   63 - 0x3f
    "00111111", --  450 - 0x1c2  :   63 - 0x3f
    "00111111", --  451 - 0x1c3  :   63 - 0x3f
    "00111111", --  452 - 0x1c4  :   63 - 0x3f
    "00111111", --  453 - 0x1c5  :   63 - 0x3f
    "00111111", --  454 - 0x1c6  :   63 - 0x3f
    "00111111", --  455 - 0x1c7  :   63 - 0x3f
    "00111111", --  456 - 0x1c8  :   63 - 0x3f
    "00111111", --  457 - 0x1c9  :   63 - 0x3f
    "00111111", --  458 - 0x1ca  :   63 - 0x3f
    "00111111", --  459 - 0x1cb  :   63 - 0x3f
    "00111111", --  460 - 0x1cc  :   63 - 0x3f
    "00111111", --  461 - 0x1cd  :   63 - 0x3f
    "00111111", --  462 - 0x1ce  :   63 - 0x3f
    "00111111", --  463 - 0x1cf  :   63 - 0x3f
    "00111111", --  464 - 0x1d0  :   63 - 0x3f
    "00111111", --  465 - 0x1d1  :   63 - 0x3f
    "00111111", --  466 - 0x1d2  :   63 - 0x3f
    "00111111", --  467 - 0x1d3  :   63 - 0x3f
    "00111111", --  468 - 0x1d4  :   63 - 0x3f
    "00111111", --  469 - 0x1d5  :   63 - 0x3f
    "00111111", --  470 - 0x1d6  :   63 - 0x3f
    "00111111", --  471 - 0x1d7  :   63 - 0x3f
    "00111111", --  472 - 0x1d8  :   63 - 0x3f
    "00111111", --  473 - 0x1d9  :   63 - 0x3f
    "00111111", --  474 - 0x1da  :   63 - 0x3f
    "00111111", --  475 - 0x1db  :   63 - 0x3f
    "00111111", --  476 - 0x1dc  :   63 - 0x3f
    "00111111", --  477 - 0x1dd  :   63 - 0x3f
    "00111111", --  478 - 0x1de  :   63 - 0x3f
    "00111111", --  479 - 0x1df  :   63 - 0x3f
    "00111111", --  480 - 0x1e0  :   63 - 0x3f -- line 0xf
    "00111111", --  481 - 0x1e1  :   63 - 0x3f
    "00111111", --  482 - 0x1e2  :   63 - 0x3f
    "00111111", --  483 - 0x1e3  :   63 - 0x3f
    "00111111", --  484 - 0x1e4  :   63 - 0x3f
    "00111111", --  485 - 0x1e5  :   63 - 0x3f
    "00111111", --  486 - 0x1e6  :   63 - 0x3f
    "00111111", --  487 - 0x1e7  :   63 - 0x3f
    "00111111", --  488 - 0x1e8  :   63 - 0x3f
    "00111111", --  489 - 0x1e9  :   63 - 0x3f
    "00111111", --  490 - 0x1ea  :   63 - 0x3f
    "00111111", --  491 - 0x1eb  :   63 - 0x3f
    "00111111", --  492 - 0x1ec  :   63 - 0x3f
    "00111111", --  493 - 0x1ed  :   63 - 0x3f
    "00111111", --  494 - 0x1ee  :   63 - 0x3f
    "00111111", --  495 - 0x1ef  :   63 - 0x3f
    "00111111", --  496 - 0x1f0  :   63 - 0x3f
    "00111111", --  497 - 0x1f1  :   63 - 0x3f
    "00111111", --  498 - 0x1f2  :   63 - 0x3f
    "00111111", --  499 - 0x1f3  :   63 - 0x3f
    "00111111", --  500 - 0x1f4  :   63 - 0x3f
    "00111111", --  501 - 0x1f5  :   63 - 0x3f
    "00111111", --  502 - 0x1f6  :   63 - 0x3f
    "00111111", --  503 - 0x1f7  :   63 - 0x3f
    "00111111", --  504 - 0x1f8  :   63 - 0x3f
    "00111111", --  505 - 0x1f9  :   63 - 0x3f
    "00111111", --  506 - 0x1fa  :   63 - 0x3f
    "00111111", --  507 - 0x1fb  :   63 - 0x3f
    "00111111", --  508 - 0x1fc  :   63 - 0x3f
    "00111111", --  509 - 0x1fd  :   63 - 0x3f
    "00111111", --  510 - 0x1fe  :   63 - 0x3f
    "00111111", --  511 - 0x1ff  :   63 - 0x3f
    "00111111", --  512 - 0x200  :   63 - 0x3f -- line 0x10
    "00111111", --  513 - 0x201  :   63 - 0x3f
    "00111111", --  514 - 0x202  :   63 - 0x3f
    "00111111", --  515 - 0x203  :   63 - 0x3f
    "00111111", --  516 - 0x204  :   63 - 0x3f
    "00111111", --  517 - 0x205  :   63 - 0x3f
    "00111111", --  518 - 0x206  :   63 - 0x3f
    "00111111", --  519 - 0x207  :   63 - 0x3f
    "00111111", --  520 - 0x208  :   63 - 0x3f
    "00111111", --  521 - 0x209  :   63 - 0x3f
    "00111111", --  522 - 0x20a  :   63 - 0x3f
    "00111111", --  523 - 0x20b  :   63 - 0x3f
    "00111111", --  524 - 0x20c  :   63 - 0x3f
    "00111111", --  525 - 0x20d  :   63 - 0x3f
    "00111111", --  526 - 0x20e  :   63 - 0x3f
    "00111111", --  527 - 0x20f  :   63 - 0x3f
    "00111111", --  528 - 0x210  :   63 - 0x3f
    "00111111", --  529 - 0x211  :   63 - 0x3f
    "00111111", --  530 - 0x212  :   63 - 0x3f
    "00111111", --  531 - 0x213  :   63 - 0x3f
    "00111111", --  532 - 0x214  :   63 - 0x3f
    "00111111", --  533 - 0x215  :   63 - 0x3f
    "00111111", --  534 - 0x216  :   63 - 0x3f
    "00111111", --  535 - 0x217  :   63 - 0x3f
    "00111111", --  536 - 0x218  :   63 - 0x3f
    "00111111", --  537 - 0x219  :   63 - 0x3f
    "00111111", --  538 - 0x21a  :   63 - 0x3f
    "00111111", --  539 - 0x21b  :   63 - 0x3f
    "00111111", --  540 - 0x21c  :   63 - 0x3f
    "00111111", --  541 - 0x21d  :   63 - 0x3f
    "00111111", --  542 - 0x21e  :   63 - 0x3f
    "00111111", --  543 - 0x21f  :   63 - 0x3f
    "00111111", --  544 - 0x220  :   63 - 0x3f -- line 0x11
    "00111111", --  545 - 0x221  :   63 - 0x3f
    "00111111", --  546 - 0x222  :   63 - 0x3f
    "00111111", --  547 - 0x223  :   63 - 0x3f
    "00111111", --  548 - 0x224  :   63 - 0x3f
    "00111111", --  549 - 0x225  :   63 - 0x3f
    "00111111", --  550 - 0x226  :   63 - 0x3f
    "00111111", --  551 - 0x227  :   63 - 0x3f
    "00111111", --  552 - 0x228  :   63 - 0x3f
    "00111111", --  553 - 0x229  :   63 - 0x3f
    "00111111", --  554 - 0x22a  :   63 - 0x3f
    "00111111", --  555 - 0x22b  :   63 - 0x3f
    "00111111", --  556 - 0x22c  :   63 - 0x3f
    "00111111", --  557 - 0x22d  :   63 - 0x3f
    "00111111", --  558 - 0x22e  :   63 - 0x3f
    "00111111", --  559 - 0x22f  :   63 - 0x3f
    "00111111", --  560 - 0x230  :   63 - 0x3f
    "00111111", --  561 - 0x231  :   63 - 0x3f
    "00111111", --  562 - 0x232  :   63 - 0x3f
    "00111111", --  563 - 0x233  :   63 - 0x3f
    "00111111", --  564 - 0x234  :   63 - 0x3f
    "00111111", --  565 - 0x235  :   63 - 0x3f
    "00111111", --  566 - 0x236  :   63 - 0x3f
    "00111111", --  567 - 0x237  :   63 - 0x3f
    "00111111", --  568 - 0x238  :   63 - 0x3f
    "00111111", --  569 - 0x239  :   63 - 0x3f
    "00111111", --  570 - 0x23a  :   63 - 0x3f
    "00111111", --  571 - 0x23b  :   63 - 0x3f
    "00111111", --  572 - 0x23c  :   63 - 0x3f
    "00111111", --  573 - 0x23d  :   63 - 0x3f
    "00111111", --  574 - 0x23e  :   63 - 0x3f
    "00111111", --  575 - 0x23f  :   63 - 0x3f
    "00111111", --  576 - 0x240  :   63 - 0x3f -- line 0x12
    "00111111", --  577 - 0x241  :   63 - 0x3f
    "00111111", --  578 - 0x242  :   63 - 0x3f
    "00111111", --  579 - 0x243  :   63 - 0x3f
    "00111111", --  580 - 0x244  :   63 - 0x3f
    "00111111", --  581 - 0x245  :   63 - 0x3f
    "00111111", --  582 - 0x246  :   63 - 0x3f
    "00111111", --  583 - 0x247  :   63 - 0x3f
    "00111111", --  584 - 0x248  :   63 - 0x3f
    "00111111", --  585 - 0x249  :   63 - 0x3f
    "00111111", --  586 - 0x24a  :   63 - 0x3f
    "00111111", --  587 - 0x24b  :   63 - 0x3f
    "00111111", --  588 - 0x24c  :   63 - 0x3f
    "00111111", --  589 - 0x24d  :   63 - 0x3f
    "00111111", --  590 - 0x24e  :   63 - 0x3f
    "00111111", --  591 - 0x24f  :   63 - 0x3f
    "00000000", --  592 - 0x250  :    0 - 0x0
    "00000010", --  593 - 0x251  :    2 - 0x2
    "00000000", --  594 - 0x252  :    0 - 0x0
    "00000010", --  595 - 0x253  :    2 - 0x2
    "00000000", --  596 - 0x254  :    0 - 0x0
    "00000010", --  597 - 0x255  :    2 - 0x2
    "00000100", --  598 - 0x256  :    4 - 0x4
    "00000110", --  599 - 0x257  :    6 - 0x6
    "00000000", --  600 - 0x258  :    0 - 0x0
    "00000010", --  601 - 0x259  :    2 - 0x2
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000010", --  603 - 0x25b  :    2 - 0x2
    "00000100", --  604 - 0x25c  :    4 - 0x4
    "00000110", --  605 - 0x25d  :    6 - 0x6
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000010", --  607 - 0x25f  :    2 - 0x2
    "00111111", --  608 - 0x260  :   63 - 0x3f -- line 0x13
    "00111111", --  609 - 0x261  :   63 - 0x3f
    "00111111", --  610 - 0x262  :   63 - 0x3f
    "00111111", --  611 - 0x263  :   63 - 0x3f
    "00111111", --  612 - 0x264  :   63 - 0x3f
    "00111111", --  613 - 0x265  :   63 - 0x3f
    "00111111", --  614 - 0x266  :   63 - 0x3f
    "00111111", --  615 - 0x267  :   63 - 0x3f
    "00111111", --  616 - 0x268  :   63 - 0x3f
    "00111111", --  617 - 0x269  :   63 - 0x3f
    "00111111", --  618 - 0x26a  :   63 - 0x3f
    "00111111", --  619 - 0x26b  :   63 - 0x3f
    "00111111", --  620 - 0x26c  :   63 - 0x3f
    "00111111", --  621 - 0x26d  :   63 - 0x3f
    "00111111", --  622 - 0x26e  :   63 - 0x3f
    "00111111", --  623 - 0x26f  :   63 - 0x3f
    "00000001", --  624 - 0x270  :    1 - 0x1
    "00000011", --  625 - 0x271  :    3 - 0x3
    "00000001", --  626 - 0x272  :    1 - 0x1
    "00000011", --  627 - 0x273  :    3 - 0x3
    "00000001", --  628 - 0x274  :    1 - 0x1
    "00000011", --  629 - 0x275  :    3 - 0x3
    "00000101", --  630 - 0x276  :    5 - 0x5
    "00000111", --  631 - 0x277  :    7 - 0x7
    "00000001", --  632 - 0x278  :    1 - 0x1
    "00000011", --  633 - 0x279  :    3 - 0x3
    "00000001", --  634 - 0x27a  :    1 - 0x1
    "00000011", --  635 - 0x27b  :    3 - 0x3
    "00000101", --  636 - 0x27c  :    5 - 0x5
    "00000111", --  637 - 0x27d  :    7 - 0x7
    "00000001", --  638 - 0x27e  :    1 - 0x1
    "00000011", --  639 - 0x27f  :    3 - 0x3
    "00111111", --  640 - 0x280  :   63 - 0x3f -- line 0x14
    "00111111", --  641 - 0x281  :   63 - 0x3f
    "00111111", --  642 - 0x282  :   63 - 0x3f
    "00111111", --  643 - 0x283  :   63 - 0x3f
    "00111111", --  644 - 0x284  :   63 - 0x3f
    "00111111", --  645 - 0x285  :   63 - 0x3f
    "00111111", --  646 - 0x286  :   63 - 0x3f
    "00111111", --  647 - 0x287  :   63 - 0x3f
    "00111111", --  648 - 0x288  :   63 - 0x3f
    "00111111", --  649 - 0x289  :   63 - 0x3f
    "00111111", --  650 - 0x28a  :   63 - 0x3f
    "00111111", --  651 - 0x28b  :   63 - 0x3f
    "00111111", --  652 - 0x28c  :   63 - 0x3f
    "00111111", --  653 - 0x28d  :   63 - 0x3f
    "00111111", --  654 - 0x28e  :   63 - 0x3f
    "00111111", --  655 - 0x28f  :   63 - 0x3f
    "00111111", --  656 - 0x290  :   63 - 0x3f
    "00111111", --  657 - 0x291  :   63 - 0x3f
    "00111111", --  658 - 0x292  :   63 - 0x3f
    "00111111", --  659 - 0x293  :   63 - 0x3f
    "00111111", --  660 - 0x294  :   63 - 0x3f
    "00111111", --  661 - 0x295  :   63 - 0x3f
    "00111111", --  662 - 0x296  :   63 - 0x3f
    "00111111", --  663 - 0x297  :   63 - 0x3f
    "00111111", --  664 - 0x298  :   63 - 0x3f
    "00111111", --  665 - 0x299  :   63 - 0x3f
    "00111111", --  666 - 0x29a  :   63 - 0x3f
    "00111111", --  667 - 0x29b  :   63 - 0x3f
    "00111111", --  668 - 0x29c  :   63 - 0x3f
    "00111111", --  669 - 0x29d  :   63 - 0x3f
    "00111111", --  670 - 0x29e  :   63 - 0x3f
    "00111111", --  671 - 0x29f  :   63 - 0x3f
    "00111111", --  672 - 0x2a0  :   63 - 0x3f -- line 0x15
    "00111111", --  673 - 0x2a1  :   63 - 0x3f
    "00111111", --  674 - 0x2a2  :   63 - 0x3f
    "00111111", --  675 - 0x2a3  :   63 - 0x3f
    "00111111", --  676 - 0x2a4  :   63 - 0x3f
    "00111111", --  677 - 0x2a5  :   63 - 0x3f
    "00111111", --  678 - 0x2a6  :   63 - 0x3f
    "00111111", --  679 - 0x2a7  :   63 - 0x3f
    "00111111", --  680 - 0x2a8  :   63 - 0x3f
    "00111111", --  681 - 0x2a9  :   63 - 0x3f
    "00111111", --  682 - 0x2aa  :   63 - 0x3f
    "00111111", --  683 - 0x2ab  :   63 - 0x3f
    "00111111", --  684 - 0x2ac  :   63 - 0x3f
    "00111111", --  685 - 0x2ad  :   63 - 0x3f
    "00111111", --  686 - 0x2ae  :   63 - 0x3f
    "00111111", --  687 - 0x2af  :   63 - 0x3f
    "00111111", --  688 - 0x2b0  :   63 - 0x3f
    "00111111", --  689 - 0x2b1  :   63 - 0x3f
    "00111111", --  690 - 0x2b2  :   63 - 0x3f
    "00111111", --  691 - 0x2b3  :   63 - 0x3f
    "00111111", --  692 - 0x2b4  :   63 - 0x3f
    "00111111", --  693 - 0x2b5  :   63 - 0x3f
    "00111111", --  694 - 0x2b6  :   63 - 0x3f
    "00111111", --  695 - 0x2b7  :   63 - 0x3f
    "00111111", --  696 - 0x2b8  :   63 - 0x3f
    "00111111", --  697 - 0x2b9  :   63 - 0x3f
    "00111111", --  698 - 0x2ba  :   63 - 0x3f
    "00111111", --  699 - 0x2bb  :   63 - 0x3f
    "00111111", --  700 - 0x2bc  :   63 - 0x3f
    "00111111", --  701 - 0x2bd  :   63 - 0x3f
    "00111111", --  702 - 0x2be  :   63 - 0x3f
    "00111111", --  703 - 0x2bf  :   63 - 0x3f
    "00111111", --  704 - 0x2c0  :   63 - 0x3f -- line 0x16
    "00111111", --  705 - 0x2c1  :   63 - 0x3f
    "00111111", --  706 - 0x2c2  :   63 - 0x3f
    "00111111", --  707 - 0x2c3  :   63 - 0x3f
    "00111111", --  708 - 0x2c4  :   63 - 0x3f
    "00111111", --  709 - 0x2c5  :   63 - 0x3f
    "00111111", --  710 - 0x2c6  :   63 - 0x3f
    "00111111", --  711 - 0x2c7  :   63 - 0x3f
    "00111111", --  712 - 0x2c8  :   63 - 0x3f
    "00111111", --  713 - 0x2c9  :   63 - 0x3f
    "00111111", --  714 - 0x2ca  :   63 - 0x3f
    "00111111", --  715 - 0x2cb  :   63 - 0x3f
    "00111111", --  716 - 0x2cc  :   63 - 0x3f
    "00111111", --  717 - 0x2cd  :   63 - 0x3f
    "00111111", --  718 - 0x2ce  :   63 - 0x3f
    "00111111", --  719 - 0x2cf  :   63 - 0x3f
    "00111111", --  720 - 0x2d0  :   63 - 0x3f
    "00111111", --  721 - 0x2d1  :   63 - 0x3f
    "00111111", --  722 - 0x2d2  :   63 - 0x3f
    "00111111", --  723 - 0x2d3  :   63 - 0x3f
    "00111111", --  724 - 0x2d4  :   63 - 0x3f
    "00111111", --  725 - 0x2d5  :   63 - 0x3f
    "00111111", --  726 - 0x2d6  :   63 - 0x3f
    "00111111", --  727 - 0x2d7  :   63 - 0x3f
    "00111111", --  728 - 0x2d8  :   63 - 0x3f
    "00111111", --  729 - 0x2d9  :   63 - 0x3f
    "00111111", --  730 - 0x2da  :   63 - 0x3f
    "00111111", --  731 - 0x2db  :   63 - 0x3f
    "00111111", --  732 - 0x2dc  :   63 - 0x3f
    "00111111", --  733 - 0x2dd  :   63 - 0x3f
    "00111111", --  734 - 0x2de  :   63 - 0x3f
    "00111111", --  735 - 0x2df  :   63 - 0x3f
    "00111111", --  736 - 0x2e0  :   63 - 0x3f -- line 0x17
    "00111111", --  737 - 0x2e1  :   63 - 0x3f
    "00111111", --  738 - 0x2e2  :   63 - 0x3f
    "00111111", --  739 - 0x2e3  :   63 - 0x3f
    "00111111", --  740 - 0x2e4  :   63 - 0x3f
    "00111111", --  741 - 0x2e5  :   63 - 0x3f
    "00111111", --  742 - 0x2e6  :   63 - 0x3f
    "00111111", --  743 - 0x2e7  :   63 - 0x3f
    "00111111", --  744 - 0x2e8  :   63 - 0x3f
    "00111111", --  745 - 0x2e9  :   63 - 0x3f
    "00111111", --  746 - 0x2ea  :   63 - 0x3f
    "00111111", --  747 - 0x2eb  :   63 - 0x3f
    "00111111", --  748 - 0x2ec  :   63 - 0x3f
    "00111111", --  749 - 0x2ed  :   63 - 0x3f
    "00111111", --  750 - 0x2ee  :   63 - 0x3f
    "00111111", --  751 - 0x2ef  :   63 - 0x3f
    "11000101", --  752 - 0x2f0  :  197 - 0xc5
    "11010110", --  753 - 0x2f1  :  214 - 0xd6
    "11000101", --  754 - 0x2f2  :  197 - 0xc5
    "11010110", --  755 - 0x2f3  :  214 - 0xd6
    "11000101", --  756 - 0x2f4  :  197 - 0xc5
    "11010110", --  757 - 0x2f5  :  214 - 0xd6
    "11000101", --  758 - 0x2f6  :  197 - 0xc5
    "11010110", --  759 - 0x2f7  :  214 - 0xd6
    "11000101", --  760 - 0x2f8  :  197 - 0xc5
    "11010110", --  761 - 0x2f9  :  214 - 0xd6
    "11000101", --  762 - 0x2fa  :  197 - 0xc5
    "11010110", --  763 - 0x2fb  :  214 - 0xd6
    "11000101", --  764 - 0x2fc  :  197 - 0xc5
    "11010110", --  765 - 0x2fd  :  214 - 0xd6
    "11000101", --  766 - 0x2fe  :  197 - 0xc5
    "11010110", --  767 - 0x2ff  :  214 - 0xd6
    "00111111", --  768 - 0x300  :   63 - 0x3f -- line 0x18
    "00111111", --  769 - 0x301  :   63 - 0x3f
    "00111111", --  770 - 0x302  :   63 - 0x3f
    "00111111", --  771 - 0x303  :   63 - 0x3f
    "00011100", --  772 - 0x304  :   28 - 0x1c
    "00011110", --  773 - 0x305  :   30 - 0x1e
    "00111111", --  774 - 0x306  :   63 - 0x3f
    "00111111", --  775 - 0x307  :   63 - 0x3f
    "00111111", --  776 - 0x308  :   63 - 0x3f
    "00111111", --  777 - 0x309  :   63 - 0x3f
    "00111111", --  778 - 0x30a  :   63 - 0x3f
    "00111111", --  779 - 0x30b  :   63 - 0x3f
    "00111111", --  780 - 0x30c  :   63 - 0x3f
    "00111111", --  781 - 0x30d  :   63 - 0x3f
    "00111111", --  782 - 0x30e  :   63 - 0x3f
    "00111111", --  783 - 0x30f  :   63 - 0x3f
    "11000111", --  784 - 0x310  :  199 - 0xc7
    "11001001", --  785 - 0x311  :  201 - 0xc9
    "11000111", --  786 - 0x312  :  199 - 0xc7
    "11001001", --  787 - 0x313  :  201 - 0xc9
    "11000111", --  788 - 0x314  :  199 - 0xc7
    "11001001", --  789 - 0x315  :  201 - 0xc9
    "11000111", --  790 - 0x316  :  199 - 0xc7
    "11001001", --  791 - 0x317  :  201 - 0xc9
    "11000111", --  792 - 0x318  :  199 - 0xc7
    "11001001", --  793 - 0x319  :  201 - 0xc9
    "11000111", --  794 - 0x31a  :  199 - 0xc7
    "11001001", --  795 - 0x31b  :  201 - 0xc9
    "11000111", --  796 - 0x31c  :  199 - 0xc7
    "11001001", --  797 - 0x31d  :  201 - 0xc9
    "11000111", --  798 - 0x31e  :  199 - 0xc7
    "11001001", --  799 - 0x31f  :  201 - 0xc9
    "00111111", --  800 - 0x320  :   63 - 0x3f -- line 0x19
    "00111111", --  801 - 0x321  :   63 - 0x3f
    "00111111", --  802 - 0x322  :   63 - 0x3f
    "00111111", --  803 - 0x323  :   63 - 0x3f
    "00011101", --  804 - 0x324  :   29 - 0x1d
    "00011111", --  805 - 0x325  :   31 - 0x1f
    "00111111", --  806 - 0x326  :   63 - 0x3f
    "00111111", --  807 - 0x327  :   63 - 0x3f
    "00111111", --  808 - 0x328  :   63 - 0x3f
    "00111111", --  809 - 0x329  :   63 - 0x3f
    "00111111", --  810 - 0x32a  :   63 - 0x3f
    "00111111", --  811 - 0x32b  :   63 - 0x3f
    "00111111", --  812 - 0x32c  :   63 - 0x3f
    "00111111", --  813 - 0x32d  :   63 - 0x3f
    "00111111", --  814 - 0x32e  :   63 - 0x3f
    "00111111", --  815 - 0x32f  :   63 - 0x3f
    "11010111", --  816 - 0x330  :  215 - 0xd7
    "11011001", --  817 - 0x331  :  217 - 0xd9
    "11010111", --  818 - 0x332  :  215 - 0xd7
    "11011001", --  819 - 0x333  :  217 - 0xd9
    "11010111", --  820 - 0x334  :  215 - 0xd7
    "11011001", --  821 - 0x335  :  217 - 0xd9
    "11010111", --  822 - 0x336  :  215 - 0xd7
    "11011001", --  823 - 0x337  :  217 - 0xd9
    "11010111", --  824 - 0x338  :  215 - 0xd7
    "11011001", --  825 - 0x339  :  217 - 0xd9
    "11010111", --  826 - 0x33a  :  215 - 0xd7
    "11011001", --  827 - 0x33b  :  217 - 0xd9
    "11010111", --  828 - 0x33c  :  215 - 0xd7
    "11011001", --  829 - 0x33d  :  217 - 0xd9
    "11010111", --  830 - 0x33e  :  215 - 0xd7
    "11011001", --  831 - 0x33f  :  217 - 0xd9
    "01110000", --  832 - 0x340  :  112 - 0x70 -- line 0x1a
    "01110001", --  833 - 0x341  :  113 - 0x71
    "01110001", --  834 - 0x342  :  113 - 0x71
    "01110001", --  835 - 0x343  :  113 - 0x71
    "01110001", --  836 - 0x344  :  113 - 0x71
    "01110001", --  837 - 0x345  :  113 - 0x71
    "01110001", --  838 - 0x346  :  113 - 0x71
    "01110001", --  839 - 0x347  :  113 - 0x71
    "01110001", --  840 - 0x348  :  113 - 0x71
    "01110001", --  841 - 0x349  :  113 - 0x71
    "01110001", --  842 - 0x34a  :  113 - 0x71
    "01110001", --  843 - 0x34b  :  113 - 0x71
    "01110001", --  844 - 0x34c  :  113 - 0x71
    "01110001", --  845 - 0x34d  :  113 - 0x71
    "01110001", --  846 - 0x34e  :  113 - 0x71
    "01110001", --  847 - 0x34f  :  113 - 0x71
    "01110001", --  848 - 0x350  :  113 - 0x71
    "01110001", --  849 - 0x351  :  113 - 0x71
    "01110001", --  850 - 0x352  :  113 - 0x71
    "01110001", --  851 - 0x353  :  113 - 0x71
    "01110001", --  852 - 0x354  :  113 - 0x71
    "01110001", --  853 - 0x355  :  113 - 0x71
    "01110001", --  854 - 0x356  :  113 - 0x71
    "01110001", --  855 - 0x357  :  113 - 0x71
    "01110001", --  856 - 0x358  :  113 - 0x71
    "01110001", --  857 - 0x359  :  113 - 0x71
    "01110001", --  858 - 0x35a  :  113 - 0x71
    "01110001", --  859 - 0x35b  :  113 - 0x71
    "01110001", --  860 - 0x35c  :  113 - 0x71
    "01110001", --  861 - 0x35d  :  113 - 0x71
    "01110001", --  862 - 0x35e  :  113 - 0x71
    "01110001", --  863 - 0x35f  :  113 - 0x71
    "01100000", --  864 - 0x360  :   96 - 0x60 -- line 0x1b
    "01110111", --  865 - 0x361  :  119 - 0x77
    "01110111", --  866 - 0x362  :  119 - 0x77
    "01110111", --  867 - 0x363  :  119 - 0x77
    "01110111", --  868 - 0x364  :  119 - 0x77
    "01110111", --  869 - 0x365  :  119 - 0x77
    "01110111", --  870 - 0x366  :  119 - 0x77
    "01110111", --  871 - 0x367  :  119 - 0x77
    "01110111", --  872 - 0x368  :  119 - 0x77
    "01110111", --  873 - 0x369  :  119 - 0x77
    "01110111", --  874 - 0x36a  :  119 - 0x77
    "01110111", --  875 - 0x36b  :  119 - 0x77
    "01110111", --  876 - 0x36c  :  119 - 0x77
    "01110111", --  877 - 0x36d  :  119 - 0x77
    "01110111", --  878 - 0x36e  :  119 - 0x77
    "01110111", --  879 - 0x36f  :  119 - 0x77
    "01110111", --  880 - 0x370  :  119 - 0x77
    "01110111", --  881 - 0x371  :  119 - 0x77
    "01110111", --  882 - 0x372  :  119 - 0x77
    "01110111", --  883 - 0x373  :  119 - 0x77
    "01110111", --  884 - 0x374  :  119 - 0x77
    "01110111", --  885 - 0x375  :  119 - 0x77
    "01110111", --  886 - 0x376  :  119 - 0x77
    "01110111", --  887 - 0x377  :  119 - 0x77
    "01110111", --  888 - 0x378  :  119 - 0x77
    "01110111", --  889 - 0x379  :  119 - 0x77
    "01110111", --  890 - 0x37a  :  119 - 0x77
    "01110111", --  891 - 0x37b  :  119 - 0x77
    "01110111", --  892 - 0x37c  :  119 - 0x77
    "01110111", --  893 - 0x37d  :  119 - 0x77
    "01110111", --  894 - 0x37e  :  119 - 0x77
    "01110111", --  895 - 0x37f  :  119 - 0x77
    "01100000", --  896 - 0x380  :   96 - 0x60 -- line 0x1c
    "01110011", --  897 - 0x381  :  115 - 0x73
    "01110011", --  898 - 0x382  :  115 - 0x73
    "01110011", --  899 - 0x383  :  115 - 0x73
    "01110011", --  900 - 0x384  :  115 - 0x73
    "01110011", --  901 - 0x385  :  115 - 0x73
    "01110011", --  902 - 0x386  :  115 - 0x73
    "01110011", --  903 - 0x387  :  115 - 0x73
    "01110011", --  904 - 0x388  :  115 - 0x73
    "01110011", --  905 - 0x389  :  115 - 0x73
    "01110011", --  906 - 0x38a  :  115 - 0x73
    "01110011", --  907 - 0x38b  :  115 - 0x73
    "01110011", --  908 - 0x38c  :  115 - 0x73
    "01110011", --  909 - 0x38d  :  115 - 0x73
    "01110011", --  910 - 0x38e  :  115 - 0x73
    "01110011", --  911 - 0x38f  :  115 - 0x73
    "01110011", --  912 - 0x390  :  115 - 0x73
    "01110011", --  913 - 0x391  :  115 - 0x73
    "01110011", --  914 - 0x392  :  115 - 0x73
    "01110011", --  915 - 0x393  :  115 - 0x73
    "01110011", --  916 - 0x394  :  115 - 0x73
    "01110011", --  917 - 0x395  :  115 - 0x73
    "01110011", --  918 - 0x396  :  115 - 0x73
    "01110011", --  919 - 0x397  :  115 - 0x73
    "01110011", --  920 - 0x398  :  115 - 0x73
    "01110011", --  921 - 0x399  :  115 - 0x73
    "01110011", --  922 - 0x39a  :  115 - 0x73
    "01110011", --  923 - 0x39b  :  115 - 0x73
    "01110011", --  924 - 0x39c  :  115 - 0x73
    "01110011", --  925 - 0x39d  :  115 - 0x73
    "01110011", --  926 - 0x39e  :  115 - 0x73
    "01110011", --  927 - 0x39f  :  115 - 0x73
    "01100000", --  928 - 0x3a0  :   96 - 0x60 -- line 0x1d
    "01110011", --  929 - 0x3a1  :  115 - 0x73
    "01110011", --  930 - 0x3a2  :  115 - 0x73
    "01110011", --  931 - 0x3a3  :  115 - 0x73
    "01110011", --  932 - 0x3a4  :  115 - 0x73
    "01110011", --  933 - 0x3a5  :  115 - 0x73
    "01110011", --  934 - 0x3a6  :  115 - 0x73
    "01110011", --  935 - 0x3a7  :  115 - 0x73
    "01110011", --  936 - 0x3a8  :  115 - 0x73
    "01110011", --  937 - 0x3a9  :  115 - 0x73
    "01110011", --  938 - 0x3aa  :  115 - 0x73
    "01110011", --  939 - 0x3ab  :  115 - 0x73
    "01110011", --  940 - 0x3ac  :  115 - 0x73
    "01110011", --  941 - 0x3ad  :  115 - 0x73
    "01110011", --  942 - 0x3ae  :  115 - 0x73
    "01110011", --  943 - 0x3af  :  115 - 0x73
    "01110011", --  944 - 0x3b0  :  115 - 0x73
    "01110011", --  945 - 0x3b1  :  115 - 0x73
    "01110011", --  946 - 0x3b2  :  115 - 0x73
    "01110011", --  947 - 0x3b3  :  115 - 0x73
    "01110011", --  948 - 0x3b4  :  115 - 0x73
    "01110011", --  949 - 0x3b5  :  115 - 0x73
    "01110011", --  950 - 0x3b6  :  115 - 0x73
    "01110011", --  951 - 0x3b7  :  115 - 0x73
    "01110011", --  952 - 0x3b8  :  115 - 0x73
    "01110011", --  953 - 0x3b9  :  115 - 0x73
    "01110011", --  954 - 0x3ba  :  115 - 0x73
    "01110011", --  955 - 0x3bb  :  115 - 0x73
    "01110011", --  956 - 0x3bc  :  115 - 0x73
    "01110011", --  957 - 0x3bd  :  115 - 0x73
    "01110011", --  958 - 0x3be  :  115 - 0x73
    "01110011", --  959 - 0x3bf  :  115 - 0x73
        ---- Attribute Table 0----
    "00000000", --  960 - 0x3c0  :    0 - 0x0
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00001000", --  974 - 0x3ce  :    8 - 0x8
    "00001000", --  975 - 0x3cf  :    8 - 0x8
    "00000000", --  976 - 0x3d0  :    0 - 0x0
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "01010001", --  981 - 0x3d5  :   81 - 0x51
    "01010000", --  982 - 0x3d6  :   80 - 0x50
    "01010000", --  983 - 0x3d7  :   80 - 0x50
    "00000000", --  984 - 0x3d8  :    0 - 0x0
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "10100000", --  996 - 0x3e4  :  160 - 0xa0
    "10100000", --  997 - 0x3e5  :  160 - 0xa0
    "10100000", --  998 - 0x3e6  :  160 - 0xa0
    "10100000", --  999 - 0x3e7  :  160 - 0xa0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0
    "00000010", -- 1009 - 0x3f1  :    2 - 0x2
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000"  -- 1023 - 0x3ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
