//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables
//- Only the first Name Table: 1KiB


//-  Original memory dump file name: pacman_ntable_start.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_NTABLE0_PACMAN_START
  (
     //input     clk,   // clock
     input      [10-1:0] addr,  //1024 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      10'h0: dout  = 8'b00100000; //    0 :  32 - 0x20 -- line 0x0
      10'h1: dout  = 8'b00100000; //    1 :  32 - 0x20
      10'h2: dout  = 8'b00100000; //    2 :  32 - 0x20
      10'h3: dout  = 8'b00100000; //    3 :  32 - 0x20
      10'h4: dout  = 8'b00100000; //    4 :  32 - 0x20
      10'h5: dout  = 8'b00100000; //    5 :  32 - 0x20
      10'h6: dout  = 8'b00100000; //    6 :  32 - 0x20
      10'h7: dout  = 8'b00100000; //    7 :  32 - 0x20
      10'h8: dout  = 8'b00100000; //    8 :  32 - 0x20
      10'h9: dout  = 8'b00100000; //    9 :  32 - 0x20
      10'hA: dout  = 8'b00100000; //   10 :  32 - 0x20
      10'hB: dout  = 8'b00100000; //   11 :  32 - 0x20
      10'hC: dout  = 8'b00100000; //   12 :  32 - 0x20
      10'hD: dout  = 8'b00100000; //   13 :  32 - 0x20
      10'hE: dout  = 8'b00100000; //   14 :  32 - 0x20
      10'hF: dout  = 8'b00100000; //   15 :  32 - 0x20
      10'h10: dout  = 8'b00100000; //   16 :  32 - 0x20
      10'h11: dout  = 8'b00100000; //   17 :  32 - 0x20
      10'h12: dout  = 8'b00100000; //   18 :  32 - 0x20
      10'h13: dout  = 8'b00100000; //   19 :  32 - 0x20
      10'h14: dout  = 8'b00100000; //   20 :  32 - 0x20
      10'h15: dout  = 8'b00100000; //   21 :  32 - 0x20
      10'h16: dout  = 8'b00100000; //   22 :  32 - 0x20
      10'h17: dout  = 8'b00100000; //   23 :  32 - 0x20
      10'h18: dout  = 8'b00100000; //   24 :  32 - 0x20
      10'h19: dout  = 8'b00100000; //   25 :  32 - 0x20
      10'h1A: dout  = 8'b00100000; //   26 :  32 - 0x20
      10'h1B: dout  = 8'b00100000; //   27 :  32 - 0x20
      10'h1C: dout  = 8'b00100000; //   28 :  32 - 0x20
      10'h1D: dout  = 8'b00100000; //   29 :  32 - 0x20
      10'h1E: dout  = 8'b00100000; //   30 :  32 - 0x20
      10'h1F: dout  = 8'b00100000; //   31 :  32 - 0x20
      10'h20: dout  = 8'b00100000; //   32 :  32 - 0x20 -- line 0x1
      10'h21: dout  = 8'b00100000; //   33 :  32 - 0x20
      10'h22: dout  = 8'b00100000; //   34 :  32 - 0x20
      10'h23: dout  = 8'b00100000; //   35 :  32 - 0x20
      10'h24: dout  = 8'b00100000; //   36 :  32 - 0x20
      10'h25: dout  = 8'b00100000; //   37 :  32 - 0x20
      10'h26: dout  = 8'b00100000; //   38 :  32 - 0x20
      10'h27: dout  = 8'b00100000; //   39 :  32 - 0x20
      10'h28: dout  = 8'b00100000; //   40 :  32 - 0x20
      10'h29: dout  = 8'b00100000; //   41 :  32 - 0x20
      10'h2A: dout  = 8'b00100000; //   42 :  32 - 0x20
      10'h2B: dout  = 8'b00100000; //   43 :  32 - 0x20
      10'h2C: dout  = 8'b00100000; //   44 :  32 - 0x20
      10'h2D: dout  = 8'b00100000; //   45 :  32 - 0x20
      10'h2E: dout  = 8'b00100000; //   46 :  32 - 0x20
      10'h2F: dout  = 8'b00100000; //   47 :  32 - 0x20
      10'h30: dout  = 8'b00100000; //   48 :  32 - 0x20
      10'h31: dout  = 8'b00100000; //   49 :  32 - 0x20
      10'h32: dout  = 8'b00100000; //   50 :  32 - 0x20
      10'h33: dout  = 8'b00100000; //   51 :  32 - 0x20
      10'h34: dout  = 8'b00100000; //   52 :  32 - 0x20
      10'h35: dout  = 8'b00100000; //   53 :  32 - 0x20
      10'h36: dout  = 8'b00100000; //   54 :  32 - 0x20
      10'h37: dout  = 8'b00100000; //   55 :  32 - 0x20
      10'h38: dout  = 8'b00100000; //   56 :  32 - 0x20
      10'h39: dout  = 8'b00100000; //   57 :  32 - 0x20
      10'h3A: dout  = 8'b00100000; //   58 :  32 - 0x20
      10'h3B: dout  = 8'b00100000; //   59 :  32 - 0x20
      10'h3C: dout  = 8'b00100000; //   60 :  32 - 0x20
      10'h3D: dout  = 8'b00100000; //   61 :  32 - 0x20
      10'h3E: dout  = 8'b00100000; //   62 :  32 - 0x20
      10'h3F: dout  = 8'b00100000; //   63 :  32 - 0x20
      10'h40: dout  = 8'b00100000; //   64 :  32 - 0x20 -- line 0x2
      10'h41: dout  = 8'b00100000; //   65 :  32 - 0x20
      10'h42: dout  = 8'b00100000; //   66 :  32 - 0x20
      10'h43: dout  = 8'b00100000; //   67 :  32 - 0x20
      10'h44: dout  = 8'b00100000; //   68 :  32 - 0x20
      10'h45: dout  = 8'b00100000; //   69 :  32 - 0x20
      10'h46: dout  = 8'b00100000; //   70 :  32 - 0x20
      10'h47: dout  = 8'b00100000; //   71 :  32 - 0x20
      10'h48: dout  = 8'b00100000; //   72 :  32 - 0x20
      10'h49: dout  = 8'b00100000; //   73 :  32 - 0x20
      10'h4A: dout  = 8'b00100000; //   74 :  32 - 0x20
      10'h4B: dout  = 8'b00100000; //   75 :  32 - 0x20
      10'h4C: dout  = 8'b00100000; //   76 :  32 - 0x20
      10'h4D: dout  = 8'b00100000; //   77 :  32 - 0x20
      10'h4E: dout  = 8'b00100000; //   78 :  32 - 0x20
      10'h4F: dout  = 8'b00100000; //   79 :  32 - 0x20
      10'h50: dout  = 8'b00100000; //   80 :  32 - 0x20
      10'h51: dout  = 8'b00100000; //   81 :  32 - 0x20
      10'h52: dout  = 8'b00100000; //   82 :  32 - 0x20
      10'h53: dout  = 8'b00100000; //   83 :  32 - 0x20
      10'h54: dout  = 8'b00100000; //   84 :  32 - 0x20
      10'h55: dout  = 8'b00100000; //   85 :  32 - 0x20
      10'h56: dout  = 8'b00100000; //   86 :  32 - 0x20
      10'h57: dout  = 8'b00100000; //   87 :  32 - 0x20
      10'h58: dout  = 8'b00100000; //   88 :  32 - 0x20
      10'h59: dout  = 8'b00100000; //   89 :  32 - 0x20
      10'h5A: dout  = 8'b00100000; //   90 :  32 - 0x20
      10'h5B: dout  = 8'b00100000; //   91 :  32 - 0x20
      10'h5C: dout  = 8'b00100000; //   92 :  32 - 0x20
      10'h5D: dout  = 8'b00100000; //   93 :  32 - 0x20
      10'h5E: dout  = 8'b00100000; //   94 :  32 - 0x20
      10'h5F: dout  = 8'b00100000; //   95 :  32 - 0x20
      10'h60: dout  = 8'b00100000; //   96 :  32 - 0x20 -- line 0x3
      10'h61: dout  = 8'b00100000; //   97 :  32 - 0x20
      10'h62: dout  = 8'b00100000; //   98 :  32 - 0x20
      10'h63: dout  = 8'b00100000; //   99 :  32 - 0x20
      10'h64: dout  = 8'b00100000; //  100 :  32 - 0x20
      10'h65: dout  = 8'b10110000; //  101 : 176 - 0xb0
      10'h66: dout  = 8'b10110011; //  102 : 179 - 0xb3
      10'h67: dout  = 8'b10110010; //  103 : 178 - 0xb2
      10'h68: dout  = 8'b00100000; //  104 :  32 - 0x20
      10'h69: dout  = 8'b00100000; //  105 :  32 - 0x20
      10'h6A: dout  = 8'b00100000; //  106 :  32 - 0x20
      10'h6B: dout  = 8'b00100000; //  107 :  32 - 0x20
      10'h6C: dout  = 8'b10110100; //  108 : 180 - 0xb4
      10'h6D: dout  = 8'b10110101; //  109 : 181 - 0xb5
      10'h6E: dout  = 8'b10110110; //  110 : 182 - 0xb6
      10'h6F: dout  = 8'b10110111; //  111 : 183 - 0xb7
      10'h70: dout  = 8'b10111000; //  112 : 184 - 0xb8
      10'h71: dout  = 8'b10111001; //  113 : 185 - 0xb9
      10'h72: dout  = 8'b10111010; //  114 : 186 - 0xba
      10'h73: dout  = 8'b10111011; //  115 : 187 - 0xbb
      10'h74: dout  = 8'b00100000; //  116 :  32 - 0x20
      10'h75: dout  = 8'b00100000; //  117 :  32 - 0x20
      10'h76: dout  = 8'b00100000; //  118 :  32 - 0x20
      10'h77: dout  = 8'b10110001; //  119 : 177 - 0xb1
      10'h78: dout  = 8'b10110011; //  120 : 179 - 0xb3
      10'h79: dout  = 8'b10110010; //  121 : 178 - 0xb2
      10'h7A: dout  = 8'b00100000; //  122 :  32 - 0x20
      10'h7B: dout  = 8'b00100000; //  123 :  32 - 0x20
      10'h7C: dout  = 8'b00100000; //  124 :  32 - 0x20
      10'h7D: dout  = 8'b00100000; //  125 :  32 - 0x20
      10'h7E: dout  = 8'b00100000; //  126 :  32 - 0x20
      10'h7F: dout  = 8'b00100000; //  127 :  32 - 0x20
      10'h80: dout  = 8'b00100000; //  128 :  32 - 0x20 -- line 0x4
      10'h81: dout  = 8'b00100000; //  129 :  32 - 0x20
      10'h82: dout  = 8'b00100000; //  130 :  32 - 0x20
      10'h83: dout  = 8'b00100000; //  131 :  32 - 0x20
      10'h84: dout  = 8'b00100000; //  132 :  32 - 0x20
      10'h85: dout  = 8'b00100000; //  133 :  32 - 0x20
      10'h86: dout  = 8'b00100000; //  134 :  32 - 0x20
      10'h87: dout  = 8'b00100000; //  135 :  32 - 0x20
      10'h88: dout  = 8'b00110101; //  136 :  53 - 0x35
      10'h89: dout  = 8'b00110000; //  137 :  48 - 0x30
      10'h8A: dout  = 8'b00100000; //  138 :  32 - 0x20
      10'h8B: dout  = 8'b00100000; //  139 :  32 - 0x20
      10'h8C: dout  = 8'b00100000; //  140 :  32 - 0x20
      10'h8D: dout  = 8'b00100000; //  141 :  32 - 0x20
      10'h8E: dout  = 8'b00110001; //  142 :  49 - 0x31
      10'h8F: dout  = 8'b00110000; //  143 :  48 - 0x30
      10'h90: dout  = 8'b00110000; //  144 :  48 - 0x30
      10'h91: dout  = 8'b00110000; //  145 :  48 - 0x30
      10'h92: dout  = 8'b00110000; //  146 :  48 - 0x30
      10'h93: dout  = 8'b00100000; //  147 :  32 - 0x20
      10'h94: dout  = 8'b00100000; //  148 :  32 - 0x20
      10'h95: dout  = 8'b00100000; //  149 :  32 - 0x20
      10'h96: dout  = 8'b00100000; //  150 :  32 - 0x20
      10'h97: dout  = 8'b00100000; //  151 :  32 - 0x20
      10'h98: dout  = 8'b00100000; //  152 :  32 - 0x20
      10'h99: dout  = 8'b00100000; //  153 :  32 - 0x20
      10'h9A: dout  = 8'b00110000; //  154 :  48 - 0x30
      10'h9B: dout  = 8'b00110000; //  155 :  48 - 0x30
      10'h9C: dout  = 8'b00100000; //  156 :  32 - 0x20
      10'h9D: dout  = 8'b00100000; //  157 :  32 - 0x20
      10'h9E: dout  = 8'b00100000; //  158 :  32 - 0x20
      10'h9F: dout  = 8'b00100000; //  159 :  32 - 0x20
      10'hA0: dout  = 8'b00100000; //  160 :  32 - 0x20 -- line 0x5
      10'hA1: dout  = 8'b00100000; //  161 :  32 - 0x20
      10'hA2: dout  = 8'b00100000; //  162 :  32 - 0x20
      10'hA3: dout  = 8'b00100000; //  163 :  32 - 0x20
      10'hA4: dout  = 8'b00100000; //  164 :  32 - 0x20
      10'hA5: dout  = 8'b00100000; //  165 :  32 - 0x20
      10'hA6: dout  = 8'b00100000; //  166 :  32 - 0x20
      10'hA7: dout  = 8'b00100000; //  167 :  32 - 0x20
      10'hA8: dout  = 8'b00100000; //  168 :  32 - 0x20
      10'hA9: dout  = 8'b00100000; //  169 :  32 - 0x20
      10'hAA: dout  = 8'b00100000; //  170 :  32 - 0x20
      10'hAB: dout  = 8'b00100000; //  171 :  32 - 0x20
      10'hAC: dout  = 8'b00100000; //  172 :  32 - 0x20
      10'hAD: dout  = 8'b00100000; //  173 :  32 - 0x20
      10'hAE: dout  = 8'b00100000; //  174 :  32 - 0x20
      10'hAF: dout  = 8'b00100000; //  175 :  32 - 0x20
      10'hB0: dout  = 8'b00100000; //  176 :  32 - 0x20
      10'hB1: dout  = 8'b00100000; //  177 :  32 - 0x20
      10'hB2: dout  = 8'b00100000; //  178 :  32 - 0x20
      10'hB3: dout  = 8'b00100000; //  179 :  32 - 0x20
      10'hB4: dout  = 8'b00100000; //  180 :  32 - 0x20
      10'hB5: dout  = 8'b00100000; //  181 :  32 - 0x20
      10'hB6: dout  = 8'b00100000; //  182 :  32 - 0x20
      10'hB7: dout  = 8'b00100000; //  183 :  32 - 0x20
      10'hB8: dout  = 8'b00100000; //  184 :  32 - 0x20
      10'hB9: dout  = 8'b00100000; //  185 :  32 - 0x20
      10'hBA: dout  = 8'b00100000; //  186 :  32 - 0x20
      10'hBB: dout  = 8'b00100000; //  187 :  32 - 0x20
      10'hBC: dout  = 8'b00100000; //  188 :  32 - 0x20
      10'hBD: dout  = 8'b00100000; //  189 :  32 - 0x20
      10'hBE: dout  = 8'b00100000; //  190 :  32 - 0x20
      10'hBF: dout  = 8'b00100000; //  191 :  32 - 0x20
      10'hC0: dout  = 8'b00100000; //  192 :  32 - 0x20 -- line 0x6
      10'hC1: dout  = 8'b00100000; //  193 :  32 - 0x20
      10'hC2: dout  = 8'b00100000; //  194 :  32 - 0x20
      10'hC3: dout  = 8'b00100000; //  195 :  32 - 0x20
      10'hC4: dout  = 8'b00100000; //  196 :  32 - 0x20
      10'hC5: dout  = 8'b00100000; //  197 :  32 - 0x20
      10'hC6: dout  = 8'b00100000; //  198 :  32 - 0x20
      10'hC7: dout  = 8'b00100000; //  199 :  32 - 0x20
      10'hC8: dout  = 8'b00100000; //  200 :  32 - 0x20
      10'hC9: dout  = 8'b00100000; //  201 :  32 - 0x20
      10'hCA: dout  = 8'b00100000; //  202 :  32 - 0x20
      10'hCB: dout  = 8'b00100000; //  203 :  32 - 0x20
      10'hCC: dout  = 8'b00100000; //  204 :  32 - 0x20
      10'hCD: dout  = 8'b00100000; //  205 :  32 - 0x20
      10'hCE: dout  = 8'b00100000; //  206 :  32 - 0x20
      10'hCF: dout  = 8'b00100000; //  207 :  32 - 0x20
      10'hD0: dout  = 8'b00100000; //  208 :  32 - 0x20
      10'hD1: dout  = 8'b00100000; //  209 :  32 - 0x20
      10'hD2: dout  = 8'b00100000; //  210 :  32 - 0x20
      10'hD3: dout  = 8'b00100000; //  211 :  32 - 0x20
      10'hD4: dout  = 8'b00100000; //  212 :  32 - 0x20
      10'hD5: dout  = 8'b00100000; //  213 :  32 - 0x20
      10'hD6: dout  = 8'b00100000; //  214 :  32 - 0x20
      10'hD7: dout  = 8'b00100000; //  215 :  32 - 0x20
      10'hD8: dout  = 8'b00100000; //  216 :  32 - 0x20
      10'hD9: dout  = 8'b00100000; //  217 :  32 - 0x20
      10'hDA: dout  = 8'b00100000; //  218 :  32 - 0x20
      10'hDB: dout  = 8'b00100000; //  219 :  32 - 0x20
      10'hDC: dout  = 8'b00100000; //  220 :  32 - 0x20
      10'hDD: dout  = 8'b00100000; //  221 :  32 - 0x20
      10'hDE: dout  = 8'b00100000; //  222 :  32 - 0x20
      10'hDF: dout  = 8'b00100000; //  223 :  32 - 0x20
      10'hE0: dout  = 8'b00100000; //  224 :  32 - 0x20 -- line 0x7
      10'hE1: dout  = 8'b00100000; //  225 :  32 - 0x20
      10'hE2: dout  = 8'b00100000; //  226 :  32 - 0x20
      10'hE3: dout  = 8'b00100000; //  227 :  32 - 0x20
      10'hE4: dout  = 8'b00100000; //  228 :  32 - 0x20
      10'hE5: dout  = 8'b11100100; //  229 : 228 - 0xe4
      10'hE6: dout  = 8'b11101000; //  230 : 232 - 0xe8
      10'hE7: dout  = 8'b11101000; //  231 : 232 - 0xe8
      10'hE8: dout  = 8'b11101000; //  232 : 232 - 0xe8
      10'hE9: dout  = 8'b11101000; //  233 : 232 - 0xe8
      10'hEA: dout  = 8'b11101000; //  234 : 232 - 0xe8
      10'hEB: dout  = 8'b11101000; //  235 : 232 - 0xe8
      10'hEC: dout  = 8'b11101000; //  236 : 232 - 0xe8
      10'hED: dout  = 8'b11101000; //  237 : 232 - 0xe8
      10'hEE: dout  = 8'b11101000; //  238 : 232 - 0xe8
      10'hEF: dout  = 8'b11101000; //  239 : 232 - 0xe8
      10'hF0: dout  = 8'b11101000; //  240 : 232 - 0xe8
      10'hF1: dout  = 8'b11101000; //  241 : 232 - 0xe8
      10'hF2: dout  = 8'b11101000; //  242 : 232 - 0xe8
      10'hF3: dout  = 8'b11101000; //  243 : 232 - 0xe8
      10'hF4: dout  = 8'b11101000; //  244 : 232 - 0xe8
      10'hF5: dout  = 8'b11101000; //  245 : 232 - 0xe8
      10'hF6: dout  = 8'b11101000; //  246 : 232 - 0xe8
      10'hF7: dout  = 8'b11101000; //  247 : 232 - 0xe8
      10'hF8: dout  = 8'b11101000; //  248 : 232 - 0xe8
      10'hF9: dout  = 8'b11101000; //  249 : 232 - 0xe8
      10'hFA: dout  = 8'b11101000; //  250 : 232 - 0xe8
      10'hFB: dout  = 8'b11100101; //  251 : 229 - 0xe5
      10'hFC: dout  = 8'b00100000; //  252 :  32 - 0x20
      10'hFD: dout  = 8'b00100000; //  253 :  32 - 0x20
      10'hFE: dout  = 8'b00100000; //  254 :  32 - 0x20
      10'hFF: dout  = 8'b00100000; //  255 :  32 - 0x20
      10'h100: dout  = 8'b00100000; //  256 :  32 - 0x20 -- line 0x8
      10'h101: dout  = 8'b00100000; //  257 :  32 - 0x20
      10'h102: dout  = 8'b00100000; //  258 :  32 - 0x20
      10'h103: dout  = 8'b00100000; //  259 :  32 - 0x20
      10'h104: dout  = 8'b00100000; //  260 :  32 - 0x20
      10'h105: dout  = 8'b11101011; //  261 : 235 - 0xeb
      10'h106: dout  = 8'b10001000; //  262 : 136 - 0x88
      10'h107: dout  = 8'b10000000; //  263 : 128 - 0x80
      10'h108: dout  = 8'b10000001; //  264 : 129 - 0x81
      10'h109: dout  = 8'b10000010; //  265 : 130 - 0x82
      10'h10A: dout  = 8'b10000011; //  266 : 131 - 0x83
      10'h10B: dout  = 8'b10000100; //  267 : 132 - 0x84
      10'h10C: dout  = 8'b10000101; //  268 : 133 - 0x85
      10'h10D: dout  = 8'b10000110; //  269 : 134 - 0x86
      10'h10E: dout  = 8'b10000111; //  270 : 135 - 0x87
      10'h10F: dout  = 8'b10001000; //  271 : 136 - 0x88
      10'h110: dout  = 8'b10001000; //  272 : 136 - 0x88
      10'h111: dout  = 8'b10001001; //  273 : 137 - 0x89
      10'h112: dout  = 8'b10001010; //  274 : 138 - 0x8a
      10'h113: dout  = 8'b10001011; //  275 : 139 - 0x8b
      10'h114: dout  = 8'b10001100; //  276 : 140 - 0x8c
      10'h115: dout  = 8'b10001101; //  277 : 141 - 0x8d
      10'h116: dout  = 8'b10001110; //  278 : 142 - 0x8e
      10'h117: dout  = 8'b10001111; //  279 : 143 - 0x8f
      10'h118: dout  = 8'b10010000; //  280 : 144 - 0x90
      10'h119: dout  = 8'b10010001; //  281 : 145 - 0x91
      10'h11A: dout  = 8'b10100011; //  282 : 163 - 0xa3
      10'h11B: dout  = 8'b11101001; //  283 : 233 - 0xe9
      10'h11C: dout  = 8'b00100000; //  284 :  32 - 0x20
      10'h11D: dout  = 8'b00100000; //  285 :  32 - 0x20
      10'h11E: dout  = 8'b00100000; //  286 :  32 - 0x20
      10'h11F: dout  = 8'b00100000; //  287 :  32 - 0x20
      10'h120: dout  = 8'b00100000; //  288 :  32 - 0x20 -- line 0x9
      10'h121: dout  = 8'b00100000; //  289 :  32 - 0x20
      10'h122: dout  = 8'b00100000; //  290 :  32 - 0x20
      10'h123: dout  = 8'b00100000; //  291 :  32 - 0x20
      10'h124: dout  = 8'b00100000; //  292 :  32 - 0x20
      10'h125: dout  = 8'b11101011; //  293 : 235 - 0xeb
      10'h126: dout  = 8'b10001000; //  294 : 136 - 0x88
      10'h127: dout  = 8'b10010010; //  295 : 146 - 0x92
      10'h128: dout  = 8'b10010011; //  296 : 147 - 0x93
      10'h129: dout  = 8'b10010100; //  297 : 148 - 0x94
      10'h12A: dout  = 8'b10010101; //  298 : 149 - 0x95
      10'h12B: dout  = 8'b10010110; //  299 : 150 - 0x96
      10'h12C: dout  = 8'b10010111; //  300 : 151 - 0x97
      10'h12D: dout  = 8'b10011000; //  301 : 152 - 0x98
      10'h12E: dout  = 8'b10011001; //  302 : 153 - 0x99
      10'h12F: dout  = 8'b10011010; //  303 : 154 - 0x9a
      10'h130: dout  = 8'b10011011; //  304 : 155 - 0x9b
      10'h131: dout  = 8'b10011100; //  305 : 156 - 0x9c
      10'h132: dout  = 8'b10011101; //  306 : 157 - 0x9d
      10'h133: dout  = 8'b10011110; //  307 : 158 - 0x9e
      10'h134: dout  = 8'b10011111; //  308 : 159 - 0x9f
      10'h135: dout  = 8'b10100000; //  309 : 160 - 0xa0
      10'h136: dout  = 8'b10100001; //  310 : 161 - 0xa1
      10'h137: dout  = 8'b10100010; //  311 : 162 - 0xa2
      10'h138: dout  = 8'b10100011; //  312 : 163 - 0xa3
      10'h139: dout  = 8'b10100100; //  313 : 164 - 0xa4
      10'h13A: dout  = 8'b10100011; //  314 : 163 - 0xa3
      10'h13B: dout  = 8'b11101001; //  315 : 233 - 0xe9
      10'h13C: dout  = 8'b00100000; //  316 :  32 - 0x20
      10'h13D: dout  = 8'b00100000; //  317 :  32 - 0x20
      10'h13E: dout  = 8'b00100000; //  318 :  32 - 0x20
      10'h13F: dout  = 8'b00100000; //  319 :  32 - 0x20
      10'h140: dout  = 8'b00100000; //  320 :  32 - 0x20 -- line 0xa
      10'h141: dout  = 8'b00100000; //  321 :  32 - 0x20
      10'h142: dout  = 8'b00100000; //  322 :  32 - 0x20
      10'h143: dout  = 8'b00100000; //  323 :  32 - 0x20
      10'h144: dout  = 8'b00100000; //  324 :  32 - 0x20
      10'h145: dout  = 8'b11101011; //  325 : 235 - 0xeb
      10'h146: dout  = 8'b10001000; //  326 : 136 - 0x88
      10'h147: dout  = 8'b10010010; //  327 : 146 - 0x92
      10'h148: dout  = 8'b10100101; //  328 : 165 - 0xa5
      10'h149: dout  = 8'b10100110; //  329 : 166 - 0xa6
      10'h14A: dout  = 8'b10100111; //  330 : 167 - 0xa7
      10'h14B: dout  = 8'b10101000; //  331 : 168 - 0xa8
      10'h14C: dout  = 8'b10101001; //  332 : 169 - 0xa9
      10'h14D: dout  = 8'b10101010; //  333 : 170 - 0xaa
      10'h14E: dout  = 8'b10101011; //  334 : 171 - 0xab
      10'h14F: dout  = 8'b10101100; //  335 : 172 - 0xac
      10'h150: dout  = 8'b10101101; //  336 : 173 - 0xad
      10'h151: dout  = 8'b10101110; //  337 : 174 - 0xae
      10'h152: dout  = 8'b10100011; //  338 : 163 - 0xa3
      10'h153: dout  = 8'b10101111; //  339 : 175 - 0xaf
      10'h154: dout  = 8'b11010000; //  340 : 208 - 0xd0
      10'h155: dout  = 8'b11010001; //  341 : 209 - 0xd1
      10'h156: dout  = 8'b11010010; //  342 : 210 - 0xd2
      10'h157: dout  = 8'b10100011; //  343 : 163 - 0xa3
      10'h158: dout  = 8'b11010011; //  344 : 211 - 0xd3
      10'h159: dout  = 8'b10100100; //  345 : 164 - 0xa4
      10'h15A: dout  = 8'b10100011; //  346 : 163 - 0xa3
      10'h15B: dout  = 8'b11101001; //  347 : 233 - 0xe9
      10'h15C: dout  = 8'b00100000; //  348 :  32 - 0x20
      10'h15D: dout  = 8'b00100000; //  349 :  32 - 0x20
      10'h15E: dout  = 8'b00100000; //  350 :  32 - 0x20
      10'h15F: dout  = 8'b00100000; //  351 :  32 - 0x20
      10'h160: dout  = 8'b00100000; //  352 :  32 - 0x20 -- line 0xb
      10'h161: dout  = 8'b00100000; //  353 :  32 - 0x20
      10'h162: dout  = 8'b00100000; //  354 :  32 - 0x20
      10'h163: dout  = 8'b00100000; //  355 :  32 - 0x20
      10'h164: dout  = 8'b00100000; //  356 :  32 - 0x20
      10'h165: dout  = 8'b11101011; //  357 : 235 - 0xeb
      10'h166: dout  = 8'b10001000; //  358 : 136 - 0x88
      10'h167: dout  = 8'b11010100; //  359 : 212 - 0xd4
      10'h168: dout  = 8'b11010101; //  360 : 213 - 0xd5
      10'h169: dout  = 8'b11010110; //  361 : 214 - 0xd6
      10'h16A: dout  = 8'b11010111; //  362 : 215 - 0xd7
      10'h16B: dout  = 8'b11011000; //  363 : 216 - 0xd8
      10'h16C: dout  = 8'b11011001; //  364 : 217 - 0xd9
      10'h16D: dout  = 8'b11011010; //  365 : 218 - 0xda
      10'h16E: dout  = 8'b11011011; //  366 : 219 - 0xdb
      10'h16F: dout  = 8'b10001000; //  367 : 136 - 0x88
      10'h170: dout  = 8'b10001000; //  368 : 136 - 0x88
      10'h171: dout  = 8'b11011100; //  369 : 220 - 0xdc
      10'h172: dout  = 8'b11010111; //  370 : 215 - 0xd7
      10'h173: dout  = 8'b11011101; //  371 : 221 - 0xdd
      10'h174: dout  = 8'b11011110; //  372 : 222 - 0xde
      10'h175: dout  = 8'b11011111; //  373 : 223 - 0xdf
      10'h176: dout  = 8'b11100000; //  374 : 224 - 0xe0
      10'h177: dout  = 8'b11100001; //  375 : 225 - 0xe1
      10'h178: dout  = 8'b11100010; //  376 : 226 - 0xe2
      10'h179: dout  = 8'b11100011; //  377 : 227 - 0xe3
      10'h17A: dout  = 8'b10100011; //  378 : 163 - 0xa3
      10'h17B: dout  = 8'b11101001; //  379 : 233 - 0xe9
      10'h17C: dout  = 8'b00100000; //  380 :  32 - 0x20
      10'h17D: dout  = 8'b00100000; //  381 :  32 - 0x20
      10'h17E: dout  = 8'b00100000; //  382 :  32 - 0x20
      10'h17F: dout  = 8'b00100000; //  383 :  32 - 0x20
      10'h180: dout  = 8'b00100000; //  384 :  32 - 0x20 -- line 0xc
      10'h181: dout  = 8'b00100000; //  385 :  32 - 0x20
      10'h182: dout  = 8'b00100000; //  386 :  32 - 0x20
      10'h183: dout  = 8'b00100000; //  387 :  32 - 0x20
      10'h184: dout  = 8'b00100000; //  388 :  32 - 0x20
      10'h185: dout  = 8'b11100111; //  389 : 231 - 0xe7
      10'h186: dout  = 8'b11101010; //  390 : 234 - 0xea
      10'h187: dout  = 8'b11101010; //  391 : 234 - 0xea
      10'h188: dout  = 8'b11101010; //  392 : 234 - 0xea
      10'h189: dout  = 8'b11101010; //  393 : 234 - 0xea
      10'h18A: dout  = 8'b11101010; //  394 : 234 - 0xea
      10'h18B: dout  = 8'b11101010; //  395 : 234 - 0xea
      10'h18C: dout  = 8'b11101010; //  396 : 234 - 0xea
      10'h18D: dout  = 8'b11101010; //  397 : 234 - 0xea
      10'h18E: dout  = 8'b11101010; //  398 : 234 - 0xea
      10'h18F: dout  = 8'b11101010; //  399 : 234 - 0xea
      10'h190: dout  = 8'b11101010; //  400 : 234 - 0xea
      10'h191: dout  = 8'b11101010; //  401 : 234 - 0xea
      10'h192: dout  = 8'b11101010; //  402 : 234 - 0xea
      10'h193: dout  = 8'b11101010; //  403 : 234 - 0xea
      10'h194: dout  = 8'b11101010; //  404 : 234 - 0xea
      10'h195: dout  = 8'b11101010; //  405 : 234 - 0xea
      10'h196: dout  = 8'b11101010; //  406 : 234 - 0xea
      10'h197: dout  = 8'b11101010; //  407 : 234 - 0xea
      10'h198: dout  = 8'b11101010; //  408 : 234 - 0xea
      10'h199: dout  = 8'b11101010; //  409 : 234 - 0xea
      10'h19A: dout  = 8'b11101010; //  410 : 234 - 0xea
      10'h19B: dout  = 8'b11100110; //  411 : 230 - 0xe6
      10'h19C: dout  = 8'b00100000; //  412 :  32 - 0x20
      10'h19D: dout  = 8'b00100000; //  413 :  32 - 0x20
      10'h19E: dout  = 8'b00100000; //  414 :  32 - 0x20
      10'h19F: dout  = 8'b00100000; //  415 :  32 - 0x20
      10'h1A0: dout  = 8'b00100000; //  416 :  32 - 0x20 -- line 0xd
      10'h1A1: dout  = 8'b00100000; //  417 :  32 - 0x20
      10'h1A2: dout  = 8'b00100000; //  418 :  32 - 0x20
      10'h1A3: dout  = 8'b00100000; //  419 :  32 - 0x20
      10'h1A4: dout  = 8'b00100000; //  420 :  32 - 0x20
      10'h1A5: dout  = 8'b00100000; //  421 :  32 - 0x20
      10'h1A6: dout  = 8'b00100000; //  422 :  32 - 0x20
      10'h1A7: dout  = 8'b00100000; //  423 :  32 - 0x20
      10'h1A8: dout  = 8'b00100000; //  424 :  32 - 0x20
      10'h1A9: dout  = 8'b00100000; //  425 :  32 - 0x20
      10'h1AA: dout  = 8'b00100000; //  426 :  32 - 0x20
      10'h1AB: dout  = 8'b00100000; //  427 :  32 - 0x20
      10'h1AC: dout  = 8'b00100000; //  428 :  32 - 0x20
      10'h1AD: dout  = 8'b00100000; //  429 :  32 - 0x20
      10'h1AE: dout  = 8'b00100000; //  430 :  32 - 0x20
      10'h1AF: dout  = 8'b00100000; //  431 :  32 - 0x20
      10'h1B0: dout  = 8'b00100000; //  432 :  32 - 0x20
      10'h1B1: dout  = 8'b00100000; //  433 :  32 - 0x20
      10'h1B2: dout  = 8'b00100000; //  434 :  32 - 0x20
      10'h1B3: dout  = 8'b00100000; //  435 :  32 - 0x20
      10'h1B4: dout  = 8'b00100000; //  436 :  32 - 0x20
      10'h1B5: dout  = 8'b00100000; //  437 :  32 - 0x20
      10'h1B6: dout  = 8'b00100000; //  438 :  32 - 0x20
      10'h1B7: dout  = 8'b00100000; //  439 :  32 - 0x20
      10'h1B8: dout  = 8'b00100000; //  440 :  32 - 0x20
      10'h1B9: dout  = 8'b00100000; //  441 :  32 - 0x20
      10'h1BA: dout  = 8'b00100000; //  442 :  32 - 0x20
      10'h1BB: dout  = 8'b00100000; //  443 :  32 - 0x20
      10'h1BC: dout  = 8'b00100000; //  444 :  32 - 0x20
      10'h1BD: dout  = 8'b00100000; //  445 :  32 - 0x20
      10'h1BE: dout  = 8'b00100000; //  446 :  32 - 0x20
      10'h1BF: dout  = 8'b00100000; //  447 :  32 - 0x20
      10'h1C0: dout  = 8'b00100000; //  448 :  32 - 0x20 -- line 0xe
      10'h1C1: dout  = 8'b00100000; //  449 :  32 - 0x20
      10'h1C2: dout  = 8'b00100000; //  450 :  32 - 0x20
      10'h1C3: dout  = 8'b00100000; //  451 :  32 - 0x20
      10'h1C4: dout  = 8'b00100000; //  452 :  32 - 0x20
      10'h1C5: dout  = 8'b00100000; //  453 :  32 - 0x20
      10'h1C6: dout  = 8'b00100000; //  454 :  32 - 0x20
      10'h1C7: dout  = 8'b00100000; //  455 :  32 - 0x20
      10'h1C8: dout  = 8'b00100000; //  456 :  32 - 0x20
      10'h1C9: dout  = 8'b00100000; //  457 :  32 - 0x20
      10'h1CA: dout  = 8'b00100000; //  458 :  32 - 0x20
      10'h1CB: dout  = 8'b00100000; //  459 :  32 - 0x20
      10'h1CC: dout  = 8'b00100000; //  460 :  32 - 0x20
      10'h1CD: dout  = 8'b00100000; //  461 :  32 - 0x20
      10'h1CE: dout  = 8'b00100000; //  462 :  32 - 0x20
      10'h1CF: dout  = 8'b00100000; //  463 :  32 - 0x20
      10'h1D0: dout  = 8'b00100000; //  464 :  32 - 0x20
      10'h1D1: dout  = 8'b00100000; //  465 :  32 - 0x20
      10'h1D2: dout  = 8'b00100000; //  466 :  32 - 0x20
      10'h1D3: dout  = 8'b00100000; //  467 :  32 - 0x20
      10'h1D4: dout  = 8'b00100000; //  468 :  32 - 0x20
      10'h1D5: dout  = 8'b00100000; //  469 :  32 - 0x20
      10'h1D6: dout  = 8'b00100000; //  470 :  32 - 0x20
      10'h1D7: dout  = 8'b00100000; //  471 :  32 - 0x20
      10'h1D8: dout  = 8'b00100000; //  472 :  32 - 0x20
      10'h1D9: dout  = 8'b00100000; //  473 :  32 - 0x20
      10'h1DA: dout  = 8'b00100000; //  474 :  32 - 0x20
      10'h1DB: dout  = 8'b00100000; //  475 :  32 - 0x20
      10'h1DC: dout  = 8'b00100000; //  476 :  32 - 0x20
      10'h1DD: dout  = 8'b00100000; //  477 :  32 - 0x20
      10'h1DE: dout  = 8'b00100000; //  478 :  32 - 0x20
      10'h1DF: dout  = 8'b00100000; //  479 :  32 - 0x20
      10'h1E0: dout  = 8'b00100000; //  480 :  32 - 0x20 -- line 0xf
      10'h1E1: dout  = 8'b00100000; //  481 :  32 - 0x20
      10'h1E2: dout  = 8'b00100000; //  482 :  32 - 0x20
      10'h1E3: dout  = 8'b00100000; //  483 :  32 - 0x20
      10'h1E4: dout  = 8'b00100000; //  484 :  32 - 0x20
      10'h1E5: dout  = 8'b00100000; //  485 :  32 - 0x20
      10'h1E6: dout  = 8'b00100000; //  486 :  32 - 0x20
      10'h1E7: dout  = 8'b00100000; //  487 :  32 - 0x20
      10'h1E8: dout  = 8'b00100000; //  488 :  32 - 0x20
      10'h1E9: dout  = 8'b00100000; //  489 :  32 - 0x20
      10'h1EA: dout  = 8'b00100000; //  490 :  32 - 0x20
      10'h1EB: dout  = 8'b00100000; //  491 :  32 - 0x20
      10'h1EC: dout  = 8'b00100000; //  492 :  32 - 0x20
      10'h1ED: dout  = 8'b00100000; //  493 :  32 - 0x20
      10'h1EE: dout  = 8'b00100000; //  494 :  32 - 0x20
      10'h1EF: dout  = 8'b00100000; //  495 :  32 - 0x20
      10'h1F0: dout  = 8'b00100000; //  496 :  32 - 0x20
      10'h1F1: dout  = 8'b00100000; //  497 :  32 - 0x20
      10'h1F2: dout  = 8'b00100000; //  498 :  32 - 0x20
      10'h1F3: dout  = 8'b00100000; //  499 :  32 - 0x20
      10'h1F4: dout  = 8'b00100000; //  500 :  32 - 0x20
      10'h1F5: dout  = 8'b00100000; //  501 :  32 - 0x20
      10'h1F6: dout  = 8'b00100000; //  502 :  32 - 0x20
      10'h1F7: dout  = 8'b00100000; //  503 :  32 - 0x20
      10'h1F8: dout  = 8'b00100000; //  504 :  32 - 0x20
      10'h1F9: dout  = 8'b00100000; //  505 :  32 - 0x20
      10'h1FA: dout  = 8'b00100000; //  506 :  32 - 0x20
      10'h1FB: dout  = 8'b00100000; //  507 :  32 - 0x20
      10'h1FC: dout  = 8'b00100000; //  508 :  32 - 0x20
      10'h1FD: dout  = 8'b00100000; //  509 :  32 - 0x20
      10'h1FE: dout  = 8'b00100000; //  510 :  32 - 0x20
      10'h1FF: dout  = 8'b00100000; //  511 :  32 - 0x20
      10'h200: dout  = 8'b00100000; //  512 :  32 - 0x20 -- line 0x10
      10'h201: dout  = 8'b00100000; //  513 :  32 - 0x20
      10'h202: dout  = 8'b00100000; //  514 :  32 - 0x20
      10'h203: dout  = 8'b00100000; //  515 :  32 - 0x20
      10'h204: dout  = 8'b00100000; //  516 :  32 - 0x20
      10'h205: dout  = 8'b00100000; //  517 :  32 - 0x20
      10'h206: dout  = 8'b00100000; //  518 :  32 - 0x20
      10'h207: dout  = 8'b00100000; //  519 :  32 - 0x20
      10'h208: dout  = 8'b00100000; //  520 :  32 - 0x20
      10'h209: dout  = 8'b00100000; //  521 :  32 - 0x20
      10'h20A: dout  = 8'b01011100; //  522 :  92 - 0x5c
      10'h20B: dout  = 8'b00100000; //  523 :  32 - 0x20
      10'h20C: dout  = 8'b00110001; //  524 :  49 - 0x31
      10'h20D: dout  = 8'b00100000; //  525 :  32 - 0x20
      10'h20E: dout  = 8'b01010000; //  526 :  80 - 0x50
      10'h20F: dout  = 8'b01001100; //  527 :  76 - 0x4c
      10'h210: dout  = 8'b01000001; //  528 :  65 - 0x41
      10'h211: dout  = 8'b01011001; //  529 :  89 - 0x59
      10'h212: dout  = 8'b01000101; //  530 :  69 - 0x45
      10'h213: dout  = 8'b01010010; //  531 :  82 - 0x52
      10'h214: dout  = 8'b00100000; //  532 :  32 - 0x20
      10'h215: dout  = 8'b00100000; //  533 :  32 - 0x20
      10'h216: dout  = 8'b00100000; //  534 :  32 - 0x20
      10'h217: dout  = 8'b00100000; //  535 :  32 - 0x20
      10'h218: dout  = 8'b00100000; //  536 :  32 - 0x20
      10'h219: dout  = 8'b00100000; //  537 :  32 - 0x20
      10'h21A: dout  = 8'b00100000; //  538 :  32 - 0x20
      10'h21B: dout  = 8'b00100000; //  539 :  32 - 0x20
      10'h21C: dout  = 8'b00100000; //  540 :  32 - 0x20
      10'h21D: dout  = 8'b00100000; //  541 :  32 - 0x20
      10'h21E: dout  = 8'b00100000; //  542 :  32 - 0x20
      10'h21F: dout  = 8'b00100000; //  543 :  32 - 0x20
      10'h220: dout  = 8'b00100000; //  544 :  32 - 0x20 -- line 0x11
      10'h221: dout  = 8'b00100000; //  545 :  32 - 0x20
      10'h222: dout  = 8'b00100000; //  546 :  32 - 0x20
      10'h223: dout  = 8'b00100000; //  547 :  32 - 0x20
      10'h224: dout  = 8'b00100000; //  548 :  32 - 0x20
      10'h225: dout  = 8'b00100000; //  549 :  32 - 0x20
      10'h226: dout  = 8'b00100000; //  550 :  32 - 0x20
      10'h227: dout  = 8'b00100000; //  551 :  32 - 0x20
      10'h228: dout  = 8'b00100000; //  552 :  32 - 0x20
      10'h229: dout  = 8'b00100000; //  553 :  32 - 0x20
      10'h22A: dout  = 8'b00100000; //  554 :  32 - 0x20
      10'h22B: dout  = 8'b00100000; //  555 :  32 - 0x20
      10'h22C: dout  = 8'b00100000; //  556 :  32 - 0x20
      10'h22D: dout  = 8'b00100000; //  557 :  32 - 0x20
      10'h22E: dout  = 8'b00100000; //  558 :  32 - 0x20
      10'h22F: dout  = 8'b00100000; //  559 :  32 - 0x20
      10'h230: dout  = 8'b00100000; //  560 :  32 - 0x20
      10'h231: dout  = 8'b00100000; //  561 :  32 - 0x20
      10'h232: dout  = 8'b00100000; //  562 :  32 - 0x20
      10'h233: dout  = 8'b00100000; //  563 :  32 - 0x20
      10'h234: dout  = 8'b00100000; //  564 :  32 - 0x20
      10'h235: dout  = 8'b00100000; //  565 :  32 - 0x20
      10'h236: dout  = 8'b00100000; //  566 :  32 - 0x20
      10'h237: dout  = 8'b00100000; //  567 :  32 - 0x20
      10'h238: dout  = 8'b00100000; //  568 :  32 - 0x20
      10'h239: dout  = 8'b00100000; //  569 :  32 - 0x20
      10'h23A: dout  = 8'b00100000; //  570 :  32 - 0x20
      10'h23B: dout  = 8'b00100000; //  571 :  32 - 0x20
      10'h23C: dout  = 8'b00100000; //  572 :  32 - 0x20
      10'h23D: dout  = 8'b00100000; //  573 :  32 - 0x20
      10'h23E: dout  = 8'b00100000; //  574 :  32 - 0x20
      10'h23F: dout  = 8'b00100000; //  575 :  32 - 0x20
      10'h240: dout  = 8'b00100000; //  576 :  32 - 0x20 -- line 0x12
      10'h241: dout  = 8'b00100000; //  577 :  32 - 0x20
      10'h242: dout  = 8'b00100000; //  578 :  32 - 0x20
      10'h243: dout  = 8'b00100000; //  579 :  32 - 0x20
      10'h244: dout  = 8'b00100000; //  580 :  32 - 0x20
      10'h245: dout  = 8'b00100000; //  581 :  32 - 0x20
      10'h246: dout  = 8'b00100000; //  582 :  32 - 0x20
      10'h247: dout  = 8'b00100000; //  583 :  32 - 0x20
      10'h248: dout  = 8'b00100000; //  584 :  32 - 0x20
      10'h249: dout  = 8'b00100000; //  585 :  32 - 0x20
      10'h24A: dout  = 8'b00100000; //  586 :  32 - 0x20
      10'h24B: dout  = 8'b00100000; //  587 :  32 - 0x20
      10'h24C: dout  = 8'b00110010; //  588 :  50 - 0x32
      10'h24D: dout  = 8'b00100000; //  589 :  32 - 0x20
      10'h24E: dout  = 8'b01010000; //  590 :  80 - 0x50
      10'h24F: dout  = 8'b01001100; //  591 :  76 - 0x4c
      10'h250: dout  = 8'b01000001; //  592 :  65 - 0x41
      10'h251: dout  = 8'b01011001; //  593 :  89 - 0x59
      10'h252: dout  = 8'b01000101; //  594 :  69 - 0x45
      10'h253: dout  = 8'b01010010; //  595 :  82 - 0x52
      10'h254: dout  = 8'b01010011; //  596 :  83 - 0x53
      10'h255: dout  = 8'b00100000; //  597 :  32 - 0x20
      10'h256: dout  = 8'b00100000; //  598 :  32 - 0x20
      10'h257: dout  = 8'b00100000; //  599 :  32 - 0x20
      10'h258: dout  = 8'b00100000; //  600 :  32 - 0x20
      10'h259: dout  = 8'b00100000; //  601 :  32 - 0x20
      10'h25A: dout  = 8'b00100000; //  602 :  32 - 0x20
      10'h25B: dout  = 8'b00100000; //  603 :  32 - 0x20
      10'h25C: dout  = 8'b00100000; //  604 :  32 - 0x20
      10'h25D: dout  = 8'b00100000; //  605 :  32 - 0x20
      10'h25E: dout  = 8'b00100000; //  606 :  32 - 0x20
      10'h25F: dout  = 8'b00100000; //  607 :  32 - 0x20
      10'h260: dout  = 8'b00100000; //  608 :  32 - 0x20 -- line 0x13
      10'h261: dout  = 8'b00100000; //  609 :  32 - 0x20
      10'h262: dout  = 8'b00100000; //  610 :  32 - 0x20
      10'h263: dout  = 8'b00100000; //  611 :  32 - 0x20
      10'h264: dout  = 8'b00100000; //  612 :  32 - 0x20
      10'h265: dout  = 8'b00100000; //  613 :  32 - 0x20
      10'h266: dout  = 8'b00100000; //  614 :  32 - 0x20
      10'h267: dout  = 8'b00100000; //  615 :  32 - 0x20
      10'h268: dout  = 8'b00100000; //  616 :  32 - 0x20
      10'h269: dout  = 8'b00100000; //  617 :  32 - 0x20
      10'h26A: dout  = 8'b00100000; //  618 :  32 - 0x20
      10'h26B: dout  = 8'b00100000; //  619 :  32 - 0x20
      10'h26C: dout  = 8'b00100000; //  620 :  32 - 0x20
      10'h26D: dout  = 8'b00100000; //  621 :  32 - 0x20
      10'h26E: dout  = 8'b00100000; //  622 :  32 - 0x20
      10'h26F: dout  = 8'b00100000; //  623 :  32 - 0x20
      10'h270: dout  = 8'b00100000; //  624 :  32 - 0x20
      10'h271: dout  = 8'b00100000; //  625 :  32 - 0x20
      10'h272: dout  = 8'b00100000; //  626 :  32 - 0x20
      10'h273: dout  = 8'b00100000; //  627 :  32 - 0x20
      10'h274: dout  = 8'b00100000; //  628 :  32 - 0x20
      10'h275: dout  = 8'b00100000; //  629 :  32 - 0x20
      10'h276: dout  = 8'b00100000; //  630 :  32 - 0x20
      10'h277: dout  = 8'b00100000; //  631 :  32 - 0x20
      10'h278: dout  = 8'b00100000; //  632 :  32 - 0x20
      10'h279: dout  = 8'b00100000; //  633 :  32 - 0x20
      10'h27A: dout  = 8'b00100000; //  634 :  32 - 0x20
      10'h27B: dout  = 8'b00100000; //  635 :  32 - 0x20
      10'h27C: dout  = 8'b00100000; //  636 :  32 - 0x20
      10'h27D: dout  = 8'b00100000; //  637 :  32 - 0x20
      10'h27E: dout  = 8'b00100000; //  638 :  32 - 0x20
      10'h27F: dout  = 8'b00100000; //  639 :  32 - 0x20
      10'h280: dout  = 8'b00100000; //  640 :  32 - 0x20 -- line 0x14
      10'h281: dout  = 8'b00100000; //  641 :  32 - 0x20
      10'h282: dout  = 8'b00100000; //  642 :  32 - 0x20
      10'h283: dout  = 8'b00100000; //  643 :  32 - 0x20
      10'h284: dout  = 8'b00100000; //  644 :  32 - 0x20
      10'h285: dout  = 8'b00100000; //  645 :  32 - 0x20
      10'h286: dout  = 8'b00100000; //  646 :  32 - 0x20
      10'h287: dout  = 8'b00100000; //  647 :  32 - 0x20
      10'h288: dout  = 8'b00100000; //  648 :  32 - 0x20
      10'h289: dout  = 8'b00100000; //  649 :  32 - 0x20
      10'h28A: dout  = 8'b00100000; //  650 :  32 - 0x20
      10'h28B: dout  = 8'b00100000; //  651 :  32 - 0x20
      10'h28C: dout  = 8'b00100000; //  652 :  32 - 0x20
      10'h28D: dout  = 8'b00100000; //  653 :  32 - 0x20
      10'h28E: dout  = 8'b00100000; //  654 :  32 - 0x20
      10'h28F: dout  = 8'b00100000; //  655 :  32 - 0x20
      10'h290: dout  = 8'b00100000; //  656 :  32 - 0x20
      10'h291: dout  = 8'b00100000; //  657 :  32 - 0x20
      10'h292: dout  = 8'b00100000; //  658 :  32 - 0x20
      10'h293: dout  = 8'b00100000; //  659 :  32 - 0x20
      10'h294: dout  = 8'b00100000; //  660 :  32 - 0x20
      10'h295: dout  = 8'b00100000; //  661 :  32 - 0x20
      10'h296: dout  = 8'b00100000; //  662 :  32 - 0x20
      10'h297: dout  = 8'b00100000; //  663 :  32 - 0x20
      10'h298: dout  = 8'b00100000; //  664 :  32 - 0x20
      10'h299: dout  = 8'b00100000; //  665 :  32 - 0x20
      10'h29A: dout  = 8'b00100000; //  666 :  32 - 0x20
      10'h29B: dout  = 8'b00100000; //  667 :  32 - 0x20
      10'h29C: dout  = 8'b00100000; //  668 :  32 - 0x20
      10'h29D: dout  = 8'b00100000; //  669 :  32 - 0x20
      10'h29E: dout  = 8'b00100000; //  670 :  32 - 0x20
      10'h29F: dout  = 8'b00100000; //  671 :  32 - 0x20
      10'h2A0: dout  = 8'b00100000; //  672 :  32 - 0x20 -- line 0x15
      10'h2A1: dout  = 8'b00100000; //  673 :  32 - 0x20
      10'h2A2: dout  = 8'b01010100; //  674 :  84 - 0x54
      10'h2A3: dout  = 8'b01001101; //  675 :  77 - 0x4d
      10'h2A4: dout  = 8'b00100000; //  676 :  32 - 0x20
      10'h2A5: dout  = 8'b01000001; //  677 :  65 - 0x41
      10'h2A6: dout  = 8'b01001110; //  678 :  78 - 0x4e
      10'h2A7: dout  = 8'b01000100; //  679 :  68 - 0x44
      10'h2A8: dout  = 8'b00100000; //  680 :  32 - 0x20
      10'h2A9: dout  = 8'b01011101; //  681 :  93 - 0x5d
      10'h2AA: dout  = 8'b00100000; //  682 :  32 - 0x20
      10'h2AB: dout  = 8'b00110001; //  683 :  49 - 0x31
      10'h2AC: dout  = 8'b00111001; //  684 :  57 - 0x39
      10'h2AD: dout  = 8'b00111000; //  685 :  56 - 0x38
      10'h2AE: dout  = 8'b00110000; //  686 :  48 - 0x30
      10'h2AF: dout  = 8'b00100000; //  687 :  32 - 0x20
      10'h2B0: dout  = 8'b00110001; //  688 :  49 - 0x31
      10'h2B1: dout  = 8'b00111001; //  689 :  57 - 0x39
      10'h2B2: dout  = 8'b00111000; //  690 :  56 - 0x38
      10'h2B3: dout  = 8'b00110100; //  691 :  52 - 0x34
      10'h2B4: dout  = 8'b00100000; //  692 :  32 - 0x20
      10'h2B5: dout  = 8'b01001110; //  693 :  78 - 0x4e
      10'h2B6: dout  = 8'b01000001; //  694 :  65 - 0x41
      10'h2B7: dout  = 8'b01001101; //  695 :  77 - 0x4d
      10'h2B8: dout  = 8'b01000011; //  696 :  67 - 0x43
      10'h2B9: dout  = 8'b01001111; //  697 :  79 - 0x4f
      10'h2BA: dout  = 8'b00100000; //  698 :  32 - 0x20
      10'h2BB: dout  = 8'b01001100; //  699 :  76 - 0x4c
      10'h2BC: dout  = 8'b01010100; //  700 :  84 - 0x54
      10'h2BD: dout  = 8'b01000100; //  701 :  68 - 0x44
      10'h2BE: dout  = 8'b01011011; //  702 :  91 - 0x5b
      10'h2BF: dout  = 8'b00100000; //  703 :  32 - 0x20
      10'h2C0: dout  = 8'b00100000; //  704 :  32 - 0x20 -- line 0x16
      10'h2C1: dout  = 8'b00100000; //  705 :  32 - 0x20
      10'h2C2: dout  = 8'b00100000; //  706 :  32 - 0x20
      10'h2C3: dout  = 8'b00100000; //  707 :  32 - 0x20
      10'h2C4: dout  = 8'b00100000; //  708 :  32 - 0x20
      10'h2C5: dout  = 8'b00100000; //  709 :  32 - 0x20
      10'h2C6: dout  = 8'b00100000; //  710 :  32 - 0x20
      10'h2C7: dout  = 8'b00100000; //  711 :  32 - 0x20
      10'h2C8: dout  = 8'b00100000; //  712 :  32 - 0x20
      10'h2C9: dout  = 8'b00100000; //  713 :  32 - 0x20
      10'h2CA: dout  = 8'b00100000; //  714 :  32 - 0x20
      10'h2CB: dout  = 8'b00100000; //  715 :  32 - 0x20
      10'h2CC: dout  = 8'b00100000; //  716 :  32 - 0x20
      10'h2CD: dout  = 8'b00100000; //  717 :  32 - 0x20
      10'h2CE: dout  = 8'b00100000; //  718 :  32 - 0x20
      10'h2CF: dout  = 8'b00100000; //  719 :  32 - 0x20
      10'h2D0: dout  = 8'b00100000; //  720 :  32 - 0x20
      10'h2D1: dout  = 8'b00100000; //  721 :  32 - 0x20
      10'h2D2: dout  = 8'b00100000; //  722 :  32 - 0x20
      10'h2D3: dout  = 8'b00100000; //  723 :  32 - 0x20
      10'h2D4: dout  = 8'b00100000; //  724 :  32 - 0x20
      10'h2D5: dout  = 8'b00100000; //  725 :  32 - 0x20
      10'h2D6: dout  = 8'b00100000; //  726 :  32 - 0x20
      10'h2D7: dout  = 8'b00100000; //  727 :  32 - 0x20
      10'h2D8: dout  = 8'b00100000; //  728 :  32 - 0x20
      10'h2D9: dout  = 8'b00100000; //  729 :  32 - 0x20
      10'h2DA: dout  = 8'b00100000; //  730 :  32 - 0x20
      10'h2DB: dout  = 8'b00100000; //  731 :  32 - 0x20
      10'h2DC: dout  = 8'b00100000; //  732 :  32 - 0x20
      10'h2DD: dout  = 8'b00100000; //  733 :  32 - 0x20
      10'h2DE: dout  = 8'b00100000; //  734 :  32 - 0x20
      10'h2DF: dout  = 8'b00100000; //  735 :  32 - 0x20
      10'h2E0: dout  = 8'b00100000; //  736 :  32 - 0x20 -- line 0x17
      10'h2E1: dout  = 8'b00100000; //  737 :  32 - 0x20
      10'h2E2: dout  = 8'b00100000; //  738 :  32 - 0x20
      10'h2E3: dout  = 8'b00100000; //  739 :  32 - 0x20
      10'h2E4: dout  = 8'b00100000; //  740 :  32 - 0x20
      10'h2E5: dout  = 8'b00100000; //  741 :  32 - 0x20
      10'h2E6: dout  = 8'b00100000; //  742 :  32 - 0x20
      10'h2E7: dout  = 8'b00100000; //  743 :  32 - 0x20
      10'h2E8: dout  = 8'b00100000; //  744 :  32 - 0x20
      10'h2E9: dout  = 8'b00100000; //  745 :  32 - 0x20
      10'h2EA: dout  = 8'b00100000; //  746 :  32 - 0x20
      10'h2EB: dout  = 8'b00100000; //  747 :  32 - 0x20
      10'h2EC: dout  = 8'b00100000; //  748 :  32 - 0x20
      10'h2ED: dout  = 8'b01010100; //  749 :  84 - 0x54
      10'h2EE: dout  = 8'b01000101; //  750 :  69 - 0x45
      10'h2EF: dout  = 8'b01001110; //  751 :  78 - 0x4e
      10'h2F0: dout  = 8'b01000111; //  752 :  71 - 0x47
      10'h2F1: dout  = 8'b01000101; //  753 :  69 - 0x45
      10'h2F2: dout  = 8'b01001110; //  754 :  78 - 0x4e
      10'h2F3: dout  = 8'b00100000; //  755 :  32 - 0x20
      10'h2F4: dout  = 8'b00100000; //  756 :  32 - 0x20
      10'h2F5: dout  = 8'b00100000; //  757 :  32 - 0x20
      10'h2F6: dout  = 8'b00100000; //  758 :  32 - 0x20
      10'h2F7: dout  = 8'b00100000; //  759 :  32 - 0x20
      10'h2F8: dout  = 8'b00100000; //  760 :  32 - 0x20
      10'h2F9: dout  = 8'b00100000; //  761 :  32 - 0x20
      10'h2FA: dout  = 8'b00100000; //  762 :  32 - 0x20
      10'h2FB: dout  = 8'b00100000; //  763 :  32 - 0x20
      10'h2FC: dout  = 8'b00100000; //  764 :  32 - 0x20
      10'h2FD: dout  = 8'b00100000; //  765 :  32 - 0x20
      10'h2FE: dout  = 8'b00100000; //  766 :  32 - 0x20
      10'h2FF: dout  = 8'b00100000; //  767 :  32 - 0x20
      10'h300: dout  = 8'b00100000; //  768 :  32 - 0x20 -- line 0x18
      10'h301: dout  = 8'b00100000; //  769 :  32 - 0x20
      10'h302: dout  = 8'b00100000; //  770 :  32 - 0x20
      10'h303: dout  = 8'b00100000; //  771 :  32 - 0x20
      10'h304: dout  = 8'b00100000; //  772 :  32 - 0x20
      10'h305: dout  = 8'b00100000; //  773 :  32 - 0x20
      10'h306: dout  = 8'b00100000; //  774 :  32 - 0x20
      10'h307: dout  = 8'b00100000; //  775 :  32 - 0x20
      10'h308: dout  = 8'b00100000; //  776 :  32 - 0x20
      10'h309: dout  = 8'b00100000; //  777 :  32 - 0x20
      10'h30A: dout  = 8'b00100000; //  778 :  32 - 0x20
      10'h30B: dout  = 8'b00100000; //  779 :  32 - 0x20
      10'h30C: dout  = 8'b00100000; //  780 :  32 - 0x20
      10'h30D: dout  = 8'b00100000; //  781 :  32 - 0x20
      10'h30E: dout  = 8'b00100000; //  782 :  32 - 0x20
      10'h30F: dout  = 8'b00100000; //  783 :  32 - 0x20
      10'h310: dout  = 8'b00100000; //  784 :  32 - 0x20
      10'h311: dout  = 8'b00100000; //  785 :  32 - 0x20
      10'h312: dout  = 8'b00100000; //  786 :  32 - 0x20
      10'h313: dout  = 8'b00100000; //  787 :  32 - 0x20
      10'h314: dout  = 8'b00100000; //  788 :  32 - 0x20
      10'h315: dout  = 8'b00100000; //  789 :  32 - 0x20
      10'h316: dout  = 8'b00100000; //  790 :  32 - 0x20
      10'h317: dout  = 8'b00100000; //  791 :  32 - 0x20
      10'h318: dout  = 8'b00100000; //  792 :  32 - 0x20
      10'h319: dout  = 8'b00100000; //  793 :  32 - 0x20
      10'h31A: dout  = 8'b00100000; //  794 :  32 - 0x20
      10'h31B: dout  = 8'b00100000; //  795 :  32 - 0x20
      10'h31C: dout  = 8'b00100000; //  796 :  32 - 0x20
      10'h31D: dout  = 8'b00100000; //  797 :  32 - 0x20
      10'h31E: dout  = 8'b00100000; //  798 :  32 - 0x20
      10'h31F: dout  = 8'b00100000; //  799 :  32 - 0x20
      10'h320: dout  = 8'b00100000; //  800 :  32 - 0x20 -- line 0x19
      10'h321: dout  = 8'b00100000; //  801 :  32 - 0x20
      10'h322: dout  = 8'b00100000; //  802 :  32 - 0x20
      10'h323: dout  = 8'b00100000; //  803 :  32 - 0x20
      10'h324: dout  = 8'b00100000; //  804 :  32 - 0x20
      10'h325: dout  = 8'b00100000; //  805 :  32 - 0x20
      10'h326: dout  = 8'b00100000; //  806 :  32 - 0x20
      10'h327: dout  = 8'b00100000; //  807 :  32 - 0x20
      10'h328: dout  = 8'b00100000; //  808 :  32 - 0x20
      10'h329: dout  = 8'b00100000; //  809 :  32 - 0x20
      10'h32A: dout  = 8'b00100000; //  810 :  32 - 0x20
      10'h32B: dout  = 8'b00100000; //  811 :  32 - 0x20
      10'h32C: dout  = 8'b00100000; //  812 :  32 - 0x20
      10'h32D: dout  = 8'b00100000; //  813 :  32 - 0x20
      10'h32E: dout  = 8'b00100000; //  814 :  32 - 0x20
      10'h32F: dout  = 8'b00100000; //  815 :  32 - 0x20
      10'h330: dout  = 8'b00100000; //  816 :  32 - 0x20
      10'h331: dout  = 8'b00100000; //  817 :  32 - 0x20
      10'h332: dout  = 8'b00100000; //  818 :  32 - 0x20
      10'h333: dout  = 8'b00100000; //  819 :  32 - 0x20
      10'h334: dout  = 8'b00100000; //  820 :  32 - 0x20
      10'h335: dout  = 8'b00100000; //  821 :  32 - 0x20
      10'h336: dout  = 8'b00100000; //  822 :  32 - 0x20
      10'h337: dout  = 8'b00100000; //  823 :  32 - 0x20
      10'h338: dout  = 8'b00100000; //  824 :  32 - 0x20
      10'h339: dout  = 8'b00100000; //  825 :  32 - 0x20
      10'h33A: dout  = 8'b00100000; //  826 :  32 - 0x20
      10'h33B: dout  = 8'b00100000; //  827 :  32 - 0x20
      10'h33C: dout  = 8'b00100000; //  828 :  32 - 0x20
      10'h33D: dout  = 8'b00100000; //  829 :  32 - 0x20
      10'h33E: dout  = 8'b00100000; //  830 :  32 - 0x20
      10'h33F: dout  = 8'b00100000; //  831 :  32 - 0x20
      10'h340: dout  = 8'b00100000; //  832 :  32 - 0x20 -- line 0x1a
      10'h341: dout  = 8'b00100000; //  833 :  32 - 0x20
      10'h342: dout  = 8'b00100000; //  834 :  32 - 0x20
      10'h343: dout  = 8'b00100000; //  835 :  32 - 0x20
      10'h344: dout  = 8'b00100000; //  836 :  32 - 0x20
      10'h345: dout  = 8'b00100000; //  837 :  32 - 0x20
      10'h346: dout  = 8'b00100000; //  838 :  32 - 0x20
      10'h347: dout  = 8'b00100000; //  839 :  32 - 0x20
      10'h348: dout  = 8'b00100000; //  840 :  32 - 0x20
      10'h349: dout  = 8'b00100000; //  841 :  32 - 0x20
      10'h34A: dout  = 8'b00100000; //  842 :  32 - 0x20
      10'h34B: dout  = 8'b00100000; //  843 :  32 - 0x20
      10'h34C: dout  = 8'b00100000; //  844 :  32 - 0x20
      10'h34D: dout  = 8'b00100000; //  845 :  32 - 0x20
      10'h34E: dout  = 8'b00100000; //  846 :  32 - 0x20
      10'h34F: dout  = 8'b00100000; //  847 :  32 - 0x20
      10'h350: dout  = 8'b00100000; //  848 :  32 - 0x20
      10'h351: dout  = 8'b00100000; //  849 :  32 - 0x20
      10'h352: dout  = 8'b00100000; //  850 :  32 - 0x20
      10'h353: dout  = 8'b00100000; //  851 :  32 - 0x20
      10'h354: dout  = 8'b00100000; //  852 :  32 - 0x20
      10'h355: dout  = 8'b00100000; //  853 :  32 - 0x20
      10'h356: dout  = 8'b00100000; //  854 :  32 - 0x20
      10'h357: dout  = 8'b00100000; //  855 :  32 - 0x20
      10'h358: dout  = 8'b00100000; //  856 :  32 - 0x20
      10'h359: dout  = 8'b00100000; //  857 :  32 - 0x20
      10'h35A: dout  = 8'b00100000; //  858 :  32 - 0x20
      10'h35B: dout  = 8'b00100000; //  859 :  32 - 0x20
      10'h35C: dout  = 8'b00100000; //  860 :  32 - 0x20
      10'h35D: dout  = 8'b00100000; //  861 :  32 - 0x20
      10'h35E: dout  = 8'b00100000; //  862 :  32 - 0x20
      10'h35F: dout  = 8'b00100000; //  863 :  32 - 0x20
      10'h360: dout  = 8'b00100000; //  864 :  32 - 0x20 -- line 0x1b
      10'h361: dout  = 8'b00100000; //  865 :  32 - 0x20
      10'h362: dout  = 8'b00100000; //  866 :  32 - 0x20
      10'h363: dout  = 8'b00100000; //  867 :  32 - 0x20
      10'h364: dout  = 8'b00100000; //  868 :  32 - 0x20
      10'h365: dout  = 8'b00100000; //  869 :  32 - 0x20
      10'h366: dout  = 8'b00100000; //  870 :  32 - 0x20
      10'h367: dout  = 8'b00100000; //  871 :  32 - 0x20
      10'h368: dout  = 8'b00100000; //  872 :  32 - 0x20
      10'h369: dout  = 8'b00100000; //  873 :  32 - 0x20
      10'h36A: dout  = 8'b00100000; //  874 :  32 - 0x20
      10'h36B: dout  = 8'b00100000; //  875 :  32 - 0x20
      10'h36C: dout  = 8'b00100000; //  876 :  32 - 0x20
      10'h36D: dout  = 8'b00100000; //  877 :  32 - 0x20
      10'h36E: dout  = 8'b00100000; //  878 :  32 - 0x20
      10'h36F: dout  = 8'b00100000; //  879 :  32 - 0x20
      10'h370: dout  = 8'b00100000; //  880 :  32 - 0x20
      10'h371: dout  = 8'b00100000; //  881 :  32 - 0x20
      10'h372: dout  = 8'b00100000; //  882 :  32 - 0x20
      10'h373: dout  = 8'b00100000; //  883 :  32 - 0x20
      10'h374: dout  = 8'b00100000; //  884 :  32 - 0x20
      10'h375: dout  = 8'b00100000; //  885 :  32 - 0x20
      10'h376: dout  = 8'b00100000; //  886 :  32 - 0x20
      10'h377: dout  = 8'b00100000; //  887 :  32 - 0x20
      10'h378: dout  = 8'b00100000; //  888 :  32 - 0x20
      10'h379: dout  = 8'b00100000; //  889 :  32 - 0x20
      10'h37A: dout  = 8'b00100000; //  890 :  32 - 0x20
      10'h37B: dout  = 8'b00100000; //  891 :  32 - 0x20
      10'h37C: dout  = 8'b00100000; //  892 :  32 - 0x20
      10'h37D: dout  = 8'b00100000; //  893 :  32 - 0x20
      10'h37E: dout  = 8'b00100000; //  894 :  32 - 0x20
      10'h37F: dout  = 8'b00100000; //  895 :  32 - 0x20
      10'h380: dout  = 8'b00100000; //  896 :  32 - 0x20 -- line 0x1c
      10'h381: dout  = 8'b00100000; //  897 :  32 - 0x20
      10'h382: dout  = 8'b00100000; //  898 :  32 - 0x20
      10'h383: dout  = 8'b00100000; //  899 :  32 - 0x20
      10'h384: dout  = 8'b00100000; //  900 :  32 - 0x20
      10'h385: dout  = 8'b00100000; //  901 :  32 - 0x20
      10'h386: dout  = 8'b00100000; //  902 :  32 - 0x20
      10'h387: dout  = 8'b00100000; //  903 :  32 - 0x20
      10'h388: dout  = 8'b00100000; //  904 :  32 - 0x20
      10'h389: dout  = 8'b00100000; //  905 :  32 - 0x20
      10'h38A: dout  = 8'b00100000; //  906 :  32 - 0x20
      10'h38B: dout  = 8'b00100000; //  907 :  32 - 0x20
      10'h38C: dout  = 8'b00100000; //  908 :  32 - 0x20
      10'h38D: dout  = 8'b00100000; //  909 :  32 - 0x20
      10'h38E: dout  = 8'b00100000; //  910 :  32 - 0x20
      10'h38F: dout  = 8'b00100000; //  911 :  32 - 0x20
      10'h390: dout  = 8'b00100000; //  912 :  32 - 0x20
      10'h391: dout  = 8'b00100000; //  913 :  32 - 0x20
      10'h392: dout  = 8'b00100000; //  914 :  32 - 0x20
      10'h393: dout  = 8'b00100000; //  915 :  32 - 0x20
      10'h394: dout  = 8'b00100000; //  916 :  32 - 0x20
      10'h395: dout  = 8'b00100000; //  917 :  32 - 0x20
      10'h396: dout  = 8'b00100000; //  918 :  32 - 0x20
      10'h397: dout  = 8'b00100000; //  919 :  32 - 0x20
      10'h398: dout  = 8'b00100000; //  920 :  32 - 0x20
      10'h399: dout  = 8'b00100000; //  921 :  32 - 0x20
      10'h39A: dout  = 8'b00100000; //  922 :  32 - 0x20
      10'h39B: dout  = 8'b00100000; //  923 :  32 - 0x20
      10'h39C: dout  = 8'b00100000; //  924 :  32 - 0x20
      10'h39D: dout  = 8'b00100000; //  925 :  32 - 0x20
      10'h39E: dout  = 8'b00100000; //  926 :  32 - 0x20
      10'h39F: dout  = 8'b00100000; //  927 :  32 - 0x20
      10'h3A0: dout  = 8'b00100000; //  928 :  32 - 0x20 -- line 0x1d
      10'h3A1: dout  = 8'b00100000; //  929 :  32 - 0x20
      10'h3A2: dout  = 8'b00100000; //  930 :  32 - 0x20
      10'h3A3: dout  = 8'b00100000; //  931 :  32 - 0x20
      10'h3A4: dout  = 8'b00100000; //  932 :  32 - 0x20
      10'h3A5: dout  = 8'b00100000; //  933 :  32 - 0x20
      10'h3A6: dout  = 8'b00100000; //  934 :  32 - 0x20
      10'h3A7: dout  = 8'b00100000; //  935 :  32 - 0x20
      10'h3A8: dout  = 8'b00100000; //  936 :  32 - 0x20
      10'h3A9: dout  = 8'b00100000; //  937 :  32 - 0x20
      10'h3AA: dout  = 8'b00100000; //  938 :  32 - 0x20
      10'h3AB: dout  = 8'b00100000; //  939 :  32 - 0x20
      10'h3AC: dout  = 8'b00100000; //  940 :  32 - 0x20
      10'h3AD: dout  = 8'b00100000; //  941 :  32 - 0x20
      10'h3AE: dout  = 8'b00100000; //  942 :  32 - 0x20
      10'h3AF: dout  = 8'b00100000; //  943 :  32 - 0x20
      10'h3B0: dout  = 8'b00100000; //  944 :  32 - 0x20
      10'h3B1: dout  = 8'b00100000; //  945 :  32 - 0x20
      10'h3B2: dout  = 8'b00100000; //  946 :  32 - 0x20
      10'h3B3: dout  = 8'b00100000; //  947 :  32 - 0x20
      10'h3B4: dout  = 8'b00100000; //  948 :  32 - 0x20
      10'h3B5: dout  = 8'b00100000; //  949 :  32 - 0x20
      10'h3B6: dout  = 8'b00100000; //  950 :  32 - 0x20
      10'h3B7: dout  = 8'b00100000; //  951 :  32 - 0x20
      10'h3B8: dout  = 8'b00100000; //  952 :  32 - 0x20
      10'h3B9: dout  = 8'b00100000; //  953 :  32 - 0x20
      10'h3BA: dout  = 8'b00100000; //  954 :  32 - 0x20
      10'h3BB: dout  = 8'b00100000; //  955 :  32 - 0x20
      10'h3BC: dout  = 8'b00100000; //  956 :  32 - 0x20
      10'h3BD: dout  = 8'b00100000; //  957 :  32 - 0x20
      10'h3BE: dout  = 8'b00100000; //  958 :  32 - 0x20
      10'h3BF: dout  = 8'b00100000; //  959 :  32 - 0x20
        //-- Attribute Table 0----
      10'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0
      10'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      10'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      10'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      10'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      10'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      10'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      10'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      10'h3C8: dout  = 8'b10000000; //  968 : 128 - 0x80
      10'h3C9: dout  = 8'b10100000; //  969 : 160 - 0xa0
      10'h3CA: dout  = 8'b10100000; //  970 : 160 - 0xa0
      10'h3CB: dout  = 8'b10100000; //  971 : 160 - 0xa0
      10'h3CC: dout  = 8'b10100000; //  972 : 160 - 0xa0
      10'h3CD: dout  = 8'b10100000; //  973 : 160 - 0xa0
      10'h3CE: dout  = 8'b10100000; //  974 : 160 - 0xa0
      10'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      10'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0
      10'h3D1: dout  = 8'b01100110; //  977 : 102 - 0x66
      10'h3D2: dout  = 8'b01010101; //  978 :  85 - 0x55
      10'h3D3: dout  = 8'b01010101; //  979 :  85 - 0x55
      10'h3D4: dout  = 8'b01010101; //  980 :  85 - 0x55
      10'h3D5: dout  = 8'b01010101; //  981 :  85 - 0x55
      10'h3D6: dout  = 8'b11011101; //  982 : 221 - 0xdd
      10'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      10'h3D8: dout  = 8'b00001000; //  984 :   8 - 0x8
      10'h3D9: dout  = 8'b00001010; //  985 :  10 - 0xa
      10'h3DA: dout  = 8'b00001010; //  986 :  10 - 0xa
      10'h3DB: dout  = 8'b00001010; //  987 :  10 - 0xa
      10'h3DC: dout  = 8'b00001010; //  988 :  10 - 0xa
      10'h3DD: dout  = 8'b00001010; //  989 :  10 - 0xa
      10'h3DE: dout  = 8'b00001010; //  990 :  10 - 0xa
      10'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      10'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0
      10'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      10'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      10'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      10'h3E4: dout  = 8'b00000000; //  996 :   0 - 0x0
      10'h3E5: dout  = 8'b00000000; //  997 :   0 - 0x0
      10'h3E6: dout  = 8'b00000000; //  998 :   0 - 0x0
      10'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      10'h3E8: dout  = 8'b11110000; // 1000 : 240 - 0xf0
      10'h3E9: dout  = 8'b11110000; // 1001 : 240 - 0xf0
      10'h3EA: dout  = 8'b11110000; // 1002 : 240 - 0xf0
      10'h3EB: dout  = 8'b11110000; // 1003 : 240 - 0xf0
      10'h3EC: dout  = 8'b11110000; // 1004 : 240 - 0xf0
      10'h3ED: dout  = 8'b11110000; // 1005 : 240 - 0xf0
      10'h3EE: dout  = 8'b11110000; // 1006 : 240 - 0xf0
      10'h3EF: dout  = 8'b11110000; // 1007 : 240 - 0xf0
      10'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0
      10'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      10'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      10'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      10'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      10'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      10'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      10'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      10'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0
      10'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      10'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      10'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      10'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      10'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      10'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      10'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
    endcase
  end

endmodule
